magic
tech sky130A
magscale 1 2
timestamp 1666360185
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 427998 1006816 428004 1006868
rect 428056 1006856 428062 1006868
rect 428056 1006828 441614 1006856
rect 428056 1006816 428062 1006828
rect 428366 1006680 428372 1006732
rect 428424 1006720 428430 1006732
rect 434438 1006720 434444 1006732
rect 428424 1006692 434444 1006720
rect 428424 1006680 428430 1006692
rect 434438 1006680 434444 1006692
rect 434496 1006680 434502 1006732
rect 357710 1006612 357716 1006664
rect 357768 1006652 357774 1006664
rect 371878 1006652 371884 1006664
rect 357768 1006624 371884 1006652
rect 357768 1006612 357774 1006624
rect 371878 1006612 371884 1006624
rect 371936 1006612 371942 1006664
rect 145558 1006544 145564 1006596
rect 145616 1006584 145622 1006596
rect 152918 1006584 152924 1006596
rect 145616 1006556 152924 1006584
rect 145616 1006544 145622 1006556
rect 152918 1006544 152924 1006556
rect 152976 1006544 152982 1006596
rect 300118 1006544 300124 1006596
rect 300176 1006584 300182 1006596
rect 308122 1006584 308128 1006596
rect 300176 1006556 308128 1006584
rect 300176 1006544 300182 1006556
rect 308122 1006544 308128 1006556
rect 308180 1006544 308186 1006596
rect 359734 1006476 359740 1006528
rect 359792 1006516 359798 1006528
rect 370498 1006516 370504 1006528
rect 359792 1006488 370504 1006516
rect 359792 1006476 359798 1006488
rect 370498 1006476 370504 1006488
rect 370556 1006476 370562 1006528
rect 422662 1006476 422668 1006528
rect 422720 1006516 422726 1006528
rect 426526 1006516 426532 1006528
rect 422720 1006488 426532 1006516
rect 422720 1006476 422726 1006488
rect 426526 1006476 426532 1006488
rect 426584 1006476 426590 1006528
rect 94498 1006408 94504 1006460
rect 94556 1006448 94562 1006460
rect 103974 1006448 103980 1006460
rect 94556 1006420 103980 1006448
rect 94556 1006408 94562 1006420
rect 103974 1006408 103980 1006420
rect 104032 1006408 104038 1006460
rect 145742 1006408 145748 1006460
rect 145800 1006448 145806 1006460
rect 152090 1006448 152096 1006460
rect 145800 1006420 152096 1006448
rect 145800 1006408 145806 1006420
rect 152090 1006408 152096 1006420
rect 152148 1006408 152154 1006460
rect 157426 1006408 157432 1006460
rect 157484 1006448 157490 1006460
rect 166258 1006448 166264 1006460
rect 157484 1006420 166264 1006448
rect 157484 1006408 157490 1006420
rect 166258 1006408 166264 1006420
rect 166316 1006408 166322 1006460
rect 171778 1006448 171784 1006460
rect 171106 1006420 171784 1006448
rect 94682 1006272 94688 1006324
rect 94740 1006312 94746 1006324
rect 101122 1006312 101128 1006324
rect 94740 1006284 101128 1006312
rect 94740 1006272 94746 1006284
rect 101122 1006272 101128 1006284
rect 101180 1006272 101186 1006324
rect 144270 1006272 144276 1006324
rect 144328 1006312 144334 1006324
rect 144328 1006284 151814 1006312
rect 144328 1006272 144334 1006284
rect 93302 1006136 93308 1006188
rect 93360 1006176 93366 1006188
rect 98270 1006176 98276 1006188
rect 93360 1006148 98276 1006176
rect 93360 1006136 93366 1006148
rect 98270 1006136 98276 1006148
rect 98328 1006136 98334 1006188
rect 107654 1006136 107660 1006188
rect 107712 1006176 107718 1006188
rect 124858 1006176 124864 1006188
rect 107712 1006148 124864 1006176
rect 107712 1006136 107718 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 144086 1006136 144092 1006188
rect 144144 1006176 144150 1006188
rect 151262 1006176 151268 1006188
rect 144144 1006148 151268 1006176
rect 144144 1006136 144150 1006148
rect 151262 1006136 151268 1006148
rect 151320 1006136 151326 1006188
rect 151786 1006176 151814 1006284
rect 158254 1006272 158260 1006324
rect 158312 1006312 158318 1006324
rect 171106 1006312 171134 1006420
rect 171778 1006408 171784 1006420
rect 171836 1006408 171842 1006460
rect 431678 1006408 431684 1006460
rect 431736 1006448 431742 1006460
rect 431736 1006420 436784 1006448
rect 431736 1006408 431742 1006420
rect 425330 1006340 425336 1006392
rect 425388 1006380 425394 1006392
rect 425388 1006352 429424 1006380
rect 425388 1006340 425394 1006352
rect 158312 1006284 171134 1006312
rect 158312 1006272 158318 1006284
rect 204898 1006272 204904 1006324
rect 204956 1006312 204962 1006324
rect 210050 1006312 210056 1006324
rect 204956 1006284 210056 1006312
rect 204956 1006272 204962 1006284
rect 210050 1006272 210056 1006284
rect 210108 1006272 210114 1006324
rect 249242 1006272 249248 1006324
rect 249300 1006312 249306 1006324
rect 254118 1006312 254124 1006324
rect 249300 1006284 254124 1006312
rect 249300 1006272 249306 1006284
rect 254118 1006272 254124 1006284
rect 254176 1006272 254182 1006324
rect 298922 1006272 298928 1006324
rect 298980 1006312 298986 1006324
rect 311802 1006312 311808 1006324
rect 298980 1006284 311808 1006312
rect 298980 1006272 298986 1006284
rect 311802 1006272 311808 1006284
rect 311860 1006272 311866 1006324
rect 358538 1006272 358544 1006324
rect 358596 1006312 358602 1006324
rect 377398 1006312 377404 1006324
rect 358596 1006284 377404 1006312
rect 358596 1006272 358602 1006284
rect 377398 1006272 377404 1006284
rect 377456 1006272 377462 1006324
rect 429396 1006244 429424 1006352
rect 431678 1006244 431684 1006256
rect 429396 1006216 431684 1006244
rect 431678 1006204 431684 1006216
rect 431736 1006204 431742 1006256
rect 153746 1006176 153752 1006188
rect 151786 1006148 153752 1006176
rect 153746 1006136 153752 1006148
rect 153804 1006136 153810 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 164878 1006176 164884 1006188
rect 160336 1006148 164884 1006176
rect 160336 1006136 160342 1006148
rect 164878 1006136 164884 1006148
rect 164936 1006136 164942 1006188
rect 166258 1006136 166264 1006188
rect 166316 1006176 166322 1006188
rect 175918 1006176 175924 1006188
rect 166316 1006148 175924 1006176
rect 166316 1006136 166322 1006148
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 210418 1006136 210424 1006188
rect 210476 1006176 210482 1006188
rect 228358 1006176 228364 1006188
rect 210476 1006148 228364 1006176
rect 210476 1006136 210482 1006148
rect 228358 1006136 228364 1006148
rect 228416 1006136 228422 1006188
rect 247034 1006136 247040 1006188
rect 247092 1006176 247098 1006188
rect 255314 1006176 255320 1006188
rect 247092 1006148 255320 1006176
rect 247092 1006136 247098 1006148
rect 255314 1006136 255320 1006148
rect 255372 1006136 255378 1006188
rect 261846 1006136 261852 1006188
rect 261904 1006176 261910 1006188
rect 279418 1006176 279424 1006188
rect 261904 1006148 279424 1006176
rect 261904 1006136 261910 1006148
rect 279418 1006136 279424 1006148
rect 279476 1006136 279482 1006188
rect 299474 1006136 299480 1006188
rect 299532 1006176 299538 1006188
rect 306098 1006176 306104 1006188
rect 299532 1006148 306104 1006176
rect 299532 1006136 299538 1006148
rect 306098 1006136 306104 1006148
rect 306156 1006136 306162 1006188
rect 361390 1006136 361396 1006188
rect 361448 1006176 361454 1006188
rect 367002 1006176 367008 1006188
rect 361448 1006148 367008 1006176
rect 361448 1006136 361454 1006148
rect 367002 1006136 367008 1006148
rect 367060 1006136 367066 1006188
rect 402238 1006136 402244 1006188
rect 402296 1006176 402302 1006188
rect 429194 1006176 429200 1006188
rect 402296 1006148 429200 1006176
rect 402296 1006136 402302 1006148
rect 429194 1006136 429200 1006148
rect 429252 1006136 429258 1006188
rect 436756 1006176 436784 1006420
rect 441586 1006312 441614 1006828
rect 504542 1006816 504548 1006868
rect 504600 1006856 504606 1006868
rect 516962 1006856 516968 1006868
rect 504600 1006828 516968 1006856
rect 504600 1006816 504606 1006828
rect 516962 1006816 516968 1006828
rect 517020 1006816 517026 1006868
rect 556982 1006816 556988 1006868
rect 557040 1006856 557046 1006868
rect 559650 1006856 559656 1006868
rect 557040 1006828 559656 1006856
rect 557040 1006816 557046 1006828
rect 559650 1006816 559656 1006828
rect 559708 1006816 559714 1006868
rect 505370 1006680 505376 1006732
rect 505428 1006720 505434 1006732
rect 515398 1006720 515404 1006732
rect 505428 1006692 515404 1006720
rect 505428 1006680 505434 1006692
rect 515398 1006680 515404 1006692
rect 515456 1006680 515462 1006732
rect 554314 1006680 554320 1006732
rect 554372 1006720 554378 1006732
rect 562318 1006720 562324 1006732
rect 554372 1006692 562324 1006720
rect 554372 1006680 554378 1006692
rect 562318 1006680 562324 1006692
rect 562376 1006680 562382 1006732
rect 506198 1006408 506204 1006460
rect 506256 1006448 506262 1006460
rect 506256 1006420 509234 1006448
rect 506256 1006408 506262 1006420
rect 464982 1006312 464988 1006324
rect 441586 1006284 464988 1006312
rect 464982 1006272 464988 1006284
rect 465040 1006272 465046 1006324
rect 509206 1006312 509234 1006420
rect 555970 1006408 555976 1006460
rect 556028 1006448 556034 1006460
rect 566458 1006448 566464 1006460
rect 556028 1006420 566464 1006448
rect 556028 1006408 556034 1006420
rect 566458 1006408 566464 1006420
rect 566516 1006408 566522 1006460
rect 520918 1006312 520924 1006324
rect 509206 1006284 520924 1006312
rect 520918 1006272 520924 1006284
rect 520976 1006272 520982 1006324
rect 471238 1006176 471244 1006188
rect 436756 1006148 471244 1006176
rect 471238 1006136 471244 1006148
rect 471296 1006136 471302 1006188
rect 508222 1006136 508228 1006188
rect 508280 1006176 508286 1006188
rect 508280 1006148 518894 1006176
rect 508280 1006136 508286 1006148
rect 93118 1006000 93124 1006052
rect 93176 1006040 93182 1006052
rect 99466 1006040 99472 1006052
rect 93176 1006012 99472 1006040
rect 93176 1006000 93182 1006012
rect 99466 1006000 99472 1006012
rect 99524 1006000 99530 1006052
rect 102778 1006000 102784 1006052
rect 102836 1006040 102842 1006052
rect 104802 1006040 104808 1006052
rect 102836 1006012 104808 1006040
rect 102836 1006000 102842 1006012
rect 104802 1006000 104808 1006012
rect 104860 1006000 104866 1006052
rect 108482 1006000 108488 1006052
rect 108540 1006040 108546 1006052
rect 126238 1006040 126244 1006052
rect 108540 1006012 126244 1006040
rect 108540 1006000 108546 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 148870 1006000 148876 1006052
rect 148928 1006040 148934 1006052
rect 150066 1006040 150072 1006052
rect 148928 1006012 150072 1006040
rect 148928 1006000 148934 1006012
rect 150066 1006000 150072 1006012
rect 150124 1006000 150130 1006052
rect 159450 1006000 159456 1006052
rect 159508 1006040 159514 1006052
rect 177298 1006040 177304 1006052
rect 159508 1006012 177304 1006040
rect 159508 1006000 159514 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 198366 1006000 198372 1006052
rect 198424 1006040 198430 1006052
rect 201034 1006040 201040 1006052
rect 198424 1006012 201040 1006040
rect 198424 1006000 198430 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 208394 1006000 208400 1006052
rect 208452 1006040 208458 1006052
rect 229738 1006040 229744 1006052
rect 208452 1006012 229744 1006040
rect 208452 1006000 208458 1006012
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 251082 1006000 251088 1006052
rect 251140 1006040 251146 1006052
rect 252462 1006040 252468 1006052
rect 251140 1006012 252468 1006040
rect 251140 1006000 251146 1006012
rect 252462 1006000 252468 1006012
rect 252520 1006000 252526 1006052
rect 260190 1006000 260196 1006052
rect 260248 1006040 260254 1006052
rect 280798 1006040 280804 1006052
rect 260248 1006012 280804 1006040
rect 260248 1006000 260254 1006012
rect 280798 1006000 280804 1006012
rect 280856 1006000 280862 1006052
rect 298738 1006000 298744 1006052
rect 298796 1006040 298802 1006052
rect 298796 1006012 299474 1006040
rect 298796 1006000 298802 1006012
rect 299446 1005836 299474 1006012
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 319438 1006040 319444 1006052
rect 314712 1006012 319444 1006040
rect 314712 1006000 314718 1006012
rect 319438 1006000 319444 1006012
rect 319496 1006000 319502 1006052
rect 382918 1006040 382924 1006052
rect 364536 1006012 382924 1006040
rect 363414 1005932 363420 1005984
rect 363472 1005972 363478 1005984
rect 364536 1005972 364564 1006012
rect 382918 1006000 382924 1006012
rect 382976 1006000 382982 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 425330 1006040 425336 1006052
rect 400916 1006012 425336 1006040
rect 400916 1006000 400922 1006012
rect 425330 1006000 425336 1006012
rect 425388 1006000 425394 1006052
rect 425514 1006000 425520 1006052
rect 425572 1006040 425578 1006052
rect 429194 1006040 429200 1006052
rect 425572 1006012 429200 1006040
rect 425572 1006000 425578 1006012
rect 429194 1006000 429200 1006012
rect 429252 1006000 429258 1006052
rect 469858 1006040 469864 1006052
rect 431926 1006012 469864 1006040
rect 363472 1005944 364564 1005972
rect 363472 1005932 363478 1005944
rect 430850 1005932 430856 1005984
rect 430908 1005972 430914 1005984
rect 431926 1005972 431954 1006012
rect 469858 1006000 469864 1006012
rect 469916 1006000 469922 1006052
rect 498102 1006000 498108 1006052
rect 498160 1006040 498166 1006052
rect 498838 1006040 498844 1006052
rect 498160 1006012 498844 1006040
rect 498160 1006000 498166 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 509050 1006000 509056 1006052
rect 509108 1006040 509114 1006052
rect 518866 1006040 518894 1006148
rect 557166 1006136 557172 1006188
rect 557224 1006176 557230 1006188
rect 567838 1006176 567844 1006188
rect 557224 1006148 567844 1006176
rect 557224 1006136 557230 1006148
rect 567838 1006136 567844 1006148
rect 567896 1006136 567902 1006188
rect 522298 1006040 522304 1006052
rect 509108 1006012 509234 1006040
rect 518866 1006012 522304 1006040
rect 509108 1006000 509114 1006012
rect 430908 1005944 431954 1005972
rect 509206 1005972 509234 1006012
rect 522298 1006000 522304 1006012
rect 522356 1006000 522362 1006052
rect 549162 1006000 549168 1006052
rect 549220 1006040 549226 1006052
rect 550266 1006040 550272 1006052
rect 549220 1006012 550272 1006040
rect 549220 1006000 549226 1006012
rect 550266 1006000 550272 1006012
rect 550324 1006000 550330 1006052
rect 553946 1006000 553952 1006052
rect 554004 1006040 554010 1006052
rect 556154 1006040 556160 1006052
rect 554004 1006012 556160 1006040
rect 554004 1006000 554010 1006012
rect 556154 1006000 556160 1006012
rect 556212 1006000 556218 1006052
rect 562318 1006000 562324 1006052
rect 562376 1006040 562382 1006052
rect 573358 1006040 573364 1006052
rect 562376 1006012 573364 1006040
rect 562376 1006000 562382 1006012
rect 573358 1006000 573364 1006012
rect 573416 1006000 573422 1006052
rect 514018 1005972 514024 1005984
rect 509206 1005944 514024 1005972
rect 430908 1005932 430914 1005944
rect 514018 1005932 514024 1005944
rect 514076 1005932 514082 1005984
rect 304074 1005836 304080 1005848
rect 299446 1005808 304080 1005836
rect 304074 1005796 304080 1005808
rect 304132 1005796 304138 1005848
rect 426342 1005728 426348 1005780
rect 426400 1005768 426406 1005780
rect 440878 1005768 440884 1005780
rect 426400 1005740 440884 1005768
rect 426400 1005728 426406 1005740
rect 440878 1005728 440884 1005740
rect 440936 1005728 440942 1005780
rect 367002 1005660 367008 1005712
rect 367060 1005700 367066 1005712
rect 380158 1005700 380164 1005712
rect 367060 1005672 380164 1005700
rect 367060 1005660 367066 1005672
rect 380158 1005660 380164 1005672
rect 380216 1005660 380222 1005712
rect 360562 1005524 360568 1005576
rect 360620 1005564 360626 1005576
rect 378778 1005564 378784 1005576
rect 360620 1005536 378784 1005564
rect 360620 1005524 360626 1005536
rect 378778 1005524 378784 1005536
rect 378836 1005524 378842 1005576
rect 426342 1005524 426348 1005576
rect 426400 1005564 426406 1005576
rect 443638 1005564 443644 1005576
rect 426400 1005536 443644 1005564
rect 426400 1005524 426406 1005536
rect 443638 1005524 443644 1005536
rect 443696 1005524 443702 1005576
rect 556154 1005524 556160 1005576
rect 556212 1005564 556218 1005576
rect 570598 1005564 570604 1005576
rect 556212 1005536 570604 1005564
rect 556212 1005524 556218 1005536
rect 570598 1005524 570604 1005536
rect 570656 1005524 570662 1005576
rect 358538 1005388 358544 1005440
rect 358596 1005428 358602 1005440
rect 373258 1005428 373264 1005440
rect 358596 1005400 373264 1005428
rect 358596 1005388 358602 1005400
rect 373258 1005388 373264 1005400
rect 373316 1005388 373322 1005440
rect 430022 1005388 430028 1005440
rect 430080 1005428 430086 1005440
rect 431954 1005428 431960 1005440
rect 430080 1005400 431960 1005428
rect 430080 1005388 430086 1005400
rect 431954 1005388 431960 1005400
rect 432012 1005388 432018 1005440
rect 434438 1005388 434444 1005440
rect 434496 1005428 434502 1005440
rect 458818 1005428 458824 1005440
rect 434496 1005400 458824 1005428
rect 434496 1005388 434502 1005400
rect 458818 1005388 458824 1005400
rect 458876 1005388 458882 1005440
rect 502150 1005388 502156 1005440
rect 502208 1005428 502214 1005440
rect 518158 1005428 518164 1005440
rect 502208 1005400 518164 1005428
rect 502208 1005388 502214 1005400
rect 518158 1005388 518164 1005400
rect 518216 1005388 518222 1005440
rect 551462 1005388 551468 1005440
rect 551520 1005428 551526 1005440
rect 569218 1005428 569224 1005440
rect 551520 1005400 569224 1005428
rect 551520 1005388 551526 1005400
rect 569218 1005388 569224 1005400
rect 569276 1005388 569282 1005440
rect 354858 1005252 354864 1005304
rect 354916 1005292 354922 1005304
rect 374638 1005292 374644 1005304
rect 354916 1005264 374644 1005292
rect 354916 1005252 354922 1005264
rect 374638 1005252 374644 1005264
rect 374696 1005252 374702 1005304
rect 423490 1005252 423496 1005304
rect 423548 1005292 423554 1005304
rect 456058 1005292 456064 1005304
rect 423548 1005264 456064 1005292
rect 423548 1005252 423554 1005264
rect 456058 1005252 456064 1005264
rect 456116 1005252 456122 1005304
rect 499666 1005252 499672 1005304
rect 499724 1005292 499730 1005304
rect 516778 1005292 516784 1005304
rect 499724 1005264 516784 1005292
rect 499724 1005252 499730 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 574738 1005292 574744 1005304
rect 557506 1005264 574744 1005292
rect 551462 1005116 551468 1005168
rect 551520 1005156 551526 1005168
rect 557506 1005156 557534 1005264
rect 574738 1005252 574744 1005264
rect 574796 1005252 574802 1005304
rect 551520 1005128 557534 1005156
rect 551520 1005116 551526 1005128
rect 149882 1005048 149888 1005100
rect 149940 1005088 149946 1005100
rect 152918 1005088 152924 1005100
rect 149940 1005060 152924 1005088
rect 149940 1005048 149946 1005060
rect 152918 1005048 152924 1005060
rect 152976 1005048 152982 1005100
rect 158622 1005048 158628 1005100
rect 158680 1005088 158686 1005100
rect 162118 1005088 162124 1005100
rect 158680 1005060 162124 1005088
rect 158680 1005048 158686 1005060
rect 162118 1005048 162124 1005060
rect 162176 1005048 162182 1005100
rect 263042 1005048 263048 1005100
rect 263100 1005088 263106 1005100
rect 268378 1005088 268384 1005100
rect 263100 1005060 268384 1005088
rect 263100 1005048 263106 1005060
rect 268378 1005048 268384 1005060
rect 268436 1005048 268442 1005100
rect 354398 1005048 354404 1005100
rect 354456 1005088 354462 1005100
rect 356514 1005088 356520 1005100
rect 354456 1005060 356520 1005088
rect 354456 1005048 354462 1005060
rect 356514 1005048 356520 1005060
rect 356572 1005048 356578 1005100
rect 361390 1005048 361396 1005100
rect 361448 1005088 361454 1005100
rect 364886 1005088 364892 1005100
rect 361448 1005060 364892 1005088
rect 361448 1005048 361454 1005060
rect 364886 1005048 364892 1005060
rect 364944 1005048 364950 1005100
rect 430022 1005048 430028 1005100
rect 430080 1005088 430086 1005100
rect 432598 1005088 432604 1005100
rect 430080 1005060 432604 1005088
rect 430080 1005048 430086 1005060
rect 432598 1005048 432604 1005060
rect 432656 1005048 432662 1005100
rect 151078 1004912 151084 1004964
rect 151136 1004952 151142 1004964
rect 153746 1004952 153752 1004964
rect 151136 1004924 153752 1004952
rect 151136 1004912 151142 1004924
rect 153746 1004912 153752 1004924
rect 153804 1004912 153810 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 313826 1004912 313832 1004964
rect 313884 1004952 313890 1004964
rect 316034 1004952 316040 1004964
rect 313884 1004924 316040 1004952
rect 313884 1004912 313890 1004924
rect 316034 1004912 316040 1004924
rect 316092 1004912 316098 1004964
rect 353202 1004912 353208 1004964
rect 353260 1004952 353266 1004964
rect 355686 1004952 355692 1004964
rect 353260 1004924 355692 1004952
rect 353260 1004912 353266 1004924
rect 355686 1004912 355692 1004924
rect 355744 1004912 355750 1004964
rect 422202 1004912 422208 1004964
rect 422260 1004952 422266 1004964
rect 423490 1004952 423496 1004964
rect 422260 1004924 423496 1004952
rect 422260 1004912 422266 1004924
rect 423490 1004912 423496 1004924
rect 423548 1004912 423554 1004964
rect 431218 1004912 431224 1004964
rect 431276 1004952 431282 1004964
rect 433518 1004952 433524 1004964
rect 431276 1004924 433524 1004952
rect 431276 1004912 431282 1004924
rect 433518 1004912 433524 1004924
rect 433576 1004912 433582 1004964
rect 507026 1004912 507032 1004964
rect 507084 1004952 507090 1004964
rect 509694 1004952 509700 1004964
rect 507084 1004924 509700 1004952
rect 507084 1004912 507090 1004924
rect 509694 1004912 509700 1004924
rect 509752 1004912 509758 1004964
rect 556798 1004912 556804 1004964
rect 556856 1004952 556862 1004964
rect 558914 1004952 558920 1004964
rect 556856 1004924 558920 1004952
rect 556856 1004912 556862 1004924
rect 558914 1004912 558920 1004924
rect 558972 1004912 558978 1004964
rect 149698 1004776 149704 1004828
rect 149756 1004816 149762 1004828
rect 151722 1004816 151728 1004828
rect 149756 1004788 151728 1004816
rect 149756 1004776 149762 1004788
rect 151722 1004776 151728 1004788
rect 151780 1004776 151786 1004828
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 207566 1004776 207572 1004828
rect 207624 1004816 207630 1004828
rect 209774 1004816 209780 1004828
rect 207624 1004788 209780 1004816
rect 207624 1004776 207630 1004788
rect 209774 1004776 209780 1004788
rect 209832 1004776 209838 1004828
rect 211246 1004776 211252 1004828
rect 211304 1004816 211310 1004828
rect 215938 1004816 215944 1004828
rect 211304 1004788 215944 1004816
rect 211304 1004776 211310 1004788
rect 215938 1004776 215944 1004788
rect 215996 1004776 216002 1004828
rect 314654 1004776 314660 1004828
rect 314712 1004816 314718 1004828
rect 316678 1004816 316684 1004828
rect 314712 1004788 316684 1004816
rect 314712 1004776 314718 1004788
rect 316678 1004776 316684 1004788
rect 316736 1004776 316742 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365254 1004816 365260 1004828
rect 362644 1004788 365260 1004816
rect 362644 1004776 362650 1004788
rect 365254 1004776 365260 1004788
rect 365312 1004776 365318 1004828
rect 420822 1004776 420828 1004828
rect 420880 1004816 420886 1004828
rect 422662 1004816 422668 1004828
rect 420880 1004788 422668 1004816
rect 420880 1004776 420886 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 507854 1004776 507860 1004828
rect 507912 1004816 507918 1004828
rect 510062 1004816 510068 1004828
rect 507912 1004788 510068 1004816
rect 507912 1004776 507918 1004788
rect 510062 1004776 510068 1004788
rect 510120 1004776 510126 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 151262 1004640 151268 1004692
rect 151320 1004680 151326 1004692
rect 154114 1004680 154120 1004692
rect 151320 1004652 154120 1004680
rect 151320 1004640 151326 1004652
rect 154114 1004640 154120 1004652
rect 154172 1004640 154178 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 212534 1004640 212540 1004692
rect 212592 1004680 212598 1004692
rect 217318 1004680 217324 1004692
rect 212592 1004652 217324 1004680
rect 212592 1004640 212598 1004652
rect 217318 1004640 217324 1004652
rect 217376 1004640 217382 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 499298 1004640 499304 1004692
rect 499356 1004680 499362 1004692
rect 501322 1004680 501328 1004692
rect 499356 1004652 501328 1004680
rect 499356 1004640 499362 1004652
rect 501322 1004640 501328 1004652
rect 501380 1004640 501386 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 505370 1004572 505376 1004624
rect 505428 1004612 505434 1004624
rect 510246 1004612 510252 1004624
rect 505428 1004584 510252 1004612
rect 505428 1004572 505434 1004584
rect 510246 1004572 510252 1004584
rect 510304 1004572 510310 1004624
rect 429194 1004028 429200 1004080
rect 429252 1004068 429258 1004080
rect 446398 1004068 446404 1004080
rect 429252 1004040 446404 1004068
rect 429252 1004028 429258 1004040
rect 446398 1004028 446404 1004040
rect 446456 1004028 446462 1004080
rect 558914 1004028 558920 1004080
rect 558972 1004068 558978 1004080
rect 571978 1004068 571984 1004080
rect 558972 1004040 571984 1004068
rect 558972 1004028 558978 1004040
rect 571978 1004028 571984 1004040
rect 572036 1004028 572042 1004080
rect 92658 1003892 92664 1003944
rect 92716 1003932 92722 1003944
rect 104802 1003932 104808 1003944
rect 92716 1003904 104808 1003932
rect 92716 1003892 92722 1003904
rect 104802 1003892 104808 1003904
rect 104860 1003892 104866 1003944
rect 356882 1003892 356888 1003944
rect 356940 1003932 356946 1003944
rect 375374 1003932 375380 1003944
rect 356940 1003904 375380 1003932
rect 356940 1003892 356946 1003904
rect 375374 1003892 375380 1003904
rect 375432 1003892 375438 1003944
rect 427170 1003892 427176 1003944
rect 427228 1003932 427234 1003944
rect 464798 1003932 464804 1003944
rect 427228 1003904 464804 1003932
rect 427228 1003892 427234 1003904
rect 464798 1003892 464804 1003904
rect 464856 1003892 464862 1003944
rect 505002 1003892 505008 1003944
rect 505060 1003932 505066 1003944
rect 517514 1003932 517520 1003944
rect 505060 1003904 517520 1003932
rect 505060 1003892 505066 1003904
rect 517514 1003892 517520 1003904
rect 517572 1003892 517578 1003944
rect 552290 1003892 552296 1003944
rect 552348 1003932 552354 1003944
rect 572622 1003932 572628 1003944
rect 552348 1003904 572628 1003932
rect 552348 1003892 552354 1003904
rect 572622 1003892 572628 1003904
rect 572680 1003892 572686 1003944
rect 464982 1003280 464988 1003332
rect 465040 1003320 465046 1003332
rect 472434 1003320 472440 1003332
rect 465040 1003292 472440 1003320
rect 465040 1003280 465046 1003292
rect 472434 1003280 472440 1003292
rect 472492 1003280 472498 1003332
rect 424318 1002804 424324 1002856
rect 424376 1002844 424382 1002856
rect 424376 1002816 441614 1002844
rect 424376 1002804 424382 1002816
rect 426526 1002668 426532 1002720
rect 426584 1002708 426590 1002720
rect 441586 1002708 441614 1002816
rect 449158 1002708 449164 1002720
rect 426584 1002680 431954 1002708
rect 441586 1002680 449164 1002708
rect 426584 1002668 426590 1002680
rect 106826 1002600 106832 1002652
rect 106884 1002640 106890 1002652
rect 109494 1002640 109500 1002652
rect 106884 1002612 109500 1002640
rect 106884 1002600 106890 1002612
rect 109494 1002600 109500 1002612
rect 109552 1002600 109558 1002652
rect 253474 1002600 253480 1002652
rect 253532 1002640 253538 1002652
rect 256142 1002640 256148 1002652
rect 253532 1002612 256148 1002640
rect 253532 1002600 253538 1002612
rect 256142 1002600 256148 1002612
rect 256200 1002600 256206 1002652
rect 261018 1002600 261024 1002652
rect 261076 1002640 261082 1002652
rect 264238 1002640 264244 1002652
rect 261076 1002612 264244 1002640
rect 261076 1002600 261082 1002612
rect 264238 1002600 264244 1002612
rect 264296 1002600 264302 1002652
rect 303246 1002600 303252 1002652
rect 303304 1002640 303310 1002652
rect 306926 1002640 306932 1002652
rect 303304 1002612 306932 1002640
rect 303304 1002600 303310 1002612
rect 306926 1002600 306932 1002612
rect 306984 1002600 306990 1002652
rect 422202 1002532 422208 1002584
rect 422260 1002572 422266 1002584
rect 427722 1002572 427728 1002584
rect 422260 1002544 427728 1002572
rect 422260 1002532 422266 1002544
rect 427722 1002532 427728 1002544
rect 427780 1002532 427786 1002584
rect 431926 1002572 431954 1002680
rect 449158 1002668 449164 1002680
rect 449216 1002668 449222 1002720
rect 504174 1002668 504180 1002720
rect 504232 1002708 504238 1002720
rect 518894 1002708 518900 1002720
rect 504232 1002680 518900 1002708
rect 504232 1002668 504238 1002680
rect 518894 1002668 518900 1002680
rect 518952 1002668 518958 1002720
rect 464982 1002572 464988 1002584
rect 431926 1002544 464988 1002572
rect 464982 1002532 464988 1002544
rect 465040 1002532 465046 1002584
rect 501690 1002532 501696 1002584
rect 501748 1002572 501754 1002584
rect 523310 1002572 523316 1002584
rect 501748 1002544 523316 1002572
rect 501748 1002532 501754 1002544
rect 523310 1002532 523316 1002544
rect 523368 1002532 523374 1002584
rect 98638 1002464 98644 1002516
rect 98696 1002504 98702 1002516
rect 101490 1002504 101496 1002516
rect 98696 1002476 101496 1002504
rect 98696 1002464 98702 1002476
rect 101490 1002464 101496 1002476
rect 101548 1002464 101554 1002516
rect 108022 1002464 108028 1002516
rect 108080 1002504 108086 1002516
rect 110690 1002504 110696 1002516
rect 108080 1002476 110696 1002504
rect 108080 1002464 108086 1002476
rect 110690 1002464 110696 1002476
rect 110748 1002464 110754 1002516
rect 251910 1002464 251916 1002516
rect 251968 1002504 251974 1002516
rect 255314 1002504 255320 1002516
rect 251968 1002476 255320 1002504
rect 251968 1002464 251974 1002476
rect 255314 1002464 255320 1002476
rect 255372 1002464 255378 1002516
rect 358722 1002464 358728 1002516
rect 358780 1002504 358786 1002516
rect 359366 1002504 359372 1002516
rect 358780 1002476 359372 1002504
rect 358780 1002464 358786 1002476
rect 359366 1002464 359372 1002476
rect 359424 1002464 359430 1002516
rect 558822 1002464 558828 1002516
rect 558880 1002504 558886 1002516
rect 562502 1002504 562508 1002516
rect 558880 1002476 562508 1002504
rect 558880 1002464 558886 1002476
rect 562502 1002464 562508 1002476
rect 562560 1002464 562566 1002516
rect 261018 1002396 261024 1002448
rect 261076 1002436 261082 1002448
rect 263686 1002436 263692 1002448
rect 261076 1002408 263692 1002436
rect 261076 1002396 261082 1002408
rect 263686 1002396 263692 1002408
rect 263744 1002396 263750 1002448
rect 97258 1002328 97264 1002380
rect 97316 1002368 97322 1002380
rect 100294 1002368 100300 1002380
rect 97316 1002340 100300 1002368
rect 97316 1002328 97322 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 100478 1002328 100484 1002380
rect 100536 1002368 100542 1002380
rect 103146 1002368 103152 1002380
rect 100536 1002340 103152 1002368
rect 100536 1002328 100542 1002340
rect 103146 1002328 103152 1002340
rect 103204 1002328 103210 1002380
rect 106826 1002328 106832 1002380
rect 106884 1002368 106890 1002380
rect 109034 1002368 109040 1002380
rect 106884 1002340 109040 1002368
rect 106884 1002328 106890 1002340
rect 109034 1002328 109040 1002340
rect 109092 1002328 109098 1002380
rect 148502 1002328 148508 1002380
rect 148560 1002368 148566 1002380
rect 150894 1002368 150900 1002380
rect 148560 1002340 150900 1002368
rect 148560 1002328 148566 1002340
rect 150894 1002328 150900 1002340
rect 150952 1002328 150958 1002380
rect 210878 1002328 210884 1002380
rect 210936 1002368 210942 1002380
rect 213178 1002368 213184 1002380
rect 210936 1002340 213184 1002368
rect 210936 1002328 210942 1002340
rect 213178 1002328 213184 1002340
rect 213236 1002328 213242 1002380
rect 253014 1002328 253020 1002380
rect 253072 1002368 253078 1002380
rect 256142 1002368 256148 1002380
rect 253072 1002340 256148 1002368
rect 253072 1002328 253078 1002340
rect 256142 1002328 256148 1002340
rect 256200 1002328 256206 1002380
rect 357342 1002328 357348 1002380
rect 357400 1002368 357406 1002380
rect 359458 1002368 359464 1002380
rect 357400 1002340 359464 1002368
rect 357400 1002328 357406 1002340
rect 359458 1002328 359464 1002340
rect 359516 1002328 359522 1002380
rect 500310 1002328 500316 1002380
rect 500368 1002368 500374 1002380
rect 503346 1002368 503352 1002380
rect 500368 1002340 503352 1002368
rect 500368 1002328 500374 1002340
rect 503346 1002328 503352 1002340
rect 503404 1002328 503410 1002380
rect 560846 1002328 560852 1002380
rect 560904 1002368 560910 1002380
rect 565262 1002368 565268 1002380
rect 560904 1002340 565268 1002368
rect 560904 1002328 560910 1002340
rect 565262 1002328 565268 1002340
rect 565320 1002328 565326 1002380
rect 262674 1002260 262680 1002312
rect 262732 1002300 262738 1002312
rect 265802 1002300 265808 1002312
rect 262732 1002272 265808 1002300
rect 262732 1002260 262738 1002272
rect 265802 1002260 265808 1002272
rect 265860 1002260 265866 1002312
rect 365070 1002260 365076 1002312
rect 365128 1002300 365134 1002312
rect 367922 1002300 367928 1002312
rect 365128 1002272 367928 1002300
rect 365128 1002260 365134 1002272
rect 367922 1002260 367928 1002272
rect 367980 1002260 367986 1002312
rect 95878 1002192 95884 1002244
rect 95936 1002232 95942 1002244
rect 99098 1002232 99104 1002244
rect 95936 1002204 99104 1002232
rect 95936 1002192 95942 1002204
rect 99098 1002192 99104 1002204
rect 99156 1002192 99162 1002244
rect 100018 1002192 100024 1002244
rect 100076 1002232 100082 1002244
rect 101950 1002232 101956 1002244
rect 100076 1002204 101956 1002232
rect 100076 1002192 100082 1002204
rect 101950 1002192 101956 1002204
rect 102008 1002192 102014 1002244
rect 105998 1002192 106004 1002244
rect 106056 1002232 106062 1002244
rect 108298 1002232 108304 1002244
rect 106056 1002204 108304 1002232
rect 106056 1002192 106062 1002204
rect 108298 1002192 108304 1002204
rect 108356 1002192 108362 1002244
rect 108850 1002192 108856 1002244
rect 108908 1002232 108914 1002244
rect 111886 1002232 111892 1002244
rect 108908 1002204 111892 1002232
rect 108908 1002192 108914 1002204
rect 111886 1002192 111892 1002204
rect 111944 1002192 111950 1002244
rect 153838 1002192 153844 1002244
rect 153896 1002232 153902 1002244
rect 155770 1002232 155776 1002244
rect 153896 1002204 155776 1002232
rect 153896 1002192 153902 1002204
rect 155770 1002192 155776 1002204
rect 155828 1002192 155834 1002244
rect 156598 1002192 156604 1002244
rect 156656 1002232 156662 1002244
rect 158714 1002232 158720 1002244
rect 156656 1002204 158720 1002232
rect 156656 1002192 156662 1002204
rect 158714 1002192 158720 1002204
rect 158772 1002192 158778 1002244
rect 203334 1002192 203340 1002244
rect 203392 1002232 203398 1002244
rect 206370 1002232 206376 1002244
rect 203392 1002204 206376 1002232
rect 203392 1002192 203398 1002204
rect 206370 1002192 206376 1002204
rect 206428 1002192 206434 1002244
rect 251450 1002192 251456 1002244
rect 251508 1002232 251514 1002244
rect 254486 1002232 254492 1002244
rect 251508 1002204 254492 1002232
rect 251508 1002192 251514 1002204
rect 254486 1002192 254492 1002204
rect 254544 1002192 254550 1002244
rect 357710 1002192 357716 1002244
rect 357768 1002232 357774 1002244
rect 360838 1002232 360844 1002244
rect 357768 1002204 360844 1002232
rect 357768 1002192 357774 1002204
rect 360838 1002192 360844 1002204
rect 360896 1002192 360902 1002244
rect 428366 1002192 428372 1002244
rect 428424 1002232 428430 1002244
rect 431402 1002232 431408 1002244
rect 428424 1002204 431408 1002232
rect 428424 1002192 428430 1002204
rect 431402 1002192 431408 1002204
rect 431460 1002192 431466 1002244
rect 432046 1002192 432052 1002244
rect 432104 1002232 432110 1002244
rect 435542 1002232 435548 1002244
rect 432104 1002204 435548 1002232
rect 432104 1002192 432110 1002204
rect 435542 1002192 435548 1002204
rect 435600 1002192 435606 1002244
rect 500494 1002192 500500 1002244
rect 500552 1002232 500558 1002244
rect 502978 1002232 502984 1002244
rect 500552 1002204 502984 1002232
rect 500552 1002192 500558 1002204
rect 502978 1002192 502984 1002204
rect 503036 1002192 503042 1002244
rect 509878 1002192 509884 1002244
rect 509936 1002232 509942 1002244
rect 512822 1002232 512828 1002244
rect 509936 1002204 512828 1002232
rect 509936 1002192 509942 1002204
rect 512822 1002192 512828 1002204
rect 512880 1002192 512886 1002244
rect 560018 1002192 560024 1002244
rect 560076 1002232 560082 1002244
rect 562318 1002232 562324 1002244
rect 560076 1002204 562324 1002232
rect 560076 1002192 560082 1002204
rect 562318 1002192 562324 1002204
rect 562376 1002192 562382 1002244
rect 263870 1002124 263876 1002176
rect 263928 1002164 263934 1002176
rect 266998 1002164 267004 1002176
rect 263928 1002136 267004 1002164
rect 263928 1002124 263934 1002136
rect 266998 1002124 267004 1002136
rect 267056 1002124 267062 1002176
rect 365898 1002124 365904 1002176
rect 365956 1002164 365962 1002176
rect 369118 1002164 369124 1002176
rect 365956 1002136 369124 1002164
rect 365956 1002124 365962 1002136
rect 369118 1002124 369124 1002136
rect 369176 1002124 369182 1002176
rect 97442 1002056 97448 1002108
rect 97500 1002096 97506 1002108
rect 100294 1002096 100300 1002108
rect 97500 1002068 100300 1002096
rect 97500 1002056 97506 1002068
rect 100294 1002056 100300 1002068
rect 100352 1002056 100358 1002108
rect 101582 1002056 101588 1002108
rect 101640 1002096 101646 1002108
rect 103146 1002096 103152 1002108
rect 101640 1002068 103152 1002096
rect 101640 1002056 101646 1002068
rect 103146 1002056 103152 1002068
rect 103204 1002056 103210 1002108
rect 105630 1002056 105636 1002108
rect 105688 1002096 105694 1002108
rect 107746 1002096 107752 1002108
rect 105688 1002068 107752 1002096
rect 105688 1002056 105694 1002068
rect 107746 1002056 107752 1002068
rect 107804 1002056 107810 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 112070 1002096 112076 1002108
rect 109736 1002068 112076 1002096
rect 109736 1002056 109742 1002068
rect 112070 1002056 112076 1002068
rect 112128 1002056 112134 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 195146 1002056 195152 1002108
rect 195204 1002096 195210 1002108
rect 203518 1002096 203524 1002108
rect 195204 1002068 203524 1002096
rect 195204 1002056 195210 1002068
rect 203518 1002056 203524 1002068
rect 203576 1002056 203582 1002108
rect 206738 1002056 206744 1002108
rect 206796 1002096 206802 1002108
rect 208394 1002096 208400 1002108
rect 206796 1002068 208400 1002096
rect 206796 1002056 206802 1002068
rect 208394 1002056 208400 1002068
rect 208452 1002056 208458 1002108
rect 210878 1002056 210884 1002108
rect 210936 1002096 210942 1002108
rect 212534 1002096 212540 1002108
rect 210936 1002068 212540 1002096
rect 210936 1002056 210942 1002068
rect 212534 1002056 212540 1002068
rect 212592 1002056 212598 1002108
rect 301498 1002056 301504 1002108
rect 301556 1002096 301562 1002108
rect 304902 1002096 304908 1002108
rect 301556 1002068 304908 1002096
rect 301556 1002056 301562 1002068
rect 304902 1002056 304908 1002068
rect 304960 1002056 304966 1002108
rect 360562 1002056 360568 1002108
rect 360620 1002096 360626 1002108
rect 363598 1002096 363604 1002108
rect 360620 1002068 363604 1002096
rect 360620 1002056 360626 1002068
rect 363598 1002056 363604 1002068
rect 363656 1002056 363662 1002108
rect 419442 1002056 419448 1002108
rect 419500 1002096 419506 1002108
rect 421466 1002096 421472 1002108
rect 419500 1002068 421472 1002096
rect 419500 1002056 419506 1002068
rect 421466 1002056 421472 1002068
rect 421524 1002056 421530 1002108
rect 427538 1002056 427544 1002108
rect 427596 1002096 427602 1002108
rect 429930 1002096 429936 1002108
rect 427596 1002068 429936 1002096
rect 427596 1002056 427602 1002068
rect 429930 1002056 429936 1002068
rect 429988 1002056 429994 1002108
rect 433334 1002056 433340 1002108
rect 433392 1002096 433398 1002108
rect 435358 1002096 435364 1002108
rect 433392 1002068 435364 1002096
rect 433392 1002056 433398 1002068
rect 435358 1002056 435364 1002068
rect 435416 1002056 435422 1002108
rect 503346 1002056 503352 1002108
rect 503404 1002096 503410 1002108
rect 505738 1002096 505744 1002108
rect 503404 1002068 505744 1002096
rect 503404 1002056 503410 1002068
rect 505738 1002056 505744 1002068
rect 505796 1002056 505802 1002108
rect 510338 1002056 510344 1002108
rect 510396 1002096 510402 1002108
rect 512638 1002096 512644 1002108
rect 510396 1002068 512644 1002096
rect 510396 1002056 510402 1002068
rect 512638 1002056 512644 1002068
rect 512696 1002056 512702 1002108
rect 552290 1002056 552296 1002108
rect 552348 1002096 552354 1002108
rect 555418 1002096 555424 1002108
rect 552348 1002068 555424 1002096
rect 552348 1002056 552354 1002068
rect 555418 1002056 555424 1002068
rect 555476 1002056 555482 1002108
rect 557994 1002056 558000 1002108
rect 558052 1002096 558058 1002108
rect 560662 1002096 560668 1002108
rect 558052 1002068 560668 1002096
rect 558052 1002056 558058 1002068
rect 560662 1002056 560668 1002068
rect 560720 1002056 560726 1002108
rect 560846 1002056 560852 1002108
rect 560904 1002096 560910 1002108
rect 565078 1002096 565084 1002108
rect 560904 1002068 565084 1002096
rect 560904 1002056 560910 1002068
rect 565078 1002056 565084 1002068
rect 565136 1002056 565142 1002108
rect 263502 1001988 263508 1002040
rect 263560 1002028 263566 1002040
rect 265618 1002028 265624 1002040
rect 263560 1002000 265624 1002028
rect 263560 1001988 263566 1002000
rect 265618 1001988 265624 1002000
rect 265676 1001988 265682 1002040
rect 365070 1001988 365076 1002040
rect 365128 1002028 365134 1002040
rect 367738 1002028 367744 1002040
rect 365128 1002000 367744 1002028
rect 365128 1001988 365134 1002000
rect 367738 1001988 367744 1002000
rect 367796 1001988 367802 1002040
rect 96062 1001920 96068 1001972
rect 96120 1001960 96126 1001972
rect 98270 1001960 98276 1001972
rect 96120 1001932 98276 1001960
rect 96120 1001920 96126 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 98822 1001920 98828 1001972
rect 98880 1001960 98886 1001972
rect 101122 1001960 101128 1001972
rect 98880 1001932 101128 1001960
rect 98880 1001920 98886 1001932
rect 101122 1001920 101128 1001932
rect 101180 1001920 101186 1001972
rect 101398 1001920 101404 1001972
rect 101456 1001960 101462 1001972
rect 102318 1001960 102324 1001972
rect 101456 1001932 102324 1001960
rect 101456 1001920 101462 1001932
rect 102318 1001920 102324 1001932
rect 102376 1001920 102382 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 108114 1001960 108120 1001972
rect 106056 1001932 108120 1001960
rect 106056 1001920 106062 1001932
rect 108114 1001920 108120 1001932
rect 108172 1001920 108178 1001972
rect 108850 1001920 108856 1001972
rect 108908 1001960 108914 1001972
rect 110506 1001960 110512 1001972
rect 108908 1001932 110512 1001960
rect 108908 1001920 108914 1001932
rect 110506 1001920 110512 1001932
rect 110564 1001920 110570 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 152458 1001920 152464 1001972
rect 152516 1001960 152522 1001972
rect 154574 1001960 154580 1001972
rect 152516 1001932 154580 1001960
rect 152516 1001920 152522 1001932
rect 154574 1001920 154580 1001932
rect 154632 1001920 154638 1001972
rect 154942 1001920 154948 1001972
rect 155000 1001960 155006 1001972
rect 157334 1001960 157340 1001972
rect 155000 1001932 157340 1001960
rect 155000 1001920 155006 1001932
rect 157334 1001920 157340 1001932
rect 157392 1001920 157398 1001972
rect 157794 1001920 157800 1001972
rect 157852 1001960 157858 1001972
rect 160094 1001960 160100 1001972
rect 157852 1001932 160100 1001960
rect 157852 1001920 157858 1001932
rect 160094 1001920 160100 1001932
rect 160152 1001920 160158 1001972
rect 202690 1001960 202696 1001972
rect 195164 1001932 202696 1001960
rect 195164 1001824 195192 1001932
rect 202690 1001920 202696 1001932
rect 202748 1001920 202754 1001972
rect 204162 1001920 204168 1001972
rect 204220 1001960 204226 1001972
rect 205542 1001960 205548 1001972
rect 204220 1001932 205548 1001960
rect 204220 1001920 204226 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 206278 1001920 206284 1001972
rect 206336 1001960 206342 1001972
rect 207566 1001960 207572 1001972
rect 206336 1001932 207572 1001960
rect 206336 1001920 206342 1001932
rect 207566 1001920 207572 1001932
rect 207624 1001920 207630 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 355686 1001920 355692 1001972
rect 355744 1001960 355750 1001972
rect 356698 1001960 356704 1001972
rect 355744 1001932 356704 1001960
rect 355744 1001920 355750 1001932
rect 356698 1001920 356704 1001932
rect 356756 1001920 356762 1001972
rect 360194 1001920 360200 1001972
rect 360252 1001960 360258 1001972
rect 362218 1001960 362224 1001972
rect 360252 1001932 362224 1001960
rect 360252 1001920 360258 1001932
rect 362218 1001920 362224 1001932
rect 362276 1001920 362282 1001972
rect 399938 1001920 399944 1001972
rect 399996 1001960 400002 1001972
rect 422294 1001960 422300 1001972
rect 399996 1001932 422300 1001960
rect 399996 1001920 400002 1001932
rect 422294 1001920 422300 1001932
rect 422352 1001920 422358 1001972
rect 423398 1001920 423404 1001972
rect 423456 1001960 423462 1001972
rect 424318 1001960 424324 1001972
rect 423456 1001932 424324 1001960
rect 423456 1001920 423462 1001932
rect 424318 1001920 424324 1001932
rect 424376 1001920 424382 1001972
rect 425514 1001920 425520 1001972
rect 425572 1001960 425578 1001972
rect 428458 1001960 428464 1001972
rect 425572 1001932 428464 1001960
rect 425572 1001920 425578 1001932
rect 428458 1001920 428464 1001932
rect 428516 1001920 428522 1001972
rect 429194 1001920 429200 1001972
rect 429252 1001960 429258 1001972
rect 431218 1001960 431224 1001972
rect 429252 1001932 431224 1001960
rect 429252 1001920 429258 1001932
rect 431218 1001920 431224 1001932
rect 431276 1001920 431282 1001972
rect 432874 1001920 432880 1001972
rect 432932 1001960 432938 1001972
rect 436738 1001960 436744 1001972
rect 432932 1001932 436744 1001960
rect 432932 1001920 432938 1001932
rect 436738 1001920 436744 1001932
rect 436796 1001920 436802 1001972
rect 496722 1001920 496728 1001972
rect 496780 1001960 496786 1001972
rect 498470 1001960 498476 1001972
rect 496780 1001932 498476 1001960
rect 496780 1001920 496786 1001932
rect 498470 1001920 498476 1001932
rect 498528 1001920 498534 1001972
rect 499574 1001920 499580 1001972
rect 499632 1001960 499638 1001972
rect 500494 1001960 500500 1001972
rect 499632 1001932 500500 1001960
rect 499632 1001920 499638 1001932
rect 500494 1001920 500500 1001932
rect 500552 1001920 500558 1001972
rect 500954 1001920 500960 1001972
rect 501012 1001960 501018 1001972
rect 502150 1001960 502156 1001972
rect 501012 1001932 502156 1001960
rect 501012 1001920 501018 1001932
rect 502150 1001920 502156 1001932
rect 502208 1001920 502214 1001972
rect 502518 1001920 502524 1001972
rect 502576 1001960 502582 1001972
rect 504358 1001960 504364 1001972
rect 502576 1001932 504364 1001960
rect 502576 1001920 502582 1001932
rect 504358 1001920 504364 1001932
rect 504416 1001920 504422 1001972
rect 553302 1001920 553308 1001972
rect 553360 1001960 553366 1001972
rect 555142 1001960 555148 1001972
rect 553360 1001932 555148 1001960
rect 553360 1001920 553366 1001932
rect 555142 1001920 555148 1001932
rect 555200 1001920 555206 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560294 1001960 560300 1001972
rect 558880 1001932 560300 1001960
rect 558880 1001920 558886 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 563698 1001960 563704 1001972
rect 561732 1001932 563704 1001960
rect 561732 1001920 561738 1001932
rect 563698 1001920 563704 1001932
rect 563756 1001920 563762 1001972
rect 195882 1001824 195888 1001836
rect 195164 1001796 195888 1001824
rect 195882 1001784 195888 1001796
rect 195940 1001784 195946 1001836
rect 510154 1001716 510160 1001768
rect 510212 1001756 510218 1001768
rect 516686 1001756 516692 1001768
rect 510212 1001728 516692 1001756
rect 510212 1001716 510218 1001728
rect 516686 1001716 516692 1001728
rect 516744 1001716 516750 1001768
rect 446398 1001580 446404 1001632
rect 446456 1001620 446462 1001632
rect 453206 1001620 453212 1001632
rect 446456 1001592 453212 1001620
rect 446456 1001580 446462 1001592
rect 453206 1001580 453212 1001592
rect 453264 1001580 453270 1001632
rect 428458 1001444 428464 1001496
rect 428516 1001484 428522 1001496
rect 446398 1001484 446404 1001496
rect 428516 1001456 446404 1001484
rect 428516 1001444 428522 1001456
rect 446398 1001444 446404 1001456
rect 446456 1001444 446462 1001496
rect 359458 1001308 359464 1001360
rect 359516 1001348 359522 1001360
rect 372706 1001348 372712 1001360
rect 359516 1001320 372712 1001348
rect 359516 1001308 359522 1001320
rect 372706 1001308 372712 1001320
rect 372764 1001308 372770 1001360
rect 431402 1001308 431408 1001360
rect 431460 1001348 431466 1001360
rect 461854 1001348 461860 1001360
rect 431460 1001320 461860 1001348
rect 431460 1001308 431466 1001320
rect 461854 1001308 461860 1001320
rect 461912 1001308 461918 1001360
rect 93486 1001172 93492 1001224
rect 93544 1001212 93550 1001224
rect 101582 1001212 101588 1001224
rect 93544 1001184 101588 1001212
rect 93544 1001172 93550 1001184
rect 101582 1001172 101588 1001184
rect 101640 1001172 101646 1001224
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 423398 1001172 423404 1001224
rect 423456 1001212 423462 1001224
rect 466454 1001212 466460 1001224
rect 423456 1001184 466460 1001212
rect 423456 1001172 423462 1001184
rect 466454 1001172 466460 1001184
rect 466512 1001172 466518 1001224
rect 496722 1001172 496728 1001224
rect 496780 1001212 496786 1001224
rect 522758 1001212 522764 1001224
rect 496780 1001184 522764 1001212
rect 496780 1001172 496786 1001184
rect 522758 1001172 522764 1001184
rect 522816 1001172 522822 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 97994 1000492 98000 1000544
rect 98052 1000532 98058 1000544
rect 100478 1000532 100484 1000544
rect 98052 1000504 100484 1000532
rect 98052 1000492 98058 1000504
rect 100478 1000492 100484 1000504
rect 100536 1000492 100542 1000544
rect 92842 999744 92848 999796
rect 92900 999784 92906 999796
rect 98822 999784 98828 999796
rect 92900 999756 98828 999784
rect 92900 999744 92906 999756
rect 98822 999744 98828 999756
rect 98880 999744 98886 999796
rect 504358 999744 504364 999796
rect 504416 999784 504422 999796
rect 519814 999784 519820 999796
rect 504416 999756 519820 999784
rect 504416 999744 504422 999756
rect 519814 999744 519820 999756
rect 519872 999744 519878 999796
rect 558178 999744 558184 999796
rect 558236 999784 558242 999796
rect 568114 999784 568120 999796
rect 558236 999756 568120 999784
rect 558236 999744 558242 999756
rect 568114 999744 568120 999756
rect 568172 999744 568178 999796
rect 518894 999200 518900 999252
rect 518952 999240 518958 999252
rect 524046 999240 524052 999252
rect 518952 999212 524052 999240
rect 518952 999200 518958 999212
rect 524046 999200 524052 999212
rect 524104 999200 524110 999252
rect 256694 999132 256700 999184
rect 256752 999172 256758 999184
rect 258166 999172 258172 999184
rect 256752 999144 258172 999172
rect 256752 999132 256758 999144
rect 258166 999132 258172 999144
rect 258224 999132 258230 999184
rect 440878 999064 440884 999116
rect 440936 999104 440942 999116
rect 444282 999104 444288 999116
rect 440936 999076 444288 999104
rect 440936 999064 440942 999076
rect 444282 999064 444288 999076
rect 444340 999064 444346 999116
rect 516962 999064 516968 999116
rect 517020 999104 517026 999116
rect 520182 999104 520188 999116
rect 517020 999076 520188 999104
rect 517020 999064 517026 999076
rect 520182 999064 520188 999076
rect 520240 999064 520246 999116
rect 370498 998792 370504 998844
rect 370556 998832 370562 998844
rect 378042 998832 378048 998844
rect 370556 998804 378048 998832
rect 370556 998792 370562 998804
rect 378042 998792 378048 998804
rect 378100 998792 378106 998844
rect 499298 998792 499304 998844
rect 499356 998832 499362 998844
rect 516870 998832 516876 998844
rect 499356 998804 516876 998832
rect 499356 998792 499362 998804
rect 516870 998792 516876 998804
rect 516928 998792 516934 998844
rect 517514 998792 517520 998844
rect 517572 998832 517578 998844
rect 523678 998832 523684 998844
rect 517572 998804 523684 998832
rect 517572 998792 517578 998804
rect 523678 998792 523684 998804
rect 523736 998792 523742 998844
rect 92474 998656 92480 998708
rect 92532 998696 92538 998708
rect 93302 998696 93308 998708
rect 92532 998668 93308 998696
rect 92532 998656 92538 998668
rect 93302 998656 93308 998668
rect 93360 998656 93366 998708
rect 196618 998656 196624 998708
rect 196676 998696 196682 998708
rect 204346 998696 204352 998708
rect 196676 998668 204352 998696
rect 196676 998656 196682 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 443638 998656 443644 998708
rect 443696 998696 443702 998708
rect 472618 998696 472624 998708
rect 443696 998668 472624 998696
rect 443696 998656 443702 998668
rect 472618 998656 472624 998668
rect 472676 998656 472682 998708
rect 499574 998656 499580 998708
rect 499632 998696 499638 998708
rect 517514 998696 517520 998708
rect 499632 998668 517520 998696
rect 499632 998656 499638 998668
rect 517514 998656 517520 998668
rect 517572 998656 517578 998708
rect 303062 998588 303068 998640
rect 303120 998628 303126 998640
rect 308950 998628 308956 998640
rect 303120 998600 308956 998628
rect 303120 998588 303126 998600
rect 308950 998588 308956 998600
rect 309008 998588 309014 998640
rect 200850 998520 200856 998572
rect 200908 998560 200914 998572
rect 203886 998560 203892 998572
rect 200908 998532 203892 998560
rect 200908 998520 200914 998532
rect 203886 998520 203892 998532
rect 203944 998520 203950 998572
rect 351822 998520 351828 998572
rect 351880 998560 351886 998572
rect 382274 998560 382280 998572
rect 351880 998532 382280 998560
rect 351880 998520 351886 998532
rect 382274 998520 382280 998532
rect 382332 998520 382338 998572
rect 427722 998520 427728 998572
rect 427780 998560 427786 998572
rect 456058 998560 456064 998572
rect 427780 998532 456064 998560
rect 427780 998520 427786 998532
rect 456058 998520 456064 998532
rect 456116 998520 456122 998572
rect 464798 998520 464804 998572
rect 464856 998560 464862 998572
rect 472250 998560 472256 998572
rect 464856 998532 472256 998560
rect 464856 998520 464862 998532
rect 472250 998520 472256 998532
rect 472308 998520 472314 998572
rect 500310 998520 500316 998572
rect 500368 998560 500374 998572
rect 522942 998560 522948 998572
rect 500368 998532 522948 998560
rect 500368 998520 500374 998532
rect 522942 998520 522948 998532
rect 523000 998520 523006 998572
rect 303246 998452 303252 998504
rect 303304 998492 303310 998504
rect 305270 998492 305276 998504
rect 303304 998464 305276 998492
rect 303304 998452 303310 998464
rect 305270 998452 305276 998464
rect 305328 998452 305334 998504
rect 92290 998384 92296 998436
rect 92348 998424 92354 998436
rect 97994 998424 98000 998436
rect 92348 998396 98000 998424
rect 92348 998384 92354 998396
rect 97994 998384 98000 998396
rect 98052 998384 98058 998436
rect 144178 998384 144184 998436
rect 144236 998424 144242 998436
rect 155218 998424 155224 998436
rect 144236 998396 155224 998424
rect 144236 998384 144242 998396
rect 155218 998384 155224 998396
rect 155276 998384 155282 998436
rect 195514 998384 195520 998436
rect 195572 998424 195578 998436
rect 204162 998424 204168 998436
rect 195572 998396 204168 998424
rect 195572 998384 195578 998396
rect 204162 998384 204168 998396
rect 204220 998384 204226 998436
rect 247402 998384 247408 998436
rect 247460 998424 247466 998436
rect 258994 998424 259000 998436
rect 247460 998396 259000 998424
rect 247460 998384 247466 998396
rect 258994 998384 259000 998396
rect 259052 998384 259058 998436
rect 354398 998384 354404 998436
rect 354456 998424 354462 998436
rect 383562 998424 383568 998436
rect 354456 998396 383568 998424
rect 354456 998384 354462 998396
rect 383562 998384 383568 998396
rect 383620 998384 383626 998436
rect 429930 998384 429936 998436
rect 429988 998424 429994 998436
rect 472066 998424 472072 998436
rect 429988 998396 472072 998424
rect 429988 998384 429994 998396
rect 472066 998384 472072 998396
rect 472124 998384 472130 998436
rect 500954 998384 500960 998436
rect 501012 998424 501018 998436
rect 523862 998424 523868 998436
rect 501012 998396 523868 998424
rect 501012 998384 501018 998396
rect 523862 998384 523868 998396
rect 523920 998384 523926 998436
rect 196802 998248 196808 998300
rect 196860 998288 196866 998300
rect 202690 998288 202696 998300
rect 196860 998260 202696 998288
rect 196860 998248 196866 998260
rect 202690 998248 202696 998260
rect 202748 998248 202754 998300
rect 247218 998248 247224 998300
rect 247276 998288 247282 998300
rect 251082 998288 251088 998300
rect 247276 998260 251088 998288
rect 247276 998248 247282 998260
rect 251082 998248 251088 998260
rect 251140 998248 251146 998300
rect 304258 998248 304264 998300
rect 304316 998288 304322 998300
rect 307294 998288 307300 998300
rect 304316 998260 307300 998288
rect 304316 998248 304322 998260
rect 307294 998248 307300 998260
rect 307352 998248 307358 998300
rect 371878 998248 371884 998300
rect 371936 998288 371942 998300
rect 372982 998288 372988 998300
rect 371936 998260 372988 998288
rect 371936 998248 371942 998260
rect 372982 998248 372988 998260
rect 373040 998248 373046 998300
rect 374638 998248 374644 998300
rect 374696 998288 374702 998300
rect 379146 998288 379152 998300
rect 374696 998260 379152 998288
rect 374696 998248 374702 998260
rect 379146 998248 379152 998260
rect 379204 998248 379210 998300
rect 456058 998248 456064 998300
rect 456116 998288 456122 998300
rect 461118 998288 461124 998300
rect 456116 998260 461124 998288
rect 456116 998248 456122 998260
rect 461118 998248 461124 998260
rect 461176 998248 461182 998300
rect 202138 998112 202144 998164
rect 202196 998152 202202 998164
rect 205542 998152 205548 998164
rect 202196 998124 205548 998152
rect 202196 998112 202202 998124
rect 205542 998112 205548 998124
rect 205600 998112 205606 998164
rect 249058 998112 249064 998164
rect 249116 998152 249122 998164
rect 253658 998152 253664 998164
rect 249116 998124 253664 998152
rect 249116 998112 249122 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 256326 998112 256332 998164
rect 256384 998152 256390 998164
rect 257338 998152 257344 998164
rect 256384 998124 257344 998152
rect 256384 998112 256390 998124
rect 257338 998112 257344 998124
rect 257396 998112 257402 998164
rect 304442 998112 304448 998164
rect 304500 998152 304506 998164
rect 306926 998152 306932 998164
rect 304500 998124 306932 998152
rect 304500 998112 304506 998124
rect 306926 998112 306932 998124
rect 306984 998112 306990 998164
rect 199378 998044 199384 998096
rect 199436 998084 199442 998096
rect 201862 998084 201868 998096
rect 199436 998056 201868 998084
rect 199436 998044 199442 998056
rect 201862 998044 201868 998056
rect 201920 998044 201926 998096
rect 555418 998044 555424 998096
rect 555476 998084 555482 998096
rect 557166 998084 557172 998096
rect 555476 998056 557172 998084
rect 555476 998044 555482 998056
rect 557166 998044 557172 998056
rect 557224 998044 557230 998096
rect 591482 998044 591488 998096
rect 591540 998084 591546 998096
rect 625706 998084 625712 998096
rect 591540 998056 625712 998084
rect 591540 998044 591546 998056
rect 625706 998044 625712 998056
rect 625764 998044 625770 998096
rect 202322 997976 202328 998028
rect 202380 998016 202386 998028
rect 204714 998016 204720 998028
rect 202380 997988 204720 998016
rect 202380 997976 202386 997988
rect 204714 997976 204720 997988
rect 204772 997976 204778 998028
rect 250438 997976 250444 998028
rect 250496 998016 250502 998028
rect 253290 998016 253296 998028
rect 250496 997988 253296 998016
rect 250496 997976 250502 997988
rect 253290 997976 253296 997988
rect 253348 997976 253354 998028
rect 302878 997976 302884 998028
rect 302936 998016 302942 998028
rect 306098 998016 306104 998028
rect 302936 997988 306104 998016
rect 302936 997976 302942 997988
rect 306098 997976 306104 997988
rect 306156 997976 306162 998028
rect 307018 997976 307024 998028
rect 307076 998016 307082 998028
rect 308950 998016 308956 998028
rect 307076 997988 308956 998016
rect 307076 997976 307082 997988
rect 308950 997976 308956 997988
rect 309008 997976 309014 998028
rect 550542 997976 550548 998028
rect 550600 998016 550606 998028
rect 553118 998016 553124 998028
rect 550600 997988 553124 998016
rect 550600 997976 550606 997988
rect 553118 997976 553124 997988
rect 553176 997976 553182 998028
rect 195330 997908 195336 997960
rect 195388 997948 195394 997960
rect 200666 997948 200672 997960
rect 195388 997920 200672 997948
rect 195388 997908 195394 997920
rect 200666 997908 200672 997920
rect 200724 997908 200730 997960
rect 254578 997908 254584 997960
rect 254636 997948 254642 997960
rect 256510 997948 256516 997960
rect 254636 997920 256516 997948
rect 254636 997908 254642 997920
rect 256510 997908 256516 997920
rect 256568 997908 256574 997960
rect 257338 997908 257344 997960
rect 257396 997948 257402 997960
rect 258994 997948 259000 997960
rect 257396 997920 259000 997948
rect 257396 997908 257402 997920
rect 258994 997908 259000 997920
rect 259052 997908 259058 997960
rect 259822 997908 259828 997960
rect 259880 997948 259886 997960
rect 262306 997948 262312 997960
rect 259880 997920 262312 997948
rect 259880 997908 259886 997920
rect 262306 997908 262312 997920
rect 262364 997908 262370 997960
rect 377398 997908 377404 997960
rect 377456 997948 377462 997960
rect 383194 997948 383200 997960
rect 377456 997920 383200 997948
rect 377456 997908 377462 997920
rect 383194 997908 383200 997920
rect 383252 997908 383258 997960
rect 591114 997908 591120 997960
rect 591172 997948 591178 997960
rect 625522 997948 625528 997960
rect 591172 997920 625528 997948
rect 591172 997908 591178 997920
rect 625522 997908 625528 997920
rect 625580 997908 625586 997960
rect 201034 997840 201040 997892
rect 201092 997880 201098 997892
rect 203518 997880 203524 997892
rect 201092 997852 203524 997880
rect 201092 997840 201098 997852
rect 203518 997840 203524 997852
rect 203576 997840 203582 997892
rect 247770 997840 247776 997892
rect 247828 997880 247834 997892
rect 252462 997880 252468 997892
rect 247828 997852 252468 997880
rect 247828 997840 247834 997852
rect 252462 997840 252468 997852
rect 252520 997840 252526 997892
rect 305638 997840 305644 997892
rect 305696 997880 305702 997892
rect 307754 997880 307760 997892
rect 305696 997852 307760 997880
rect 305696 997840 305702 997852
rect 307754 997840 307760 997852
rect 307812 997840 307818 997892
rect 308398 997840 308404 997892
rect 308456 997880 308462 997892
rect 310606 997880 310612 997892
rect 308456 997852 310612 997880
rect 308456 997840 308462 997852
rect 310606 997840 310612 997852
rect 310664 997840 310670 997892
rect 461854 997840 461860 997892
rect 461912 997880 461918 997892
rect 463878 997880 463884 997892
rect 461912 997852 463884 997880
rect 461912 997840 461918 997852
rect 463878 997840 463884 997852
rect 463936 997840 463942 997892
rect 196066 997772 196072 997824
rect 196124 997812 196130 997824
rect 198366 997812 198372 997824
rect 196124 997784 198372 997812
rect 196124 997772 196130 997784
rect 198366 997772 198372 997784
rect 198424 997772 198430 997824
rect 254946 997772 254952 997824
rect 255004 997812 255010 997824
rect 256970 997812 256976 997824
rect 255004 997784 256976 997812
rect 255004 997772 255010 997784
rect 256970 997772 256976 997784
rect 257028 997772 257034 997824
rect 258166 997772 258172 997824
rect 258224 997812 258230 997824
rect 259454 997812 259460 997824
rect 258224 997784 259460 997812
rect 258224 997772 258230 997784
rect 259454 997772 259460 997784
rect 259512 997772 259518 997824
rect 260190 997772 260196 997824
rect 260248 997812 260254 997824
rect 262490 997812 262496 997824
rect 260248 997784 262496 997812
rect 260248 997772 260254 997784
rect 262490 997772 262496 997784
rect 262548 997772 262554 997824
rect 378778 997772 378784 997824
rect 378836 997812 378842 997824
rect 383378 997812 383384 997824
rect 378836 997784 383384 997812
rect 378836 997772 378842 997784
rect 383378 997772 383384 997784
rect 383436 997772 383442 997824
rect 551738 997772 551744 997824
rect 551796 997812 551802 997824
rect 553118 997812 553124 997824
rect 551796 997784 553124 997812
rect 551796 997772 551802 997784
rect 553118 997772 553124 997784
rect 553176 997772 553182 997824
rect 591298 997772 591304 997824
rect 591356 997812 591362 997824
rect 625338 997812 625344 997824
rect 591356 997784 625344 997812
rect 591356 997772 591362 997784
rect 625338 997772 625344 997784
rect 625396 997772 625402 997824
rect 93302 997704 93308 997756
rect 93360 997744 93366 997756
rect 103514 997744 103520 997756
rect 93360 997716 103520 997744
rect 93360 997704 93366 997716
rect 103514 997704 103520 997716
rect 103572 997704 103578 997756
rect 109494 997704 109500 997756
rect 109552 997744 109558 997756
rect 116302 997744 116308 997756
rect 109552 997716 116308 997744
rect 109552 997704 109558 997716
rect 116302 997704 116308 997716
rect 116360 997704 116366 997756
rect 143994 997704 144000 997756
rect 144052 997744 144058 997756
rect 160094 997744 160100 997756
rect 144052 997716 160100 997744
rect 144052 997704 144058 997716
rect 160094 997704 160100 997716
rect 160152 997704 160158 997756
rect 162118 997704 162124 997756
rect 162176 997744 162182 997756
rect 170306 997744 170312 997756
rect 162176 997716 170312 997744
rect 162176 997704 162182 997716
rect 170306 997704 170312 997716
rect 170364 997704 170370 997756
rect 209774 997744 209780 997756
rect 200086 997716 209780 997744
rect 195698 997636 195704 997688
rect 195756 997676 195762 997688
rect 200086 997676 200114 997716
rect 209774 997704 209780 997716
rect 209832 997704 209838 997756
rect 246574 997704 246580 997756
rect 246632 997744 246638 997756
rect 254762 997744 254768 997756
rect 246632 997716 254768 997744
rect 246632 997704 246638 997716
rect 254762 997704 254768 997716
rect 254820 997704 254826 997756
rect 299106 997704 299112 997756
rect 299164 997744 299170 997756
rect 311894 997744 311900 997756
rect 299164 997716 311900 997744
rect 299164 997704 299170 997716
rect 311894 997704 311900 997716
rect 311952 997704 311958 997756
rect 365254 997704 365260 997756
rect 365312 997744 365318 997756
rect 372522 997744 372528 997756
rect 365312 997716 372528 997744
rect 365312 997704 365318 997716
rect 372522 997704 372528 997716
rect 372580 997704 372586 997756
rect 399938 997704 399944 997756
rect 399996 997744 400002 997756
rect 431954 997744 431960 997756
rect 399996 997716 431960 997744
rect 399996 997704 400002 997716
rect 431954 997704 431960 997716
rect 432012 997704 432018 997756
rect 432598 997704 432604 997756
rect 432656 997744 432662 997756
rect 439866 997744 439872 997756
rect 432656 997716 439872 997744
rect 432656 997704 432662 997716
rect 439866 997704 439872 997716
rect 439924 997704 439930 997756
rect 464982 997704 464988 997756
rect 465040 997744 465046 997756
rect 471054 997744 471060 997756
rect 465040 997716 471060 997744
rect 465040 997704 465046 997716
rect 471054 997704 471060 997716
rect 471112 997704 471118 997756
rect 488902 997704 488908 997756
rect 488960 997744 488966 997756
rect 507854 997744 507860 997756
rect 488960 997716 507860 997744
rect 488960 997704 488966 997716
rect 507854 997704 507860 997716
rect 507912 997704 507918 997756
rect 509694 997704 509700 997756
rect 509752 997744 509758 997756
rect 516686 997744 516692 997756
rect 509752 997716 516692 997744
rect 509752 997704 509758 997716
rect 516686 997704 516692 997716
rect 516744 997704 516750 997756
rect 195756 997648 200114 997676
rect 195756 997636 195762 997648
rect 540514 997636 540520 997688
rect 540572 997676 540578 997688
rect 556982 997676 556988 997688
rect 540572 997648 556988 997676
rect 540572 997636 540578 997648
rect 556982 997636 556988 997648
rect 557040 997636 557046 997688
rect 566458 997636 566464 997688
rect 566516 997676 566522 997688
rect 591482 997676 591488 997688
rect 566516 997648 591488 997676
rect 566516 997636 566522 997648
rect 591482 997636 591488 997648
rect 591540 997636 591546 997688
rect 108298 997568 108304 997620
rect 108356 997608 108362 997620
rect 117222 997608 117228 997620
rect 108356 997580 117228 997608
rect 108356 997568 108362 997580
rect 117222 997568 117228 997580
rect 117280 997568 117286 997620
rect 144822 997568 144828 997620
rect 144880 997608 144886 997620
rect 158714 997608 158720 997620
rect 144880 997580 158720 997608
rect 144880 997568 144886 997580
rect 158714 997568 158720 997580
rect 158772 997568 158778 997620
rect 360838 997568 360844 997620
rect 360896 997608 360902 997620
rect 372338 997608 372344 997620
rect 360896 997580 372344 997608
rect 360896 997568 360902 997580
rect 372338 997568 372344 997580
rect 372396 997568 372402 997620
rect 422294 997568 422300 997620
rect 422352 997608 422358 997620
rect 426250 997608 426256 997620
rect 422352 997580 426256 997608
rect 422352 997568 422358 997580
rect 426250 997568 426256 997580
rect 426308 997568 426314 997620
rect 431218 997568 431224 997620
rect 431276 997608 431282 997620
rect 439682 997608 439688 997620
rect 431276 997580 439688 997608
rect 431276 997568 431282 997580
rect 439682 997568 439688 997580
rect 439740 997568 439746 997620
rect 489086 997568 489092 997620
rect 489144 997608 489150 997620
rect 506474 997608 506480 997620
rect 489144 997580 506480 997608
rect 489144 997568 489150 997580
rect 506474 997568 506480 997580
rect 506532 997568 506538 997620
rect 509970 997568 509976 997620
rect 510028 997608 510034 997620
rect 517054 997608 517060 997620
rect 510028 997580 517060 997608
rect 510028 997568 510034 997580
rect 517054 997568 517060 997580
rect 517112 997568 517118 997620
rect 554498 997500 554504 997552
rect 554556 997540 554562 997552
rect 591114 997540 591120 997552
rect 554556 997512 591120 997540
rect 554556 997500 554562 997512
rect 591114 997500 591120 997512
rect 591172 997500 591178 997552
rect 540330 997364 540336 997416
rect 540388 997404 540394 997416
rect 560294 997404 560300 997416
rect 540388 997376 560300 997404
rect 540388 997364 540394 997376
rect 560294 997364 560300 997376
rect 560352 997364 560358 997416
rect 573358 997364 573364 997416
rect 573416 997404 573422 997416
rect 591298 997404 591304 997416
rect 573416 997376 591304 997404
rect 573416 997364 573422 997376
rect 591298 997364 591304 997376
rect 591356 997364 591362 997416
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 204898 997268 204904 997280
rect 200264 997240 204904 997268
rect 200264 997228 200270 997240
rect 204898 997228 204904 997240
rect 204956 997228 204962 997280
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 554682 997160 554688 997212
rect 554740 997200 554746 997212
rect 568942 997200 568948 997212
rect 554740 997172 568948 997200
rect 554740 997160 554746 997172
rect 568942 997160 568948 997172
rect 569000 997160 569006 997212
rect 572622 997160 572628 997212
rect 572680 997200 572686 997212
rect 623682 997200 623688 997212
rect 572680 997172 623688 997200
rect 572680 997160 572686 997172
rect 623682 997160 623688 997172
rect 623740 997160 623746 997212
rect 444282 997024 444288 997076
rect 444340 997064 444346 997076
rect 470502 997064 470508 997076
rect 444340 997036 470508 997064
rect 444340 997024 444346 997036
rect 470502 997024 470508 997036
rect 470560 997024 470566 997076
rect 505738 997024 505744 997076
rect 505796 997064 505802 997076
rect 519998 997064 520004 997076
rect 505796 997036 520004 997064
rect 505796 997024 505802 997036
rect 519998 997024 520004 997036
rect 520056 997024 520062 997076
rect 550542 997024 550548 997076
rect 550600 997064 550606 997076
rect 620094 997064 620100 997076
rect 550600 997036 620100 997064
rect 550600 997024 550606 997036
rect 620094 997024 620100 997036
rect 620152 997024 620158 997076
rect 197354 996888 197360 996940
rect 197412 996928 197418 996940
rect 200942 996928 200948 996940
rect 197412 996900 200948 996928
rect 197412 996888 197418 996900
rect 200942 996888 200948 996900
rect 201000 996888 201006 996940
rect 570598 996888 570604 996940
rect 570656 996928 570662 996940
rect 590562 996928 590568 996940
rect 570656 996900 590568 996928
rect 570656 996888 570662 996900
rect 590562 996888 590568 996900
rect 590620 996888 590626 996940
rect 106918 996752 106924 996804
rect 106976 996792 106982 996804
rect 110506 996792 110512 996804
rect 106976 996764 110512 996792
rect 106976 996752 106982 996764
rect 110506 996752 110512 996764
rect 110564 996752 110570 996804
rect 303246 996684 303252 996736
rect 303304 996724 303310 996736
rect 304442 996724 304448 996736
rect 303304 996696 304448 996724
rect 303304 996684 303310 996696
rect 304442 996684 304448 996696
rect 304500 996684 304506 996736
rect 144822 996480 144828 996532
rect 144880 996520 144886 996532
rect 150434 996520 150440 996532
rect 144880 996492 150440 996520
rect 144880 996480 144886 996492
rect 150434 996480 150440 996492
rect 150492 996480 150498 996532
rect 103882 996384 103888 996396
rect 93320 996356 103888 996384
rect 93320 996260 93348 996356
rect 103882 996344 103888 996356
rect 103940 996344 103946 996396
rect 143994 996344 144000 996396
rect 144052 996384 144058 996396
rect 151262 996384 151268 996396
rect 144052 996356 151268 996384
rect 144052 996344 144058 996356
rect 151262 996344 151268 996356
rect 151320 996344 151326 996396
rect 199378 996384 199384 996396
rect 195716 996356 199384 996384
rect 195716 996260 195744 996356
rect 199378 996344 199384 996356
rect 199436 996344 199442 996396
rect 299382 996344 299388 996396
rect 299440 996384 299446 996396
rect 360194 996384 360200 996396
rect 299440 996356 360200 996384
rect 299440 996344 299446 996356
rect 360194 996344 360200 996356
rect 360252 996344 360258 996396
rect 200942 996276 200948 996328
rect 201000 996316 201006 996328
rect 206278 996316 206284 996328
rect 201000 996288 206284 996316
rect 201000 996276 201006 996288
rect 206278 996276 206284 996288
rect 206336 996276 206342 996328
rect 553302 996276 553308 996328
rect 553360 996316 553366 996328
rect 553360 996288 605834 996316
rect 553360 996276 553366 996288
rect 93302 996208 93308 996260
rect 93360 996208 93366 996260
rect 195698 996208 195704 996260
rect 195756 996208 195762 996260
rect 247586 996208 247592 996260
rect 247644 996248 247650 996260
rect 263686 996248 263692 996260
rect 247644 996220 263692 996248
rect 247644 996208 247650 996220
rect 263686 996208 263692 996220
rect 263744 996208 263750 996260
rect 605806 996248 605834 996288
rect 618162 996248 618168 996260
rect 605806 996220 618168 996248
rect 618162 996208 618168 996220
rect 618220 996208 618226 996260
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 211154 996112 211160 996124
rect 171836 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 211798 996072 211804 996124
rect 211856 996112 211862 996124
rect 262490 996112 262496 996124
rect 211856 996084 262496 996112
rect 211856 996072 211862 996084
rect 262490 996072 262496 996084
rect 262548 996072 262554 996124
rect 265802 996072 265808 996124
rect 265860 996112 265866 996124
rect 316034 996112 316040 996124
rect 265860 996084 316040 996112
rect 265860 996072 265866 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 382918 996072 382924 996124
rect 382976 996112 382982 996124
rect 433518 996112 433524 996124
rect 382976 996084 433524 996112
rect 382976 996072 382982 996084
rect 433518 996072 433524 996084
rect 433576 996072 433582 996124
rect 169386 995936 169392 995988
rect 169444 995976 169450 995988
rect 171502 995976 171508 995988
rect 169444 995948 171508 995976
rect 169444 995936 169450 995948
rect 171502 995936 171508 995948
rect 171560 995936 171566 995988
rect 177298 995936 177304 995988
rect 177356 995976 177362 995988
rect 212534 995976 212540 995988
rect 177356 995948 212540 995976
rect 177356 995936 177362 995948
rect 212534 995936 212540 995948
rect 212592 995936 212598 995988
rect 229738 995936 229744 995988
rect 229796 995976 229802 995988
rect 262306 995976 262312 995988
rect 229796 995948 262312 995976
rect 229796 995936 229802 995948
rect 262306 995936 262312 995948
rect 262364 995936 262370 995988
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 299290 995976 299296 995988
rect 264296 995948 299296 995976
rect 264296 995936 264302 995948
rect 299290 995936 299296 995948
rect 299348 995936 299354 995988
rect 366358 995936 366364 995988
rect 366416 995976 366422 995988
rect 400858 995976 400864 995988
rect 366416 995948 400864 995976
rect 366416 995936 366422 995948
rect 400858 995936 400864 995948
rect 400916 995936 400922 995988
rect 136450 995800 136456 995852
rect 136508 995840 136514 995852
rect 143810 995840 143816 995852
rect 136508 995812 143816 995840
rect 136508 995800 136514 995812
rect 143810 995800 143816 995812
rect 143868 995800 143874 995852
rect 170674 995800 170680 995852
rect 170732 995840 170738 995852
rect 171686 995840 171692 995852
rect 170732 995812 171692 995840
rect 170732 995800 170738 995812
rect 171686 995800 171692 995812
rect 171744 995800 171750 995852
rect 213178 995800 213184 995852
rect 213236 995840 213242 995852
rect 261294 995840 261300 995852
rect 213236 995812 261300 995840
rect 213236 995800 213242 995812
rect 261294 995800 261300 995812
rect 261352 995800 261358 995852
rect 364886 995800 364892 995852
rect 364944 995840 364950 995852
rect 402238 995840 402244 995852
rect 364944 995812 402244 995840
rect 364944 995800 364950 995812
rect 402238 995800 402244 995812
rect 402296 995800 402302 995852
rect 518158 995800 518164 995852
rect 518216 995840 518222 995852
rect 524046 995840 524052 995852
rect 518216 995812 524052 995840
rect 518216 995800 518222 995812
rect 524046 995800 524052 995812
rect 524104 995800 524110 995852
rect 92658 995528 92664 995580
rect 92716 995568 92722 995580
rect 97442 995568 97448 995580
rect 92716 995540 97448 995568
rect 92716 995528 92722 995540
rect 97442 995528 97448 995540
rect 97500 995528 97506 995580
rect 171042 995528 171048 995580
rect 171100 995568 171106 995580
rect 171100 995540 171916 995568
rect 171100 995528 171106 995540
rect 171888 995415 171916 995540
rect 246206 995528 246212 995580
rect 246264 995568 246270 995580
rect 256326 995568 256332 995580
rect 246264 995540 256332 995568
rect 246264 995528 246270 995540
rect 256326 995528 256332 995540
rect 256384 995528 256390 995580
rect 383194 995528 383200 995580
rect 383252 995568 383258 995580
rect 385034 995568 385040 995580
rect 383252 995540 385040 995568
rect 383252 995528 383258 995540
rect 385034 995528 385040 995540
rect 385092 995528 385098 995580
rect 415946 995528 415952 995580
rect 416004 995528 416010 995580
rect 472618 995528 472624 995580
rect 472676 995568 472682 995580
rect 473354 995568 473360 995580
rect 472676 995540 473360 995568
rect 472676 995528 472682 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 494698 995528 494704 995580
rect 494756 995568 494762 995580
rect 511074 995568 511080 995580
rect 494756 995540 511080 995568
rect 494756 995528 494762 995540
rect 511074 995528 511080 995540
rect 511132 995528 511138 995580
rect 523678 995528 523684 995580
rect 523736 995568 523742 995580
rect 524782 995568 524788 995580
rect 523736 995540 524788 995568
rect 523736 995528 523742 995540
rect 524782 995528 524788 995540
rect 524840 995528 524846 995580
rect 625706 995528 625712 995580
rect 625764 995568 625770 995580
rect 626534 995568 626540 995580
rect 625764 995540 626540 995568
rect 625764 995528 625770 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 194870 995460 194876 995512
rect 194928 995500 194934 995512
rect 197354 995500 197360 995512
rect 194928 995472 197360 995500
rect 194928 995460 194934 995472
rect 197354 995460 197360 995472
rect 197412 995460 197418 995512
rect 246758 995392 246764 995444
rect 246816 995432 246822 995444
rect 253474 995432 253480 995444
rect 246816 995404 253480 995432
rect 246816 995392 246822 995404
rect 253474 995392 253480 995404
rect 253532 995392 253538 995444
rect 383470 995392 383476 995444
rect 383528 995432 383534 995444
rect 385678 995432 385684 995444
rect 383528 995404 385684 995432
rect 383528 995392 383534 995404
rect 385678 995392 385684 995404
rect 385736 995392 385742 995444
rect 171686 995277 171692 995329
rect 171744 995277 171750 995329
rect 189442 995324 189448 995376
rect 189500 995364 189506 995376
rect 192938 995364 192944 995376
rect 189500 995336 192944 995364
rect 189500 995324 189506 995336
rect 192938 995324 192944 995336
rect 192996 995324 193002 995376
rect 193122 995324 193128 995376
rect 193180 995364 193186 995376
rect 196066 995364 196072 995376
rect 193180 995336 196072 995364
rect 193180 995324 193186 995336
rect 196066 995324 196072 995336
rect 196124 995324 196130 995376
rect 228358 995324 228364 995376
rect 228416 995364 228422 995376
rect 245286 995364 245292 995376
rect 228416 995336 245292 995364
rect 228416 995324 228422 995336
rect 245286 995324 245292 995336
rect 245344 995324 245350 995376
rect 245562 995324 245568 995376
rect 245620 995364 245626 995376
rect 246574 995364 246580 995376
rect 245620 995336 246580 995364
rect 245620 995324 245626 995336
rect 246574 995324 246580 995336
rect 246632 995324 246638 995376
rect 292298 995324 292304 995376
rect 292356 995364 292362 995376
rect 295978 995364 295984 995376
rect 292356 995336 295984 995364
rect 292356 995324 292362 995336
rect 295978 995324 295984 995336
rect 296036 995324 296042 995376
rect 296162 995324 296168 995376
rect 296220 995364 296226 995376
rect 298462 995364 298468 995376
rect 296220 995336 298468 995364
rect 296220 995324 296226 995336
rect 298462 995324 298468 995336
rect 298520 995324 298526 995376
rect 396626 995324 396632 995376
rect 396684 995364 396690 995376
rect 400122 995364 400128 995376
rect 396684 995336 400128 995364
rect 396684 995324 396690 995336
rect 400122 995324 400128 995336
rect 400180 995324 400186 995376
rect 415964 995373 415992 995528
rect 362218 995256 362224 995308
rect 362276 995296 362282 995308
rect 387794 995296 387800 995308
rect 362276 995268 387800 995296
rect 362276 995256 362282 995268
rect 387794 995256 387800 995268
rect 387852 995256 387858 995308
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 184796 995188 184802 995240
rect 184854 995228 184860 995240
rect 194134 995228 194140 995240
rect 184854 995200 194140 995228
rect 184854 995188 184860 995200
rect 194134 995188 194140 995200
rect 194192 995188 194198 995240
rect 194318 995188 194324 995240
rect 194376 995228 194382 995240
rect 195514 995228 195520 995240
rect 194376 995200 195520 995228
rect 194376 995188 194382 995200
rect 195514 995188 195520 995200
rect 195572 995188 195578 995240
rect 244228 995188 244234 995240
rect 244286 995228 244292 995240
rect 247218 995228 247224 995240
rect 244286 995200 247224 995228
rect 244286 995188 244292 995200
rect 247218 995188 247224 995200
rect 247276 995188 247282 995240
rect 283466 995188 283472 995240
rect 283524 995228 283530 995240
rect 300118 995228 300124 995240
rect 283524 995200 300124 995228
rect 283524 995188 283530 995200
rect 300118 995188 300124 995200
rect 300176 995188 300182 995240
rect 380894 995120 380900 995172
rect 380952 995160 380958 995172
rect 416148 995160 416176 995261
rect 380952 995132 416176 995160
rect 380952 995120 380958 995132
rect 489730 995120 489736 995172
rect 489788 995160 489794 995172
rect 489914 995160 489920 995172
rect 489788 995132 489920 995160
rect 489788 995120 489794 995132
rect 489914 995120 489920 995132
rect 489972 995120 489978 995172
rect 172330 995092 172336 995104
rect 171428 995064 172336 995092
rect 172330 995052 172336 995064
rect 172388 995052 172394 995104
rect 180610 995052 180616 995104
rect 180668 995092 180674 995104
rect 202138 995092 202144 995104
rect 180668 995064 202144 995092
rect 180668 995052 180674 995064
rect 202138 995052 202144 995064
rect 202196 995052 202202 995104
rect 232866 995052 232872 995104
rect 232924 995092 232930 995104
rect 257338 995092 257344 995104
rect 232924 995064 257344 995092
rect 232924 995052 232930 995064
rect 257338 995052 257344 995064
rect 257396 995052 257402 995104
rect 285950 995052 285956 995104
rect 286008 995092 286014 995104
rect 309134 995092 309140 995104
rect 286008 995064 309140 995092
rect 286008 995052 286014 995064
rect 309134 995052 309140 995064
rect 309192 995052 309198 995104
rect 425146 995052 425152 995104
rect 425204 995092 425210 995104
rect 484118 995092 484124 995104
rect 425204 995064 484124 995092
rect 425204 995052 425210 995064
rect 484118 995052 484124 995064
rect 484176 995052 484182 995104
rect 515398 995052 515404 995104
rect 515456 995092 515462 995104
rect 537386 995092 537392 995104
rect 515456 995064 537392 995092
rect 515456 995052 515462 995064
rect 537386 995052 537392 995064
rect 537444 995052 537450 995104
rect 568114 995052 568120 995104
rect 568172 995092 568178 995104
rect 629662 995092 629668 995104
rect 568172 995064 629668 995092
rect 568172 995052 568178 995064
rect 629662 995052 629668 995064
rect 629720 995052 629726 995104
rect 358722 994984 358728 995036
rect 358780 995024 358786 995036
rect 398834 995024 398840 995036
rect 358780 994996 398840 995024
rect 358780 994984 358786 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 638862 994984 638868 995036
rect 638920 995024 638926 995036
rect 640794 995024 640800 995036
rect 638920 994996 640800 995024
rect 638920 994984 638926 994996
rect 640794 994984 640800 994996
rect 640852 994984 640858 995036
rect 641714 994984 641720 995036
rect 641772 995024 641778 995036
rect 660408 995024 660436 995121
rect 641772 994996 660436 995024
rect 641772 994984 641778 994996
rect 660574 994983 660580 995035
rect 660632 994983 660638 995035
rect 171244 994881 171272 994967
rect 181438 994916 181444 994968
rect 181496 994956 181502 994968
rect 200942 994956 200948 994968
rect 181496 994928 200948 994956
rect 181496 994916 181502 994928
rect 200942 994916 200948 994928
rect 201000 994916 201006 994968
rect 229002 994916 229008 994968
rect 229060 994956 229066 994968
rect 246206 994956 246212 994968
rect 229060 994928 246212 994956
rect 229060 994916 229066 994928
rect 246206 994916 246212 994928
rect 246264 994916 246270 994968
rect 284110 994916 284116 994968
rect 284168 994956 284174 994968
rect 308398 994956 308404 994968
rect 284168 994928 308404 994956
rect 284168 994916 284174 994928
rect 308398 994916 308404 994928
rect 308456 994916 308462 994968
rect 419442 994916 419448 994968
rect 419500 994956 419506 994968
rect 568206 994956 568212 994968
rect 419500 994928 568212 994956
rect 419500 994916 419506 994928
rect 568206 994916 568212 994928
rect 568264 994916 568270 994968
rect 568942 994916 568948 994968
rect 569000 994956 569006 994968
rect 569000 994928 636056 994956
rect 569000 994916 569006 994928
rect 78306 994780 78312 994832
rect 78364 994820 78370 994832
rect 102778 994820 102784 994832
rect 78364 994792 102784 994820
rect 78364 994780 78370 994792
rect 102778 994780 102784 994792
rect 102836 994780 102842 994832
rect 129734 994780 129740 994832
rect 129792 994820 129798 994832
rect 155954 994820 155960 994832
rect 129792 994792 155960 994820
rect 129792 994780 129798 994792
rect 155954 994780 155960 994792
rect 156012 994780 156018 994832
rect 170858 994829 170864 994881
rect 170916 994829 170922 994881
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 363598 994848 363604 994900
rect 363656 994888 363662 994900
rect 396994 994888 397000 994900
rect 363656 994860 397000 994888
rect 363656 994848 363662 994860
rect 396994 994848 397000 994860
rect 397052 994848 397058 994900
rect 636028 994888 636056 994928
rect 640978 994888 640984 994900
rect 636028 994860 640984 994888
rect 640978 994848 640984 994860
rect 641036 994848 641042 994900
rect 245286 994780 245292 994832
rect 245344 994820 245350 994832
rect 247586 994820 247592 994832
rect 245344 994792 247592 994820
rect 245344 994780 245350 994792
rect 247586 994780 247592 994792
rect 247644 994780 247650 994832
rect 287146 994780 287152 994832
rect 287204 994820 287210 994832
rect 296714 994820 296720 994832
rect 287204 994792 296720 994820
rect 287204 994780 287210 994792
rect 296714 994780 296720 994792
rect 296772 994780 296778 994832
rect 456242 994780 456248 994832
rect 456300 994820 456306 994832
rect 471238 994820 471244 994832
rect 456300 994792 471244 994820
rect 456300 994780 456306 994792
rect 471238 994780 471244 994792
rect 471296 994780 471302 994832
rect 472434 994780 472440 994832
rect 472492 994820 472498 994832
rect 475930 994820 475936 994832
rect 472492 994792 475936 994820
rect 472492 994780 472498 994792
rect 475930 994780 475936 994792
rect 475988 994780 475994 994832
rect 476114 994780 476120 994832
rect 476172 994820 476178 994832
rect 485222 994820 485228 994832
rect 476172 994792 485228 994820
rect 476172 994780 476178 994792
rect 485222 994780 485228 994792
rect 485280 994780 485286 994832
rect 486602 994780 486608 994832
rect 486660 994820 486666 994832
rect 489730 994820 489736 994832
rect 486660 994792 489736 994820
rect 486660 994780 486666 994792
rect 489730 994780 489736 994792
rect 489788 994780 489794 994832
rect 502978 994780 502984 994832
rect 503036 994820 503042 994832
rect 534350 994820 534356 994832
rect 503036 994792 534356 994820
rect 503036 994780 503042 994792
rect 534350 994780 534356 994792
rect 534408 994780 534414 994832
rect 569218 994780 569224 994832
rect 569276 994820 569282 994832
rect 635826 994820 635832 994832
rect 569276 994792 635832 994820
rect 569276 994780 569282 994792
rect 635826 994780 635832 994792
rect 635884 994780 635890 994832
rect 169386 994712 169392 994764
rect 169444 994752 169450 994764
rect 243170 994752 243176 994764
rect 169444 994724 243176 994752
rect 169444 994712 169450 994724
rect 243170 994712 243176 994724
rect 243228 994712 243234 994764
rect 253198 994712 253204 994764
rect 253256 994752 253262 994764
rect 259454 994752 259460 994764
rect 253256 994724 259460 994752
rect 253256 994712 253262 994724
rect 259454 994712 259460 994724
rect 259512 994712 259518 994764
rect 379146 994712 379152 994764
rect 379204 994752 379210 994764
rect 397638 994752 397644 994764
rect 379204 994724 397644 994752
rect 379204 994712 379210 994724
rect 397638 994712 397644 994724
rect 397696 994712 397702 994764
rect 74626 994644 74632 994696
rect 74684 994684 74690 994696
rect 81986 994684 81992 994696
rect 74684 994656 81992 994684
rect 74684 994644 74690 994656
rect 81986 994644 81992 994656
rect 82044 994644 82050 994696
rect 85482 994644 85488 994696
rect 85540 994684 85546 994696
rect 98638 994684 98644 994696
rect 85540 994656 98644 994684
rect 85540 994644 85546 994656
rect 98638 994644 98644 994656
rect 98696 994644 98702 994696
rect 128446 994644 128452 994696
rect 128504 994684 128510 994696
rect 153838 994684 153844 994696
rect 128504 994656 153844 994684
rect 128504 994644 128510 994656
rect 153838 994644 153844 994656
rect 153896 994644 153902 994696
rect 289538 994644 289544 994696
rect 289596 994684 289602 994696
rect 305638 994684 305644 994696
rect 289596 994656 305644 994684
rect 289596 994644 289602 994656
rect 305638 994644 305644 994656
rect 305696 994644 305702 994696
rect 420822 994644 420828 994696
rect 420880 994684 420886 994696
rect 590562 994684 590568 994696
rect 420880 994656 590568 994684
rect 420880 994644 420886 994656
rect 590562 994644 590568 994656
rect 590620 994644 590626 994696
rect 625338 994644 625344 994696
rect 625396 994684 625402 994696
rect 630214 994684 630220 994696
rect 625396 994656 630220 994684
rect 625396 994644 625402 994656
rect 630214 994644 630220 994656
rect 630272 994644 630278 994696
rect 660776 994628 660804 994897
rect 171042 994576 171048 994628
rect 171100 994616 171106 994628
rect 287698 994616 287704 994628
rect 171100 994588 287704 994616
rect 171100 994576 171106 994588
rect 287698 994576 287704 994588
rect 287756 994576 287762 994628
rect 372706 994576 372712 994628
rect 372764 994616 372770 994628
rect 393314 994616 393320 994628
rect 372764 994588 393320 994616
rect 372764 994576 372770 994588
rect 393314 994576 393320 994588
rect 393372 994576 393378 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 74442 994508 74448 994560
rect 74500 994548 74506 994560
rect 97258 994548 97264 994560
rect 74500 994520 97264 994548
rect 74500 994508 74506 994520
rect 97258 994508 97264 994520
rect 97316 994508 97322 994560
rect 132402 994508 132408 994560
rect 132460 994548 132466 994560
rect 149698 994548 149704 994560
rect 132460 994520 149704 994548
rect 132460 994508 132466 994520
rect 149698 994508 149704 994520
rect 149756 994508 149762 994560
rect 301314 994548 301320 994560
rect 296686 994520 301320 994548
rect 170674 994440 170680 994492
rect 170732 994480 170738 994492
rect 296686 994480 296714 994520
rect 301314 994508 301320 994520
rect 301372 994508 301378 994560
rect 470502 994508 470508 994560
rect 470560 994548 470566 994560
rect 475654 994548 475660 994560
rect 470560 994520 475660 994548
rect 470560 994508 470566 994520
rect 475654 994508 475660 994520
rect 475712 994508 475718 994560
rect 475930 994508 475936 994560
rect 475988 994548 475994 994560
rect 490098 994548 490104 994560
rect 475988 994520 490104 994548
rect 475988 994508 475994 994520
rect 490098 994508 490104 994520
rect 490156 994508 490162 994560
rect 519998 994508 520004 994560
rect 520056 994548 520062 994560
rect 539226 994548 539232 994560
rect 520056 994520 539232 994548
rect 520056 994508 520062 994520
rect 539226 994508 539232 994520
rect 539284 994508 539290 994560
rect 567838 994508 567844 994560
rect 567896 994548 567902 994560
rect 591298 994548 591304 994560
rect 567896 994520 591304 994548
rect 567896 994508 567902 994520
rect 591298 994508 591304 994520
rect 591356 994508 591362 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 170732 994452 296714 994480
rect 170732 994440 170738 994452
rect 356698 994440 356704 994492
rect 356756 994480 356762 994492
rect 393958 994480 393964 994492
rect 356756 994452 393964 994480
rect 356756 994440 356762 994452
rect 393958 994440 393964 994452
rect 394016 994440 394022 994492
rect 81342 994372 81348 994424
rect 81400 994412 81406 994424
rect 85482 994412 85488 994424
rect 81400 994384 85488 994412
rect 81400 994372 81406 994384
rect 85482 994372 85488 994384
rect 85540 994372 85546 994424
rect 85666 994372 85672 994424
rect 85724 994412 85730 994424
rect 100018 994412 100024 994424
rect 85724 994384 100024 994412
rect 85724 994372 85730 994384
rect 100018 994372 100024 994384
rect 100076 994372 100082 994424
rect 103882 994372 103888 994424
rect 103940 994412 103946 994424
rect 121730 994412 121736 994424
rect 103940 994384 121736 994412
rect 103940 994372 103946 994384
rect 121730 994372 121736 994384
rect 121788 994372 121794 994424
rect 129090 994372 129096 994424
rect 129148 994412 129154 994424
rect 151078 994412 151084 994424
rect 129148 994384 151084 994412
rect 129148 994372 129154 994384
rect 151078 994372 151084 994384
rect 151136 994372 151142 994424
rect 296806 994372 296812 994424
rect 296864 994412 296870 994424
rect 304258 994412 304264 994424
rect 296864 994384 304264 994412
rect 296864 994372 296870 994384
rect 304258 994372 304264 994384
rect 304316 994372 304322 994424
rect 463878 994372 463884 994424
rect 463936 994412 463942 994424
rect 463936 994384 466454 994412
rect 463936 994372 463942 994384
rect 191742 994304 191748 994356
rect 191800 994344 191806 994356
rect 197354 994344 197360 994356
rect 191800 994316 197360 994344
rect 191800 994304 191806 994316
rect 197354 994304 197360 994316
rect 197412 994304 197418 994356
rect 229186 994304 229192 994356
rect 229244 994344 229250 994356
rect 234062 994344 234068 994356
rect 229244 994316 234068 994344
rect 229244 994304 229250 994316
rect 234062 994304 234068 994316
rect 234120 994304 234126 994356
rect 256694 994344 256700 994356
rect 237300 994316 256700 994344
rect 73154 994236 73160 994288
rect 73212 994276 73218 994288
rect 111886 994276 111892 994288
rect 73212 994248 111892 994276
rect 73212 994236 73218 994248
rect 111886 994236 111892 994248
rect 111944 994236 111950 994288
rect 150434 994236 150440 994288
rect 150492 994276 150498 994288
rect 186498 994276 186504 994288
rect 150492 994248 186504 994276
rect 150492 994236 150498 994248
rect 186498 994236 186504 994248
rect 186556 994236 186562 994288
rect 139210 994168 139216 994220
rect 139268 994208 139274 994220
rect 144546 994208 144552 994220
rect 139268 994180 144552 994208
rect 139268 994168 139274 994180
rect 144546 994168 144552 994180
rect 144604 994168 144610 994220
rect 231578 994168 231584 994220
rect 231636 994208 231642 994220
rect 237300 994208 237328 994316
rect 256694 994304 256700 994316
rect 256752 994304 256758 994356
rect 287698 994304 287704 994356
rect 287756 994344 287762 994356
rect 287756 994316 296714 994344
rect 287756 994304 287762 994316
rect 296686 994276 296714 994316
rect 298830 994276 298836 994288
rect 296686 994248 298836 994276
rect 298830 994236 298836 994248
rect 298888 994236 298894 994288
rect 360194 994236 360200 994288
rect 360252 994276 360258 994288
rect 381170 994276 381176 994288
rect 360252 994248 381176 994276
rect 360252 994236 360258 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 426250 994236 426256 994288
rect 426308 994276 426314 994288
rect 446122 994276 446128 994288
rect 426308 994248 446128 994276
rect 426308 994236 426314 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 466426 994276 466454 994384
rect 466546 994372 466552 994424
rect 466604 994412 466610 994424
rect 475746 994412 475752 994424
rect 466604 994384 475752 994412
rect 466604 994372 466610 994384
rect 475746 994372 475752 994384
rect 475804 994372 475810 994424
rect 476068 994372 476074 994424
rect 476126 994412 476132 994424
rect 476126 994384 485084 994412
rect 476126 994372 476132 994384
rect 485056 994276 485084 994384
rect 485222 994372 485228 994424
rect 485280 994412 485286 994424
rect 487798 994412 487804 994424
rect 485280 994384 487804 994412
rect 485280 994372 485286 994384
rect 487798 994372 487804 994384
rect 487856 994372 487862 994424
rect 498102 994372 498108 994424
rect 498160 994412 498166 994424
rect 538030 994412 538036 994424
rect 498160 994384 538036 994412
rect 498160 994372 498166 994384
rect 538030 994372 538036 994384
rect 538088 994372 538094 994424
rect 571978 994372 571984 994424
rect 572036 994412 572042 994424
rect 639046 994412 639052 994424
rect 572036 994384 639052 994412
rect 572036 994372 572042 994384
rect 639046 994372 639052 994384
rect 639104 994372 639110 994424
rect 489914 994276 489920 994288
rect 466426 994248 482140 994276
rect 485056 994248 489920 994276
rect 231636 994180 237328 994208
rect 231636 994168 231642 994180
rect 237466 994168 237472 994220
rect 237524 994208 237530 994220
rect 254578 994208 254584 994220
rect 237524 994180 254584 994208
rect 237524 994168 237530 994180
rect 254578 994168 254584 994180
rect 254636 994168 254642 994220
rect 286502 994168 286508 994220
rect 286560 994208 286566 994220
rect 289538 994208 289544 994220
rect 286560 994180 289544 994208
rect 286560 994168 286566 994180
rect 289538 994168 289544 994180
rect 289596 994168 289602 994220
rect 80698 994100 80704 994152
rect 80756 994140 80762 994152
rect 85666 994140 85672 994152
rect 80756 994112 85672 994140
rect 80756 994100 80762 994112
rect 85666 994100 85672 994112
rect 85724 994100 85730 994152
rect 184934 994100 184940 994152
rect 184992 994140 184998 994152
rect 196618 994140 196624 994152
rect 184992 994112 196624 994140
rect 184992 994100 184998 994112
rect 196618 994100 196624 994112
rect 196676 994100 196682 994152
rect 471054 994100 471060 994152
rect 471112 994140 471118 994152
rect 476022 994140 476028 994152
rect 471112 994112 476028 994140
rect 471112 994100 471118 994112
rect 476022 994100 476028 994112
rect 476080 994100 476086 994152
rect 481634 994140 481640 994152
rect 480226 994112 481640 994140
rect 137554 994032 137560 994084
rect 137612 994072 137618 994084
rect 141786 994072 141792 994084
rect 137612 994044 141792 994072
rect 137612 994032 137618 994044
rect 141786 994032 141792 994044
rect 141844 994032 141850 994084
rect 235902 994032 235908 994084
rect 235960 994072 235966 994084
rect 253014 994072 253020 994084
rect 235960 994044 253020 994072
rect 235960 994032 235966 994044
rect 253014 994032 253020 994044
rect 253072 994032 253078 994084
rect 471238 993964 471244 994016
rect 471296 994004 471302 994016
rect 480226 994004 480254 994112
rect 481634 994100 481640 994112
rect 481692 994100 481698 994152
rect 471296 993976 480254 994004
rect 482112 994004 482140 994248
rect 489914 994236 489920 994248
rect 489972 994236 489978 994288
rect 524046 994236 524052 994288
rect 524104 994276 524110 994288
rect 535546 994276 535552 994288
rect 524104 994248 535552 994276
rect 524104 994236 524110 994248
rect 535546 994236 535552 994248
rect 535604 994236 535610 994288
rect 482278 994100 482284 994152
rect 482336 994140 482342 994152
rect 489546 994140 489552 994152
rect 482336 994112 489552 994140
rect 482336 994100 482342 994112
rect 489546 994100 489552 994112
rect 489604 994100 489610 994152
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 485958 994004 485964 994016
rect 482112 993976 485964 994004
rect 471296 993964 471302 993976
rect 485958 993964 485964 993976
rect 486016 993964 486022 994016
rect 228818 993896 228824 993948
rect 228876 993936 228882 993948
rect 253198 993936 253204 993948
rect 228876 993908 253204 993936
rect 228876 993896 228882 993908
rect 253198 993896 253204 993908
rect 253256 993896 253262 993948
rect 574738 993896 574744 993948
rect 574796 993936 574802 993948
rect 661328 993936 661356 994561
rect 574796 993908 661356 993936
rect 574796 993896 574802 993908
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 195146 993800 195152 993812
rect 171284 993772 195152 993800
rect 171284 993760 171290 993772
rect 195146 993760 195152 993772
rect 195204 993760 195210 993812
rect 232222 993760 232228 993812
rect 232280 993800 232286 993812
rect 237466 993800 237472 993812
rect 232280 993772 237472 993800
rect 232280 993760 232286 993772
rect 237466 993760 237472 993772
rect 237524 993760 237530 993812
rect 243170 993760 243176 993812
rect 243228 993800 243234 993812
rect 247770 993800 247776 993812
rect 243228 993772 247776 993800
rect 243228 993760 243234 993772
rect 247770 993760 247776 993772
rect 247828 993760 247834 993812
rect 522758 993760 522764 993812
rect 522816 993800 522822 993812
rect 660758 993800 660764 993812
rect 522816 993772 660764 993800
rect 522816 993760 522822 993772
rect 660758 993760 660764 993772
rect 660816 993760 660822 993812
rect 170858 993624 170864 993676
rect 170916 993664 170922 993676
rect 195698 993664 195704 993676
rect 170916 993636 195704 993664
rect 170916 993624 170922 993636
rect 195698 993624 195704 993636
rect 195756 993624 195762 993676
rect 229370 993624 229376 993676
rect 229428 993664 229434 993676
rect 238386 993664 238392 993676
rect 229428 993636 238392 993664
rect 229428 993624 229434 993636
rect 238386 993624 238392 993636
rect 238444 993624 238450 993676
rect 516502 993624 516508 993676
rect 516560 993664 516566 993676
rect 660942 993664 660948 993676
rect 516560 993636 660948 993664
rect 516560 993624 516566 993636
rect 660942 993624 660948 993636
rect 661000 993624 661006 993676
rect 549162 993488 549168 993540
rect 549220 993528 549226 993540
rect 639506 993528 639512 993540
rect 549220 993500 639512 993528
rect 549220 993488 549226 993500
rect 639506 993488 639512 993500
rect 639564 993488 639570 993540
rect 551738 993352 551744 993404
rect 551796 993392 551802 993404
rect 637022 993392 637028 993404
rect 551796 993364 637028 993392
rect 551796 993352 551802 993364
rect 637022 993352 637028 993364
rect 637080 993352 637086 993404
rect 51718 993148 51724 993200
rect 51776 993188 51782 993200
rect 107746 993188 107752 993200
rect 51776 993160 107752 993188
rect 51776 993148 51782 993160
rect 107746 993148 107752 993160
rect 107804 993148 107810 993200
rect 50338 993012 50344 993064
rect 50396 993052 50402 993064
rect 108114 993052 108120 993064
rect 50396 993024 108120 993052
rect 50396 993012 50402 993024
rect 108114 993012 108120 993024
rect 108172 993012 108178 993064
rect 202874 993012 202880 993064
rect 202932 993052 202938 993064
rect 213914 993052 213920 993064
rect 202932 993024 213920 993052
rect 202932 993012 202938 993024
rect 213914 993012 213920 993024
rect 213972 993012 213978 993064
rect 563698 993012 563704 993064
rect 563756 993052 563762 993064
rect 608594 993052 608600 993064
rect 563756 993024 608600 993052
rect 563756 993012 563762 993024
rect 608594 993012 608600 993024
rect 608652 993012 608658 993064
rect 55858 992876 55864 992928
rect 55916 992916 55922 992928
rect 146938 992916 146944 992928
rect 55916 992888 146944 992916
rect 55916 992876 55922 992888
rect 146938 992876 146944 992888
rect 146996 992876 147002 992928
rect 197354 992876 197360 992928
rect 197412 992916 197418 992928
rect 251450 992916 251456 992928
rect 197412 992888 251456 992916
rect 197412 992876 197418 992888
rect 251450 992876 251456 992888
rect 251508 992876 251514 992928
rect 316678 992876 316684 992928
rect 316736 992916 316742 992928
rect 364978 992916 364984 992928
rect 316736 992888 364984 992916
rect 316736 992876 316742 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 367922 992876 367928 992928
rect 367980 992916 367986 992928
rect 429930 992916 429936 992928
rect 367980 992888 429936 992916
rect 367980 992876 367986 992888
rect 429930 992876 429936 992888
rect 429988 992876 429994 992928
rect 435542 992876 435548 992928
rect 435600 992916 435606 992928
rect 494698 992916 494704 992928
rect 435600 992888 494704 992916
rect 435600 992876 435606 992888
rect 494698 992876 494704 992888
rect 494756 992876 494762 992928
rect 512822 992876 512828 992928
rect 512880 992916 512886 992928
rect 527266 992916 527272 992928
rect 512880 992888 527272 992916
rect 512880 992876 512886 992888
rect 527266 992876 527272 992888
rect 527324 992876 527330 992928
rect 562502 992876 562508 992928
rect 562560 992916 562566 992928
rect 660298 992916 660304 992928
rect 562560 992888 660304 992916
rect 562560 992876 562566 992888
rect 660298 992876 660304 992888
rect 660356 992876 660362 992928
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 48958 991584 48964 991636
rect 49016 991624 49022 991636
rect 110690 991624 110696 991636
rect 49016 991596 110696 991624
rect 49016 991584 49022 991596
rect 110690 991584 110696 991596
rect 110748 991584 110754 991636
rect 138290 991584 138296 991636
rect 138348 991624 138354 991636
rect 163130 991624 163136 991636
rect 138348 991596 163136 991624
rect 138348 991584 138354 991596
rect 163130 991584 163136 991596
rect 163188 991584 163194 991636
rect 54478 991448 54484 991500
rect 54536 991488 54542 991500
rect 148318 991488 148324 991500
rect 54536 991460 148324 991488
rect 54536 991448 54542 991460
rect 148318 991448 148324 991460
rect 148376 991448 148382 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 318058 991448 318064 991500
rect 318116 991488 318122 991500
rect 349154 991488 349160 991500
rect 318116 991460 349160 991488
rect 318116 991448 318122 991460
rect 349154 991448 349160 991460
rect 349212 991448 349218 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 397822 991488 397828 991500
rect 367796 991460 397828 991488
rect 367796 991448 367802 991460
rect 397822 991448 397828 991460
rect 397880 991448 397886 991500
rect 435358 991448 435364 991500
rect 435416 991488 435422 991500
rect 478966 991488 478972 991500
rect 435416 991460 478972 991488
rect 435416 991448 435422 991460
rect 478966 991448 478972 991460
rect 479024 991448 479030 991500
rect 512638 991448 512644 991500
rect 512696 991488 512702 991500
rect 543826 991488 543832 991500
rect 512696 991460 543832 991488
rect 512696 991448 512702 991460
rect 543826 991448 543832 991460
rect 543884 991448 543890 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 164878 990836 164884 990888
rect 164936 990876 164942 990888
rect 170766 990876 170772 990888
rect 164936 990848 170772 990876
rect 164936 990836 164942 990848
rect 170766 990836 170772 990848
rect 170824 990836 170830 990888
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 89714 990224 89720 990276
rect 89772 990264 89778 990276
rect 112070 990264 112076 990276
rect 89772 990236 112076 990264
rect 89772 990224 89778 990236
rect 112070 990224 112076 990236
rect 112128 990224 112134 990276
rect 560938 990224 560944 990276
rect 560996 990264 561002 990276
rect 668578 990264 668584 990276
rect 560996 990236 668584 990264
rect 560996 990224 561002 990236
rect 668578 990224 668584 990236
rect 668636 990224 668642 990276
rect 44818 990088 44824 990140
rect 44876 990128 44882 990140
rect 109034 990128 109040 990140
rect 44876 990100 109040 990128
rect 44876 990088 44882 990100
rect 109034 990088 109040 990100
rect 109092 990088 109098 990140
rect 319438 990088 319444 990140
rect 319496 990128 319502 990140
rect 332962 990128 332968 990140
rect 319496 990100 332968 990128
rect 319496 990088 319502 990100
rect 332962 990088 332968 990100
rect 333020 990088 333026 990140
rect 369118 990088 369124 990140
rect 369176 990128 369182 990140
rect 414106 990128 414112 990140
rect 369176 990100 414112 990128
rect 369176 990088 369182 990100
rect 414106 990088 414112 990100
rect 414164 990088 414170 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 669958 990128 669964 990140
rect 562376 990100 669964 990128
rect 562376 990088 562382 990100
rect 669958 990088 669964 990100
rect 670016 990088 670022 990140
rect 53282 988728 53288 988780
rect 53340 988768 53346 988780
rect 95878 988768 95884 988780
rect 53340 988740 95884 988768
rect 53340 988728 53346 988740
rect 95878 988728 95884 988740
rect 95936 988728 95942 988780
rect 217318 986620 217324 986672
rect 217376 986660 217382 986672
rect 219434 986660 219440 986672
rect 217376 986632 219440 986660
rect 217376 986620 217382 986632
rect 219434 986620 219440 986632
rect 219492 986620 219498 986672
rect 105814 986552 105820 986604
rect 105872 986592 105878 986604
rect 106918 986592 106924 986604
rect 105872 986564 106924 986592
rect 105872 986552 105878 986564
rect 106918 986552 106924 986564
rect 106976 986552 106982 986604
rect 565078 986076 565084 986128
rect 565136 986116 565142 986128
rect 592494 986116 592500 986128
rect 565136 986088 592500 986116
rect 565136 986076 565142 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 462774 985980 462780 985992
rect 436796 985952 462780 985980
rect 436796 985940 436802 985952
rect 462774 985940 462780 985952
rect 462832 985940 462838 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565262 985940 565268 985992
rect 565320 985980 565326 985992
rect 624970 985980 624976 985992
rect 565320 985952 624976 985980
rect 565320 985940 565326 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 667198 975712 667204 975724
rect 651708 975684 667204 975712
rect 651708 975672 651714 975684
rect 667198 975672 667204 975684
rect 667256 975672 667262 975724
rect 43438 961868 43444 961920
rect 43496 961908 43502 961920
rect 62114 961908 62120 961920
rect 43496 961880 62120 961908
rect 43496 961868 43502 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952416 36544 952468
rect 36596 952456 36602 952468
rect 41690 952456 41696 952468
rect 36596 952428 41696 952456
rect 36596 952416 36602 952428
rect 41690 952416 41696 952428
rect 41748 952416 41754 952468
rect 37918 952212 37924 952264
rect 37976 952252 37982 952264
rect 41690 952252 41696 952264
rect 37976 952224 41696 952252
rect 37976 952212 37982 952224
rect 41690 952212 41696 952224
rect 41748 952212 41754 952264
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 663058 948104 663064 948116
rect 652260 948076 663064 948104
rect 652260 948064 652266 948076
rect 663058 948064 663064 948076
rect 663116 948064 663122 948116
rect 46290 945956 46296 946008
rect 46348 945996 46354 946008
rect 62114 945996 62120 946008
rect 46348 945968 62120 945996
rect 46348 945956 46354 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 35802 942692 35808 942744
rect 35860 942732 35866 942744
rect 40402 942732 40408 942744
rect 35860 942704 40408 942732
rect 35860 942692 35866 942704
rect 40402 942692 40408 942704
rect 40460 942692 40466 942744
rect 35802 941332 35808 941384
rect 35860 941372 35866 941384
rect 38470 941372 38476 941384
rect 35860 941344 38476 941372
rect 35860 941332 35866 941344
rect 38470 941332 38476 941344
rect 38528 941332 38534 941384
rect 35802 939836 35808 939888
rect 35860 939876 35866 939888
rect 39482 939876 39488 939888
rect 35860 939848 39488 939876
rect 35860 939836 35866 939848
rect 39482 939836 39488 939848
rect 39540 939836 39546 939888
rect 39482 938136 39488 938188
rect 39540 938176 39546 938188
rect 41690 938176 41696 938188
rect 39540 938148 41696 938176
rect 39540 938136 39546 938148
rect 41690 938136 41696 938148
rect 41748 938136 41754 938188
rect 38470 937524 38476 937576
rect 38528 937564 38534 937576
rect 41690 937564 41696 937576
rect 38528 937536 41696 937564
rect 38528 937524 38534 937536
rect 41690 937524 41696 937536
rect 41748 937524 41754 937576
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 41322 934328 41328 934380
rect 41380 934368 41386 934380
rect 41690 934368 41696 934380
rect 41380 934340 41696 934368
rect 41380 934328 41386 934340
rect 41690 934328 41696 934340
rect 41748 934328 41754 934380
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 663058 921856 663064 921868
rect 651524 921828 663064 921856
rect 651524 921816 651530 921828
rect 663058 921816 663064 921828
rect 663116 921816 663122 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 665818 909480 665824 909492
rect 652444 909452 665824 909480
rect 652444 909440 652450 909452
rect 665818 909440 665824 909452
rect 665876 909440 665882 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 670970 895676 670976 895688
rect 651524 895648 670976 895676
rect 651524 895636 651530 895648
rect 670970 895636 670976 895648
rect 671028 895636 671034 895688
rect 44082 892752 44088 892764
rect 42858 892724 44088 892752
rect 42858 892466 42886 892724
rect 44082 892712 44088 892724
rect 44140 892712 44146 892764
rect 42938 892254 42990 892260
rect 42938 892196 42990 892202
rect 43076 891948 43128 891954
rect 43076 891890 43128 891896
rect 44082 891868 44088 891880
rect 43194 891840 44088 891868
rect 44082 891828 44088 891840
rect 44140 891828 44146 891880
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 651466 852116 651472 852168
rect 651524 852156 651530 852168
rect 664438 852156 664444 852168
rect 651524 852128 664444 852156
rect 651524 852116 651530 852128
rect 664438 852116 664444 852128
rect 664496 852116 664502 852168
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651834 841780 651840 841832
rect 651892 841820 651898 841832
rect 669958 841820 669964 841832
rect 651892 841792 669964 841820
rect 651892 841780 651898 841792
rect 669958 841780 669964 841792
rect 670016 841780 670022 841832
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817028 35808 817080
rect 35860 817068 35866 817080
rect 41690 817068 41696 817080
rect 35860 817040 41696 817068
rect 35860 817028 35866 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 41598 815640 41604 815652
rect 35860 815612 41604 815640
rect 35860 815600 35866 815612
rect 41598 815600 41604 815612
rect 41656 815600 41662 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 661678 815640 661684 815652
rect 651524 815612 661684 815640
rect 651524 815600 651530 815612
rect 661678 815600 661684 815612
rect 661736 815600 661742 815652
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 41414 814280 41420 814292
rect 35860 814252 41420 814280
rect 35860 814240 35866 814252
rect 41414 814240 41420 814252
rect 41472 814240 41478 814292
rect 41322 810704 41328 810756
rect 41380 810744 41386 810756
rect 41690 810744 41696 810756
rect 41380 810716 41696 810744
rect 41380 810704 41386 810716
rect 41690 810704 41696 810716
rect 41748 810704 41754 810756
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 33042 802408 33048 802460
rect 33100 802448 33106 802460
rect 41690 802448 41696 802460
rect 33100 802420 41696 802448
rect 33100 802408 33106 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 39298 801660 39304 801712
rect 39356 801700 39362 801712
rect 41598 801700 41604 801712
rect 39356 801672 41604 801700
rect 39356 801660 39362 801672
rect 41598 801660 41604 801672
rect 41656 801660 41662 801712
rect 44818 793568 44824 793620
rect 44876 793608 44882 793620
rect 62114 793608 62120 793620
rect 44876 793580 62120 793608
rect 44876 793568 44882 793580
rect 62114 793568 62120 793580
rect 62172 793568 62178 793620
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 652386 775548 652392 775600
rect 652444 775588 652450 775600
rect 668394 775588 668400 775600
rect 652444 775560 668400 775588
rect 652444 775548 652450 775560
rect 668394 775548 668400 775560
rect 668452 775548 668458 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35526 768952 35532 769004
rect 35584 768992 35590 769004
rect 39298 768992 39304 769004
rect 35584 768964 39304 768992
rect 35584 768952 35590 768964
rect 39298 768952 39304 768964
rect 39356 768952 39362 769004
rect 35342 768816 35348 768868
rect 35400 768856 35406 768868
rect 40402 768856 40408 768868
rect 35400 768828 40408 768856
rect 35400 768816 35406 768828
rect 40402 768816 40408 768828
rect 40460 768816 40466 768868
rect 35802 768680 35808 768732
rect 35860 768720 35866 768732
rect 40586 768720 40592 768732
rect 35860 768692 40592 768720
rect 35860 768680 35866 768692
rect 40586 768680 40592 768692
rect 40644 768680 40650 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 35618 767320 35624 767372
rect 35676 767360 35682 767372
rect 41322 767360 41328 767372
rect 35676 767332 41328 767360
rect 35676 767320 35682 767332
rect 41322 767320 41328 767332
rect 41380 767320 41386 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 35802 763240 35808 763292
rect 35860 763280 35866 763292
rect 37918 763280 37924 763292
rect 35860 763252 37924 763280
rect 35860 763240 35866 763252
rect 37918 763240 37924 763252
rect 37976 763240 37982 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 31018 759636 31024 759688
rect 31076 759676 31082 759688
rect 41506 759676 41512 759688
rect 31076 759648 41512 759676
rect 31076 759636 31082 759648
rect 41506 759636 41512 759648
rect 41564 759636 41570 759688
rect 40586 758384 40592 758396
rect 38626 758356 40592 758384
rect 35158 758276 35164 758328
rect 35216 758316 35222 758328
rect 38626 758316 38654 758356
rect 40586 758344 40592 758356
rect 40644 758344 40650 758396
rect 35216 758288 38654 758316
rect 35216 758276 35222 758288
rect 37918 757732 37924 757784
rect 37976 757772 37982 757784
rect 41598 757772 41604 757784
rect 37976 757744 41604 757772
rect 37976 757732 37982 757744
rect 41598 757732 41604 757744
rect 41656 757732 41662 757784
rect 675846 754264 675852 754316
rect 675904 754304 675910 754316
rect 683114 754304 683120 754316
rect 675904 754276 683120 754304
rect 675904 754264 675910 754276
rect 683114 754264 683120 754276
rect 683172 754264 683178 754316
rect 676030 753584 676036 753636
rect 676088 753624 676094 753636
rect 676582 753624 676588 753636
rect 676088 753596 676588 753624
rect 676088 753584 676094 753596
rect 676582 753584 676588 753596
rect 676640 753584 676646 753636
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 672902 734000 672908 734052
rect 672960 734040 672966 734052
rect 673546 734040 673552 734052
rect 672960 734012 673552 734040
rect 672960 734000 672966 734012
rect 673546 734000 673552 734012
rect 673604 734000 673610 734052
rect 35802 730056 35808 730108
rect 35860 730096 35866 730108
rect 41690 730096 41696 730108
rect 35860 730068 41696 730096
rect 35860 730056 35866 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 674098 728628 674104 728680
rect 674156 728668 674162 728680
rect 674156 728640 674406 728668
rect 674156 728628 674162 728640
rect 673086 728424 673092 728476
rect 673144 728464 673150 728476
rect 673144 728436 674268 728464
rect 673144 728424 673150 728436
rect 673914 728152 673920 728204
rect 673972 728192 673978 728204
rect 673972 728164 674072 728192
rect 673972 728152 673978 728164
rect 674044 728110 674072 728164
rect 674150 728136 674202 728142
rect 674150 728078 674202 728084
rect 41322 725908 41328 725960
rect 41380 725948 41386 725960
rect 41690 725948 41696 725960
rect 41380 725920 41696 725948
rect 41380 725908 41386 725920
rect 41690 725908 41696 725920
rect 41748 725908 41754 725960
rect 41322 724480 41328 724532
rect 41380 724520 41386 724532
rect 41690 724520 41696 724532
rect 41380 724492 41696 724520
rect 41380 724480 41386 724492
rect 41690 724480 41696 724492
rect 41748 724480 41754 724532
rect 677318 724208 677324 724260
rect 677376 724248 677382 724260
rect 683850 724248 683856 724260
rect 677376 724220 683856 724248
rect 677376 724208 677382 724220
rect 683850 724208 683856 724220
rect 683908 724208 683914 724260
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 36538 717340 36544 717392
rect 36596 717380 36602 717392
rect 41414 717380 41420 717392
rect 36596 717352 41420 717380
rect 36596 717340 36602 717352
rect 41414 717340 41420 717352
rect 41472 717340 41478 717392
rect 34514 715640 34520 715692
rect 34572 715680 34578 715692
rect 41690 715680 41696 715692
rect 34572 715652 41696 715680
rect 34572 715640 34578 715652
rect 41690 715640 41696 715652
rect 41748 715640 41754 715692
rect 33778 715504 33784 715556
rect 33836 715544 33842 715556
rect 40310 715544 40316 715556
rect 33836 715516 40316 715544
rect 33836 715504 33842 715516
rect 40310 715504 40316 715516
rect 40368 715504 40374 715556
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 651466 709316 651472 709368
rect 651524 709356 651530 709368
rect 664438 709356 664444 709368
rect 651524 709328 664444 709356
rect 651524 709316 651530 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 672534 707208 672540 707260
rect 672592 707248 672598 707260
rect 673270 707248 673276 707260
rect 672592 707220 673276 707248
rect 672592 707208 672598 707220
rect 673270 707208 673276 707220
rect 673328 707208 673334 707260
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 651466 696940 651472 696992
rect 651524 696980 651530 696992
rect 669958 696980 669964 696992
rect 651524 696952 669964 696980
rect 651524 696940 651530 696952
rect 669958 696940 669964 696952
rect 670016 696940 670022 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 35802 687216 35808 687268
rect 35860 687256 35866 687268
rect 41414 687256 41420 687268
rect 35860 687228 41420 687256
rect 35860 687216 35866 687228
rect 41414 687216 41420 687228
rect 41472 687216 41478 687268
rect 35802 683340 35808 683392
rect 35860 683380 35866 683392
rect 35860 683340 35894 683380
rect 35866 683312 35894 683340
rect 41506 683312 41512 683324
rect 35866 683284 41512 683312
rect 41506 683272 41512 683284
rect 41564 683272 41570 683324
rect 35802 683136 35808 683188
rect 35860 683176 35866 683188
rect 41690 683176 41696 683188
rect 35860 683148 41696 683176
rect 35860 683136 35866 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 651650 683136 651656 683188
rect 651708 683176 651714 683188
rect 658918 683176 658924 683188
rect 651708 683148 658924 683176
rect 651708 683136 651714 683148
rect 658918 683136 658924 683148
rect 658976 683136 658982 683188
rect 35802 681980 35808 682032
rect 35860 682020 35866 682032
rect 36538 682020 36544 682032
rect 35860 681992 36544 682020
rect 35860 681980 35866 681992
rect 36538 681980 36544 681992
rect 36596 681980 36602 682032
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35434 681708 35440 681760
rect 35492 681748 35498 681760
rect 40954 681748 40960 681760
rect 35492 681720 40960 681748
rect 35492 681708 35498 681720
rect 40954 681708 40960 681720
rect 41012 681708 41018 681760
rect 35618 674092 35624 674144
rect 35676 674132 35682 674144
rect 39666 674132 39672 674144
rect 35676 674104 39672 674132
rect 35676 674092 35682 674104
rect 39666 674092 39672 674104
rect 39724 674092 39730 674144
rect 36538 673140 36544 673192
rect 36596 673180 36602 673192
rect 40586 673180 40592 673192
rect 36596 673152 40592 673180
rect 36596 673140 36602 673152
rect 40586 673140 40592 673152
rect 40644 673140 40650 673192
rect 32398 672732 32404 672784
rect 32456 672772 32462 672784
rect 41690 672772 41696 672784
rect 32456 672744 41696 672772
rect 32456 672732 32462 672744
rect 41690 672732 41696 672744
rect 41748 672732 41754 672784
rect 37182 670964 37188 671016
rect 37240 671004 37246 671016
rect 40126 671004 40132 671016
rect 37240 670976 40132 671004
rect 37240 670964 37246 670976
rect 40126 670964 40132 670976
rect 40184 670964 40190 671016
rect 651466 669332 651472 669384
rect 651524 669372 651530 669384
rect 661678 669372 661684 669384
rect 651524 669344 661684 669372
rect 651524 669332 651530 669344
rect 661678 669332 661684 669344
rect 661736 669332 661742 669384
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651466 656888 651472 656940
rect 651524 656928 651530 656940
rect 663058 656928 663064 656940
rect 651524 656900 663064 656928
rect 651524 656888 651530 656900
rect 663058 656888 663064 656900
rect 663116 656888 663122 656940
rect 54478 647844 54484 647896
rect 54536 647884 54542 647896
rect 62114 647884 62120 647896
rect 54536 647856 62120 647884
rect 54536 647844 54542 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 41690 644484 41696 644496
rect 35860 644456 41696 644484
rect 35860 644444 35866 644456
rect 41690 644444 41696 644456
rect 41748 644444 41754 644496
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639208 35808 639260
rect 35860 639248 35866 639260
rect 40034 639248 40040 639260
rect 35860 639220 40040 639248
rect 35860 639208 35866 639220
rect 40034 639208 40040 639220
rect 40092 639208 40098 639260
rect 35342 639072 35348 639124
rect 35400 639112 35406 639124
rect 41690 639112 41696 639124
rect 35400 639084 41696 639112
rect 35400 639072 35406 639084
rect 41690 639072 41696 639084
rect 41748 639072 41754 639124
rect 35526 638936 35532 638988
rect 35584 638976 35590 638988
rect 36538 638976 36544 638988
rect 35584 638948 36544 638976
rect 35584 638936 35590 638948
rect 36538 638936 36544 638948
rect 36596 638936 36602 638988
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 41322 637616 41328 637628
rect 35860 637588 41328 637616
rect 35860 637576 35866 637588
rect 41322 637576 41328 637588
rect 41380 637576 41386 637628
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 33778 629892 33784 629944
rect 33836 629932 33842 629944
rect 41690 629932 41696 629944
rect 33836 629904 41696 629932
rect 33836 629892 33842 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651558 628532 651564 628584
rect 651616 628572 651622 628584
rect 667198 628572 667204 628584
rect 651616 628544 667204 628572
rect 651616 628532 651622 628544
rect 667198 628532 667204 628544
rect 667256 628532 667262 628584
rect 48958 623772 48964 623824
rect 49016 623812 49022 623824
rect 62114 623812 62120 623824
rect 49016 623784 62120 623812
rect 49016 623772 49022 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 671062 616156 671068 616208
rect 671120 616196 671126 616208
rect 671706 616196 671712 616208
rect 671120 616168 671712 616196
rect 671120 616156 671126 616168
rect 671706 616156 671712 616168
rect 671764 616156 671770 616208
rect 43286 612904 43971 612932
rect 43622 612728 43628 612740
rect 43397 612700 43628 612728
rect 43622 612688 43628 612700
rect 43680 612688 43686 612740
rect 43806 612620 43812 612672
rect 43864 612660 43870 612672
rect 43943 612660 43971 612904
rect 43864 612632 43971 612660
rect 43864 612620 43870 612632
rect 43990 612524 43996 612536
rect 43516 612496 43996 612524
rect 43990 612484 43996 612496
rect 44048 612484 44054 612536
rect 43582 612332 43634 612338
rect 43714 612280 43720 612332
rect 43772 612280 43778 612332
rect 43582 612274 43634 612280
rect 43732 612102 43760 612280
rect 46934 611912 46940 611924
rect 43838 611884 46940 611912
rect 46934 611872 46940 611884
rect 46992 611872 46998 611924
rect 46106 611708 46112 611720
rect 43957 611680 46112 611708
rect 46106 611668 46112 611680
rect 46164 611668 46170 611720
rect 45554 611504 45560 611516
rect 44068 611476 45560 611504
rect 45554 611464 45560 611476
rect 45612 611464 45618 611516
rect 45738 611300 45744 611312
rect 44181 611272 45744 611300
rect 45738 611260 45744 611272
rect 45796 611260 45802 611312
rect 44272 610972 44324 610978
rect 44272 610914 44324 610920
rect 44379 610836 44431 610842
rect 44379 610778 44431 610784
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 661678 603140 661684 603152
rect 651524 603112 661684 603140
rect 651524 603100 651530 603112
rect 661678 603100 661684 603112
rect 661736 603100 661742 603152
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 41322 596028 41328 596080
rect 41380 596068 41386 596080
rect 41598 596068 41604 596080
rect 41380 596040 41604 596068
rect 41380 596028 41386 596040
rect 41598 596028 41604 596040
rect 41656 596028 41662 596080
rect 41138 594736 41144 594788
rect 41196 594776 41202 594788
rect 41690 594776 41696 594788
rect 41196 594748 41696 594776
rect 41196 594736 41202 594748
rect 41690 594736 41696 594748
rect 41748 594736 41754 594788
rect 40862 593240 40868 593292
rect 40920 593280 40926 593292
rect 41598 593280 41604 593292
rect 40920 593252 41604 593280
rect 40920 593240 40926 593252
rect 41598 593240 41604 593252
rect 41656 593240 41662 593292
rect 40494 592288 40500 592340
rect 40552 592328 40558 592340
rect 41598 592328 41604 592340
rect 40552 592300 41604 592328
rect 40552 592288 40558 592300
rect 41598 592288 41604 592300
rect 41656 592288 41662 592340
rect 675846 591336 675852 591388
rect 675904 591376 675910 591388
rect 682378 591376 682384 591388
rect 675904 591348 682384 591376
rect 675904 591336 675910 591348
rect 682378 591336 682384 591348
rect 682436 591336 682442 591388
rect 652386 590656 652392 590708
rect 652444 590696 652450 590708
rect 665818 590696 665824 590708
rect 652444 590668 665824 590696
rect 652444 590656 652450 590668
rect 665818 590656 665824 590668
rect 665876 590656 665882 590708
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 40126 587160 40132 587172
rect 33100 587132 40132 587160
rect 33100 587120 33106 587132
rect 40126 587120 40132 587132
rect 40184 587120 40190 587172
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 41690 585936 41696 585948
rect 35216 585908 41696 585936
rect 35216 585896 35222 585908
rect 41690 585896 41696 585908
rect 41748 585896 41754 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 39390 585800 39396 585812
rect 31076 585772 39396 585800
rect 31076 585760 31082 585772
rect 39390 585760 39396 585772
rect 39448 585760 39454 585812
rect 40862 584536 40868 584588
rect 40920 584576 40926 584588
rect 41598 584576 41604 584588
rect 40920 584548 41604 584576
rect 40920 584536 40926 584548
rect 41598 584536 41604 584548
rect 41656 584536 41662 584588
rect 50338 583720 50344 583772
rect 50396 583760 50402 583772
rect 62114 583760 62120 583772
rect 50396 583732 62120 583760
rect 50396 583720 50402 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 671614 578252 671620 578264
rect 671448 578224 671620 578252
rect 671448 577992 671476 578224
rect 671614 578212 671620 578224
rect 671672 578212 671678 578264
rect 671430 577940 671436 577992
rect 671488 577940 671494 577992
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 664438 576892 664444 576904
rect 651524 576864 664444 576892
rect 651524 576852 651530 576864
rect 664438 576852 664444 576864
rect 664496 576852 664502 576904
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 41322 557540 41328 557592
rect 41380 557580 41386 557592
rect 41506 557580 41512 557592
rect 41380 557552 41512 557580
rect 41380 557540 41386 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 41322 554752 41328 554804
rect 41380 554792 41386 554804
rect 41690 554792 41696 554804
rect 41380 554764 41696 554792
rect 41380 554752 41386 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 41138 552100 41144 552152
rect 41196 552140 41202 552152
rect 41598 552140 41604 552152
rect 41196 552112 41604 552140
rect 41196 552100 41202 552112
rect 41598 552100 41604 552112
rect 41656 552100 41662 552152
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 40586 549380 40592 549432
rect 40644 549420 40650 549432
rect 41598 549420 41604 549432
rect 40644 549392 41604 549420
rect 40644 549380 40650 549392
rect 41598 549380 41604 549392
rect 41656 549380 41662 549432
rect 41230 549244 41236 549296
rect 41288 549284 41294 549296
rect 41690 549284 41696 549296
rect 41288 549256 41696 549284
rect 41288 549244 41294 549256
rect 41690 549244 41696 549256
rect 41748 549244 41754 549296
rect 41230 548088 41236 548140
rect 41288 548128 41294 548140
rect 41690 548128 41696 548140
rect 41288 548100 41696 548128
rect 41288 548088 41294 548100
rect 41690 548088 41696 548100
rect 41748 548088 41754 548140
rect 31754 547816 31760 547868
rect 31812 547856 31818 547868
rect 38286 547856 38292 547868
rect 31812 547828 38292 547856
rect 31812 547816 31818 547828
rect 38286 547816 38292 547828
rect 38344 547816 38350 547868
rect 675938 547612 675944 547664
rect 675996 547652 676002 547664
rect 678238 547652 678244 547664
rect 675996 547624 678244 547652
rect 675996 547612 676002 547624
rect 678238 547612 678244 547624
rect 678296 547612 678302 547664
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 32398 542988 32404 543040
rect 32456 543028 32462 543040
rect 41506 543028 41512 543040
rect 32456 543000 41512 543028
rect 32456 542988 32462 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 38286 542308 38292 542360
rect 38344 542348 38350 542360
rect 41690 542348 41696 542360
rect 38344 542320 41696 542348
rect 38344 542308 38350 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669958 536840 669964 536852
rect 651524 536812 669964 536840
rect 651524 536800 651530 536812
rect 669958 536800 669964 536812
rect 670016 536800 670022 536852
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 676858 520276 676864 520328
rect 676916 520316 676922 520328
rect 683114 520316 683120 520328
rect 676916 520288 683120 520316
rect 676916 520276 676922 520288
rect 683114 520276 683120 520288
rect 683172 520276 683178 520328
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 676030 518780 676036 518832
rect 676088 518820 676094 518832
rect 677870 518820 677876 518832
rect 676088 518792 677876 518820
rect 676088 518780 676094 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675846 503616 675852 503668
rect 675904 503656 675910 503668
rect 679618 503656 679624 503668
rect 675904 503628 679624 503656
rect 675904 503616 675910 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 675846 500896 675852 500948
rect 675904 500936 675910 500948
rect 680998 500936 681004 500948
rect 675904 500908 681004 500936
rect 675904 500896 675910 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 652570 494708 652576 494760
rect 652628 494748 652634 494760
rect 663242 494748 663248 494760
rect 652628 494720 663248 494748
rect 652628 494708 652634 494720
rect 663242 494708 663248 494720
rect 663300 494708 663306 494760
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 677410 489880 677416 489932
rect 677468 489920 677474 489932
rect 683114 489920 683120 489932
rect 677468 489892 683120 489920
rect 677468 489880 677474 489892
rect 683114 489880 683120 489892
rect 683172 489880 683178 489932
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 667198 484412 667204 484424
rect 654106 484384 667204 484412
rect 667198 484372 667204 484384
rect 667256 484372 667262 484424
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 665818 470608 665824 470620
rect 651524 470580 665824 470608
rect 651524 470568 651530 470580
rect 665818 470568 665824 470580
rect 665876 470568 665882 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 661678 456804 661684 456816
rect 652444 456776 661684 456804
rect 652444 456764 652450 456776
rect 661678 456764 661684 456776
rect 661736 456764 661742 456816
rect 673454 456560 673460 456612
rect 673512 456600 673518 456612
rect 673512 456572 673988 456600
rect 673512 456560 673518 456572
rect 673960 456246 673988 456572
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673736 455796 673788 455802
rect 673736 455738 673788 455744
rect 673598 455592 673650 455598
rect 675846 455540 675852 455592
rect 675904 455580 675910 455592
rect 677042 455580 677048 455592
rect 675904 455552 677048 455580
rect 675904 455540 675910 455552
rect 677042 455540 677048 455552
rect 677100 455540 677106 455592
rect 673598 455534 673650 455540
rect 672258 455336 672264 455388
rect 672316 455376 672322 455388
rect 672316 455348 673532 455376
rect 672316 455336 672322 455348
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 671798 454996 671804 455048
rect 671856 455036 671862 455048
rect 671856 455008 673302 455036
rect 671856 454996 671862 455008
rect 673040 454860 673046 454912
rect 673098 454860 673104 454912
rect 672902 454656 672908 454708
rect 672960 454696 672966 454708
rect 672960 454656 672994 454696
rect 672966 454410 672994 454656
rect 673058 454614 673086 454860
rect 673164 454640 673216 454646
rect 673164 454582 673216 454588
rect 672816 454232 672868 454238
rect 672816 454174 672868 454180
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 671338 430624 671344 430636
rect 651524 430596 671344 430624
rect 651524 430584 651530 430596
rect 671338 430584 671344 430596
rect 671396 430584 671402 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41322 425008 41328 425060
rect 41380 425048 41386 425060
rect 41690 425048 41696 425060
rect 41380 425020 41696 425048
rect 41380 425008 41386 425020
rect 41690 425008 41696 425020
rect 41748 425008 41754 425060
rect 41322 423784 41328 423836
rect 41380 423824 41386 423836
rect 41598 423824 41604 423836
rect 41380 423796 41604 423824
rect 41380 423784 41386 423796
rect 41598 423784 41604 423796
rect 41656 423784 41662 423836
rect 41322 422288 41328 422340
rect 41380 422328 41386 422340
rect 41598 422328 41604 422340
rect 41380 422300 41604 422328
rect 41380 422288 41386 422300
rect 41598 422288 41604 422300
rect 41656 422288 41662 422340
rect 41322 420928 41328 420980
rect 41380 420968 41386 420980
rect 41598 420968 41604 420980
rect 41380 420940 41604 420968
rect 41380 420928 41386 420940
rect 41598 420928 41604 420940
rect 41656 420928 41662 420980
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 663058 416820 663064 416832
rect 651892 416792 663064 416820
rect 651892 416780 651898 416792
rect 663058 416780 663064 416792
rect 663116 416780 663122 416832
rect 33686 416168 33692 416220
rect 33744 416208 33750 416220
rect 41690 416208 41696 416220
rect 33744 416180 41696 416208
rect 33744 416168 33750 416180
rect 41690 416168 41696 416180
rect 41748 416168 41754 416220
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 41138 387064 41144 387116
rect 41196 387104 41202 387116
rect 41690 387104 41696 387116
rect 41196 387076 41696 387104
rect 41196 387064 41202 387076
rect 41690 387064 41696 387076
rect 41748 387064 41754 387116
rect 44634 385432 44640 385484
rect 44692 385472 44698 385484
rect 45002 385472 45008 385484
rect 44692 385444 45008 385472
rect 44692 385432 44698 385444
rect 45002 385432 45008 385444
rect 45060 385432 45066 385484
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41690 382412 41696 382424
rect 41380 382384 41696 382412
rect 41380 382372 41386 382384
rect 41690 382372 41696 382384
rect 41748 382372 41754 382424
rect 41138 382236 41144 382288
rect 41196 382276 41202 382288
rect 41690 382276 41696 382288
rect 41196 382248 41696 382276
rect 41196 382236 41202 382248
rect 41690 382236 41696 382248
rect 41748 382236 41754 382288
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 41690 379556 41696 379568
rect 35860 379528 41696 379556
rect 35860 379516 35866 379528
rect 41690 379516 41696 379528
rect 41748 379516 41754 379568
rect 35802 375980 35808 376032
rect 35860 376020 35866 376032
rect 39574 376020 39580 376032
rect 35860 375992 39580 376020
rect 35860 375980 35866 375992
rect 39574 375980 39580 375992
rect 39632 375980 39638 376032
rect 51718 375368 51724 375420
rect 51776 375408 51782 375420
rect 62114 375408 62120 375420
rect 51776 375380 62120 375408
rect 51776 375368 51782 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 28902 371832 28908 371884
rect 28960 371872 28966 371884
rect 41690 371872 41696 371884
rect 28960 371844 41696 371872
rect 28960 371832 28966 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 651834 364352 651840 364404
rect 651892 364392 651898 364404
rect 661862 364392 661868 364404
rect 651892 364364 661868 364392
rect 651892 364352 651898 364364
rect 661862 364352 661868 364364
rect 661920 364352 661926 364404
rect 46382 362924 46388 362976
rect 46440 362964 46446 362976
rect 62114 362964 62120 362976
rect 46440 362936 62120 362964
rect 46440 362924 46446 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 45002 355784 45008 355836
rect 45060 355824 45066 355836
rect 45646 355824 45652 355836
rect 45060 355796 45652 355824
rect 45060 355784 45066 355796
rect 45646 355784 45652 355796
rect 45704 355784 45710 355836
rect 44634 355648 44640 355700
rect 44692 355688 44698 355700
rect 44692 355660 45048 355688
rect 44692 355648 44698 355660
rect 44569 354832 44575 354884
rect 44627 354872 44633 354884
rect 44627 354844 44839 354872
rect 44627 354832 44633 354844
rect 44575 354680 44627 354686
rect 44575 354622 44627 354628
rect 44811 354600 44839 354844
rect 45020 354600 45048 355660
rect 44811 354572 44956 354600
rect 45020 354572 45063 354600
rect 44793 354424 44799 354476
rect 44851 354424 44857 354476
rect 44686 354340 44738 354346
rect 44811 354314 44839 354424
rect 44686 354282 44738 354288
rect 44928 354110 44956 354572
rect 45035 353906 45063 354572
rect 45646 354056 45652 354068
rect 45158 354028 45652 354056
rect 45158 353702 45186 354028
rect 45646 354016 45652 354028
rect 45704 354016 45710 354068
rect 45922 353784 45928 353796
rect 45250 353756 45928 353784
rect 45250 353498 45278 353756
rect 45922 353744 45928 353756
rect 45980 353744 45986 353796
rect 45554 353240 45560 353252
rect 45385 353212 45560 353240
rect 45554 353200 45560 353212
rect 45612 353200 45618 353252
rect 652386 350548 652392 350600
rect 652444 350588 652450 350600
rect 667382 350588 667388 350600
rect 652444 350560 667388 350588
rect 652444 350548 652450 350560
rect 667382 350548 667388 350560
rect 667440 350548 667446 350600
rect 35802 343612 35808 343664
rect 35860 343652 35866 343664
rect 40218 343652 40224 343664
rect 35860 343624 40224 343652
rect 35860 343612 35866 343624
rect 40218 343612 40224 343624
rect 40276 343612 40282 343664
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 36630 339504 36636 339516
rect 35860 339476 36636 339504
rect 35860 339464 35866 339476
rect 36630 339464 36636 339476
rect 36688 339464 36694 339516
rect 46198 336744 46204 336796
rect 46256 336784 46262 336796
rect 62114 336784 62120 336796
rect 46256 336756 62120 336784
rect 46256 336744 46262 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 667750 324340 667756 324352
rect 651524 324312 667756 324340
rect 651524 324300 651530 324312
rect 667750 324300 667756 324312
rect 667808 324300 667814 324352
rect 53282 322940 53288 322992
rect 53340 322980 53346 322992
rect 62114 322980 62120 322992
rect 53340 322952 62120 322980
rect 53340 322940 53346 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 54478 310496 54484 310548
rect 54536 310536 54542 310548
rect 62114 310536 62120 310548
rect 54536 310508 62120 310536
rect 54536 310496 54542 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667198 310536 667204 310548
rect 651524 310508 667204 310536
rect 651524 310496 651530 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 678974 298092 678980 298104
rect 675904 298064 678980 298092
rect 675904 298052 675910 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676030 297916 676036 297968
rect 676088 297956 676094 297968
rect 680998 297956 681004 297968
rect 676088 297928 681004 297956
rect 676088 297916 676094 297928
rect 680998 297916 681004 297928
rect 681056 297916 681062 297968
rect 41322 284928 41328 284980
rect 41380 284968 41386 284980
rect 41690 284968 41696 284980
rect 41380 284940 41696 284968
rect 41380 284928 41386 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 37918 284724 37924 284776
rect 37976 284764 37982 284776
rect 41690 284764 41696 284776
rect 37976 284736 41696 284764
rect 37976 284724 37982 284736
rect 41690 284724 41696 284736
rect 41748 284724 41754 284776
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667566 284356 667572 284368
rect 651524 284328 667572 284356
rect 651524 284316 651530 284328
rect 667566 284316 667572 284328
rect 667624 284316 667630 284368
rect 464798 276768 464804 276820
rect 464856 276808 464862 276820
rect 532786 276808 532792 276820
rect 464856 276780 532792 276808
rect 464856 276768 464862 276780
rect 532786 276768 532792 276780
rect 532844 276768 532850 276820
rect 482830 276632 482836 276684
rect 482888 276672 482894 276684
rect 558822 276672 558828 276684
rect 482888 276644 558828 276672
rect 482888 276632 482894 276644
rect 558822 276632 558828 276644
rect 558880 276632 558886 276684
rect 103698 275952 103704 276004
rect 103756 275992 103762 276004
rect 160738 275992 160744 276004
rect 103756 275964 160744 275992
rect 103756 275952 103762 275964
rect 160738 275952 160744 275964
rect 160796 275952 160802 276004
rect 166350 275952 166356 276004
rect 166408 275992 166414 276004
rect 182082 275992 182088 276004
rect 166408 275964 182088 275992
rect 166408 275952 166414 275964
rect 182082 275952 182088 275964
rect 182140 275952 182146 276004
rect 188798 275952 188804 276004
rect 188856 275992 188862 276004
rect 222838 275992 222844 276004
rect 188856 275964 222844 275992
rect 188856 275952 188862 275964
rect 222838 275952 222844 275964
rect 222896 275952 222902 276004
rect 385954 275952 385960 276004
rect 386012 275992 386018 276004
rect 401594 275992 401600 276004
rect 386012 275964 401600 275992
rect 386012 275952 386018 275964
rect 401594 275952 401600 275964
rect 401652 275952 401658 276004
rect 432966 275952 432972 276004
rect 433024 275992 433030 276004
rect 487890 275992 487896 276004
rect 433024 275964 487896 275992
rect 433024 275952 433030 275964
rect 487890 275952 487896 275964
rect 487948 275952 487954 276004
rect 512546 275952 512552 276004
rect 512604 275992 512610 276004
rect 526898 275992 526904 276004
rect 512604 275964 526904 275992
rect 512604 275952 512610 275964
rect 526898 275952 526904 275964
rect 526956 275952 526962 276004
rect 527358 275952 527364 276004
rect 527416 275992 527422 276004
rect 607306 275992 607312 276004
rect 527416 275964 607312 275992
rect 527416 275952 527422 275964
rect 607306 275952 607312 275964
rect 607364 275952 607370 276004
rect 88334 275816 88340 275868
rect 88392 275856 88398 275868
rect 146938 275856 146944 275868
rect 88392 275828 146944 275856
rect 88392 275816 88398 275828
rect 146938 275816 146944 275828
rect 146996 275816 147002 275868
rect 149790 275816 149796 275868
rect 149848 275856 149854 275868
rect 187878 275856 187884 275868
rect 149848 275828 187884 275856
rect 149848 275816 149854 275828
rect 187878 275816 187884 275828
rect 187936 275816 187942 275868
rect 393866 275816 393872 275868
rect 393924 275856 393930 275868
rect 411070 275856 411076 275868
rect 393924 275828 411076 275856
rect 393924 275816 393930 275828
rect 411070 275816 411076 275828
rect 411128 275816 411134 275868
rect 411254 275816 411260 275868
rect 411312 275856 411318 275868
rect 415762 275856 415768 275868
rect 411312 275828 415768 275856
rect 411312 275816 411318 275828
rect 415762 275816 415768 275828
rect 415820 275816 415826 275868
rect 423582 275816 423588 275868
rect 423640 275856 423646 275868
rect 439406 275856 439412 275868
rect 423640 275828 439412 275856
rect 423640 275816 423646 275828
rect 439406 275816 439412 275828
rect 439464 275816 439470 275868
rect 443638 275816 443644 275868
rect 443696 275856 443702 275868
rect 498562 275856 498568 275868
rect 443696 275828 498568 275856
rect 443696 275816 443702 275828
rect 498562 275816 498568 275828
rect 498620 275816 498626 275868
rect 504726 275816 504732 275868
rect 504784 275856 504790 275868
rect 590746 275856 590752 275868
rect 504784 275828 590752 275856
rect 504784 275816 504790 275828
rect 590746 275816 590752 275828
rect 590804 275816 590810 275868
rect 260926 275748 260932 275800
rect 260984 275788 260990 275800
rect 263502 275788 263508 275800
rect 260984 275760 263508 275788
rect 260984 275748 260990 275760
rect 263502 275748 263508 275760
rect 263560 275748 263566 275800
rect 96614 275680 96620 275732
rect 96672 275720 96678 275732
rect 156598 275720 156604 275732
rect 96672 275692 156604 275720
rect 96672 275680 96678 275692
rect 156598 275680 156604 275692
rect 156656 275680 156662 275732
rect 174630 275680 174636 275732
rect 174688 275720 174694 275732
rect 208670 275720 208676 275732
rect 174688 275692 208676 275720
rect 174688 275680 174694 275692
rect 208670 275680 208676 275692
rect 208728 275680 208734 275732
rect 212442 275680 212448 275732
rect 212500 275720 212506 275732
rect 220538 275720 220544 275732
rect 212500 275692 220544 275720
rect 212500 275680 212506 275692
rect 220538 275680 220544 275692
rect 220596 275680 220602 275732
rect 232498 275680 232504 275732
rect 232556 275720 232562 275732
rect 232556 275692 243584 275720
rect 232556 275680 232562 275692
rect 220722 275612 220728 275664
rect 220780 275652 220786 275664
rect 224954 275652 224960 275664
rect 220780 275624 224960 275652
rect 220780 275612 220786 275624
rect 224954 275612 224960 275624
rect 225012 275612 225018 275664
rect 85942 275544 85948 275596
rect 86000 275584 86006 275596
rect 150802 275584 150808 275596
rect 86000 275556 150808 275584
rect 86000 275544 86006 275556
rect 150802 275544 150808 275556
rect 150860 275544 150866 275596
rect 160462 275544 160468 275596
rect 160520 275584 160526 275596
rect 172422 275584 172428 275596
rect 160520 275556 172428 275584
rect 160520 275544 160526 275556
rect 172422 275544 172428 275556
rect 172480 275544 172486 275596
rect 181714 275544 181720 275596
rect 181772 275584 181778 275596
rect 218606 275584 218612 275596
rect 181772 275556 218612 275584
rect 181772 275544 181778 275556
rect 218606 275544 218612 275556
rect 218664 275544 218670 275596
rect 225414 275544 225420 275596
rect 225472 275584 225478 275596
rect 242250 275584 242256 275596
rect 225472 275556 242256 275584
rect 225472 275544 225478 275556
rect 242250 275544 242256 275556
rect 242308 275544 242314 275596
rect 243556 275584 243584 275692
rect 244366 275680 244372 275732
rect 244424 275720 244430 275732
rect 247034 275720 247040 275732
rect 244424 275692 247040 275720
rect 244424 275680 244430 275692
rect 247034 275680 247040 275692
rect 247092 275680 247098 275732
rect 268010 275680 268016 275732
rect 268068 275720 268074 275732
rect 269114 275720 269120 275732
rect 268068 275692 269120 275720
rect 268068 275680 268074 275692
rect 269114 275680 269120 275692
rect 269172 275680 269178 275732
rect 365898 275680 365904 275732
rect 365956 275720 365962 275732
rect 369670 275720 369676 275732
rect 365956 275692 369676 275720
rect 365956 275680 365962 275692
rect 369670 275680 369676 275692
rect 369728 275680 369734 275732
rect 373074 275680 373080 275732
rect 373132 275720 373138 275732
rect 385034 275720 385040 275732
rect 373132 275692 385040 275720
rect 373132 275680 373138 275692
rect 385034 275680 385040 275692
rect 385092 275680 385098 275732
rect 400214 275680 400220 275732
rect 400272 275720 400278 275732
rect 418154 275720 418160 275732
rect 400272 275692 418160 275720
rect 400272 275680 400278 275692
rect 418154 275680 418160 275692
rect 418212 275680 418218 275732
rect 418338 275680 418344 275732
rect 418396 275720 418402 275732
rect 435910 275720 435916 275732
rect 418396 275692 435916 275720
rect 418396 275680 418402 275692
rect 435910 275680 435916 275692
rect 435968 275680 435974 275732
rect 457438 275680 457444 275732
rect 457496 275720 457502 275732
rect 516226 275720 516232 275732
rect 457496 275692 516232 275720
rect 457496 275680 457502 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 516686 275680 516692 275732
rect 516744 275720 516750 275732
rect 604914 275720 604920 275732
rect 516744 275692 604920 275720
rect 516744 275680 516750 275692
rect 604914 275680 604920 275692
rect 604972 275680 604978 275732
rect 605098 275680 605104 275732
rect 605156 275720 605162 275732
rect 616782 275720 616788 275732
rect 605156 275692 616788 275720
rect 605156 275680 605162 275692
rect 616782 275680 616788 275692
rect 616840 275680 616846 275732
rect 245654 275584 245660 275596
rect 243556 275556 245660 275584
rect 245654 275544 245660 275556
rect 245712 275544 245718 275596
rect 347406 275544 347412 275596
rect 347464 275584 347470 275596
rect 349614 275584 349620 275596
rect 347464 275556 349620 275584
rect 347464 275544 347470 275556
rect 349614 275544 349620 275556
rect 349672 275544 349678 275596
rect 352374 275544 352380 275596
rect 352432 275584 352438 275596
rect 360194 275584 360200 275596
rect 352432 275556 360200 275584
rect 352432 275544 352438 275556
rect 360194 275544 360200 275556
rect 360252 275544 360258 275596
rect 376570 275544 376576 275596
rect 376628 275584 376634 275596
rect 393314 275584 393320 275596
rect 376628 275556 393320 275584
rect 376628 275544 376634 275556
rect 393314 275544 393320 275556
rect 393372 275544 393378 275596
rect 395062 275544 395068 275596
rect 395120 275584 395126 275596
rect 403986 275584 403992 275596
rect 395120 275556 403992 275584
rect 395120 275544 395126 275556
rect 403986 275544 403992 275556
rect 404044 275544 404050 275596
rect 407666 275544 407672 275596
rect 407724 275584 407730 275596
rect 432322 275584 432328 275596
rect 407724 275556 432328 275584
rect 407724 275544 407730 275556
rect 432322 275544 432328 275556
rect 432380 275544 432386 275596
rect 438854 275544 438860 275596
rect 438912 275584 438918 275596
rect 446490 275584 446496 275596
rect 438912 275556 446496 275584
rect 438912 275544 438918 275556
rect 446490 275544 446496 275556
rect 446548 275544 446554 275596
rect 453942 275544 453948 275596
rect 454000 275584 454006 275596
rect 464246 275584 464252 275596
rect 454000 275556 464252 275584
rect 454000 275544 454006 275556
rect 464246 275544 464252 275556
rect 464304 275544 464310 275596
rect 464430 275544 464436 275596
rect 464488 275584 464494 275596
rect 523402 275584 523408 275596
rect 464488 275556 523408 275584
rect 464488 275544 464494 275556
rect 523402 275544 523408 275556
rect 523460 275544 523466 275596
rect 525794 275544 525800 275596
rect 525852 275584 525858 275596
rect 527358 275584 527364 275596
rect 525852 275556 527364 275584
rect 525852 275544 525858 275556
rect 527358 275544 527364 275556
rect 527416 275544 527422 275596
rect 532694 275544 532700 275596
rect 532752 275584 532758 275596
rect 626166 275584 626172 275596
rect 532752 275556 626172 275584
rect 532752 275544 532758 275556
rect 626166 275544 626172 275556
rect 626224 275544 626230 275596
rect 76466 275408 76472 275460
rect 76524 275448 76530 275460
rect 143258 275448 143264 275460
rect 76524 275420 143264 275448
rect 76524 275408 76530 275420
rect 143258 275408 143264 275420
rect 143316 275408 143322 275460
rect 148594 275408 148600 275460
rect 148652 275448 148658 275460
rect 164142 275448 164148 275460
rect 148652 275420 164148 275448
rect 148652 275408 148658 275420
rect 164142 275408 164148 275420
rect 164200 275408 164206 275460
rect 167546 275408 167552 275460
rect 167604 275448 167610 275460
rect 209038 275448 209044 275460
rect 167604 275420 209044 275448
rect 167604 275408 167610 275420
rect 209038 275408 209044 275420
rect 209096 275408 209102 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 239398 275448 239404 275460
rect 218388 275420 239404 275448
rect 218388 275408 218394 275420
rect 239398 275408 239404 275420
rect 239456 275408 239462 275460
rect 253842 275408 253848 275460
rect 253900 275448 253906 275460
rect 261478 275448 261484 275460
rect 253900 275420 261484 275448
rect 253900 275408 253906 275420
rect 261478 275408 261484 275420
rect 261536 275408 261542 275460
rect 349706 275408 349712 275460
rect 349764 275448 349770 275460
rect 361390 275448 361396 275460
rect 349764 275420 361396 275448
rect 349764 275408 349770 275420
rect 361390 275408 361396 275420
rect 361448 275408 361454 275460
rect 362954 275408 362960 275460
rect 363012 275448 363018 275460
rect 367278 275448 367284 275460
rect 363012 275420 367284 275448
rect 363012 275408 363018 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 367830 275408 367836 275460
rect 367888 275448 367894 275460
rect 377950 275448 377956 275460
rect 367888 275420 377956 275448
rect 367888 275408 367894 275420
rect 377950 275408 377956 275420
rect 378008 275408 378014 275460
rect 382458 275408 382464 275460
rect 382516 275448 382522 275460
rect 400398 275448 400404 275460
rect 382516 275420 400404 275448
rect 382516 275408 382522 275420
rect 400398 275408 400404 275420
rect 400456 275408 400462 275460
rect 403618 275408 403624 275460
rect 403676 275448 403682 275460
rect 428826 275448 428832 275460
rect 403676 275420 428832 275448
rect 403676 275408 403682 275420
rect 428826 275408 428832 275420
rect 428884 275408 428890 275460
rect 435726 275408 435732 275460
rect 435784 275448 435790 275460
rect 491478 275448 491484 275460
rect 435784 275420 491484 275448
rect 435784 275408 435790 275420
rect 491478 275408 491484 275420
rect 491536 275408 491542 275460
rect 494054 275408 494060 275460
rect 494112 275448 494118 275460
rect 502058 275448 502064 275460
rect 494112 275420 502064 275448
rect 494112 275408 494118 275420
rect 502058 275408 502064 275420
rect 502116 275408 502122 275460
rect 505830 275408 505836 275460
rect 505888 275448 505894 275460
rect 512730 275448 512736 275460
rect 505888 275420 512736 275448
rect 505888 275408 505894 275420
rect 512730 275408 512736 275420
rect 512788 275408 512794 275460
rect 525610 275408 525616 275460
rect 525668 275448 525674 275460
rect 619082 275448 619088 275460
rect 525668 275420 619088 275448
rect 525668 275408 525674 275420
rect 619082 275408 619088 275420
rect 619140 275408 619146 275460
rect 626442 275408 626448 275460
rect 626500 275448 626506 275460
rect 640426 275448 640432 275460
rect 626500 275420 640432 275448
rect 626500 275408 626506 275420
rect 640426 275408 640432 275420
rect 640484 275408 640490 275460
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 156874 275272 156880 275324
rect 156932 275312 156938 275324
rect 199286 275312 199292 275324
rect 156932 275284 199292 275312
rect 156932 275272 156938 275284
rect 199286 275272 199292 275284
rect 199344 275272 199350 275324
rect 211246 275272 211252 275324
rect 211304 275312 211310 275324
rect 232682 275312 232688 275324
rect 211304 275284 232688 275312
rect 211304 275272 211310 275284
rect 232682 275272 232688 275284
rect 232740 275272 232746 275324
rect 259730 275272 259736 275324
rect 259788 275312 259794 275324
rect 268838 275312 268844 275324
rect 259788 275284 268844 275312
rect 259788 275272 259794 275284
rect 268838 275272 268844 275284
rect 268896 275272 268902 275324
rect 276290 275272 276296 275324
rect 276348 275312 276354 275324
rect 284294 275312 284300 275324
rect 276348 275284 284300 275312
rect 276348 275272 276354 275284
rect 284294 275272 284300 275284
rect 284352 275272 284358 275324
rect 284570 275272 284576 275324
rect 284628 275312 284634 275324
rect 290090 275312 290096 275324
rect 284628 275284 290096 275312
rect 284628 275272 284634 275284
rect 290090 275272 290096 275284
rect 290148 275272 290154 275324
rect 339126 275272 339132 275324
rect 339184 275312 339190 275324
rect 353110 275312 353116 275324
rect 339184 275284 353116 275312
rect 339184 275272 339190 275284
rect 353110 275272 353116 275284
rect 353168 275272 353174 275324
rect 359458 275272 359464 275324
rect 359516 275312 359522 275324
rect 370866 275312 370872 275324
rect 359516 275284 370872 275312
rect 359516 275272 359522 275284
rect 370866 275272 370872 275284
rect 370924 275272 370930 275324
rect 377398 275272 377404 275324
rect 377456 275312 377462 275324
rect 396902 275312 396908 275324
rect 377456 275284 396908 275312
rect 377456 275272 377462 275284
rect 396902 275272 396908 275284
rect 396960 275272 396966 275324
rect 400398 275272 400404 275324
rect 400456 275312 400462 275324
rect 425238 275312 425244 275324
rect 400456 275284 425244 275312
rect 400456 275272 400462 275284
rect 425238 275272 425244 275284
rect 425296 275272 425302 275324
rect 427814 275272 427820 275324
rect 427872 275312 427878 275324
rect 442994 275312 443000 275324
rect 427872 275284 443000 275312
rect 427872 275272 427878 275284
rect 442994 275272 443000 275284
rect 443052 275272 443058 275324
rect 448238 275272 448244 275324
rect 448296 275312 448302 275324
rect 509142 275312 509148 275324
rect 448296 275284 509148 275312
rect 448296 275272 448302 275284
rect 509142 275272 509148 275284
rect 509200 275272 509206 275324
rect 513742 275272 513748 275324
rect 513800 275312 513806 275324
rect 533982 275312 533988 275324
rect 513800 275284 533988 275312
rect 513800 275272 513806 275284
rect 533982 275272 533988 275284
rect 534040 275272 534046 275324
rect 539502 275272 539508 275324
rect 539560 275312 539566 275324
rect 542262 275312 542268 275324
rect 539560 275284 542268 275312
rect 539560 275272 539566 275284
rect 542262 275272 542268 275284
rect 542320 275272 542326 275324
rect 543274 275272 543280 275324
rect 543332 275312 543338 275324
rect 645118 275312 645124 275324
rect 543332 275284 645124 275312
rect 543332 275272 543338 275284
rect 645118 275272 645124 275284
rect 645176 275272 645182 275324
rect 249058 275204 249064 275256
rect 249116 275244 249122 275256
rect 253566 275244 253572 275256
rect 249116 275216 253572 275244
rect 249116 275204 249122 275216
rect 253566 275204 253572 275216
rect 253624 275204 253630 275256
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 164970 275176 164976 275188
rect 110840 275148 164976 275176
rect 110840 275136 110846 275148
rect 164970 275136 164976 275148
rect 165028 275136 165034 275188
rect 171042 275136 171048 275188
rect 171100 275176 171106 275188
rect 191098 275176 191104 275188
rect 171100 275148 191104 275176
rect 171100 275136 171106 275148
rect 191098 275136 191104 275148
rect 191156 275136 191162 275188
rect 429194 275136 429200 275188
rect 429252 275176 429258 275188
rect 480806 275176 480812 275188
rect 429252 275148 480812 275176
rect 429252 275136 429258 275148
rect 480806 275136 480812 275148
rect 480864 275136 480870 275188
rect 487154 275136 487160 275188
rect 487212 275176 487218 275188
rect 544654 275176 544660 275188
rect 487212 275148 544660 275176
rect 487212 275136 487218 275148
rect 544654 275136 544660 275148
rect 544712 275136 544718 275188
rect 552566 275136 552572 275188
rect 552624 275176 552630 275188
rect 560018 275176 560024 275188
rect 552624 275148 560024 275176
rect 552624 275136 552630 275148
rect 560018 275136 560024 275148
rect 560076 275136 560082 275188
rect 246758 275068 246764 275120
rect 246816 275108 246822 275120
rect 256694 275108 256700 275120
rect 246816 275080 256700 275108
rect 246816 275068 246822 275080
rect 256694 275068 256700 275080
rect 256752 275068 256758 275120
rect 270402 275068 270408 275120
rect 270460 275108 270466 275120
rect 276198 275108 276204 275120
rect 270460 275080 276204 275108
rect 270460 275068 270466 275080
rect 276198 275068 276204 275080
rect 276256 275068 276262 275120
rect 580258 275068 580264 275120
rect 580316 275108 580322 275120
rect 583662 275108 583668 275120
rect 580316 275080 583668 275108
rect 580316 275068 580322 275080
rect 583662 275068 583668 275080
rect 583720 275068 583726 275120
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 167638 275040 167644 275052
rect 135680 275012 167644 275040
rect 135680 275000 135686 275012
rect 167638 275000 167644 275012
rect 167696 275000 167702 275052
rect 426250 275000 426256 275052
rect 426308 275040 426314 275052
rect 477218 275040 477224 275052
rect 426308 275012 477224 275040
rect 426308 275000 426314 275012
rect 477218 275000 477224 275012
rect 477276 275000 477282 275052
rect 485038 275000 485044 275052
rect 485096 275040 485102 275052
rect 494054 275040 494060 275052
rect 485096 275012 494060 275040
rect 485096 275000 485102 275012
rect 494054 275000 494060 275012
rect 494112 275000 494118 275052
rect 494422 275000 494428 275052
rect 494480 275040 494486 275052
rect 537294 275040 537300 275052
rect 494480 275012 537300 275040
rect 494480 275000 494486 275012
rect 537294 275000 537300 275012
rect 537352 275000 537358 275052
rect 537662 275000 537668 275052
rect 537720 275040 537726 275052
rect 538766 275040 538772 275052
rect 537720 275012 538772 275040
rect 537720 275000 537726 275012
rect 538766 275000 538772 275012
rect 538824 275000 538830 275052
rect 541986 275000 541992 275052
rect 542044 275040 542050 275052
rect 549346 275040 549352 275052
rect 542044 275012 549352 275040
rect 542044 275000 542050 275012
rect 549346 275000 549352 275012
rect 549404 275000 549410 275052
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 86218 274972 86224 274984
rect 81308 274944 86224 274972
rect 81308 274932 81314 274944
rect 86218 274932 86224 274944
rect 86276 274932 86282 274984
rect 241974 274932 241980 274984
rect 242032 274972 242038 274984
rect 244090 274972 244096 274984
rect 242032 274944 244096 274972
rect 242032 274932 242038 274944
rect 244090 274932 244096 274944
rect 244148 274932 244154 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136082 274904 136088 274916
rect 129700 274876 136088 274904
rect 129700 274864 129706 274876
rect 136082 274864 136088 274876
rect 136140 274864 136146 274916
rect 142706 274864 142712 274916
rect 142764 274904 142770 274916
rect 166258 274904 166264 274916
rect 142764 274876 166264 274904
rect 142764 274864 142770 274876
rect 166258 274864 166264 274876
rect 166316 274864 166322 274916
rect 210050 274864 210056 274916
rect 210108 274904 210114 274916
rect 212442 274904 212448 274916
rect 210108 274876 212448 274904
rect 210108 274864 210114 274876
rect 212442 274864 212448 274876
rect 212500 274864 212506 274916
rect 418522 274864 418528 274916
rect 418580 274904 418586 274916
rect 422846 274904 422852 274916
rect 418580 274876 422852 274904
rect 418580 274864 418586 274876
rect 422846 274864 422852 274876
rect 422904 274864 422910 274916
rect 478966 274864 478972 274916
rect 479024 274904 479030 274916
rect 482002 274904 482008 274916
rect 479024 274876 482008 274904
rect 479024 274864 479030 274876
rect 482002 274864 482008 274876
rect 482060 274864 482066 274916
rect 487798 274864 487804 274916
rect 487856 274904 487862 274916
rect 530486 274904 530492 274916
rect 487856 274876 530492 274904
rect 487856 274864 487862 274876
rect 530486 274864 530492 274876
rect 530544 274864 530550 274916
rect 530670 274864 530676 274916
rect 530728 274904 530734 274916
rect 541066 274904 541072 274916
rect 530728 274876 541072 274904
rect 530728 274864 530734 274876
rect 541066 274864 541072 274876
rect 541124 274864 541130 274916
rect 545114 274864 545120 274916
rect 545172 274904 545178 274916
rect 552934 274904 552940 274916
rect 545172 274876 552940 274904
rect 545172 274864 545178 274876
rect 552934 274864 552940 274876
rect 552992 274864 552998 274916
rect 559190 274864 559196 274916
rect 559248 274904 559254 274916
rect 567010 274904 567016 274916
rect 559248 274876 567016 274904
rect 559248 274864 559254 274876
rect 567010 274864 567016 274876
rect 567068 274864 567074 274916
rect 199470 274796 199476 274848
rect 199528 274836 199534 274848
rect 202782 274836 202788 274848
rect 199528 274808 202788 274836
rect 199528 274796 199534 274808
rect 202782 274796 202788 274808
rect 202840 274796 202846 274848
rect 243170 274796 243176 274848
rect 243228 274836 243234 274848
rect 249058 274836 249064 274848
rect 243228 274808 249064 274836
rect 243228 274796 243234 274808
rect 249058 274796 249064 274808
rect 249116 274796 249122 274848
rect 263226 274796 263232 274848
rect 263284 274836 263290 274848
rect 266446 274836 266452 274848
rect 263284 274808 266452 274836
rect 263284 274796 263290 274808
rect 266446 274796 266452 274808
rect 266504 274796 266510 274848
rect 277486 274796 277492 274848
rect 277544 274836 277550 274848
rect 283190 274836 283196 274848
rect 277544 274808 283196 274836
rect 277544 274796 277550 274808
rect 283190 274796 283196 274808
rect 283248 274796 283254 274848
rect 289262 274796 289268 274848
rect 289320 274836 289326 274848
rect 293402 274836 293408 274848
rect 289320 274808 293408 274836
rect 289320 274796 289326 274808
rect 293402 274796 293408 274808
rect 293460 274796 293466 274848
rect 336642 274796 336648 274848
rect 336700 274836 336706 274848
rect 343634 274836 343640 274848
rect 336700 274808 343640 274836
rect 336700 274796 336706 274808
rect 343634 274796 343640 274808
rect 343692 274796 343698 274848
rect 369854 274796 369860 274848
rect 369912 274836 369918 274848
rect 375558 274836 375564 274848
rect 369912 274808 375564 274836
rect 369912 274796 369918 274808
rect 375558 274796 375564 274808
rect 375616 274796 375622 274848
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149698 274768 149704 274780
rect 146260 274740 149704 274768
rect 146260 274728 146266 274740
rect 149698 274728 149704 274740
rect 149756 274728 149762 274780
rect 150986 274728 150992 274780
rect 151044 274768 151050 274780
rect 152734 274768 152740 274780
rect 151044 274740 152740 274768
rect 151044 274728 151050 274740
rect 152734 274728 152740 274740
rect 152792 274728 152798 274780
rect 163958 274728 163964 274780
rect 164016 274768 164022 274780
rect 170398 274768 170404 274780
rect 164016 274740 170404 274768
rect 164016 274728 164022 274740
rect 170398 274728 170404 274740
rect 170456 274728 170462 274780
rect 172238 274728 172244 274780
rect 172296 274768 172302 274780
rect 174906 274768 174912 274780
rect 172296 274740 174912 274768
rect 172296 274728 172302 274740
rect 174906 274728 174912 274740
rect 174964 274728 174970 274780
rect 208854 274728 208860 274780
rect 208912 274768 208918 274780
rect 210602 274768 210608 274780
rect 208912 274740 210608 274768
rect 208912 274728 208918 274740
rect 210602 274728 210608 274740
rect 210660 274728 210666 274780
rect 415302 274728 415308 274780
rect 415360 274768 415366 274780
rect 419350 274768 419356 274780
rect 415360 274740 419356 274768
rect 415360 274728 415366 274740
rect 419350 274728 419356 274740
rect 419408 274728 419414 274780
rect 423030 274728 423036 274780
rect 423088 274768 423094 274780
rect 424042 274768 424048 274780
rect 423088 274740 424048 274768
rect 423088 274728 423094 274740
rect 424042 274728 424048 274740
rect 424100 274728 424106 274780
rect 471882 274728 471888 274780
rect 471940 274768 471946 274780
rect 496170 274768 496176 274780
rect 471940 274740 496176 274768
rect 471940 274728 471946 274740
rect 496170 274728 496176 274740
rect 496228 274728 496234 274780
rect 510522 274728 510528 274780
rect 510580 274768 510586 274780
rect 519814 274768 519820 274780
rect 510580 274740 519820 274768
rect 510580 274728 510586 274740
rect 519814 274728 519820 274740
rect 519872 274728 519878 274780
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 545850 274768 545856 274780
rect 523736 274740 545856 274768
rect 523736 274728 523742 274740
rect 545850 274728 545856 274740
rect 545908 274728 545914 274780
rect 551278 274728 551284 274780
rect 551336 274768 551342 274780
rect 574186 274768 574192 274780
rect 551336 274740 574192 274768
rect 551336 274728 551342 274740
rect 574186 274728 574192 274740
rect 574244 274728 574250 274780
rect 71774 274660 71780 274712
rect 71832 274700 71838 274712
rect 73798 274700 73804 274712
rect 71832 274672 73804 274700
rect 71832 274660 71838 274672
rect 73798 274660 73804 274672
rect 73856 274660 73862 274712
rect 74074 274660 74080 274712
rect 74132 274700 74138 274712
rect 77202 274700 77208 274712
rect 74132 274672 77208 274700
rect 74132 274660 74138 274672
rect 77202 274660 77208 274672
rect 77260 274660 77266 274712
rect 257338 274660 257344 274712
rect 257396 274700 257402 274712
rect 260190 274700 260196 274712
rect 257396 274672 260196 274700
rect 257396 274660 257402 274672
rect 260190 274660 260196 274672
rect 260248 274660 260254 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294322 274700 294328 274712
rect 290516 274672 294328 274700
rect 290516 274660 290522 274672
rect 294322 274660 294328 274672
rect 294380 274660 294386 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 298738 274660 298744 274712
rect 298796 274700 298802 274712
rect 300118 274700 300124 274712
rect 298796 274672 300124 274700
rect 298796 274660 298802 274672
rect 300118 274660 300124 274672
rect 300176 274660 300182 274712
rect 324958 274660 324964 274712
rect 325016 274700 325022 274712
rect 327074 274700 327080 274712
rect 325016 274672 327080 274700
rect 325016 274660 325022 274672
rect 327074 274660 327080 274672
rect 327132 274660 327138 274712
rect 331398 274660 331404 274712
rect 331456 274700 331462 274712
rect 335354 274700 335360 274712
rect 331456 274672 335360 274700
rect 331456 274660 331462 274672
rect 335354 274660 335360 274672
rect 335412 274660 335418 274712
rect 337102 274660 337108 274712
rect 337160 274700 337166 274712
rect 338942 274700 338948 274712
rect 337160 274672 338948 274700
rect 337160 274660 337166 274672
rect 338942 274660 338948 274672
rect 339000 274660 339006 274712
rect 344278 274660 344284 274712
rect 344336 274700 344342 274712
rect 347222 274700 347228 274712
rect 344336 274672 347228 274700
rect 344336 274660 344342 274672
rect 347222 274660 347228 274672
rect 347280 274660 347286 274712
rect 360194 274660 360200 274712
rect 360252 274700 360258 274712
rect 363782 274700 363788 274712
rect 360252 274672 363788 274700
rect 360252 274660 360258 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 368750 274660 368756 274712
rect 368808 274700 368814 274712
rect 373258 274700 373264 274712
rect 368808 274672 373264 274700
rect 368808 274660 368814 274672
rect 373258 274660 373264 274672
rect 373316 274660 373322 274712
rect 453574 274700 453580 274712
rect 446416 274672 453580 274700
rect 120258 274592 120264 274644
rect 120316 274632 120322 274644
rect 175274 274632 175280 274644
rect 120316 274604 175280 274632
rect 120316 274592 120322 274604
rect 175274 274592 175280 274604
rect 175332 274592 175338 274644
rect 204714 274592 204720 274644
rect 204772 274632 204778 274644
rect 218790 274632 218796 274644
rect 204772 274604 218796 274632
rect 204772 274592 204778 274604
rect 218790 274592 218796 274604
rect 218848 274592 218854 274644
rect 403986 274592 403992 274644
rect 404044 274632 404050 274644
rect 438854 274632 438860 274644
rect 404044 274604 438860 274632
rect 404044 274592 404050 274604
rect 438854 274592 438860 274604
rect 438912 274592 438918 274644
rect 114278 274456 114284 274508
rect 114336 274496 114342 274508
rect 171594 274496 171600 274508
rect 114336 274468 171600 274496
rect 114336 274456 114342 274468
rect 171594 274456 171600 274468
rect 171652 274456 171658 274508
rect 179322 274456 179328 274508
rect 179380 274496 179386 274508
rect 213178 274496 213184 274508
rect 179380 274468 213184 274496
rect 179380 274456 179386 274468
rect 213178 274456 213184 274468
rect 213236 274456 213242 274508
rect 378778 274456 378784 274508
rect 378836 274496 378842 274508
rect 395706 274496 395712 274508
rect 378836 274468 395712 274496
rect 378836 274456 378842 274468
rect 395706 274456 395712 274468
rect 395764 274456 395770 274508
rect 409230 274456 409236 274508
rect 409288 274496 409294 274508
rect 446416 274496 446444 274672
rect 453574 274660 453580 274672
rect 453632 274660 453638 274712
rect 498470 274660 498476 274712
rect 498528 274700 498534 274712
rect 499758 274700 499764 274712
rect 498528 274672 499764 274700
rect 498528 274660 498534 274672
rect 499758 274660 499764 274672
rect 499816 274660 499822 274712
rect 501598 274660 501604 274712
rect 501656 274700 501662 274712
rect 505646 274700 505652 274712
rect 501656 274672 505652 274700
rect 501656 274660 501662 274672
rect 505646 274660 505652 274672
rect 505704 274660 505710 274712
rect 506474 274660 506480 274712
rect 506532 274700 506538 274712
rect 510338 274700 510344 274712
rect 506532 274672 510344 274700
rect 506532 274660 506538 274672
rect 510338 274660 510344 274672
rect 510396 274660 510402 274712
rect 619174 274660 619180 274712
rect 619232 274700 619238 274712
rect 623866 274700 623872 274712
rect 619232 274672 623872 274700
rect 619232 274660 619238 274672
rect 623866 274660 623872 274672
rect 623924 274660 623930 274712
rect 458818 274592 458824 274644
rect 458876 274632 458882 274644
rect 484302 274632 484308 274644
rect 458876 274604 484308 274632
rect 458876 274592 458882 274604
rect 484302 274592 484308 274604
rect 484360 274592 484366 274644
rect 493134 274592 493140 274644
rect 493192 274632 493198 274644
rect 494422 274632 494428 274644
rect 493192 274604 494428 274632
rect 493192 274592 493198 274604
rect 494422 274592 494428 274604
rect 494480 274592 494486 274644
rect 522390 274592 522396 274644
rect 522448 274632 522454 274644
rect 595438 274632 595444 274644
rect 522448 274604 595444 274632
rect 522448 274592 522454 274604
rect 595438 274592 595444 274604
rect 595496 274592 595502 274644
rect 409288 274468 446444 274496
rect 409288 274456 409294 274468
rect 453298 274456 453304 274508
rect 453356 274496 453362 274508
rect 478414 274496 478420 274508
rect 453356 274468 478420 274496
rect 453356 274456 453362 274468
rect 478414 274456 478420 274468
rect 478472 274456 478478 274508
rect 481358 274456 481364 274508
rect 481416 274496 481422 274508
rect 556430 274496 556436 274508
rect 481416 274468 556436 274496
rect 481416 274456 481422 274468
rect 556430 274456 556436 274468
rect 556488 274456 556494 274508
rect 559558 274456 559564 274508
rect 559616 274496 559622 274508
rect 587158 274496 587164 274508
rect 559616 274468 587164 274496
rect 559616 274456 559622 274468
rect 587158 274456 587164 274468
rect 587216 274456 587222 274508
rect 93026 274320 93032 274372
rect 93084 274360 93090 274372
rect 95878 274360 95884 274372
rect 93084 274332 95884 274360
rect 93084 274320 93090 274332
rect 95878 274320 95884 274332
rect 95936 274320 95942 274372
rect 97718 274320 97724 274372
rect 97776 274360 97782 274372
rect 158806 274360 158812 274372
rect 97776 274332 158812 274360
rect 97776 274320 97782 274332
rect 158806 274320 158812 274332
rect 158864 274320 158870 274372
rect 180518 274320 180524 274372
rect 180576 274360 180582 274372
rect 216950 274360 216956 274372
rect 180576 274332 216956 274360
rect 180576 274320 180582 274332
rect 216950 274320 216956 274332
rect 217008 274320 217014 274372
rect 223114 274320 223120 274372
rect 223172 274360 223178 274372
rect 247218 274360 247224 274372
rect 223172 274332 247224 274360
rect 223172 274320 223178 274332
rect 247218 274320 247224 274332
rect 247276 274320 247282 274372
rect 384942 274320 384948 274372
rect 385000 274360 385006 274372
rect 400214 274360 400220 274372
rect 385000 274332 400220 274360
rect 385000 274320 385006 274332
rect 400214 274320 400220 274332
rect 400272 274320 400278 274372
rect 416590 274320 416596 274372
rect 416648 274360 416654 274372
rect 453942 274360 453948 274372
rect 416648 274332 453948 274360
rect 416648 274320 416654 274332
rect 453942 274320 453948 274332
rect 454000 274320 454006 274372
rect 474366 274320 474372 274372
rect 474424 274360 474430 274372
rect 523678 274360 523684 274372
rect 474424 274332 523684 274360
rect 474424 274320 474430 274332
rect 523678 274320 523684 274332
rect 523736 274320 523742 274372
rect 537478 274320 537484 274372
rect 537536 274360 537542 274372
rect 613194 274360 613200 274372
rect 537536 274332 613200 274360
rect 537536 274320 537542 274332
rect 613194 274320 613200 274332
rect 613252 274320 613258 274372
rect 95418 274184 95424 274236
rect 95476 274224 95482 274236
rect 157610 274224 157616 274236
rect 95476 274196 157616 274224
rect 95476 274184 95482 274196
rect 157610 274184 157616 274196
rect 157668 274184 157674 274236
rect 165614 274184 165620 274236
rect 165672 274224 165678 274236
rect 205726 274224 205732 274236
rect 165672 274196 205732 274224
rect 165672 274184 165678 274196
rect 205726 274184 205732 274196
rect 205784 274184 205790 274236
rect 213638 274184 213644 274236
rect 213696 274224 213702 274236
rect 240410 274224 240416 274236
rect 213696 274196 240416 274224
rect 213696 274184 213702 274196
rect 240410 274184 240416 274196
rect 240468 274184 240474 274236
rect 362770 274184 362776 274236
rect 362828 274224 362834 274236
rect 386230 274224 386236 274236
rect 362828 274196 386236 274224
rect 362828 274184 362834 274196
rect 386230 274184 386236 274196
rect 386288 274184 386294 274236
rect 400122 274184 400128 274236
rect 400180 274224 400186 274236
rect 423582 274224 423588 274236
rect 400180 274196 423588 274224
rect 400180 274184 400186 274196
rect 423582 274184 423588 274196
rect 423640 274184 423646 274236
rect 427446 274184 427452 274236
rect 427504 274224 427510 274236
rect 479334 274224 479340 274236
rect 427504 274196 479340 274224
rect 427504 274184 427510 274196
rect 479334 274184 479340 274196
rect 479392 274184 479398 274236
rect 486970 274184 486976 274236
rect 487028 274224 487034 274236
rect 563514 274224 563520 274236
rect 487028 274196 563520 274224
rect 487028 274184 487034 274196
rect 563514 274184 563520 274196
rect 563572 274184 563578 274236
rect 563698 274184 563704 274236
rect 563756 274224 563762 274236
rect 611998 274224 612004 274236
rect 563756 274196 612004 274224
rect 563756 274184 563762 274196
rect 611998 274184 612004 274196
rect 612056 274184 612062 274236
rect 75270 274048 75276 274100
rect 75328 274088 75334 274100
rect 142154 274088 142160 274100
rect 75328 274060 142160 274088
rect 75328 274048 75334 274060
rect 142154 274048 142160 274060
rect 142212 274048 142218 274100
rect 147398 274048 147404 274100
rect 147456 274088 147462 274100
rect 193306 274088 193312 274100
rect 147456 274060 193312 274088
rect 147456 274048 147462 274060
rect 193306 274048 193312 274060
rect 193364 274048 193370 274100
rect 193490 274048 193496 274100
rect 193548 274088 193554 274100
rect 204714 274088 204720 274100
rect 193548 274060 204720 274088
rect 193548 274048 193554 274060
rect 204714 274048 204720 274060
rect 204772 274048 204778 274100
rect 206554 274048 206560 274100
rect 206612 274088 206618 274100
rect 234614 274088 234620 274100
rect 206612 274060 234620 274088
rect 206612 274048 206618 274060
rect 234614 274048 234620 274060
rect 234672 274048 234678 274100
rect 245654 274048 245660 274100
rect 245712 274088 245718 274100
rect 254026 274088 254032 274100
rect 245712 274060 254032 274088
rect 245712 274048 245718 274060
rect 254026 274048 254032 274060
rect 254084 274048 254090 274100
rect 269114 274048 269120 274100
rect 269172 274088 269178 274100
rect 278774 274088 278780 274100
rect 269172 274060 278780 274088
rect 269172 274048 269178 274060
rect 278774 274048 278780 274060
rect 278832 274048 278838 274100
rect 349890 274048 349896 274100
rect 349948 274088 349954 274100
rect 362586 274088 362592 274100
rect 349948 274060 362592 274088
rect 349948 274048 349954 274060
rect 362586 274048 362592 274060
rect 362644 274048 362650 274100
rect 368290 274048 368296 274100
rect 368348 274088 368354 274100
rect 394510 274088 394516 274100
rect 368348 274060 394516 274088
rect 368348 274048 368354 274060
rect 394510 274048 394516 274060
rect 394568 274048 394574 274100
rect 395338 274048 395344 274100
rect 395396 274088 395402 274100
rect 426434 274088 426440 274100
rect 395396 274060 426440 274088
rect 395396 274048 395402 274060
rect 426434 274048 426440 274060
rect 426492 274048 426498 274100
rect 431678 274048 431684 274100
rect 431736 274088 431742 274100
rect 485498 274088 485504 274100
rect 431736 274060 485504 274088
rect 431736 274048 431742 274060
rect 485498 274048 485504 274060
rect 485556 274048 485562 274100
rect 529842 274048 529848 274100
rect 529900 274088 529906 274100
rect 532694 274088 532700 274100
rect 529900 274060 532700 274088
rect 529900 274048 529906 274060
rect 532694 274048 532700 274060
rect 532752 274048 532758 274100
rect 540882 274048 540888 274100
rect 540940 274088 540946 274100
rect 626442 274088 626448 274100
rect 540940 274060 626448 274088
rect 540940 274048 540946 274060
rect 626442 274048 626448 274060
rect 626500 274048 626506 274100
rect 77662 273912 77668 273964
rect 77720 273952 77726 273964
rect 145098 273952 145104 273964
rect 77720 273924 145104 273952
rect 77720 273912 77726 273924
rect 145098 273912 145104 273924
rect 145156 273912 145162 273964
rect 145282 273912 145288 273964
rect 145340 273952 145346 273964
rect 145340 273924 190454 273952
rect 145340 273912 145346 273924
rect 130838 273776 130844 273828
rect 130896 273816 130902 273828
rect 181438 273816 181444 273828
rect 130896 273788 181444 273816
rect 130896 273776 130902 273788
rect 181438 273776 181444 273788
rect 181496 273776 181502 273828
rect 190426 273816 190454 273924
rect 191834 273912 191840 273964
rect 191892 273952 191898 273964
rect 191892 273924 219434 273952
rect 191892 273912 191898 273924
rect 191834 273816 191840 273828
rect 190426 273788 191840 273816
rect 191834 273776 191840 273788
rect 191892 273776 191898 273828
rect 219406 273816 219434 273924
rect 224954 273912 224960 273964
rect 225012 273952 225018 273964
rect 245746 273952 245752 273964
rect 225012 273924 245752 273952
rect 225012 273912 225018 273924
rect 245746 273912 245752 273924
rect 245804 273912 245810 273964
rect 247034 273912 247040 273964
rect 247092 273952 247098 273964
rect 262214 273952 262220 273964
rect 247092 273924 262220 273952
rect 247092 273912 247098 273924
rect 262214 273912 262220 273924
rect 262272 273912 262278 273964
rect 263502 273912 263508 273964
rect 263560 273952 263566 273964
rect 273530 273952 273536 273964
rect 263560 273924 273536 273952
rect 263560 273912 263566 273924
rect 273530 273912 273536 273924
rect 273588 273912 273594 273964
rect 279786 273912 279792 273964
rect 279844 273952 279850 273964
rect 287146 273952 287152 273964
rect 279844 273924 287152 273952
rect 279844 273912 279850 273924
rect 287146 273912 287152 273924
rect 287204 273912 287210 273964
rect 333790 273912 333796 273964
rect 333848 273952 333854 273964
rect 344462 273952 344468 273964
rect 333848 273924 344468 273952
rect 333848 273912 333854 273924
rect 344462 273912 344468 273924
rect 344520 273912 344526 273964
rect 344646 273912 344652 273964
rect 344704 273952 344710 273964
rect 349706 273952 349712 273964
rect 344704 273924 349712 273952
rect 344704 273912 344710 273924
rect 349706 273912 349712 273924
rect 349764 273912 349770 273964
rect 365898 273952 365904 273964
rect 354646 273924 365904 273952
rect 224954 273816 224960 273828
rect 219406 273788 224960 273816
rect 224954 273776 224960 273788
rect 225012 273776 225018 273828
rect 350350 273776 350356 273828
rect 350408 273816 350414 273828
rect 354646 273816 354674 273924
rect 365898 273912 365904 273924
rect 365956 273912 365962 273964
rect 367002 273912 367008 273964
rect 367060 273952 367066 273964
rect 376570 273952 376576 273964
rect 367060 273924 376576 273952
rect 367060 273912 367066 273924
rect 376570 273912 376576 273924
rect 376628 273912 376634 273964
rect 407482 273952 407488 273964
rect 383626 273924 407488 273952
rect 350408 273788 354674 273816
rect 350408 273776 350414 273788
rect 376570 273776 376576 273828
rect 376628 273816 376634 273828
rect 383626 273816 383654 273924
rect 407482 273912 407488 273924
rect 407540 273912 407546 273964
rect 420730 273912 420736 273964
rect 420788 273952 420794 273964
rect 470134 273952 470140 273964
rect 420788 273924 470140 273952
rect 420788 273912 420794 273924
rect 470134 273912 470140 273924
rect 470192 273912 470198 273964
rect 470410 273912 470416 273964
rect 470468 273952 470474 273964
rect 539870 273952 539876 273964
rect 470468 273924 539876 273952
rect 470468 273912 470474 273924
rect 539870 273912 539876 273924
rect 539928 273912 539934 273964
rect 542170 273912 542176 273964
rect 542228 273952 542234 273964
rect 642726 273952 642732 273964
rect 542228 273924 642732 273952
rect 542228 273912 542234 273924
rect 642726 273912 642732 273924
rect 642784 273912 642790 273964
rect 376628 273788 383654 273816
rect 376628 273776 376634 273788
rect 397270 273776 397276 273828
rect 397328 273816 397334 273828
rect 418338 273816 418344 273828
rect 397328 273788 418344 273816
rect 397328 273776 397334 273788
rect 418338 273776 418344 273788
rect 418396 273776 418402 273828
rect 439314 273776 439320 273828
rect 439372 273816 439378 273828
rect 471330 273816 471336 273828
rect 439372 273788 471336 273816
rect 439372 273776 439378 273788
rect 471330 273776 471336 273788
rect 471388 273776 471394 273828
rect 473078 273776 473084 273828
rect 473136 273816 473142 273828
rect 487154 273816 487160 273828
rect 473136 273788 487160 273816
rect 473136 273776 473142 273788
rect 487154 273776 487160 273788
rect 487212 273776 487218 273828
rect 488350 273776 488356 273828
rect 488408 273816 488414 273828
rect 559190 273816 559196 273828
rect 488408 273788 559196 273816
rect 488408 273776 488414 273788
rect 559190 273776 559196 273788
rect 559248 273776 559254 273828
rect 124950 273640 124956 273692
rect 125008 273680 125014 273692
rect 148410 273680 148416 273692
rect 125008 273652 148416 273680
rect 125008 273640 125014 273652
rect 148410 273640 148416 273652
rect 148468 273640 148474 273692
rect 155678 273640 155684 273692
rect 155736 273680 155742 273692
rect 198090 273680 198096 273692
rect 155736 273652 198096 273680
rect 155736 273640 155742 273652
rect 198090 273640 198096 273652
rect 198148 273640 198154 273692
rect 438118 273640 438124 273692
rect 438176 273680 438182 273692
rect 467834 273680 467840 273692
rect 438176 273652 467840 273680
rect 438176 273640 438182 273652
rect 467834 273640 467840 273652
rect 467892 273640 467898 273692
rect 484302 273640 484308 273692
rect 484360 273680 484366 273692
rect 552566 273680 552572 273692
rect 484360 273652 552572 273680
rect 484360 273640 484366 273652
rect 552566 273640 552572 273652
rect 552624 273640 552630 273692
rect 446398 273504 446404 273556
rect 446456 273544 446462 273556
rect 468938 273544 468944 273556
rect 446456 273516 468944 273544
rect 446456 273504 446462 273516
rect 468938 273504 468944 273516
rect 468996 273504 469002 273556
rect 478782 273504 478788 273556
rect 478840 273544 478846 273556
rect 545114 273544 545120 273556
rect 478840 273516 545120 273544
rect 478840 273504 478846 273516
rect 545114 273504 545120 273516
rect 545172 273504 545178 273556
rect 552658 273504 552664 273556
rect 552716 273544 552722 273556
rect 580074 273544 580080 273556
rect 552716 273516 580080 273544
rect 552716 273504 552722 273516
rect 580074 273504 580080 273516
rect 580132 273504 580138 273556
rect 475746 273368 475752 273420
rect 475804 273408 475810 273420
rect 541986 273408 541992 273420
rect 475804 273380 541992 273408
rect 475804 273368 475810 273380
rect 541986 273368 541992 273380
rect 542044 273368 542050 273420
rect 330478 273232 330484 273284
rect 330536 273272 330542 273284
rect 333054 273272 333060 273284
rect 330536 273244 333060 273272
rect 330536 273232 330542 273244
rect 333054 273232 333060 273244
rect 333112 273232 333118 273284
rect 128538 273164 128544 273216
rect 128596 273204 128602 273216
rect 181254 273204 181260 273216
rect 128596 273176 181260 273204
rect 128596 273164 128602 273176
rect 181254 273164 181260 273176
rect 181312 273164 181318 273216
rect 268838 273164 268844 273216
rect 268896 273204 268902 273216
rect 272610 273204 272616 273216
rect 268896 273176 272616 273204
rect 268896 273164 268902 273176
rect 272610 273164 272616 273176
rect 272668 273164 272674 273216
rect 401502 273164 401508 273216
rect 401560 273204 401566 273216
rect 427814 273204 427820 273216
rect 401560 273176 427820 273204
rect 401560 273164 401566 273176
rect 427814 273164 427820 273176
rect 427872 273164 427878 273216
rect 438762 273164 438768 273216
rect 438820 273204 438826 273216
rect 471882 273204 471888 273216
rect 438820 273176 471888 273204
rect 438820 273164 438826 273176
rect 471882 273164 471888 273176
rect 471940 273164 471946 273216
rect 475930 273164 475936 273216
rect 475988 273204 475994 273216
rect 548150 273204 548156 273216
rect 475988 273176 548156 273204
rect 475988 273164 475994 273176
rect 548150 273164 548156 273176
rect 548208 273164 548214 273216
rect 111978 273028 111984 273080
rect 112036 273068 112042 273080
rect 168374 273068 168380 273080
rect 112036 273040 168380 273068
rect 112036 273028 112042 273040
rect 168374 273028 168380 273040
rect 168432 273028 168438 273080
rect 182082 273028 182088 273080
rect 182140 273068 182146 273080
rect 207290 273068 207296 273080
rect 182140 273040 207296 273068
rect 182140 273028 182146 273040
rect 207290 273028 207296 273040
rect 207348 273028 207354 273080
rect 217410 273068 217416 273080
rect 209746 273040 217416 273068
rect 102502 272892 102508 272944
rect 102560 272932 102566 272944
rect 162118 272932 162124 272944
rect 102560 272904 162124 272932
rect 102560 272892 102566 272904
rect 162118 272892 162124 272904
rect 162176 272892 162182 272944
rect 189994 272892 190000 272944
rect 190052 272932 190058 272944
rect 209746 272932 209774 273040
rect 217410 273028 217416 273040
rect 217468 273028 217474 273080
rect 381998 273028 382004 273080
rect 382056 273068 382062 273080
rect 414566 273068 414572 273080
rect 382056 273040 414572 273068
rect 382056 273028 382062 273040
rect 414566 273028 414572 273040
rect 414624 273028 414630 273080
rect 424962 273028 424968 273080
rect 425020 273068 425026 273080
rect 474918 273068 474924 273080
rect 425020 273040 474924 273068
rect 425020 273028 425026 273040
rect 474918 273028 474924 273040
rect 474976 273028 474982 273080
rect 500862 273028 500868 273080
rect 500920 273068 500926 273080
rect 580258 273068 580264 273080
rect 500920 273040 580264 273068
rect 500920 273028 500926 273040
rect 580258 273028 580264 273040
rect 580316 273028 580322 273080
rect 190052 272904 209774 272932
rect 190052 272892 190058 272904
rect 217134 272892 217140 272944
rect 217192 272932 217198 272944
rect 242894 272932 242900 272944
rect 217192 272904 242900 272932
rect 217192 272892 217198 272904
rect 242894 272892 242900 272904
rect 242952 272892 242958 272944
rect 388806 272892 388812 272944
rect 388864 272932 388870 272944
rect 400398 272932 400404 272944
rect 388864 272904 400404 272932
rect 388864 272892 388870 272904
rect 400398 272892 400404 272904
rect 400456 272892 400462 272944
rect 406838 272892 406844 272944
rect 406896 272932 406902 272944
rect 450078 272932 450084 272944
rect 406896 272904 450084 272932
rect 406896 272892 406902 272904
rect 450078 272892 450084 272904
rect 450136 272892 450142 272944
rect 451090 272892 451096 272944
rect 451148 272932 451154 272944
rect 513926 272932 513932 272944
rect 451148 272904 513932 272932
rect 451148 272892 451154 272904
rect 513926 272892 513932 272904
rect 513984 272892 513990 272944
rect 520090 272892 520096 272944
rect 520148 272932 520154 272944
rect 610802 272932 610808 272944
rect 520148 272904 610808 272932
rect 520148 272892 520154 272904
rect 610802 272892 610808 272904
rect 610860 272892 610866 272944
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 155954 272796 155960 272808
rect 94280 272768 155960 272796
rect 94280 272756 94286 272768
rect 155954 272756 155960 272768
rect 156012 272756 156018 272808
rect 187602 272756 187608 272808
rect 187660 272796 187666 272808
rect 220078 272796 220084 272808
rect 187660 272768 220084 272796
rect 187660 272756 187666 272768
rect 220078 272756 220084 272768
rect 220136 272756 220142 272808
rect 220538 272756 220544 272808
rect 220596 272796 220602 272808
rect 239214 272796 239220 272808
rect 220596 272768 239220 272796
rect 220596 272756 220602 272768
rect 239214 272756 239220 272768
rect 239272 272756 239278 272808
rect 343542 272756 343548 272808
rect 343600 272796 343606 272808
rect 358998 272796 359004 272808
rect 343600 272768 359004 272796
rect 343600 272756 343606 272768
rect 358998 272756 359004 272768
rect 359056 272756 359062 272808
rect 360838 272756 360844 272808
rect 360896 272796 360902 272808
rect 381538 272796 381544 272808
rect 360896 272768 381544 272796
rect 360896 272756 360902 272768
rect 381538 272756 381544 272768
rect 381596 272756 381602 272808
rect 394326 272756 394332 272808
rect 394384 272796 394390 272808
rect 407666 272796 407672 272808
rect 394384 272768 407672 272796
rect 394384 272756 394390 272768
rect 407666 272756 407672 272768
rect 407724 272756 407730 272808
rect 408126 272756 408132 272808
rect 408184 272796 408190 272808
rect 452102 272796 452108 272808
rect 408184 272768 452108 272796
rect 408184 272756 408190 272768
rect 452102 272756 452108 272768
rect 452160 272756 452166 272808
rect 452286 272756 452292 272808
rect 452344 272796 452350 272808
rect 515122 272796 515128 272808
rect 452344 272768 515128 272796
rect 452344 272756 452350 272768
rect 515122 272756 515128 272768
rect 515180 272756 515186 272808
rect 524046 272756 524052 272808
rect 524104 272796 524110 272808
rect 617978 272796 617984 272808
rect 524104 272768 617984 272796
rect 524104 272756 524110 272768
rect 617978 272756 617984 272768
rect 618036 272756 618042 272808
rect 82354 272620 82360 272672
rect 82412 272660 82418 272672
rect 148226 272660 148232 272672
rect 82412 272632 148232 272660
rect 82412 272620 82418 272632
rect 148226 272620 148232 272632
rect 148284 272620 148290 272672
rect 161566 272620 161572 272672
rect 161624 272660 161630 272672
rect 203058 272660 203064 272672
rect 161624 272632 203064 272660
rect 161624 272620 161630 272632
rect 203058 272620 203064 272632
rect 203116 272620 203122 272672
rect 203242 272620 203248 272672
rect 203300 272660 203306 272672
rect 233234 272660 233240 272672
rect 203300 272632 233240 272660
rect 203300 272620 203306 272632
rect 233234 272620 233240 272632
rect 233292 272620 233298 272672
rect 239582 272620 239588 272672
rect 239640 272660 239646 272672
rect 251818 272660 251824 272672
rect 239640 272632 251824 272660
rect 239640 272620 239646 272632
rect 251818 272620 251824 272632
rect 251876 272620 251882 272672
rect 252646 272620 252652 272672
rect 252704 272660 252710 272672
rect 252704 272632 267734 272660
rect 252704 272620 252710 272632
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 187694 272524 187700 272536
rect 137980 272496 187700 272524
rect 137980 272484 137986 272496
rect 187694 272484 187700 272496
rect 187752 272484 187758 272536
rect 192294 272484 192300 272536
rect 192352 272524 192358 272536
rect 225506 272524 225512 272536
rect 192352 272496 225512 272524
rect 192352 272484 192358 272496
rect 225506 272484 225512 272496
rect 225564 272484 225570 272536
rect 228818 272484 228824 272536
rect 228876 272524 228882 272536
rect 238018 272524 238024 272536
rect 228876 272496 238024 272524
rect 228876 272484 228882 272496
rect 238018 272484 238024 272496
rect 238076 272484 238082 272536
rect 238478 272484 238484 272536
rect 238536 272524 238542 272536
rect 258074 272524 258080 272536
rect 238536 272496 258080 272524
rect 238536 272484 238542 272496
rect 258074 272484 258080 272496
rect 258132 272484 258138 272536
rect 267706 272524 267734 272632
rect 347590 272620 347596 272672
rect 347648 272660 347654 272672
rect 366082 272660 366088 272672
rect 347648 272632 366088 272660
rect 347648 272620 347654 272632
rect 366082 272620 366088 272632
rect 366140 272620 366146 272672
rect 370958 272620 370964 272672
rect 371016 272660 371022 272672
rect 399202 272660 399208 272672
rect 371016 272632 399208 272660
rect 371016 272620 371022 272632
rect 399202 272620 399208 272632
rect 399260 272620 399266 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 457162 272660 457168 272672
rect 412324 272632 457168 272660
rect 412324 272620 412330 272632
rect 457162 272620 457168 272632
rect 457220 272620 457226 272672
rect 457990 272620 457996 272672
rect 458048 272660 458054 272672
rect 522206 272660 522212 272672
rect 458048 272632 522212 272660
rect 458048 272620 458054 272632
rect 522206 272620 522212 272632
rect 522264 272620 522270 272672
rect 526806 272620 526812 272672
rect 526864 272660 526870 272672
rect 621474 272660 621480 272672
rect 526864 272632 621480 272660
rect 526864 272620 526870 272632
rect 621474 272620 621480 272632
rect 621532 272620 621538 272672
rect 267826 272524 267832 272536
rect 267706 272496 267832 272524
rect 267826 272484 267832 272496
rect 267884 272484 267890 272536
rect 273898 272484 273904 272536
rect 273956 272524 273962 272536
rect 283006 272524 283012 272536
rect 273956 272496 283012 272524
rect 273956 272484 273962 272496
rect 283006 272484 283012 272496
rect 283064 272484 283070 272536
rect 322750 272484 322756 272536
rect 322808 272524 322814 272536
rect 330662 272524 330668 272536
rect 322808 272496 330668 272524
rect 322808 272484 322814 272496
rect 330662 272484 330668 272496
rect 330720 272484 330726 272536
rect 331030 272484 331036 272536
rect 331088 272524 331094 272536
rect 342438 272524 342444 272536
rect 331088 272496 342444 272524
rect 331088 272484 331094 272496
rect 342438 272484 342444 272496
rect 342496 272484 342502 272536
rect 356698 272484 356704 272536
rect 356756 272524 356762 272536
rect 376754 272524 376760 272536
rect 356756 272496 376760 272524
rect 356756 272484 356762 272496
rect 376754 272484 376760 272496
rect 376812 272484 376818 272536
rect 380802 272484 380808 272536
rect 380860 272524 380866 272536
rect 411990 272524 411996 272536
rect 380860 272496 411996 272524
rect 380860 272484 380866 272496
rect 411990 272484 411996 272496
rect 412048 272484 412054 272536
rect 413830 272484 413836 272536
rect 413888 272524 413894 272536
rect 460658 272524 460664 272536
rect 413888 272496 460664 272524
rect 413888 272484 413894 272496
rect 460658 272484 460664 272496
rect 460716 272484 460722 272536
rect 461946 272484 461952 272536
rect 462004 272524 462010 272536
rect 529290 272524 529296 272536
rect 462004 272496 529296 272524
rect 462004 272484 462010 272496
rect 529290 272484 529296 272496
rect 529348 272484 529354 272536
rect 529474 272484 529480 272536
rect 529532 272524 529538 272536
rect 624694 272524 624700 272536
rect 529532 272496 624700 272524
rect 529532 272484 529538 272496
rect 624694 272484 624700 272496
rect 624752 272484 624758 272536
rect 127342 272348 127348 272400
rect 127400 272388 127406 272400
rect 179874 272388 179880 272400
rect 127400 272360 179880 272388
rect 127400 272348 127406 272360
rect 179874 272348 179880 272360
rect 179932 272348 179938 272400
rect 258534 272348 258540 272400
rect 258592 272388 258598 272400
rect 269758 272388 269764 272400
rect 258592 272360 269764 272388
rect 258592 272348 258598 272360
rect 269758 272348 269764 272360
rect 269816 272348 269822 272400
rect 429838 272348 429844 272400
rect 429896 272388 429902 272400
rect 447686 272388 447692 272400
rect 429896 272360 447692 272388
rect 429896 272348 429902 272360
rect 447686 272348 447692 272360
rect 447744 272348 447750 272400
rect 471606 272348 471612 272400
rect 471664 272388 471670 272400
rect 543458 272388 543464 272400
rect 471664 272360 543464 272388
rect 471664 272348 471670 272360
rect 543458 272348 543464 272360
rect 543516 272348 543522 272400
rect 116670 272212 116676 272264
rect 116728 272252 116734 272264
rect 166074 272252 166080 272264
rect 116728 272224 166080 272252
rect 116728 272212 116734 272224
rect 166074 272212 166080 272224
rect 166132 272212 166138 272264
rect 166258 272212 166264 272264
rect 166316 272252 166322 272264
rect 192018 272252 192024 272264
rect 166316 272224 192024 272252
rect 166316 272212 166322 272224
rect 192018 272212 192024 272224
rect 192076 272212 192082 272264
rect 467742 272212 467748 272264
rect 467800 272252 467806 272264
rect 536374 272252 536380 272264
rect 467800 272224 536380 272252
rect 467800 272212 467806 272224
rect 536374 272212 536380 272224
rect 536432 272212 536438 272264
rect 541618 272212 541624 272264
rect 541676 272252 541682 272264
rect 603718 272252 603724 272264
rect 541676 272224 603724 272252
rect 541676 272212 541682 272224
rect 603718 272212 603724 272224
rect 603776 272212 603782 272264
rect 152182 272076 152188 272128
rect 152240 272116 152246 272128
rect 189810 272116 189816 272128
rect 152240 272088 189816 272116
rect 152240 272076 152246 272088
rect 189810 272076 189816 272088
rect 189868 272076 189874 272128
rect 447778 272076 447784 272128
rect 447836 272116 447842 272128
rect 506842 272116 506848 272128
rect 447836 272088 506848 272116
rect 447836 272076 447842 272088
rect 506842 272076 506848 272088
rect 506900 272076 506906 272128
rect 507302 272076 507308 272128
rect 507360 272116 507366 272128
rect 565906 272116 565912 272128
rect 507360 272088 565912 272116
rect 507360 272076 507366 272088
rect 565906 272076 565912 272088
rect 565964 272076 565970 272128
rect 516042 271940 516048 271992
rect 516100 271980 516106 271992
rect 516686 271980 516692 271992
rect 516100 271952 516692 271980
rect 516100 271940 516106 271952
rect 516686 271940 516692 271952
rect 516744 271940 516750 271992
rect 517330 271940 517336 271992
rect 517388 271980 517394 271992
rect 525794 271980 525800 271992
rect 517388 271952 525800 271980
rect 517388 271940 517394 271952
rect 525794 271940 525800 271952
rect 525852 271940 525858 271992
rect 121362 271804 121368 271856
rect 121420 271844 121426 271856
rect 176746 271844 176752 271856
rect 121420 271816 176752 271844
rect 121420 271804 121426 271816
rect 176746 271804 176752 271816
rect 176804 271804 176810 271856
rect 187878 271804 187884 271856
rect 187936 271844 187942 271856
rect 196434 271844 196440 271856
rect 187936 271816 196440 271844
rect 187936 271804 187942 271816
rect 196434 271804 196440 271816
rect 196492 271804 196498 271856
rect 283190 271804 283196 271856
rect 283248 271844 283254 271856
rect 285122 271844 285128 271856
rect 283248 271816 285128 271844
rect 283248 271804 283254 271816
rect 285122 271804 285128 271816
rect 285180 271804 285186 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 395062 271844 395068 271856
rect 375340 271816 395068 271844
rect 375340 271804 375346 271816
rect 395062 271804 395068 271816
rect 395120 271804 395126 271856
rect 433150 271804 433156 271856
rect 433208 271844 433214 271856
rect 486694 271844 486700 271856
rect 433208 271816 486700 271844
rect 433208 271804 433214 271816
rect 486694 271804 486700 271816
rect 486752 271804 486758 271856
rect 496538 271804 496544 271856
rect 496596 271844 496602 271856
rect 578878 271844 578884 271856
rect 496596 271816 578884 271844
rect 496596 271804 496602 271816
rect 578878 271804 578884 271816
rect 578936 271804 578942 271856
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 104894 271668 104900 271720
rect 104952 271708 104958 271720
rect 163314 271708 163320 271720
rect 104952 271680 163320 271708
rect 104952 271668 104958 271680
rect 163314 271668 163320 271680
rect 163372 271668 163378 271720
rect 164142 271668 164148 271720
rect 164200 271708 164206 271720
rect 194778 271708 194784 271720
rect 164200 271680 194784 271708
rect 164200 271668 164206 271680
rect 194778 271668 194784 271680
rect 194836 271668 194842 271720
rect 197078 271668 197084 271720
rect 197136 271708 197142 271720
rect 224218 271708 224224 271720
rect 197136 271680 224224 271708
rect 197136 271668 197142 271680
rect 224218 271668 224224 271680
rect 224276 271668 224282 271720
rect 224586 271668 224592 271720
rect 224644 271708 224650 271720
rect 247770 271708 247776 271720
rect 224644 271680 247776 271708
rect 224644 271668 224650 271680
rect 247770 271668 247776 271680
rect 247828 271668 247834 271720
rect 363598 271668 363604 271720
rect 363656 271708 363662 271720
rect 374362 271708 374368 271720
rect 363656 271680 374368 271708
rect 363656 271668 363662 271680
rect 374362 271668 374368 271680
rect 374420 271668 374426 271720
rect 384758 271668 384764 271720
rect 384816 271708 384822 271720
rect 415302 271708 415308 271720
rect 384816 271680 415308 271708
rect 384816 271668 384822 271680
rect 415302 271668 415308 271680
rect 415360 271668 415366 271720
rect 437198 271668 437204 271720
rect 437256 271708 437262 271720
rect 493778 271708 493784 271720
rect 437256 271680 493784 271708
rect 437256 271668 437262 271680
rect 493778 271668 493784 271680
rect 493836 271668 493842 271720
rect 499482 271668 499488 271720
rect 499540 271708 499546 271720
rect 582466 271708 582472 271720
rect 499540 271680 582472 271708
rect 499540 271668 499546 271680
rect 582466 271668 582472 271680
rect 582524 271668 582530 271720
rect 105998 271532 106004 271584
rect 106056 271572 106062 271584
rect 164786 271572 164792 271584
rect 106056 271544 164792 271572
rect 106056 271532 106062 271544
rect 164786 271532 164792 271544
rect 164844 271532 164850 271584
rect 178126 271532 178132 271584
rect 178184 271572 178190 271584
rect 184198 271572 184204 271584
rect 178184 271544 184204 271572
rect 178184 271532 178190 271544
rect 184198 271532 184204 271544
rect 184256 271532 184262 271584
rect 184474 271532 184480 271584
rect 184532 271572 184538 271584
rect 215938 271572 215944 271584
rect 184532 271544 215944 271572
rect 184532 271532 184538 271544
rect 215938 271532 215944 271544
rect 215996 271532 216002 271584
rect 216306 271532 216312 271584
rect 216364 271572 216370 271584
rect 242066 271572 242072 271584
rect 216364 271544 242072 271572
rect 216364 271532 216370 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 340598 271532 340604 271584
rect 340656 271572 340662 271584
rect 355134 271572 355140 271584
rect 340656 271544 355140 271572
rect 340656 271532 340662 271544
rect 355134 271532 355140 271544
rect 355192 271532 355198 271584
rect 355318 271532 355324 271584
rect 355376 271572 355382 271584
rect 368474 271572 368480 271584
rect 355376 271544 368480 271572
rect 355376 271532 355382 271544
rect 368474 271532 368480 271544
rect 368532 271532 368538 271584
rect 369486 271532 369492 271584
rect 369544 271572 369550 271584
rect 377398 271572 377404 271584
rect 369544 271544 377404 271572
rect 369544 271532 369550 271544
rect 377398 271532 377404 271544
rect 377456 271532 377462 271584
rect 379330 271532 379336 271584
rect 379388 271572 379394 271584
rect 393866 271572 393872 271584
rect 379388 271544 393872 271572
rect 379388 271532 379394 271544
rect 393866 271532 393872 271544
rect 393924 271532 393930 271584
rect 395522 271532 395528 271584
rect 395580 271572 395586 271584
rect 427630 271572 427636 271584
rect 395580 271544 427636 271572
rect 395580 271532 395586 271544
rect 427630 271532 427636 271544
rect 427688 271532 427694 271584
rect 434438 271532 434444 271584
rect 434496 271572 434502 271584
rect 490282 271572 490288 271584
rect 434496 271544 490288 271572
rect 434496 271532 434502 271544
rect 490282 271532 490288 271544
rect 490340 271532 490346 271584
rect 494698 271532 494704 271584
rect 494756 271572 494762 271584
rect 500494 271572 500500 271584
rect 494756 271544 500500 271572
rect 494756 271532 494762 271544
rect 500494 271532 500500 271544
rect 500552 271532 500558 271584
rect 501966 271532 501972 271584
rect 502024 271572 502030 271584
rect 585594 271572 585600 271584
rect 502024 271544 585600 271572
rect 502024 271532 502030 271544
rect 585594 271532 585600 271544
rect 585652 271532 585658 271584
rect 585778 271532 585784 271584
rect 585836 271572 585842 271584
rect 608502 271572 608508 271584
rect 585836 271544 608508 271572
rect 585836 271532 585842 271544
rect 608502 271532 608508 271544
rect 608560 271532 608566 271584
rect 89530 271396 89536 271448
rect 89588 271436 89594 271448
rect 152366 271436 152372 271448
rect 89588 271408 152372 271436
rect 89588 271396 89594 271408
rect 152366 271396 152372 271408
rect 152424 271396 152430 271448
rect 162762 271396 162768 271448
rect 162820 271436 162826 271448
rect 204714 271436 204720 271448
rect 162820 271408 204720 271436
rect 162820 271396 162826 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 205358 271396 205364 271448
rect 205416 271436 205422 271448
rect 234982 271436 234988 271448
rect 205416 271408 234988 271436
rect 205416 271396 205422 271408
rect 234982 271396 234988 271408
rect 235040 271396 235046 271448
rect 248414 271396 248420 271448
rect 248472 271436 248478 271448
rect 264330 271436 264336 271448
rect 248472 271408 264336 271436
rect 248472 271396 248478 271408
rect 264330 271396 264336 271408
rect 264388 271396 264394 271448
rect 348878 271396 348884 271448
rect 348936 271436 348942 271448
rect 362954 271436 362960 271448
rect 348936 271408 362960 271436
rect 348936 271396 348942 271408
rect 362954 271396 362960 271408
rect 363012 271396 363018 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 379146 271436 379152 271448
rect 366416 271408 379152 271436
rect 366416 271396 366422 271408
rect 379146 271396 379152 271408
rect 379204 271396 379210 271448
rect 383378 271396 383384 271448
rect 383436 271436 383442 271448
rect 416958 271436 416964 271448
rect 383436 271408 416964 271436
rect 383436 271396 383442 271408
rect 416958 271396 416964 271408
rect 417016 271396 417022 271448
rect 418982 271396 418988 271448
rect 419040 271436 419046 271448
rect 429654 271436 429660 271448
rect 419040 271408 429660 271436
rect 419040 271396 419046 271408
rect 429654 271396 429660 271408
rect 429712 271396 429718 271448
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 497366 271436 497372 271448
rect 440016 271408 497372 271436
rect 440016 271396 440022 271408
rect 497366 271396 497372 271408
rect 497424 271396 497430 271448
rect 504910 271396 504916 271448
rect 504968 271436 504974 271448
rect 589550 271436 589556 271448
rect 504968 271408 589556 271436
rect 504968 271396 504974 271408
rect 589550 271396 589556 271408
rect 589608 271396 589614 271448
rect 592678 271396 592684 271448
rect 592736 271436 592742 271448
rect 622670 271436 622676 271448
rect 592736 271408 622676 271436
rect 592736 271396 592742 271408
rect 622670 271396 622676 271408
rect 622728 271396 622734 271448
rect 68186 271260 68192 271312
rect 68244 271300 68250 271312
rect 138474 271300 138480 271312
rect 68244 271272 138480 271300
rect 68244 271260 68250 271272
rect 138474 271260 138480 271272
rect 138532 271260 138538 271312
rect 139118 271260 139124 271312
rect 139176 271300 139182 271312
rect 141602 271300 141608 271312
rect 139176 271272 141608 271300
rect 139176 271260 139182 271272
rect 141602 271260 141608 271272
rect 141660 271260 141666 271312
rect 141786 271260 141792 271312
rect 141844 271300 141850 271312
rect 189626 271300 189632 271312
rect 141844 271272 189632 271300
rect 141844 271260 141850 271272
rect 189626 271260 189632 271272
rect 189684 271260 189690 271312
rect 195698 271260 195704 271312
rect 195756 271300 195762 271312
rect 227898 271300 227904 271312
rect 195756 271272 227904 271300
rect 195756 271260 195762 271272
rect 227898 271260 227904 271272
rect 227956 271260 227962 271312
rect 237282 271260 237288 271312
rect 237340 271300 237346 271312
rect 256970 271300 256976 271312
rect 237340 271272 256976 271300
rect 237340 271260 237346 271272
rect 256970 271260 256976 271272
rect 257028 271260 257034 271312
rect 260190 271260 260196 271312
rect 260248 271300 260254 271312
rect 270954 271300 270960 271312
rect 260248 271272 270960 271300
rect 260248 271260 260254 271272
rect 270954 271260 270960 271272
rect 271012 271260 271018 271312
rect 271506 271260 271512 271312
rect 271564 271300 271570 271312
rect 280890 271300 280896 271312
rect 271564 271272 280896 271300
rect 271564 271260 271570 271272
rect 280890 271260 280896 271272
rect 280948 271260 280954 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 325510 271260 325516 271312
rect 325568 271300 325574 271312
rect 334158 271300 334164 271312
rect 325568 271272 334164 271300
rect 325568 271260 325574 271272
rect 334158 271260 334164 271272
rect 334216 271260 334222 271312
rect 334618 271260 334624 271312
rect 334676 271300 334682 271312
rect 341334 271300 341340 271312
rect 334676 271272 341340 271300
rect 334676 271260 334682 271272
rect 341334 271260 341340 271272
rect 341392 271260 341398 271312
rect 354582 271260 354588 271312
rect 354640 271300 354646 271312
rect 369854 271300 369860 271312
rect 354640 271272 369860 271300
rect 354640 271260 354646 271272
rect 369854 271260 369860 271272
rect 369912 271260 369918 271312
rect 372522 271260 372528 271312
rect 372580 271300 372586 271312
rect 382458 271300 382464 271312
rect 372580 271272 382464 271300
rect 372580 271260 372586 271272
rect 382458 271260 382464 271272
rect 382516 271260 382522 271312
rect 387518 271260 387524 271312
rect 387576 271300 387582 271312
rect 421374 271300 421380 271312
rect 387576 271272 421380 271300
rect 387576 271260 387582 271272
rect 421374 271260 421380 271272
rect 421432 271260 421438 271312
rect 421558 271260 421564 271312
rect 421616 271300 421622 271312
rect 437014 271300 437020 271312
rect 421616 271272 437020 271300
rect 421616 271260 421622 271272
rect 437014 271260 437020 271272
rect 437072 271260 437078 271312
rect 445662 271260 445668 271312
rect 445720 271300 445726 271312
rect 455782 271300 455788 271312
rect 445720 271272 455788 271300
rect 445720 271260 445726 271272
rect 455782 271260 455788 271272
rect 455840 271260 455846 271312
rect 465718 271300 465724 271312
rect 456168 271272 465724 271300
rect 456168 271232 456196 271272
rect 465718 271260 465724 271272
rect 465776 271260 465782 271312
rect 465902 271260 465908 271312
rect 465960 271300 465966 271312
rect 507946 271300 507952 271312
rect 465960 271272 507952 271300
rect 465960 271260 465966 271272
rect 507946 271260 507952 271272
rect 508004 271260 508010 271312
rect 509142 271260 509148 271312
rect 509200 271300 509206 271312
rect 596634 271300 596640 271312
rect 509200 271272 596640 271300
rect 509200 271260 509206 271272
rect 596634 271260 596640 271272
rect 596692 271260 596698 271312
rect 596818 271260 596824 271312
rect 596876 271300 596882 271312
rect 629754 271300 629760 271312
rect 596876 271272 629760 271300
rect 596876 271260 596882 271272
rect 629754 271260 629760 271272
rect 629812 271260 629818 271312
rect 455984 271204 456196 271232
rect 72970 271124 72976 271176
rect 73028 271164 73034 271176
rect 142338 271164 142344 271176
rect 73028 271136 142344 271164
rect 73028 271124 73034 271136
rect 142338 271124 142344 271136
rect 142396 271124 142402 271176
rect 143258 271124 143264 271176
rect 143316 271164 143322 271176
rect 144362 271164 144368 271176
rect 143316 271136 144368 271164
rect 143316 271124 143322 271136
rect 144362 271124 144368 271136
rect 144420 271124 144426 271176
rect 154298 271124 154304 271176
rect 154356 271164 154362 271176
rect 197906 271164 197912 271176
rect 154356 271136 197912 271164
rect 154356 271124 154362 271136
rect 197906 271124 197912 271136
rect 197964 271124 197970 271176
rect 198274 271124 198280 271176
rect 198332 271164 198338 271176
rect 229554 271164 229560 271176
rect 198332 271136 229560 271164
rect 198332 271124 198338 271136
rect 229554 271124 229560 271136
rect 229612 271124 229618 271176
rect 231394 271124 231400 271176
rect 231452 271164 231458 271176
rect 252738 271164 252744 271176
rect 231452 271136 252744 271164
rect 231452 271124 231458 271136
rect 252738 271124 252744 271136
rect 252796 271124 252802 271176
rect 253566 271124 253572 271176
rect 253624 271164 253630 271176
rect 265250 271164 265256 271176
rect 253624 271136 265256 271164
rect 253624 271124 253630 271136
rect 265250 271124 265256 271136
rect 265308 271124 265314 271176
rect 269482 271124 269488 271176
rect 269540 271164 269546 271176
rect 279234 271164 279240 271176
rect 269540 271136 279240 271164
rect 269540 271124 269546 271136
rect 279234 271124 279240 271136
rect 279292 271124 279298 271176
rect 285766 271124 285772 271176
rect 285824 271164 285830 271176
rect 291194 271164 291200 271176
rect 285824 271136 291200 271164
rect 285824 271124 285830 271136
rect 291194 271124 291200 271136
rect 291252 271124 291258 271176
rect 328086 271124 328092 271176
rect 328144 271164 328150 271176
rect 337746 271164 337752 271176
rect 328144 271136 337752 271164
rect 328144 271124 328150 271136
rect 337746 271124 337752 271136
rect 337804 271124 337810 271176
rect 339310 271124 339316 271176
rect 339368 271164 339374 271176
rect 354306 271164 354312 271176
rect 339368 271136 354312 271164
rect 339368 271124 339374 271136
rect 354306 271124 354312 271136
rect 354364 271124 354370 271176
rect 362678 271124 362684 271176
rect 362736 271164 362742 271176
rect 387150 271164 387156 271176
rect 362736 271136 387156 271164
rect 362736 271124 362742 271136
rect 387150 271124 387156 271136
rect 387208 271124 387214 271176
rect 391750 271124 391756 271176
rect 391808 271164 391814 271176
rect 403618 271164 403624 271176
rect 391808 271136 403624 271164
rect 391808 271124 391814 271136
rect 403618 271124 403624 271136
rect 403676 271124 403682 271176
rect 404170 271124 404176 271176
rect 404228 271164 404234 271176
rect 445294 271164 445300 271176
rect 404228 271136 445300 271164
rect 404228 271124 404234 271136
rect 445294 271124 445300 271136
rect 445352 271124 445358 271176
rect 449802 271124 449808 271176
rect 449860 271164 449866 271176
rect 455984 271164 456012 271204
rect 449860 271136 456012 271164
rect 449860 271124 449866 271136
rect 456334 271124 456340 271176
rect 456392 271164 456398 271176
rect 504174 271164 504180 271176
rect 456392 271136 504180 271164
rect 456392 271124 456398 271136
rect 504174 271124 504180 271136
rect 504232 271124 504238 271176
rect 511534 271164 511540 271176
rect 504376 271136 511540 271164
rect 83550 270988 83556 271040
rect 83608 271028 83614 271040
rect 123478 271028 123484 271040
rect 83608 271000 123484 271028
rect 83608 270988 83614 271000
rect 123478 270988 123484 271000
rect 123536 270988 123542 271040
rect 123754 270988 123760 271040
rect 123812 271028 123818 271040
rect 177482 271028 177488 271040
rect 123812 271000 177488 271028
rect 123812 270988 123818 271000
rect 177482 270988 177488 271000
rect 177540 270988 177546 271040
rect 418062 270988 418068 271040
rect 418120 271028 418126 271040
rect 463786 271028 463792 271040
rect 418120 271000 463792 271028
rect 418120 270988 418126 271000
rect 463786 270988 463792 271000
rect 463844 270988 463850 271040
rect 465718 270988 465724 271040
rect 465776 271028 465782 271040
rect 504376 271028 504404 271136
rect 511534 271124 511540 271136
rect 511592 271124 511598 271176
rect 511902 271124 511908 271176
rect 511960 271164 511966 271176
rect 600222 271164 600228 271176
rect 511960 271136 600228 271164
rect 511960 271124 511966 271136
rect 600222 271124 600228 271136
rect 600280 271124 600286 271176
rect 623038 271124 623044 271176
rect 623096 271164 623102 271176
rect 643922 271164 643928 271176
rect 623096 271136 643928 271164
rect 623096 271124 623102 271136
rect 643922 271124 643928 271136
rect 643980 271124 643986 271176
rect 465776 271000 504404 271028
rect 465776 270988 465782 271000
rect 504542 270988 504548 271040
rect 504600 271028 504606 271040
rect 575382 271028 575388 271040
rect 504600 271000 575388 271028
rect 504600 270988 504606 271000
rect 575382 270988 575388 271000
rect 575440 270988 575446 271040
rect 576118 270988 576124 271040
rect 576176 271028 576182 271040
rect 594334 271028 594340 271040
rect 576176 271000 594340 271028
rect 576176 270988 576182 271000
rect 594334 270988 594340 271000
rect 594392 270988 594398 271040
rect 134426 270852 134432 270904
rect 134484 270892 134490 270904
rect 184934 270892 184940 270904
rect 134484 270864 184940 270892
rect 134484 270852 134490 270864
rect 184934 270852 184940 270864
rect 184992 270852 184998 270904
rect 404998 270852 405004 270904
rect 405056 270892 405062 270904
rect 434714 270892 434720 270904
rect 405056 270864 434720 270892
rect 405056 270852 405062 270864
rect 434714 270852 434720 270864
rect 434772 270852 434778 270904
rect 456058 270852 456064 270904
rect 456116 270892 456122 270904
rect 465902 270892 465908 270904
rect 456116 270864 465908 270892
rect 456116 270852 456122 270864
rect 465902 270852 465908 270864
rect 465960 270852 465966 270904
rect 492030 270852 492036 270904
rect 492088 270892 492094 270904
rect 571794 270892 571800 270904
rect 492088 270864 571800 270892
rect 492088 270852 492094 270864
rect 571794 270852 571800 270864
rect 571852 270852 571858 270904
rect 113174 270716 113180 270768
rect 113232 270756 113238 270768
rect 154022 270756 154028 270768
rect 113232 270728 154028 270756
rect 113232 270716 113238 270728
rect 154022 270716 154028 270728
rect 154080 270716 154086 270768
rect 175826 270716 175832 270768
rect 175884 270756 175890 270768
rect 206278 270756 206284 270768
rect 175884 270728 206284 270756
rect 175884 270716 175890 270728
rect 206278 270716 206284 270728
rect 206336 270716 206342 270768
rect 425698 270716 425704 270768
rect 425756 270756 425762 270768
rect 448882 270756 448888 270768
rect 425756 270728 448888 270756
rect 425756 270716 425762 270728
rect 448882 270716 448888 270728
rect 448940 270716 448946 270768
rect 463786 270716 463792 270768
rect 463844 270756 463850 270768
rect 466638 270756 466644 270768
rect 463844 270728 466644 270756
rect 463844 270716 463850 270728
rect 466638 270716 466644 270728
rect 466696 270716 466702 270768
rect 467098 270716 467104 270768
rect 467156 270756 467162 270768
rect 525334 270756 525340 270768
rect 467156 270728 525340 270756
rect 467156 270716 467162 270728
rect 525334 270716 525340 270728
rect 525392 270716 525398 270768
rect 526438 270716 526444 270768
rect 526496 270756 526502 270768
rect 576578 270756 576584 270768
rect 526496 270728 576584 270756
rect 526496 270716 526502 270728
rect 576578 270716 576584 270728
rect 576636 270716 576642 270768
rect 414474 270580 414480 270632
rect 414532 270620 414538 270632
rect 437934 270620 437940 270632
rect 414532 270592 437940 270620
rect 414532 270580 414538 270592
rect 437934 270580 437940 270592
rect 437992 270580 437998 270632
rect 445018 270580 445024 270632
rect 445076 270620 445082 270632
rect 494698 270620 494704 270632
rect 445076 270592 494704 270620
rect 445076 270580 445082 270592
rect 494698 270580 494704 270592
rect 494756 270580 494762 270632
rect 495342 270580 495348 270632
rect 495400 270620 495406 270632
rect 504542 270620 504548 270632
rect 495400 270592 504548 270620
rect 495400 270580 495406 270592
rect 504542 270580 504548 270592
rect 504600 270580 504606 270632
rect 100662 270444 100668 270496
rect 100720 270484 100726 270496
rect 119798 270484 119804 270496
rect 100720 270456 119804 270484
rect 100720 270444 100726 270456
rect 119798 270444 119804 270456
rect 119856 270444 119862 270496
rect 122742 270444 122748 270496
rect 122800 270484 122806 270496
rect 176194 270484 176200 270496
rect 122800 270456 176200 270484
rect 122800 270444 122806 270456
rect 176194 270444 176200 270456
rect 176252 270444 176258 270496
rect 176930 270444 176936 270496
rect 176988 270484 176994 270496
rect 214742 270484 214748 270496
rect 176988 270456 214748 270484
rect 176988 270444 176994 270456
rect 214742 270444 214748 270456
rect 214800 270444 214806 270496
rect 230382 270444 230388 270496
rect 230440 270484 230446 270496
rect 252094 270484 252100 270496
rect 230440 270456 252100 270484
rect 230440 270444 230446 270456
rect 252094 270444 252100 270456
rect 252152 270444 252158 270496
rect 275094 270444 275100 270496
rect 275152 270484 275158 270496
rect 276014 270484 276020 270496
rect 275152 270456 276020 270484
rect 275152 270444 275158 270456
rect 276014 270444 276020 270456
rect 276072 270444 276078 270496
rect 281442 270444 281448 270496
rect 281500 270484 281506 270496
rect 285674 270484 285680 270496
rect 281500 270456 285680 270484
rect 281500 270444 281506 270456
rect 285674 270444 285680 270456
rect 285732 270444 285738 270496
rect 292850 270444 292856 270496
rect 292908 270484 292914 270496
rect 293954 270484 293960 270496
rect 292908 270456 293960 270484
rect 292908 270444 292914 270456
rect 293954 270444 293960 270456
rect 294012 270444 294018 270496
rect 297910 270444 297916 270496
rect 297968 270484 297974 270496
rect 299566 270484 299572 270496
rect 297968 270456 299572 270484
rect 297968 270444 297974 270456
rect 299566 270444 299572 270456
rect 299624 270444 299630 270496
rect 299934 270444 299940 270496
rect 299992 270484 299998 270496
rect 300854 270484 300860 270496
rect 299992 270456 300860 270484
rect 299992 270444 299998 270456
rect 300854 270444 300860 270456
rect 300912 270444 300918 270496
rect 327074 270444 327080 270496
rect 327132 270484 327138 270496
rect 328454 270484 328460 270496
rect 327132 270456 328460 270484
rect 327132 270444 327138 270456
rect 328454 270444 328460 270456
rect 328512 270444 328518 270496
rect 360194 270484 360200 270496
rect 354646 270456 360200 270484
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132586 270348 132592 270360
rect 78916 270320 132592 270348
rect 78916 270308 78922 270320
rect 132586 270308 132592 270320
rect 132644 270308 132650 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 183646 270348 183652 270360
rect 133840 270320 183652 270348
rect 133840 270308 133846 270320
rect 183646 270308 183652 270320
rect 183704 270308 183710 270360
rect 185210 270308 185216 270360
rect 185268 270348 185274 270360
rect 186314 270348 186320 270360
rect 185268 270320 186320 270348
rect 185268 270308 185274 270320
rect 186314 270308 186320 270320
rect 186372 270308 186378 270360
rect 186498 270308 186504 270360
rect 186556 270348 186562 270360
rect 202322 270348 202328 270360
rect 186556 270320 202328 270348
rect 186556 270308 186562 270320
rect 202322 270308 202328 270320
rect 202380 270308 202386 270360
rect 202782 270308 202788 270360
rect 202840 270348 202846 270360
rect 205910 270348 205916 270360
rect 202840 270320 205916 270348
rect 202840 270308 202846 270320
rect 205910 270308 205916 270320
rect 205968 270308 205974 270360
rect 219526 270308 219532 270360
rect 219584 270348 219590 270360
rect 244918 270348 244924 270360
rect 219584 270320 244924 270348
rect 219584 270308 219590 270320
rect 244918 270308 244924 270320
rect 244976 270308 244982 270360
rect 278590 270308 278596 270360
rect 278648 270348 278654 270360
rect 286318 270348 286324 270360
rect 278648 270320 286324 270348
rect 278648 270308 278654 270320
rect 286318 270308 286324 270320
rect 286376 270308 286382 270360
rect 291654 270308 291660 270360
rect 291712 270348 291718 270360
rect 295518 270348 295524 270360
rect 291712 270320 295524 270348
rect 291712 270308 291718 270320
rect 295518 270308 295524 270320
rect 295576 270308 295582 270360
rect 85482 270172 85488 270224
rect 85540 270212 85546 270224
rect 149422 270212 149428 270224
rect 85540 270184 149428 270212
rect 85540 270172 85546 270184
rect 149422 270172 149428 270184
rect 149480 270172 149486 270224
rect 153286 270172 153292 270224
rect 153344 270212 153350 270224
rect 169846 270212 169852 270224
rect 153344 270184 169852 270212
rect 153344 270172 153350 270184
rect 169846 270172 169852 270184
rect 169904 270172 169910 270224
rect 170030 270172 170036 270224
rect 170088 270212 170094 270224
rect 210142 270212 210148 270224
rect 170088 270184 210148 270212
rect 170088 270172 170094 270184
rect 210142 270172 210148 270184
rect 210200 270172 210206 270224
rect 210602 270172 210608 270224
rect 210660 270212 210666 270224
rect 237466 270212 237472 270224
rect 210660 270184 237472 270212
rect 210660 270172 210666 270184
rect 237466 270172 237472 270184
rect 237524 270172 237530 270224
rect 255222 270172 255228 270224
rect 255280 270212 255286 270224
rect 269390 270212 269396 270224
rect 255280 270184 269396 270212
rect 255280 270172 255286 270184
rect 269390 270172 269396 270184
rect 269448 270172 269454 270224
rect 288250 270172 288256 270224
rect 288308 270212 288314 270224
rect 292942 270212 292948 270224
rect 288308 270184 292948 270212
rect 288308 270172 288314 270184
rect 292942 270172 292948 270184
rect 293000 270172 293006 270224
rect 321094 270172 321100 270224
rect 321152 270212 321158 270224
rect 327442 270212 327448 270224
rect 321152 270184 327448 270212
rect 321152 270172 321158 270184
rect 327442 270172 327448 270184
rect 327500 270172 327506 270224
rect 329374 270172 329380 270224
rect 329432 270212 329438 270224
rect 339494 270212 339500 270224
rect 329432 270184 339500 270212
rect 329432 270172 329438 270184
rect 339494 270172 339500 270184
rect 339552 270172 339558 270224
rect 345934 270172 345940 270224
rect 345992 270212 345998 270224
rect 354646 270212 354674 270456
rect 360194 270444 360200 270456
rect 360252 270444 360258 270496
rect 382274 270484 382280 270496
rect 373966 270456 382280 270484
rect 359182 270308 359188 270360
rect 359240 270348 359246 270360
rect 373966 270348 373994 270456
rect 382274 270444 382280 270456
rect 382332 270444 382338 270496
rect 383838 270444 383844 270496
rect 383896 270484 383902 270496
rect 391934 270484 391940 270496
rect 383896 270456 391940 270484
rect 383896 270444 383902 270456
rect 391934 270444 391940 270456
rect 391992 270444 391998 270496
rect 400582 270444 400588 270496
rect 400640 270484 400646 270496
rect 441614 270484 441620 270496
rect 400640 270456 441620 270484
rect 400640 270444 400646 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 453574 270444 453580 270496
rect 453632 270484 453638 270496
rect 516502 270484 516508 270496
rect 453632 270456 516508 270484
rect 453632 270444 453638 270456
rect 516502 270444 516508 270456
rect 516560 270444 516566 270496
rect 517790 270444 517796 270496
rect 517848 270484 517854 270496
rect 597554 270484 597560 270496
rect 517848 270456 597560 270484
rect 517848 270444 517854 270456
rect 597554 270444 597560 270456
rect 597612 270444 597618 270496
rect 359240 270320 373994 270348
rect 359240 270308 359246 270320
rect 377950 270308 377956 270360
rect 378008 270348 378014 270360
rect 387794 270348 387800 270360
rect 378008 270320 387800 270348
rect 378008 270308 378014 270320
rect 387794 270308 387800 270320
rect 387852 270308 387858 270360
rect 407206 270308 407212 270360
rect 407264 270348 407270 270360
rect 451458 270348 451464 270360
rect 407264 270320 451464 270348
rect 407264 270308 407270 270320
rect 451458 270308 451464 270320
rect 451516 270308 451522 270360
rect 456426 270308 456432 270360
rect 456484 270348 456490 270360
rect 520274 270348 520280 270360
rect 456484 270320 520280 270348
rect 456484 270308 456490 270320
rect 520274 270308 520280 270320
rect 520332 270308 520338 270360
rect 523126 270308 523132 270360
rect 523184 270348 523190 270360
rect 605098 270348 605104 270360
rect 523184 270320 605104 270348
rect 523184 270308 523190 270320
rect 605098 270308 605104 270320
rect 605156 270308 605162 270360
rect 345992 270184 354674 270212
rect 345992 270172 345998 270184
rect 360194 270172 360200 270224
rect 360252 270212 360258 270224
rect 383654 270212 383660 270224
rect 360252 270184 383660 270212
rect 360252 270172 360258 270184
rect 383654 270172 383660 270184
rect 383712 270172 383718 270224
rect 387702 270172 387708 270224
rect 387760 270212 387766 270224
rect 401778 270212 401784 270224
rect 387760 270184 401784 270212
rect 387760 270172 387766 270184
rect 401778 270172 401784 270184
rect 401836 270172 401842 270224
rect 410518 270172 410524 270224
rect 410576 270212 410582 270224
rect 455414 270212 455420 270224
rect 410576 270184 455420 270212
rect 410576 270172 410582 270184
rect 455414 270172 455420 270184
rect 455472 270172 455478 270224
rect 461394 270172 461400 270224
rect 461452 270212 461458 270224
rect 527174 270212 527180 270224
rect 461452 270184 527180 270212
rect 461452 270172 461458 270184
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528094 270172 528100 270224
rect 528152 270212 528158 270224
rect 619174 270212 619180 270224
rect 528152 270184 619180 270212
rect 528152 270172 528158 270184
rect 619174 270172 619180 270184
rect 619232 270172 619238 270224
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 67542 270036 67548 270088
rect 67600 270076 67606 270088
rect 75914 270076 75920 270088
rect 67600 270048 75920 270076
rect 67600 270036 67606 270048
rect 75914 270036 75920 270048
rect 75972 270036 75978 270088
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 158622 270036 158628 270088
rect 158680 270076 158686 270088
rect 201034 270076 201040 270088
rect 158680 270048 201040 270076
rect 158680 270036 158686 270048
rect 201034 270036 201040 270048
rect 201092 270036 201098 270088
rect 201770 270036 201776 270088
rect 201828 270076 201834 270088
rect 201828 270048 205772 270076
rect 201828 270036 201834 270048
rect 77202 269900 77208 269952
rect 77260 269940 77266 269952
rect 143902 269940 143908 269952
rect 77260 269912 143908 269940
rect 77260 269900 77266 269912
rect 143902 269900 143908 269912
rect 143960 269900 143966 269952
rect 144086 269900 144092 269952
rect 144144 269940 144150 269952
rect 190822 269940 190828 269952
rect 144144 269912 190828 269940
rect 144144 269900 144150 269912
rect 190822 269900 190828 269912
rect 190880 269900 190886 269952
rect 204162 269900 204168 269952
rect 204220 269940 204226 269952
rect 205082 269940 205088 269952
rect 204220 269912 205088 269940
rect 204220 269900 204226 269912
rect 205082 269900 205088 269912
rect 205140 269900 205146 269952
rect 205744 269940 205772 270048
rect 205910 270036 205916 270088
rect 205968 270076 205974 270088
rect 230842 270076 230848 270088
rect 205968 270048 230848 270076
rect 205968 270036 205974 270048
rect 230842 270036 230848 270048
rect 230900 270036 230906 270088
rect 244090 270036 244096 270088
rect 244148 270076 244154 270088
rect 260650 270076 260656 270088
rect 244148 270048 260656 270076
rect 244148 270036 244154 270048
rect 260650 270036 260656 270048
rect 260708 270036 260714 270088
rect 262030 270036 262036 270088
rect 262088 270076 262094 270088
rect 274726 270076 274732 270088
rect 262088 270048 274732 270076
rect 262088 270036 262094 270048
rect 274726 270036 274732 270048
rect 274784 270036 274790 270088
rect 316954 270036 316960 270088
rect 317012 270076 317018 270088
rect 321554 270076 321560 270088
rect 317012 270048 321560 270076
rect 317012 270036 317018 270048
rect 321554 270036 321560 270048
rect 321612 270036 321618 270088
rect 332226 270036 332232 270088
rect 332284 270076 332290 270088
rect 336642 270076 336648 270088
rect 332284 270048 336648 270076
rect 332284 270036 332290 270048
rect 336642 270036 336648 270048
rect 336700 270036 336706 270088
rect 347406 270076 347412 270088
rect 344986 270048 347412 270076
rect 232498 269940 232504 269952
rect 205744 269912 232504 269940
rect 232498 269900 232504 269912
rect 232556 269900 232562 269952
rect 233694 269900 233700 269952
rect 233752 269940 233758 269952
rect 243906 269940 243912 269952
rect 233752 269912 243912 269940
rect 233752 269900 233758 269912
rect 243906 269900 243912 269912
rect 243964 269900 243970 269952
rect 245470 269900 245476 269952
rect 245528 269940 245534 269952
rect 263134 269940 263140 269952
rect 245528 269912 263140 269940
rect 245528 269900 245534 269912
rect 263134 269900 263140 269912
rect 263192 269900 263198 269952
rect 266262 269900 266268 269952
rect 266320 269940 266326 269952
rect 272886 269940 272892 269952
rect 266320 269912 272892 269940
rect 266320 269900 266326 269912
rect 272886 269900 272892 269912
rect 272944 269900 272950 269952
rect 286962 269900 286968 269952
rect 287020 269940 287026 269952
rect 292114 269940 292120 269952
rect 287020 269912 292120 269940
rect 287020 269900 287026 269912
rect 292114 269900 292120 269912
rect 292172 269900 292178 269952
rect 323578 269900 323584 269952
rect 323636 269940 323642 269952
rect 331214 269940 331220 269952
rect 323636 269912 331220 269940
rect 323636 269900 323642 269912
rect 331214 269900 331220 269912
rect 331272 269900 331278 269952
rect 335998 269900 336004 269952
rect 336056 269940 336062 269952
rect 344986 269940 345014 270048
rect 347406 270036 347412 270048
rect 347464 270036 347470 270088
rect 349706 270036 349712 270088
rect 349764 270076 349770 270088
rect 357434 270076 357440 270088
rect 349764 270048 357440 270076
rect 349764 270036 349770 270048
rect 357434 270036 357440 270048
rect 357492 270036 357498 270088
rect 364150 270036 364156 270088
rect 364208 270076 364214 270088
rect 389174 270076 389180 270088
rect 364208 270048 389180 270076
rect 364208 270036 364214 270048
rect 389174 270036 389180 270048
rect 389232 270036 389238 270088
rect 389634 270036 389640 270088
rect 389692 270076 389698 270088
rect 405734 270076 405740 270088
rect 389692 270048 405740 270076
rect 389692 270036 389698 270048
rect 405734 270036 405740 270048
rect 405792 270036 405798 270088
rect 409690 270036 409696 270088
rect 409748 270076 409754 270088
rect 454126 270076 454132 270088
rect 409748 270048 454132 270076
rect 409748 270036 409754 270048
rect 454126 270036 454132 270048
rect 454184 270036 454190 270088
rect 454494 270036 454500 270088
rect 454552 270076 454558 270088
rect 473354 270076 473360 270088
rect 454552 270048 473360 270076
rect 454552 270036 454558 270048
rect 473354 270036 473360 270048
rect 473412 270036 473418 270088
rect 525518 270036 525524 270088
rect 525576 270076 525582 270088
rect 619634 270076 619640 270088
rect 525576 270048 619640 270076
rect 525576 270036 525582 270048
rect 619634 270036 619640 270048
rect 619692 270036 619698 270088
rect 336056 269912 345014 269940
rect 336056 269900 336062 269912
rect 346762 269900 346768 269952
rect 346820 269940 346826 269952
rect 364334 269940 364340 269952
rect 346820 269912 364340 269940
rect 346820 269900 346826 269912
rect 364334 269900 364340 269912
rect 364392 269900 364398 269952
rect 364978 269900 364984 269952
rect 365036 269940 365042 269952
rect 390554 269940 390560 269952
rect 365036 269912 390560 269940
rect 365036 269900 365042 269912
rect 390554 269900 390560 269912
rect 390612 269900 390618 269952
rect 391934 269900 391940 269952
rect 391992 269940 391998 269952
rect 409874 269940 409880 269952
rect 391992 269912 409880 269940
rect 391992 269900 391998 269912
rect 409874 269900 409880 269912
rect 409932 269900 409938 269952
rect 412450 269900 412456 269952
rect 412508 269940 412514 269952
rect 458174 269940 458180 269952
rect 412508 269912 458180 269940
rect 412508 269900 412514 269912
rect 458174 269900 458180 269912
rect 458232 269900 458238 269952
rect 458542 269900 458548 269952
rect 458600 269940 458606 269952
rect 524414 269940 524420 269952
rect 458600 269912 524420 269940
rect 458600 269900 458606 269912
rect 524414 269900 524420 269912
rect 524472 269900 524478 269952
rect 531682 269900 531688 269952
rect 531740 269940 531746 269952
rect 627914 269940 627920 269952
rect 531740 269912 627920 269940
rect 531740 269900 531746 269912
rect 627914 269900 627920 269912
rect 627972 269900 627978 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 140682 269764 140688 269816
rect 140740 269804 140746 269816
rect 188614 269804 188620 269816
rect 140740 269776 188620 269804
rect 140740 269764 140746 269776
rect 188614 269764 188620 269776
rect 188672 269764 188678 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 119062 269628 119068 269680
rect 119120 269668 119126 269680
rect 173342 269668 173348 269680
rect 119120 269640 173348 269668
rect 119120 269628 119126 269640
rect 173342 269628 173348 269640
rect 173400 269628 173406 269680
rect 174906 269628 174912 269680
rect 174964 269668 174970 269680
rect 174964 269640 204944 269668
rect 174964 269628 174970 269640
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 204162 269532 204168 269544
rect 183520 269504 204168 269532
rect 183520 269492 183526 269504
rect 204162 269492 204168 269504
rect 204220 269492 204226 269544
rect 136082 269356 136088 269408
rect 136140 269396 136146 269408
rect 180886 269396 180892 269408
rect 136140 269368 180892 269396
rect 136140 269356 136146 269368
rect 180886 269356 180892 269368
rect 180944 269356 180950 269408
rect 204916 269396 204944 269640
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 250254 269764 250260 269816
rect 250312 269804 250318 269816
rect 266630 269804 266636 269816
rect 250312 269776 266636 269804
rect 250312 269764 250318 269776
rect 266630 269764 266636 269776
rect 266688 269764 266694 269816
rect 266814 269764 266820 269816
rect 266872 269804 266878 269816
rect 278038 269804 278044 269816
rect 266872 269776 278044 269804
rect 266872 269764 266878 269776
rect 278038 269764 278044 269776
rect 278096 269764 278102 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318978 269804 318984 269816
rect 314528 269776 318984 269804
rect 314528 269764 314534 269776
rect 318978 269764 318984 269776
rect 319036 269764 319042 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 336826 269764 336832 269816
rect 336884 269804 336890 269816
rect 350534 269804 350540 269816
rect 336884 269776 350540 269804
rect 336884 269764 336890 269776
rect 350534 269764 350540 269776
rect 350592 269764 350598 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 374914 269764 374920 269816
rect 374972 269804 374978 269816
rect 404354 269804 404360 269816
rect 374972 269776 404360 269804
rect 374972 269764 374978 269776
rect 404354 269764 404360 269776
rect 404412 269764 404418 269816
rect 417142 269764 417148 269816
rect 417200 269804 417206 269816
rect 465074 269804 465080 269816
rect 417200 269776 465080 269804
rect 417200 269764 417206 269776
rect 465074 269764 465080 269776
rect 465132 269764 465138 269816
rect 465994 269764 466000 269816
rect 466052 269804 466058 269816
rect 534350 269804 534356 269816
rect 466052 269776 534356 269804
rect 466052 269764 466058 269776
rect 534350 269764 534356 269776
rect 534408 269764 534414 269816
rect 535546 269764 535552 269816
rect 535604 269804 535610 269816
rect 633526 269804 633532 269816
rect 535604 269776 633532 269804
rect 535604 269764 535610 269776
rect 633526 269764 633532 269776
rect 633584 269764 633590 269816
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 236086 269628 236092 269680
rect 236144 269668 236150 269680
rect 253750 269668 253756 269680
rect 236144 269640 253756 269668
rect 236144 269628 236150 269640
rect 253750 269628 253756 269640
rect 253808 269628 253814 269680
rect 341794 269628 341800 269680
rect 341852 269668 341858 269680
rect 349706 269668 349712 269680
rect 341852 269640 349712 269668
rect 341852 269628 341858 269640
rect 349706 269628 349712 269640
rect 349764 269628 349770 269680
rect 393314 269628 393320 269680
rect 393372 269668 393378 269680
rect 412634 269668 412640 269680
rect 393372 269640 412640 269668
rect 393372 269628 393378 269640
rect 412634 269628 412640 269640
rect 412692 269628 412698 269680
rect 422110 269628 422116 269680
rect 422168 269668 422174 269680
rect 472066 269668 472072 269680
rect 422168 269640 472072 269668
rect 422168 269628 422174 269640
rect 472066 269628 472072 269640
rect 472124 269628 472130 269680
rect 474642 269628 474648 269680
rect 474700 269668 474706 269680
rect 546494 269668 546500 269680
rect 474700 269640 546500 269668
rect 474700 269628 474706 269640
rect 546494 269628 546500 269640
rect 546552 269628 546558 269680
rect 205082 269492 205088 269544
rect 205140 269532 205146 269544
rect 223482 269532 223488 269544
rect 205140 269504 223488 269532
rect 205140 269492 205146 269504
rect 223482 269492 223488 269504
rect 223540 269492 223546 269544
rect 388162 269492 388168 269544
rect 388220 269532 388226 269544
rect 423030 269532 423036 269544
rect 388220 269504 423036 269532
rect 388220 269492 388226 269504
rect 423030 269492 423036 269504
rect 423088 269492 423094 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 476114 269532 476120 269544
rect 424652 269504 476120 269532
rect 424652 269492 424658 269504
rect 476114 269492 476120 269504
rect 476172 269492 476178 269544
rect 476758 269492 476764 269544
rect 476816 269532 476822 269544
rect 549898 269532 549904 269544
rect 476816 269504 549904 269532
rect 476816 269492 476822 269504
rect 549898 269492 549904 269504
rect 549956 269492 549962 269544
rect 210970 269396 210976 269408
rect 204916 269368 210976 269396
rect 210970 269356 210976 269368
rect 211028 269356 211034 269408
rect 273070 269356 273076 269408
rect 273128 269396 273134 269408
rect 277394 269396 277400 269408
rect 273128 269368 277400 269396
rect 273128 269356 273134 269368
rect 277394 269356 277400 269368
rect 277452 269356 277458 269408
rect 401686 269356 401692 269408
rect 401744 269396 401750 269408
rect 419534 269396 419540 269408
rect 401744 269368 419540 269396
rect 401744 269356 401750 269368
rect 419534 269356 419540 269368
rect 419592 269356 419598 269408
rect 419810 269356 419816 269408
rect 419868 269396 419874 269408
rect 462314 269396 462320 269408
rect 419868 269368 462320 269396
rect 419868 269356 419874 269368
rect 462314 269356 462320 269368
rect 462372 269356 462378 269408
rect 507946 269356 507952 269408
rect 508004 269396 508010 269408
rect 560294 269396 560300 269408
rect 508004 269368 560300 269396
rect 508004 269356 508010 269368
rect 560294 269356 560300 269368
rect 560352 269356 560358 269408
rect 251450 269220 251456 269272
rect 251508 269260 251514 269272
rect 258258 269260 258264 269272
rect 251508 269232 258264 269260
rect 251508 269220 251514 269232
rect 258258 269220 258264 269232
rect 258316 269220 258322 269272
rect 295334 269220 295340 269272
rect 295392 269260 295398 269272
rect 297910 269260 297916 269272
rect 295392 269232 297916 269260
rect 295392 269220 295398 269232
rect 297910 269220 297916 269232
rect 297968 269220 297974 269272
rect 441614 269220 441620 269272
rect 441672 269260 441678 269272
rect 460934 269260 460940 269272
rect 441672 269232 460940 269260
rect 441672 269220 441678 269232
rect 460934 269220 460940 269232
rect 460992 269220 460998 269272
rect 463510 269220 463516 269272
rect 463568 269260 463574 269272
rect 531314 269260 531320 269272
rect 463568 269232 531320 269260
rect 463568 269220 463574 269232
rect 531314 269220 531320 269232
rect 531372 269220 531378 269272
rect 146938 269152 146944 269204
rect 146996 269192 147002 269204
rect 153838 269192 153844 269204
rect 146996 269164 153844 269192
rect 146996 269152 147002 269164
rect 153838 269152 153844 269164
rect 153896 269152 153902 269204
rect 294138 269084 294144 269136
rect 294196 269124 294202 269136
rect 297082 269124 297088 269136
rect 294196 269096 297088 269124
rect 294196 269084 294202 269096
rect 297082 269084 297088 269096
rect 297140 269084 297146 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 342254 269084 342260 269136
rect 342312 269124 342318 269136
rect 345106 269124 345112 269136
rect 342312 269096 345112 269124
rect 342312 269084 342318 269096
rect 345106 269084 345112 269096
rect 345164 269084 345170 269136
rect 115842 269016 115848 269068
rect 115900 269056 115906 269068
rect 171226 269056 171232 269068
rect 115900 269028 171232 269056
rect 115900 269016 115906 269028
rect 171226 269016 171232 269028
rect 171284 269016 171290 269068
rect 428734 269016 428740 269068
rect 428792 269056 428798 269068
rect 475194 269056 475200 269068
rect 428792 269028 475200 269056
rect 428792 269016 428798 269028
rect 475194 269016 475200 269028
rect 475252 269016 475258 269068
rect 475378 269016 475384 269068
rect 475436 269056 475442 269068
rect 494238 269056 494244 269068
rect 475436 269028 494244 269056
rect 475436 269016 475442 269028
rect 494238 269016 494244 269028
rect 494296 269016 494302 269068
rect 495802 269016 495808 269068
rect 495860 269056 495866 269068
rect 576854 269056 576860 269068
rect 495860 269028 576860 269056
rect 495860 269016 495866 269028
rect 576854 269016 576860 269028
rect 576912 269016 576918 269068
rect 108942 268880 108948 268932
rect 109000 268920 109006 268932
rect 166258 268920 166264 268932
rect 109000 268892 166264 268920
rect 109000 268880 109006 268892
rect 166258 268880 166264 268892
rect 166316 268880 166322 268932
rect 172422 268880 172428 268932
rect 172480 268920 172486 268932
rect 204346 268920 204352 268932
rect 172480 268892 204352 268920
rect 172480 268880 172486 268892
rect 204346 268880 204352 268892
rect 204404 268880 204410 268932
rect 208210 268880 208216 268932
rect 208268 268920 208274 268932
rect 227714 268920 227720 268932
rect 208268 268892 227720 268920
rect 208268 268880 208274 268892
rect 227714 268880 227720 268892
rect 227772 268880 227778 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 411254 268920 411260 268932
rect 382424 268892 411260 268920
rect 382424 268880 382430 268892
rect 411254 268880 411260 268892
rect 411312 268880 411318 268932
rect 429562 268880 429568 268932
rect 429620 268920 429626 268932
rect 483106 268920 483112 268932
rect 429620 268892 483112 268920
rect 429620 268880 429626 268892
rect 483106 268880 483112 268892
rect 483164 268880 483170 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 582282 268880 582288 268932
rect 582340 268920 582346 268932
rect 600590 268920 600596 268932
rect 582340 268892 600596 268920
rect 582340 268880 582346 268892
rect 600590 268880 600596 268892
rect 600648 268880 600654 268932
rect 99282 268744 99288 268796
rect 99340 268784 99346 268796
rect 99340 268756 103514 268784
rect 99340 268744 99346 268756
rect 91002 268608 91008 268660
rect 91060 268648 91066 268660
rect 99282 268648 99288 268660
rect 91060 268620 99288 268648
rect 91060 268608 91066 268620
rect 99282 268608 99288 268620
rect 99340 268608 99346 268660
rect 103486 268648 103514 268756
rect 110230 268744 110236 268796
rect 110288 268784 110294 268796
rect 167914 268784 167920 268796
rect 110288 268756 167920 268784
rect 110288 268744 110294 268756
rect 167914 268744 167920 268756
rect 167972 268744 167978 268796
rect 173802 268744 173808 268796
rect 173860 268784 173866 268796
rect 212626 268784 212632 268796
rect 173860 268756 212632 268784
rect 173860 268744 173866 268756
rect 212626 268744 212632 268756
rect 212684 268744 212690 268796
rect 215202 268744 215208 268796
rect 215260 268784 215266 268796
rect 220814 268784 220820 268796
rect 215260 268756 220820 268784
rect 215260 268744 215266 268756
rect 220814 268744 220820 268756
rect 220872 268744 220878 268796
rect 377398 268744 377404 268796
rect 377456 268784 377462 268796
rect 408494 268784 408500 268796
rect 377456 268756 408500 268784
rect 377456 268744 377462 268756
rect 408494 268744 408500 268756
rect 408552 268744 408558 268796
rect 416406 268744 416412 268796
rect 416464 268784 416470 268796
rect 433334 268784 433340 268796
rect 416464 268756 433340 268784
rect 416464 268744 416470 268756
rect 433334 268744 433340 268756
rect 433392 268744 433398 268796
rect 441154 268744 441160 268796
rect 441212 268784 441218 268796
rect 498470 268784 498476 268796
rect 441212 268756 498476 268784
rect 441212 268744 441218 268756
rect 498470 268744 498476 268756
rect 498528 268744 498534 268796
rect 500678 268744 500684 268796
rect 500736 268784 500742 268796
rect 583846 268784 583852 268796
rect 500736 268756 583852 268784
rect 500736 268744 500742 268756
rect 583846 268744 583852 268756
rect 583904 268744 583910 268796
rect 160462 268648 160468 268660
rect 103486 268620 160468 268648
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 168650 268608 168656 268660
rect 168708 268648 168714 268660
rect 208486 268648 208492 268660
rect 168708 268620 208492 268648
rect 168708 268608 168714 268620
rect 208486 268608 208492 268620
rect 208544 268608 208550 268660
rect 208670 268608 208676 268660
rect 208728 268648 208734 268660
rect 214282 268648 214288 268660
rect 208728 268620 214288 268648
rect 208728 268608 208734 268620
rect 214282 268608 214288 268620
rect 214340 268608 214346 268660
rect 228082 268608 228088 268660
rect 228140 268648 228146 268660
rect 250714 268648 250720 268660
rect 228140 268620 250720 268648
rect 228140 268608 228146 268620
rect 250714 268608 250720 268620
rect 250772 268608 250778 268660
rect 256694 268608 256700 268660
rect 256752 268648 256758 268660
rect 263962 268648 263968 268660
rect 256752 268620 263968 268648
rect 256752 268608 256758 268620
rect 263962 268608 263968 268620
rect 264020 268608 264026 268660
rect 355870 268608 355876 268660
rect 355928 268648 355934 268660
rect 367830 268648 367836 268660
rect 355928 268620 367836 268648
rect 355928 268608 355934 268620
rect 367830 268608 367836 268620
rect 367888 268608 367894 268660
rect 372338 268608 372344 268660
rect 372396 268648 372402 268660
rect 385954 268648 385960 268660
rect 372396 268620 385960 268648
rect 372396 268608 372402 268620
rect 385954 268608 385960 268620
rect 386012 268608 386018 268660
rect 387334 268608 387340 268660
rect 387392 268648 387398 268660
rect 418522 268648 418528 268660
rect 387392 268620 418528 268648
rect 387392 268608 387398 268620
rect 418522 268608 418528 268620
rect 418580 268608 418586 268660
rect 443914 268608 443920 268660
rect 443972 268648 443978 268660
rect 502334 268648 502340 268660
rect 443972 268620 502340 268648
rect 443972 268608 443978 268620
rect 502334 268608 502340 268620
rect 502392 268608 502398 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 160002 268472 160008 268524
rect 160060 268512 160066 268524
rect 200390 268512 200396 268524
rect 160060 268484 200396 268512
rect 160060 268472 160066 268484
rect 200390 268472 200396 268484
rect 200448 268472 200454 268524
rect 212442 268472 212448 268524
rect 212500 268512 212506 268524
rect 238294 268512 238300 268524
rect 212500 268484 238300 268512
rect 212500 268472 212506 268484
rect 238294 268472 238300 268484
rect 238352 268472 238358 268524
rect 241330 268472 241336 268524
rect 241388 268512 241394 268524
rect 256694 268512 256700 268524
rect 241388 268484 256700 268512
rect 241388 268472 241394 268484
rect 256694 268472 256700 268484
rect 256752 268472 256758 268524
rect 266446 268472 266452 268524
rect 266504 268512 266510 268524
rect 275554 268512 275560 268524
rect 266504 268484 275560 268512
rect 266504 268472 266510 268484
rect 275554 268472 275560 268484
rect 275612 268472 275618 268524
rect 326062 268472 326068 268524
rect 326120 268512 326126 268524
rect 331398 268512 331404 268524
rect 326120 268484 331404 268512
rect 326120 268472 326126 268484
rect 331398 268472 331404 268484
rect 331456 268472 331462 268524
rect 335170 268472 335176 268524
rect 335228 268512 335234 268524
rect 347774 268512 347780 268524
rect 335228 268484 347780 268512
rect 335228 268472 335234 268484
rect 347774 268472 347780 268484
rect 347832 268472 347838 268524
rect 357526 268472 357532 268524
rect 357584 268512 357590 268524
rect 379514 268512 379520 268524
rect 357584 268484 379520 268512
rect 357584 268472 357590 268484
rect 379514 268472 379520 268484
rect 379572 268472 379578 268524
rect 398742 268472 398748 268524
rect 398800 268512 398806 268524
rect 430574 268512 430580 268524
rect 398800 268484 430580 268512
rect 398800 268472 398806 268484
rect 430574 268472 430580 268484
rect 430632 268472 430638 268524
rect 433702 268472 433708 268524
rect 433760 268512 433766 268524
rect 488534 268512 488540 268524
rect 433760 268484 488540 268512
rect 433760 268472 433766 268484
rect 488534 268472 488540 268484
rect 488592 268472 488598 268524
rect 510706 268472 510712 268524
rect 510764 268512 510770 268524
rect 598934 268512 598940 268524
rect 510764 268484 598940 268512
rect 510764 268472 510770 268484
rect 598934 268472 598940 268484
rect 598992 268472 598998 268524
rect 87138 268336 87144 268388
rect 87196 268376 87202 268388
rect 152182 268376 152188 268388
rect 87196 268348 152188 268376
rect 87196 268336 87202 268348
rect 152182 268336 152188 268348
rect 152240 268336 152246 268388
rect 152734 268336 152740 268388
rect 152792 268376 152798 268388
rect 196066 268376 196072 268388
rect 152792 268348 196072 268376
rect 152792 268336 152798 268348
rect 196066 268336 196072 268348
rect 196124 268336 196130 268388
rect 200574 268336 200580 268388
rect 200632 268376 200638 268388
rect 231670 268376 231676 268388
rect 200632 268348 231676 268376
rect 200632 268336 200638 268348
rect 231670 268336 231676 268348
rect 231728 268336 231734 268388
rect 234798 268336 234804 268388
rect 234856 268376 234862 268388
rect 255682 268376 255688 268388
rect 234856 268348 255688 268376
rect 234856 268336 234862 268348
rect 255682 268336 255688 268348
rect 255740 268336 255746 268388
rect 256510 268336 256516 268388
rect 256568 268376 256574 268388
rect 270586 268376 270592 268388
rect 256568 268348 270592 268376
rect 256568 268336 256574 268348
rect 270586 268336 270592 268348
rect 270644 268336 270650 268388
rect 276198 268336 276204 268388
rect 276256 268376 276262 268388
rect 280522 268376 280528 268388
rect 276256 268348 280528 268376
rect 276256 268336 276262 268348
rect 280522 268336 280528 268348
rect 280580 268336 280586 268388
rect 337654 268336 337660 268388
rect 337712 268376 337718 268388
rect 351914 268376 351920 268388
rect 337712 268348 351920 268376
rect 337712 268336 337718 268348
rect 351914 268336 351920 268348
rect 351972 268336 351978 268388
rect 352558 268336 352564 268388
rect 352616 268376 352622 268388
rect 368750 268376 368756 268388
rect 352616 268348 368756 268376
rect 352616 268336 352622 268348
rect 368750 268336 368756 268348
rect 368808 268336 368814 268388
rect 369946 268336 369952 268388
rect 370004 268376 370010 268388
rect 397454 268376 397460 268388
rect 370004 268348 397460 268376
rect 370004 268336 370010 268348
rect 397454 268336 397460 268348
rect 397512 268336 397518 268388
rect 399754 268336 399760 268388
rect 399812 268376 399818 268388
rect 440234 268376 440240 268388
rect 399812 268348 440240 268376
rect 399812 268336 399818 268348
rect 440234 268336 440240 268348
rect 440292 268336 440298 268388
rect 459554 268336 459560 268388
rect 459612 268376 459618 268388
rect 517606 268376 517612 268388
rect 459612 268348 517612 268376
rect 459612 268336 459618 268348
rect 517606 268336 517612 268348
rect 517664 268336 517670 268388
rect 534718 268336 534724 268388
rect 534776 268376 534782 268388
rect 535730 268376 535736 268388
rect 534776 268348 535736 268376
rect 534776 268336 534782 268348
rect 535730 268336 535736 268348
rect 535788 268336 535794 268388
rect 536374 268336 536380 268388
rect 536432 268376 536438 268388
rect 634814 268376 634820 268388
rect 536432 268348 634820 268376
rect 536432 268336 536438 268348
rect 634814 268336 634820 268348
rect 634872 268336 634878 268388
rect 118602 268200 118608 268252
rect 118660 268240 118666 268252
rect 174538 268240 174544 268252
rect 118660 268212 174544 268240
rect 118660 268200 118666 268212
rect 174538 268200 174544 268212
rect 174596 268200 174602 268252
rect 413002 268200 413008 268252
rect 413060 268240 413066 268252
rect 459738 268240 459744 268252
rect 413060 268212 459744 268240
rect 413060 268200 413066 268212
rect 459738 268200 459744 268212
rect 459796 268200 459802 268252
rect 469490 268200 469496 268252
rect 469548 268240 469554 268252
rect 475378 268240 475384 268252
rect 469548 268212 475384 268240
rect 469548 268200 469554 268212
rect 475378 268200 475384 268212
rect 475436 268200 475442 268252
rect 490834 268200 490840 268252
rect 490892 268240 490898 268252
rect 569954 268240 569960 268252
rect 490892 268212 569960 268240
rect 490892 268200 490898 268212
rect 569954 268200 569960 268212
rect 570012 268200 570018 268252
rect 137002 268064 137008 268116
rect 137060 268104 137066 268116
rect 182174 268104 182180 268116
rect 137060 268076 182180 268104
rect 137060 268064 137066 268076
rect 182174 268064 182180 268076
rect 182232 268064 182238 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 443270 268104 443276 268116
rect 422352 268076 443276 268104
rect 422352 268064 422358 268076
rect 443270 268064 443276 268076
rect 443328 268064 443334 268116
rect 475194 268064 475200 268116
rect 475252 268104 475258 268116
rect 478966 268104 478972 268116
rect 475252 268076 478972 268104
rect 475252 268064 475258 268076
rect 478966 268064 478972 268076
rect 479024 268064 479030 268116
rect 489178 268064 489184 268116
rect 489236 268104 489242 268116
rect 567286 268104 567292 268116
rect 489236 268076 567292 268104
rect 489236 268064 489242 268076
rect 567286 268064 567292 268076
rect 567344 268064 567350 268116
rect 448606 267928 448612 267980
rect 448664 267968 448670 267980
rect 506474 267968 506480 267980
rect 448664 267940 506480 267968
rect 448664 267928 448670 267940
rect 506474 267928 506480 267940
rect 506532 267928 506538 267980
rect 436186 267792 436192 267844
rect 436244 267832 436250 267844
rect 491846 267832 491852 267844
rect 436244 267804 491852 267832
rect 436244 267792 436250 267804
rect 491846 267792 491852 267804
rect 491904 267792 491910 267844
rect 493318 267792 493324 267844
rect 493376 267832 493382 267844
rect 551278 267832 551284 267844
rect 493376 267804 551284 267832
rect 493376 267792 493382 267804
rect 551278 267792 551284 267804
rect 551336 267792 551342 267844
rect 328546 267724 328552 267776
rect 328604 267764 328610 267776
rect 337102 267764 337108 267776
rect 328604 267736 337108 267764
rect 328604 267724 328610 267736
rect 337102 267724 337108 267736
rect 337160 267724 337166 267776
rect 356054 267764 356060 267776
rect 347746 267736 356060 267764
rect 132402 267656 132408 267708
rect 132460 267696 132466 267708
rect 184474 267696 184480 267708
rect 132460 267668 184480 267696
rect 132460 267656 132466 267668
rect 184474 267656 184480 267668
rect 184532 267656 184538 267708
rect 189810 267656 189816 267708
rect 189868 267696 189874 267708
rect 197722 267696 197728 267708
rect 189868 267668 197728 267696
rect 189868 267656 189874 267668
rect 197722 267656 197728 267668
rect 197780 267656 197786 267708
rect 204162 267656 204168 267708
rect 204220 267696 204226 267708
rect 218422 267696 218428 267708
rect 204220 267668 218428 267696
rect 204220 267656 204226 267668
rect 218422 267656 218428 267668
rect 218480 267656 218486 267708
rect 224218 267656 224224 267708
rect 224276 267696 224282 267708
rect 229186 267696 229192 267708
rect 224276 267668 229192 267696
rect 224276 267656 224282 267668
rect 229186 267656 229192 267668
rect 229244 267656 229250 267708
rect 99282 267520 99288 267572
rect 99340 267560 99346 267572
rect 154666 267560 154672 267572
rect 99340 267532 154672 267560
rect 99340 267520 99346 267532
rect 154666 267520 154672 267532
rect 154724 267520 154730 267572
rect 167638 267520 167644 267572
rect 167696 267560 167702 267572
rect 186958 267560 186964 267572
rect 167696 267532 186964 267560
rect 167696 267520 167702 267532
rect 186958 267520 186964 267532
rect 187016 267520 187022 267572
rect 195238 267520 195244 267572
rect 195296 267560 195302 267572
rect 216766 267560 216772 267572
rect 195296 267532 216772 267560
rect 195296 267520 195302 267532
rect 216766 267520 216772 267532
rect 216824 267520 216830 267572
rect 218790 267520 218796 267572
rect 218848 267560 218854 267572
rect 226702 267560 226708 267572
rect 218848 267532 226708 267560
rect 218848 267520 218854 267532
rect 226702 267520 226708 267532
rect 226760 267520 226766 267572
rect 107654 267384 107660 267436
rect 107712 267424 107718 267436
rect 167086 267424 167092 267436
rect 107712 267396 167092 267424
rect 107712 267384 107718 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 170398 267384 170404 267436
rect 170456 267424 170462 267436
rect 170456 267396 173756 267424
rect 170456 267384 170462 267396
rect 95878 267248 95884 267300
rect 95936 267288 95942 267300
rect 156414 267288 156420 267300
rect 95936 267260 156420 267288
rect 95936 267248 95942 267260
rect 156414 267248 156420 267260
rect 156472 267248 156478 267300
rect 156598 267248 156604 267300
rect 156656 267288 156662 267300
rect 159634 267288 159640 267300
rect 156656 267260 159640 267288
rect 156656 267248 156662 267260
rect 159634 267248 159640 267260
rect 159692 267248 159698 267300
rect 160738 267248 160744 267300
rect 160796 267288 160802 267300
rect 164602 267288 164608 267300
rect 160796 267260 164608 267288
rect 160796 267248 160802 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 166442 267248 166448 267300
rect 166500 267288 166506 267300
rect 172882 267288 172888 267300
rect 166500 267260 172888 267288
rect 166500 267248 166506 267260
rect 172882 267248 172888 267260
rect 172940 267248 172946 267300
rect 173728 267288 173756 267396
rect 186314 267384 186320 267436
rect 186372 267424 186378 267436
rect 221734 267424 221740 267436
rect 186372 267396 221740 267424
rect 186372 267384 186378 267396
rect 221734 267384 221740 267396
rect 221792 267384 221798 267436
rect 227714 267384 227720 267436
rect 227772 267424 227778 267436
rect 236638 267424 236644 267436
rect 227772 267396 236644 267424
rect 227772 267384 227778 267396
rect 236638 267384 236644 267396
rect 236696 267384 236702 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 347746 267424 347774 267736
rect 356054 267724 356060 267736
rect 356112 267724 356118 267776
rect 368106 267656 368112 267708
rect 368164 267696 368170 267708
rect 378778 267696 378784 267708
rect 368164 267668 378784 267696
rect 368164 267656 368170 267668
rect 378778 267656 378784 267668
rect 378836 267656 378842 267708
rect 380618 267656 380624 267708
rect 380676 267696 380682 267708
rect 393314 267696 393320 267708
rect 380676 267668 393320 267696
rect 380676 267656 380682 267668
rect 393314 267656 393320 267668
rect 393372 267656 393378 267708
rect 402238 267656 402244 267708
rect 402296 267696 402302 267708
rect 422294 267696 422300 267708
rect 402296 267668 422300 267696
rect 402296 267656 402302 267668
rect 422294 267656 422300 267668
rect 422352 267656 422358 267708
rect 430390 267656 430396 267708
rect 430448 267696 430454 267708
rect 458818 267696 458824 267708
rect 430448 267668 458824 267696
rect 430448 267656 430454 267668
rect 458818 267656 458824 267668
rect 458876 267656 458882 267708
rect 460198 267656 460204 267708
rect 460256 267696 460262 267708
rect 512546 267696 512552 267708
rect 460256 267668 512552 267696
rect 460256 267656 460262 267668
rect 512546 267656 512552 267668
rect 512604 267656 512610 267708
rect 514386 267656 514392 267708
rect 514444 267696 514450 267708
rect 541618 267696 541624 267708
rect 514444 267668 541624 267696
rect 514444 267656 514450 267668
rect 541618 267656 541624 267668
rect 541676 267656 541682 267708
rect 357066 267520 357072 267572
rect 357124 267560 357130 267572
rect 357124 267532 364334 267560
rect 357124 267520 357130 267532
rect 341024 267396 347774 267424
rect 341024 267384 341030 267396
rect 358354 267384 358360 267436
rect 358412 267424 358418 267436
rect 360838 267424 360844 267436
rect 358412 267396 360844 267424
rect 358412 267384 358418 267396
rect 360838 267384 360844 267396
rect 360896 267384 360902 267436
rect 364306 267424 364334 267532
rect 373258 267520 373264 267572
rect 373316 267560 373322 267572
rect 387702 267560 387708 267572
rect 373316 267532 387708 267560
rect 373316 267520 373322 267532
rect 387702 267520 387708 267532
rect 387760 267520 387766 267572
rect 404722 267520 404728 267572
rect 404780 267560 404786 267572
rect 429838 267560 429844 267572
rect 404780 267532 429844 267560
rect 404780 267520 404786 267532
rect 429838 267520 429844 267532
rect 429896 267520 429902 267572
rect 436738 267520 436744 267572
rect 436796 267560 436802 267572
rect 441614 267560 441620 267572
rect 436796 267532 441620 267560
rect 436796 267520 436802 267532
rect 441614 267520 441620 267532
rect 441672 267520 441678 267572
rect 442810 267520 442816 267572
rect 442868 267560 442874 267572
rect 485038 267560 485044 267572
rect 442868 267532 485044 267560
rect 442868 267520 442874 267532
rect 485038 267520 485044 267532
rect 485096 267520 485102 267572
rect 487154 267520 487160 267572
rect 487212 267560 487218 267572
rect 487798 267560 487804 267572
rect 487212 267532 487804 267560
rect 487212 267520 487218 267532
rect 487798 267520 487804 267532
rect 487856 267520 487862 267572
rect 494698 267520 494704 267572
rect 494756 267560 494762 267572
rect 501598 267560 501604 267572
rect 494756 267532 501604 267560
rect 494756 267520 494762 267532
rect 501598 267520 501604 267532
rect 501656 267520 501662 267572
rect 502426 267520 502432 267572
rect 502484 267560 502490 267572
rect 502484 267532 506060 267560
rect 502484 267520 502490 267532
rect 366358 267424 366364 267436
rect 364306 267396 366364 267424
rect 366358 267384 366364 267396
rect 366416 267384 366422 267436
rect 375742 267384 375748 267436
rect 375800 267424 375806 267436
rect 389634 267424 389640 267436
rect 375800 267396 389640 267424
rect 375800 267384 375806 267396
rect 389634 267384 389640 267396
rect 389692 267384 389698 267436
rect 394786 267384 394792 267436
rect 394844 267424 394850 267436
rect 416406 267424 416412 267436
rect 394844 267396 416412 267424
rect 394844 267384 394850 267396
rect 416406 267384 416412 267396
rect 416464 267384 416470 267436
rect 419626 267384 419632 267436
rect 419684 267424 419690 267436
rect 446398 267424 446404 267436
rect 419684 267396 446404 267424
rect 419684 267384 419690 267396
rect 446398 267384 446404 267396
rect 446456 267384 446462 267436
rect 450262 267384 450268 267436
rect 450320 267424 450326 267436
rect 505830 267424 505836 267436
rect 450320 267396 505836 267424
rect 450320 267384 450326 267396
rect 505830 267384 505836 267396
rect 505888 267384 505894 267436
rect 506032 267424 506060 267532
rect 507578 267520 507584 267572
rect 507636 267560 507642 267572
rect 576118 267560 576124 267572
rect 507636 267532 576124 267560
rect 507636 267520 507642 267532
rect 576118 267520 576124 267532
rect 576176 267520 576182 267572
rect 508406 267424 508412 267436
rect 506032 267396 508412 267424
rect 508406 267384 508412 267396
rect 508464 267384 508470 267436
rect 509878 267384 509884 267436
rect 509936 267424 509942 267436
rect 517790 267424 517796 267436
rect 509936 267396 517796 267424
rect 509936 267384 509942 267396
rect 517790 267384 517796 267396
rect 517848 267384 517854 267436
rect 582282 267424 582288 267436
rect 518866 267396 582288 267424
rect 173728 267260 206140 267288
rect 86218 267112 86224 267164
rect 86276 267152 86282 267164
rect 148042 267152 148048 267164
rect 86276 267124 148048 267152
rect 86276 267112 86282 267124
rect 148042 267112 148048 267124
rect 148100 267112 148106 267164
rect 149698 267112 149704 267164
rect 149756 267152 149762 267164
rect 194410 267152 194416 267164
rect 149756 267124 194416 267152
rect 149756 267112 149762 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 199286 267112 199292 267164
rect 199344 267152 199350 267164
rect 201862 267152 201868 267164
rect 199344 267124 201868 267152
rect 199344 267112 199350 267124
rect 201862 267112 201868 267124
rect 201920 267112 201926 267164
rect 206112 267152 206140 267260
rect 206278 267248 206284 267300
rect 206336 267288 206342 267300
rect 213454 267288 213460 267300
rect 206336 267260 213460 267288
rect 206336 267248 206342 267260
rect 213454 267248 213460 267260
rect 213512 267248 213518 267300
rect 217410 267248 217416 267300
rect 217468 267288 217474 267300
rect 219894 267288 219900 267300
rect 217468 267260 219900 267288
rect 217468 267248 217474 267260
rect 219894 267248 219900 267260
rect 219952 267248 219958 267300
rect 220078 267248 220084 267300
rect 220136 267288 220142 267300
rect 222562 267288 222568 267300
rect 220136 267260 222568 267288
rect 220136 267248 220142 267260
rect 222562 267248 222568 267260
rect 222620 267248 222626 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 234154 267288 234160 267300
rect 223540 267260 234160 267288
rect 223540 267248 223546 267260
rect 234154 267248 234160 267260
rect 234212 267248 234218 267300
rect 238018 267248 238024 267300
rect 238076 267288 238082 267300
rect 251542 267288 251548 267300
rect 238076 267260 251548 267288
rect 238076 267248 238082 267260
rect 251542 267248 251548 267260
rect 251600 267248 251606 267300
rect 261478 267248 261484 267300
rect 261536 267288 261542 267300
rect 268930 267288 268936 267300
rect 261536 267260 268936 267288
rect 261536 267248 261542 267260
rect 268930 267248 268936 267260
rect 268988 267248 268994 267300
rect 334342 267248 334348 267300
rect 334400 267288 334406 267300
rect 344278 267288 344284 267300
rect 334400 267260 344284 267288
rect 334400 267248 334406 267260
rect 344278 267248 344284 267260
rect 344336 267248 344342 267300
rect 360838 267248 360844 267300
rect 360896 267288 360902 267300
rect 373074 267288 373080 267300
rect 360896 267260 373080 267288
rect 360896 267248 360902 267260
rect 373074 267248 373080 267260
rect 373132 267248 373138 267300
rect 378226 267248 378232 267300
rect 378284 267288 378290 267300
rect 378284 267260 385540 267288
rect 378284 267248 378290 267260
rect 206830 267152 206836 267164
rect 206112 267124 206836 267152
rect 206830 267112 206836 267124
rect 206888 267112 206894 267164
rect 207014 267112 207020 267164
rect 207072 267152 207078 267164
rect 207072 267124 214604 267152
rect 207072 267112 207078 267124
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 141418 267016 141424 267028
rect 73856 266988 141424 267016
rect 73856 266976 73862 266988
rect 141418 266976 141424 266988
rect 141476 266976 141482 267028
rect 146938 266976 146944 267028
rect 146996 267016 147002 267028
rect 189442 267016 189448 267028
rect 146996 266988 189448 267016
rect 146996 266976 147002 266988
rect 189442 266976 189448 266988
rect 189500 266976 189506 267028
rect 191098 266976 191104 267028
rect 191156 267016 191162 267028
rect 211798 267016 211804 267028
rect 191156 266988 211804 267016
rect 191156 266976 191162 266988
rect 211798 266976 211804 266988
rect 211856 266976 211862 267028
rect 214576 267016 214604 267124
rect 215938 267112 215944 267164
rect 215996 267152 216002 267164
rect 220078 267152 220084 267164
rect 215996 267124 220084 267152
rect 215996 267112 216002 267124
rect 220078 267112 220084 267124
rect 220136 267112 220142 267164
rect 220814 267112 220820 267164
rect 220872 267152 220878 267164
rect 241606 267152 241612 267164
rect 220872 267124 241612 267152
rect 220872 267112 220878 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 243906 267112 243912 267164
rect 243964 267152 243970 267164
rect 254854 267152 254860 267164
rect 243964 267124 254860 267152
rect 243964 267112 243970 267124
rect 254854 267112 254860 267124
rect 254912 267112 254918 267164
rect 282822 267112 282828 267164
rect 282880 267152 282886 267164
rect 288802 267152 288808 267164
rect 282880 267124 288808 267152
rect 282880 267112 282886 267124
rect 288802 267112 288808 267124
rect 288860 267112 288866 267164
rect 324406 267112 324412 267164
rect 324464 267152 324470 267164
rect 330478 267152 330484 267164
rect 324464 267124 330484 267152
rect 324464 267112 324470 267124
rect 330478 267112 330484 267124
rect 330536 267112 330542 267164
rect 333514 267112 333520 267164
rect 333572 267152 333578 267164
rect 342254 267152 342260 267164
rect 333572 267124 342260 267152
rect 333572 267112 333578 267124
rect 342254 267112 342260 267124
rect 342312 267112 342318 267164
rect 350902 267112 350908 267164
rect 350960 267152 350966 267164
rect 359458 267152 359464 267164
rect 350960 267124 359464 267152
rect 350960 267112 350966 267124
rect 359458 267112 359464 267124
rect 359516 267112 359522 267164
rect 363322 267112 363328 267164
rect 363380 267152 363386 267164
rect 377950 267152 377956 267164
rect 363380 267124 377956 267152
rect 363380 267112 363386 267124
rect 377950 267112 377956 267124
rect 378008 267112 378014 267164
rect 383838 267152 383844 267164
rect 383626 267124 383844 267152
rect 220906 267016 220912 267028
rect 214576 266988 220912 267016
rect 220906 266976 220912 266988
rect 220964 266976 220970 267028
rect 222010 266976 222016 267028
rect 222068 267016 222074 267028
rect 246574 267016 246580 267028
rect 222068 266988 246580 267016
rect 222068 266976 222074 266988
rect 246574 266976 246580 266988
rect 246632 266976 246638 267028
rect 249058 266976 249064 267028
rect 249116 267016 249122 267028
rect 261478 267016 261484 267028
rect 249116 266988 261484 267016
rect 249116 266976 249122 266988
rect 261478 266976 261484 266988
rect 261536 266976 261542 267028
rect 276014 266976 276020 267028
rect 276072 267016 276078 267028
rect 283834 267016 283840 267028
rect 276072 266988 283840 267016
rect 276072 266976 276078 266988
rect 283834 266976 283840 266988
rect 283892 266976 283898 267028
rect 343358 266976 343364 267028
rect 343416 267016 343422 267028
rect 352374 267016 352380 267028
rect 343416 266988 352380 267016
rect 343416 266976 343422 266988
rect 352374 266976 352380 266988
rect 352432 266976 352438 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 363598 267016 363604 267028
rect 353444 266988 363604 267016
rect 353444 266976 353450 266988
rect 363598 266976 363604 266988
rect 363656 266976 363662 267028
rect 365806 266976 365812 267028
rect 365864 267016 365870 267028
rect 383626 267016 383654 267124
rect 383838 267112 383844 267124
rect 383896 267112 383902 267164
rect 365864 266988 383654 267016
rect 385512 267016 385540 267260
rect 389818 267248 389824 267300
rect 389876 267288 389882 267300
rect 395338 267288 395344 267300
rect 389876 267260 395344 267288
rect 389876 267248 389882 267260
rect 395338 267248 395344 267260
rect 395396 267248 395402 267300
rect 397086 267248 397092 267300
rect 397144 267288 397150 267300
rect 421558 267288 421564 267300
rect 397144 267260 421564 267288
rect 397144 267248 397150 267260
rect 421558 267248 421564 267260
rect 421616 267248 421622 267300
rect 426066 267248 426072 267300
rect 426124 267288 426130 267300
rect 453298 267288 453304 267300
rect 426124 267260 453304 267288
rect 426124 267248 426130 267260
rect 453298 267248 453304 267260
rect 453356 267248 453362 267300
rect 455230 267248 455236 267300
rect 455288 267288 455294 267300
rect 510522 267288 510528 267300
rect 455288 267260 510528 267288
rect 455288 267248 455294 267260
rect 510522 267248 510528 267260
rect 510580 267248 510586 267300
rect 512362 267248 512368 267300
rect 512420 267288 512426 267300
rect 518866 267288 518894 267396
rect 582282 267384 582288 267396
rect 582340 267384 582346 267436
rect 512420 267260 518894 267288
rect 512420 267248 512426 267260
rect 520642 267248 520648 267300
rect 520700 267288 520706 267300
rect 537478 267288 537484 267300
rect 520700 267260 537484 267288
rect 520700 267248 520706 267260
rect 537478 267248 537484 267260
rect 537536 267248 537542 267300
rect 539686 267248 539692 267300
rect 539744 267288 539750 267300
rect 540882 267288 540888 267300
rect 539744 267260 540888 267288
rect 539744 267248 539750 267260
rect 540882 267248 540888 267260
rect 540940 267248 540946 267300
rect 541342 267248 541348 267300
rect 541400 267288 541406 267300
rect 542170 267288 542176 267300
rect 541400 267260 542176 267288
rect 541400 267248 541406 267260
rect 542170 267248 542176 267260
rect 542228 267248 542234 267300
rect 542354 267248 542360 267300
rect 542412 267288 542418 267300
rect 623038 267288 623044 267300
rect 542412 267260 623044 267288
rect 542412 267248 542418 267260
rect 623038 267248 623044 267260
rect 623096 267248 623102 267300
rect 385678 267112 385684 267164
rect 385736 267152 385742 267164
rect 401686 267152 401692 267164
rect 385736 267124 401692 267152
rect 385736 267112 385742 267124
rect 401686 267112 401692 267124
rect 401744 267112 401750 267164
rect 414658 267112 414664 267164
rect 414716 267152 414722 267164
rect 436738 267152 436744 267164
rect 414716 267124 436744 267152
rect 414716 267112 414722 267124
rect 436738 267112 436744 267124
rect 436796 267112 436802 267164
rect 440326 267112 440332 267164
rect 440384 267152 440390 267164
rect 443638 267152 443644 267164
rect 440384 267124 443644 267152
rect 440384 267112 440390 267124
rect 443638 267112 443644 267124
rect 443696 267112 443702 267164
rect 445294 267112 445300 267164
rect 445352 267152 445358 267164
rect 494698 267152 494704 267164
rect 445352 267124 494704 267152
rect 445352 267112 445358 267124
rect 494698 267112 494704 267124
rect 494756 267112 494762 267164
rect 494882 267112 494888 267164
rect 494940 267152 494946 267164
rect 507302 267152 507308 267164
rect 494940 267124 507308 267152
rect 494940 267112 494946 267124
rect 507302 267112 507308 267124
rect 507360 267112 507366 267164
rect 508222 267112 508228 267164
rect 508280 267152 508286 267164
rect 522390 267152 522396 267164
rect 508280 267124 522396 267152
rect 508280 267112 508286 267124
rect 522390 267112 522396 267124
rect 522448 267112 522454 267164
rect 522666 267112 522672 267164
rect 522724 267152 522730 267164
rect 526622 267152 526628 267164
rect 522724 267124 526628 267152
rect 522724 267112 522730 267124
rect 526622 267112 526628 267124
rect 526680 267112 526686 267164
rect 532234 267112 532240 267164
rect 532292 267152 532298 267164
rect 596818 267152 596824 267164
rect 532292 267124 596824 267152
rect 532292 267112 532298 267124
rect 596818 267112 596824 267124
rect 596876 267112 596882 267164
rect 391934 267016 391940 267028
rect 385512 266988 391940 267016
rect 365864 266976 365870 266988
rect 391934 266976 391940 266988
rect 391992 266976 391998 267028
rect 392302 266976 392308 267028
rect 392360 267016 392366 267028
rect 418982 267016 418988 267028
rect 392360 266988 418988 267016
rect 392360 266976 392366 266988
rect 418982 266976 418988 266988
rect 419040 266976 419046 267028
rect 422938 266976 422944 267028
rect 422996 267016 423002 267028
rect 454494 267016 454500 267028
rect 422996 266988 454500 267016
rect 422996 266976 423002 266988
rect 454494 266976 454500 266988
rect 454552 266976 454558 267028
rect 454770 266976 454776 267028
rect 454828 267016 454834 267028
rect 459186 267016 459192 267028
rect 454828 266988 459192 267016
rect 454828 266976 454834 266988
rect 459186 266976 459192 266988
rect 459244 266976 459250 267028
rect 459370 266976 459376 267028
rect 459428 267016 459434 267028
rect 467098 267016 467104 267028
rect 459428 266988 467104 267016
rect 459428 266976 459434 266988
rect 467098 266976 467104 266988
rect 467156 266976 467162 267028
rect 467282 266976 467288 267028
rect 467340 267016 467346 267028
rect 469490 267016 469496 267028
rect 467340 266988 469496 267016
rect 467340 266976 467346 266988
rect 469490 266976 469496 266988
rect 469548 266976 469554 267028
rect 530670 267016 530676 267028
rect 470566 266988 530676 267016
rect 119798 266840 119804 266892
rect 119856 266880 119862 266892
rect 156598 266880 156604 266892
rect 119856 266852 156604 266880
rect 119856 266840 119862 266852
rect 156598 266840 156604 266852
rect 156656 266840 156662 266892
rect 169846 266840 169852 266892
rect 169904 266880 169910 266892
rect 169904 266852 180794 266880
rect 169904 266840 169910 266852
rect 132586 266704 132592 266756
rect 132644 266744 132650 266756
rect 147214 266744 147220 266756
rect 132644 266716 147220 266744
rect 132644 266704 132650 266716
rect 147214 266704 147220 266716
rect 147272 266704 147278 266756
rect 148502 266704 148508 266756
rect 148560 266744 148566 266756
rect 179506 266744 179512 266756
rect 148560 266716 179512 266744
rect 148560 266704 148566 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 180766 266744 180794 266852
rect 198182 266840 198188 266892
rect 198240 266880 198246 266892
rect 200206 266880 200212 266892
rect 198240 266852 200212 266880
rect 198240 266840 198246 266852
rect 200206 266840 200212 266852
rect 200264 266840 200270 266892
rect 202322 266840 202328 266892
rect 202380 266880 202386 266892
rect 207014 266880 207020 266892
rect 202380 266852 207020 266880
rect 202380 266840 202386 266852
rect 207014 266840 207020 266852
rect 207072 266840 207078 266892
rect 219894 266840 219900 266892
rect 219952 266880 219958 266892
rect 223390 266880 223396 266892
rect 219952 266852 223396 266880
rect 219952 266840 219958 266852
rect 223390 266840 223396 266852
rect 223448 266840 223454 266892
rect 242250 266840 242256 266892
rect 242308 266880 242314 266892
rect 249058 266880 249064 266892
rect 242308 266852 249064 266880
rect 242308 266840 242314 266852
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 251818 266840 251824 266892
rect 251876 266880 251882 266892
rect 258994 266880 259000 266892
rect 251876 266852 259000 266880
rect 251876 266840 251882 266852
rect 258994 266840 259000 266852
rect 259052 266840 259058 266892
rect 264974 266840 264980 266892
rect 265032 266880 265038 266892
rect 276382 266880 276388 266892
rect 265032 266852 276388 266880
rect 265032 266840 265038 266852
rect 276382 266840 276388 266852
rect 276440 266840 276446 266892
rect 285674 266840 285680 266892
rect 285732 266880 285738 266892
rect 287974 266880 287980 266892
rect 285732 266852 287980 266880
rect 285732 266840 285738 266852
rect 287974 266840 287980 266852
rect 288032 266840 288038 266892
rect 312814 266840 312820 266892
rect 312872 266880 312878 266892
rect 316402 266880 316408 266892
rect 312872 266852 316408 266880
rect 312872 266840 312878 266852
rect 316402 266840 316408 266852
rect 316460 266840 316466 266892
rect 321922 266840 321928 266892
rect 321980 266880 321986 266892
rect 327074 266880 327080 266892
rect 321980 266852 327080 266880
rect 321980 266840 321986 266852
rect 327074 266840 327080 266852
rect 327132 266840 327138 266892
rect 349246 266840 349252 266892
rect 349304 266880 349310 266892
rect 355318 266880 355324 266892
rect 349304 266852 355324 266880
rect 349304 266840 349310 266852
rect 355318 266840 355324 266852
rect 355376 266840 355382 266892
rect 393130 266840 393136 266892
rect 393188 266880 393194 266892
rect 398742 266880 398748 266892
rect 393188 266852 398748 266880
rect 393188 266840 393194 266852
rect 398742 266840 398748 266852
rect 398800 266840 398806 266892
rect 403066 266840 403072 266892
rect 403124 266880 403130 266892
rect 404170 266880 404176 266892
rect 403124 266852 404176 266880
rect 403124 266840 403130 266852
rect 404170 266840 404176 266852
rect 404228 266840 404234 266892
rect 405550 266840 405556 266892
rect 405608 266880 405614 266892
rect 425698 266880 425704 266892
rect 405608 266852 425704 266880
rect 405608 266840 405614 266852
rect 425698 266840 425704 266852
rect 425756 266840 425762 266892
rect 438118 266880 438124 266892
rect 431926 266852 438124 266880
rect 199378 266744 199384 266756
rect 180766 266716 199384 266744
rect 199378 266704 199384 266716
rect 199436 266704 199442 266756
rect 232682 266704 232688 266756
rect 232740 266744 232746 266756
rect 239122 266744 239128 266756
rect 232740 266716 239128 266744
rect 232740 266704 232746 266716
rect 239122 266704 239128 266716
rect 239180 266704 239186 266756
rect 317782 266704 317788 266756
rect 317840 266744 317846 266756
rect 322934 266744 322940 266756
rect 317840 266716 322940 266744
rect 317840 266704 317846 266716
rect 322934 266704 322940 266716
rect 322992 266704 322998 266756
rect 390646 266704 390652 266756
rect 390704 266744 390710 266756
rect 395522 266744 395528 266756
rect 390704 266716 395528 266744
rect 390704 266704 390710 266716
rect 395522 266704 395528 266716
rect 395580 266704 395586 266756
rect 398098 266704 398104 266756
rect 398156 266744 398162 266756
rect 414474 266744 414480 266756
rect 398156 266716 414480 266744
rect 398156 266704 398162 266716
rect 414474 266704 414480 266716
rect 414532 266704 414538 266756
rect 423766 266704 423772 266756
rect 423824 266744 423830 266756
rect 424962 266744 424968 266756
rect 423824 266716 424968 266744
rect 423824 266704 423830 266716
rect 424962 266704 424968 266716
rect 425020 266704 425026 266756
rect 425422 266704 425428 266756
rect 425480 266744 425486 266756
rect 426250 266744 426256 266756
rect 425480 266716 426256 266744
rect 425480 266704 425486 266716
rect 426250 266704 426256 266716
rect 426308 266704 426314 266756
rect 427906 266704 427912 266756
rect 427964 266744 427970 266756
rect 428918 266744 428924 266756
rect 427964 266716 428924 266744
rect 427964 266704 427970 266716
rect 428918 266704 428924 266716
rect 428976 266704 428982 266756
rect 312354 266636 312360 266688
rect 312412 266676 312418 266688
rect 314654 266676 314660 266688
rect 312412 266648 314660 266676
rect 312412 266636 312418 266648
rect 314654 266636 314660 266648
rect 314712 266636 314718 266688
rect 123478 266568 123484 266620
rect 123536 266608 123542 266620
rect 150526 266608 150532 266620
rect 123536 266580 150532 266608
rect 123536 266568 123542 266580
rect 150526 266568 150532 266580
rect 150584 266568 150590 266620
rect 154022 266568 154028 266620
rect 154080 266608 154086 266620
rect 161934 266608 161940 266620
rect 154080 266580 161940 266608
rect 154080 266568 154086 266580
rect 161934 266568 161940 266580
rect 161992 266568 161998 266620
rect 162118 266568 162124 266620
rect 162176 266608 162182 266620
rect 162946 266608 162952 266620
rect 162176 266580 162952 266608
rect 162176 266568 162182 266580
rect 162946 266568 162952 266580
rect 163004 266568 163010 266620
rect 195238 266608 195244 266620
rect 190426 266580 195244 266608
rect 170398 266540 170404 266552
rect 164896 266512 170404 266540
rect 141602 266432 141608 266484
rect 141660 266472 141666 266484
rect 146938 266472 146944 266484
rect 141660 266444 146944 266472
rect 141660 266432 141666 266444
rect 146938 266432 146944 266444
rect 146996 266432 147002 266484
rect 156598 266432 156604 266484
rect 156656 266472 156662 266484
rect 162118 266472 162124 266484
rect 156656 266444 162124 266472
rect 156656 266432 156662 266444
rect 162118 266432 162124 266444
rect 162176 266432 162182 266484
rect 164896 266472 164924 266512
rect 170398 266500 170404 266512
rect 170456 266500 170462 266552
rect 182174 266500 182180 266552
rect 182232 266540 182238 266552
rect 186130 266540 186136 266552
rect 182232 266512 186136 266540
rect 182232 266500 182238 266512
rect 186130 266500 186136 266512
rect 186188 266500 186194 266552
rect 162320 266444 164924 266472
rect 161934 266296 161940 266348
rect 161992 266336 161998 266348
rect 162320 266336 162348 266444
rect 165062 266364 165068 266416
rect 165120 266404 165126 266416
rect 169570 266404 169576 266416
rect 165120 266376 169576 266404
rect 165120 266364 165126 266376
rect 169570 266364 169576 266376
rect 169628 266364 169634 266416
rect 181530 266364 181536 266416
rect 181588 266404 181594 266416
rect 182818 266404 182824 266416
rect 181588 266376 182824 266404
rect 181588 266364 181594 266376
rect 182818 266364 182824 266376
rect 182876 266364 182882 266416
rect 184198 266364 184204 266416
rect 184256 266404 184262 266416
rect 190426 266404 190454 266580
rect 195238 266568 195244 266580
rect 195296 266568 195302 266620
rect 316126 266568 316132 266620
rect 316184 266608 316190 266620
rect 320542 266608 320548 266620
rect 316184 266580 320548 266608
rect 316184 266568 316190 266580
rect 320542 266568 320548 266580
rect 320600 266568 320606 266620
rect 418798 266568 418804 266620
rect 418856 266608 418862 266620
rect 431926 266608 431954 266852
rect 438118 266840 438124 266852
rect 438176 266840 438182 266892
rect 446950 266840 446956 266892
rect 447008 266880 447014 266892
rect 456058 266880 456064 266892
rect 447008 266852 456064 266880
rect 447008 266840 447014 266852
rect 456058 266840 456064 266852
rect 456116 266840 456122 266892
rect 457714 266840 457720 266892
rect 457772 266880 457778 266892
rect 464430 266880 464436 266892
rect 457772 266852 464436 266880
rect 457772 266840 457778 266852
rect 464430 266840 464436 266852
rect 464488 266840 464494 266892
rect 469950 266880 469956 266892
rect 464632 266852 469956 266880
rect 437842 266704 437848 266756
rect 437900 266744 437906 266756
rect 437900 266716 451274 266744
rect 437900 266704 437906 266716
rect 418856 266580 431954 266608
rect 451246 266608 451274 266716
rect 452746 266704 452752 266756
rect 452804 266744 452810 266756
rect 457438 266744 457444 266756
rect 452804 266716 457444 266744
rect 452804 266704 452810 266716
rect 457438 266704 457444 266716
rect 457496 266704 457502 266756
rect 462682 266704 462688 266756
rect 462740 266744 462746 266756
rect 464632 266744 464660 266852
rect 469950 266840 469956 266852
rect 470008 266840 470014 266892
rect 470134 266840 470140 266892
rect 470192 266880 470198 266892
rect 470566 266880 470594 266988
rect 530670 266976 530676 266988
rect 530728 266976 530734 267028
rect 537202 266976 537208 267028
rect 537260 267016 537266 267028
rect 636194 267016 636200 267028
rect 537260 266988 636200 267016
rect 537260 266976 537266 266988
rect 636194 266976 636200 266988
rect 636252 266976 636258 267028
rect 470192 266852 470594 266880
rect 470192 266840 470198 266852
rect 473446 266840 473452 266892
rect 473504 266880 473510 266892
rect 474366 266880 474372 266892
rect 473504 266852 474372 266880
rect 473504 266840 473510 266852
rect 474366 266840 474372 266852
rect 474424 266840 474430 266892
rect 475102 266840 475108 266892
rect 475160 266880 475166 266892
rect 475930 266880 475936 266892
rect 475160 266852 475936 266880
rect 475160 266840 475166 266852
rect 475930 266840 475936 266852
rect 475988 266840 475994 266892
rect 513742 266880 513748 266892
rect 480226 266852 513748 266880
rect 462740 266716 464660 266744
rect 462740 266704 462746 266716
rect 465166 266704 465172 266756
rect 465224 266744 465230 266756
rect 480226 266744 480254 266852
rect 513742 266840 513748 266852
rect 513800 266840 513806 266892
rect 514018 266840 514024 266892
rect 514076 266880 514082 266892
rect 518710 266880 518716 266892
rect 514076 266852 518716 266880
rect 514076 266840 514082 266852
rect 518710 266840 518716 266852
rect 518768 266840 518774 266892
rect 518894 266840 518900 266892
rect 518952 266880 518958 266892
rect 526438 266880 526444 266892
rect 518952 266852 526444 266880
rect 518952 266840 518958 266852
rect 526438 266840 526444 266852
rect 526496 266840 526502 266892
rect 526622 266840 526628 266892
rect 526680 266880 526686 266892
rect 615494 266880 615500 266892
rect 526680 266852 615500 266880
rect 526680 266840 526686 266852
rect 615494 266840 615500 266852
rect 615552 266840 615558 266892
rect 465224 266716 480254 266744
rect 465224 266704 465230 266716
rect 483198 266704 483204 266756
rect 483256 266744 483262 266756
rect 487154 266744 487160 266756
rect 483256 266716 487160 266744
rect 483256 266704 483262 266716
rect 487154 266704 487160 266716
rect 487212 266704 487218 266756
rect 487522 266704 487528 266756
rect 487580 266744 487586 266756
rect 494698 266744 494704 266756
rect 487580 266716 494704 266744
rect 487580 266704 487586 266716
rect 494698 266704 494704 266716
rect 494756 266704 494762 266756
rect 497458 266744 497464 266756
rect 494900 266716 497464 266744
rect 467282 266608 467288 266620
rect 451246 266580 467288 266608
rect 418856 266568 418862 266580
rect 467282 266568 467288 266580
rect 467340 266568 467346 266620
rect 467558 266568 467564 266620
rect 467616 266608 467622 266620
rect 493134 266608 493140 266620
rect 467616 266580 493140 266608
rect 467616 266568 467622 266580
rect 493134 266568 493140 266580
rect 493192 266568 493198 266620
rect 494900 266608 494928 266716
rect 497458 266704 497464 266716
rect 497516 266704 497522 266756
rect 499942 266704 499948 266756
rect 500000 266744 500006 266756
rect 500862 266744 500868 266756
rect 500000 266716 500868 266744
rect 500000 266704 500006 266716
rect 500862 266704 500868 266716
rect 500920 266704 500926 266756
rect 504082 266704 504088 266756
rect 504140 266744 504146 266756
rect 504910 266744 504916 266756
rect 504140 266716 504916 266744
rect 504140 266704 504146 266716
rect 504910 266704 504916 266716
rect 504968 266704 504974 266756
rect 506566 266704 506572 266756
rect 506624 266744 506630 266756
rect 507762 266744 507768 266756
rect 506624 266716 507768 266744
rect 506624 266704 506630 266716
rect 507762 266704 507768 266716
rect 507820 266704 507826 266756
rect 508406 266704 508412 266756
rect 508464 266744 508470 266756
rect 559558 266744 559564 266756
rect 508464 266716 559564 266744
rect 508464 266704 508470 266716
rect 559558 266704 559564 266716
rect 559616 266704 559622 266756
rect 493336 266580 494928 266608
rect 258258 266500 258264 266552
rect 258316 266540 258322 266552
rect 267274 266540 267280 266552
rect 258316 266512 267280 266540
rect 258316 266500 258322 266512
rect 267274 266500 267280 266512
rect 267332 266500 267338 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 330202 266500 330208 266552
rect 330260 266540 330266 266552
rect 334618 266540 334624 266552
rect 330260 266512 334624 266540
rect 330260 266500 330266 266512
rect 334618 266500 334624 266512
rect 334676 266500 334682 266552
rect 395614 266500 395620 266552
rect 395672 266540 395678 266552
rect 404998 266540 405004 266552
rect 395672 266512 402974 266540
rect 395672 266500 395678 266512
rect 313642 266432 313648 266484
rect 313700 266472 313706 266484
rect 317414 266472 317420 266484
rect 313700 266444 317420 266472
rect 313700 266432 313706 266444
rect 317414 266432 317420 266444
rect 317472 266432 317478 266484
rect 184256 266376 190454 266404
rect 184256 266364 184262 266376
rect 200390 266364 200396 266416
rect 200448 266404 200454 266416
rect 202690 266404 202696 266416
rect 200448 266376 202696 266404
rect 200448 266364 200454 266376
rect 202690 266364 202696 266376
rect 202748 266364 202754 266416
rect 213178 266364 213184 266416
rect 213236 266404 213242 266416
rect 215938 266404 215944 266416
rect 213236 266376 215944 266404
rect 213236 266364 213242 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 222838 266364 222844 266416
rect 222896 266404 222902 266416
rect 224218 266404 224224 266416
rect 222896 266376 224224 266404
rect 222896 266364 222902 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 239490 266364 239496 266416
rect 239548 266404 239554 266416
rect 244090 266404 244096 266416
rect 239548 266376 244096 266404
rect 239548 266364 239554 266376
rect 244090 266364 244096 266376
rect 244148 266364 244154 266416
rect 253750 266364 253756 266416
rect 253808 266404 253814 266416
rect 256510 266404 256516 266416
rect 253808 266376 256516 266404
rect 253808 266364 253814 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 256694 266364 256700 266416
rect 256752 266404 256758 266416
rect 259822 266404 259828 266416
rect 256752 266376 259828 266404
rect 256752 266364 256758 266376
rect 259822 266364 259828 266376
rect 259880 266364 259886 266416
rect 269758 266364 269764 266416
rect 269816 266404 269822 266416
rect 272242 266404 272248 266416
rect 269816 266376 272248 266404
rect 269816 266364 269822 266376
rect 272242 266364 272248 266376
rect 272300 266364 272306 266416
rect 272886 266364 272892 266416
rect 272944 266404 272950 266416
rect 277210 266404 277216 266416
rect 272944 266376 277216 266404
rect 272944 266364 272950 266376
rect 277210 266364 277216 266376
rect 277268 266364 277274 266416
rect 277394 266364 277400 266416
rect 277452 266404 277458 266416
rect 282178 266404 282184 266416
rect 277452 266376 282184 266404
rect 277452 266364 277458 266376
rect 282178 266364 282184 266376
rect 282236 266364 282242 266416
rect 293954 266364 293960 266416
rect 294012 266404 294018 266416
rect 296254 266404 296260 266416
rect 294012 266376 296260 266404
rect 294012 266364 294018 266376
rect 296254 266364 296260 266376
rect 296312 266364 296318 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 324958 266404 324964 266416
rect 320324 266376 324964 266404
rect 320324 266364 320330 266376
rect 324958 266364 324964 266376
rect 325016 266364 325022 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333790 266404 333796 266416
rect 332744 266376 333796 266404
rect 332744 266364 332750 266376
rect 333790 266364 333796 266376
rect 333848 266364 333854 266416
rect 342622 266364 342628 266416
rect 342680 266404 342686 266416
rect 343542 266404 343548 266416
rect 342680 266376 343548 266404
rect 342680 266364 342686 266376
rect 343542 266364 343548 266376
rect 343600 266364 343606 266416
rect 345106 266364 345112 266416
rect 345164 266404 345170 266416
rect 349890 266404 349896 266416
rect 345164 266376 349896 266404
rect 345164 266364 345170 266376
rect 349890 266364 349896 266376
rect 349948 266364 349954 266416
rect 355042 266364 355048 266416
rect 355100 266404 355106 266416
rect 356698 266404 356704 266416
rect 355100 266376 356704 266404
rect 355100 266364 355106 266376
rect 356698 266364 356704 266376
rect 356756 266364 356762 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362862 266404 362868 266416
rect 361724 266376 362868 266404
rect 361724 266364 361730 266376
rect 362862 266364 362868 266376
rect 362920 266364 362926 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368290 266404 368296 266416
rect 367520 266376 368296 266404
rect 367520 266364 367526 266376
rect 368290 266364 368296 266376
rect 368348 266364 368354 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 380802 266404 380808 266416
rect 379940 266376 380808 266404
rect 379940 266364 379946 266376
rect 380802 266364 380808 266376
rect 380860 266364 380866 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387518 266404 387524 266416
rect 386564 266376 387524 266404
rect 386564 266364 386570 266376
rect 387518 266364 387524 266376
rect 387576 266364 387582 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 402946 266404 402974 266512
rect 403084 266512 405004 266540
rect 403084 266404 403112 266512
rect 404998 266500 405004 266512
rect 405056 266500 405062 266552
rect 441982 266500 441988 266552
rect 442040 266540 442046 266552
rect 445018 266540 445024 266552
rect 442040 266512 445024 266540
rect 442040 266500 442046 266512
rect 445018 266500 445024 266512
rect 445076 266500 445082 266552
rect 421282 266432 421288 266484
rect 421340 266472 421346 266484
rect 483198 266472 483204 266484
rect 421340 266444 431954 266472
rect 421340 266432 421346 266444
rect 402946 266376 403112 266404
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 419810 266404 419816 266416
rect 415544 266376 419816 266404
rect 415544 266364 415550 266376
rect 419810 266364 419816 266376
rect 419868 266364 419874 266416
rect 161992 266308 162348 266336
rect 161992 266296 161998 266308
rect 431926 266268 431954 266444
rect 470566 266444 483204 266472
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 439314 266404 439320 266416
rect 433352 266376 439320 266404
rect 433352 266268 433380 266376
rect 439314 266364 439320 266376
rect 439372 266364 439378 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 446122 266364 446128 266416
rect 446180 266404 446186 266416
rect 447778 266404 447784 266416
rect 446180 266376 447784 266404
rect 446180 266364 446186 266376
rect 447778 266364 447784 266376
rect 447836 266364 447842 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 457990 266404 457996 266416
rect 456944 266376 457996 266404
rect 456944 266364 456950 266376
rect 457990 266364 457996 266376
rect 458048 266364 458054 266416
rect 466822 266364 466828 266416
rect 466880 266404 466886 266416
rect 467742 266404 467748 266416
rect 466880 266376 467748 266404
rect 466880 266364 466886 266376
rect 467742 266364 467748 266376
rect 467800 266364 467806 266416
rect 469306 266364 469312 266416
rect 469364 266404 469370 266416
rect 470410 266404 470416 266416
rect 469364 266376 470416 266404
rect 469364 266364 469370 266376
rect 470410 266364 470416 266376
rect 470468 266364 470474 266416
rect 431926 266240 433380 266268
rect 469950 266228 469956 266280
rect 470008 266268 470014 266280
rect 470566 266268 470594 266444
rect 483198 266432 483204 266444
rect 483256 266432 483262 266484
rect 483382 266432 483388 266484
rect 483440 266472 483446 266484
rect 484302 266472 484308 266484
rect 483440 266444 484308 266472
rect 483440 266432 483446 266444
rect 484302 266432 484308 266444
rect 484360 266432 484366 266484
rect 485866 266432 485872 266484
rect 485924 266472 485930 266484
rect 486970 266472 486976 266484
rect 485924 266444 486976 266472
rect 485924 266432 485930 266444
rect 486970 266432 486976 266444
rect 487028 266432 487034 266484
rect 490006 266432 490012 266484
rect 490064 266472 490070 266484
rect 493336 266472 493364 266580
rect 495158 266568 495164 266620
rect 495216 266608 495222 266620
rect 495216 266580 495572 266608
rect 495216 266568 495222 266580
rect 490064 266444 493364 266472
rect 490064 266432 490070 266444
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495342 266472 495348 266484
rect 494204 266444 495348 266472
rect 494204 266432 494210 266444
rect 495342 266432 495348 266444
rect 495400 266432 495406 266484
rect 495544 266472 495572 266580
rect 497458 266568 497464 266620
rect 497516 266608 497522 266620
rect 552658 266608 552664 266620
rect 497516 266580 552664 266608
rect 497516 266568 497522 266580
rect 552658 266568 552664 266580
rect 552716 266568 552722 266620
rect 514018 266472 514024 266484
rect 495544 266444 514024 266472
rect 514018 266432 514024 266444
rect 514076 266432 514082 266484
rect 514846 266432 514852 266484
rect 514904 266472 514910 266484
rect 516042 266472 516048 266484
rect 514904 266444 516048 266472
rect 514904 266432 514910 266444
rect 516042 266432 516048 266444
rect 516100 266432 516106 266484
rect 516502 266432 516508 266484
rect 516560 266472 516566 266484
rect 517330 266472 517336 266484
rect 516560 266444 517336 266472
rect 516560 266432 516566 266444
rect 517330 266432 517336 266444
rect 517388 266432 517394 266484
rect 518986 266432 518992 266484
rect 519044 266472 519050 266484
rect 520090 266472 520096 266484
rect 519044 266444 520096 266472
rect 519044 266432 519050 266444
rect 520090 266432 520096 266444
rect 520148 266432 520154 266484
rect 524782 266432 524788 266484
rect 524840 266472 524846 266484
rect 525702 266472 525708 266484
rect 524840 266444 525708 266472
rect 524840 266432 524846 266444
rect 525702 266432 525708 266444
rect 525760 266432 525766 266484
rect 527266 266432 527272 266484
rect 527324 266472 527330 266484
rect 592678 266472 592684 266484
rect 527324 266444 592684 266472
rect 527324 266432 527330 266444
rect 592678 266432 592684 266444
rect 592736 266432 592742 266484
rect 480070 266296 480076 266348
rect 480128 266336 480134 266348
rect 554774 266336 554780 266348
rect 480128 266308 554780 266336
rect 480128 266296 480134 266308
rect 554774 266296 554780 266308
rect 554832 266296 554838 266348
rect 470008 266240 470594 266268
rect 470008 266228 470014 266240
rect 485038 266160 485044 266212
rect 485096 266200 485102 266212
rect 561674 266200 561680 266212
rect 485096 266172 561680 266200
rect 485096 266160 485102 266172
rect 561674 266160 561680 266172
rect 561732 266160 561738 266212
rect 486694 266024 486700 266076
rect 486752 266064 486758 266076
rect 564434 266064 564440 266076
rect 486752 266036 564440 266064
rect 486752 266024 486758 266036
rect 564434 266024 564440 266036
rect 564492 266024 564498 266076
rect 492490 265888 492496 265940
rect 492548 265928 492554 265940
rect 572714 265928 572720 265940
rect 492548 265900 572720 265928
rect 492548 265888 492554 265900
rect 572714 265888 572720 265900
rect 572772 265888 572778 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 142154 265616 142160 265668
rect 142212 265656 142218 265668
rect 142798 265656 142804 265668
rect 142212 265628 142804 265656
rect 142212 265616 142218 265628
rect 142798 265616 142804 265628
rect 142856 265616 142862 265668
rect 191834 265616 191840 265668
rect 191892 265656 191898 265668
rect 192478 265656 192484 265668
rect 191892 265628 192484 265656
rect 191892 265616 191898 265628
rect 192478 265616 192484 265628
rect 192536 265616 192542 265668
rect 234614 265616 234620 265668
rect 234672 265656 234678 265668
rect 235534 265656 235540 265668
rect 234672 265628 235540 265656
rect 234672 265616 234678 265628
rect 235534 265616 235540 265628
rect 235592 265616 235598 265668
rect 518158 265616 518164 265668
rect 518216 265656 518222 265668
rect 608686 265656 608692 265668
rect 518216 265628 608692 265656
rect 518216 265616 518222 265628
rect 608686 265616 608692 265628
rect 608744 265616 608750 265668
rect 481726 265480 481732 265532
rect 481784 265520 481790 265532
rect 557534 265520 557540 265532
rect 481784 265492 557540 265520
rect 481784 265480 481790 265492
rect 557534 265480 557540 265492
rect 557592 265480 557598 265532
rect 479242 265344 479248 265396
rect 479300 265384 479306 265396
rect 553394 265384 553400 265396
rect 479300 265356 553400 265384
rect 479300 265344 479306 265356
rect 553394 265344 553400 265356
rect 553452 265344 553458 265396
rect 571978 261468 571984 261520
rect 572036 261508 572042 261520
rect 645854 261508 645860 261520
rect 572036 261480 645860 261508
rect 572036 261468 572042 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 563698 259468 563704 259480
rect 554372 259440 563704 259468
rect 554372 259428 554378 259440
rect 563698 259428 563704 259440
rect 563756 259428 563762 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 560938 256748 560944 256760
rect 554004 256720 560944 256748
rect 554004 256708 554010 256720
rect 560938 256708 560944 256720
rect 560996 256708 561002 256760
rect 553762 255280 553768 255332
rect 553820 255320 553826 255332
rect 556798 255320 556804 255332
rect 553820 255292 556804 255320
rect 553820 255280 553826 255292
rect 556798 255280 556804 255292
rect 556856 255280 556862 255332
rect 35802 252832 35808 252884
rect 35860 252872 35866 252884
rect 41322 252872 41328 252884
rect 35860 252844 41328 252872
rect 35860 252832 35866 252844
rect 41322 252832 41328 252844
rect 41380 252832 41386 252884
rect 35618 252696 35624 252748
rect 35676 252736 35682 252748
rect 41690 252736 41696 252748
rect 35676 252708 41696 252736
rect 35676 252696 35682 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35802 252560 35808 252612
rect 35860 252600 35866 252612
rect 40678 252600 40684 252612
rect 35860 252572 40684 252600
rect 35860 252560 35866 252572
rect 40678 252560 40684 252572
rect 40736 252560 40742 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 676030 252356 676036 252408
rect 676088 252396 676094 252408
rect 679618 252396 679624 252408
rect 676088 252368 679624 252396
rect 676088 252356 676094 252368
rect 679618 252356 679624 252368
rect 679676 252356 679682 252408
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 37918 251240 37924 251252
rect 35860 251212 37924 251240
rect 35860 251200 35866 251212
rect 37918 251200 37924 251212
rect 37976 251200 37982 251252
rect 553486 251200 553492 251252
rect 553544 251240 553550 251252
rect 555418 251240 555424 251252
rect 553544 251212 555424 251240
rect 553544 251200 553550 251212
rect 555418 251200 555424 251212
rect 555476 251200 555482 251252
rect 558178 246304 558184 246356
rect 558236 246344 558242 246356
rect 647234 246344 647240 246356
rect 558236 246316 647240 246344
rect 558236 246304 558242 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 606478 245664 606484 245676
rect 553912 245636 606484 245664
rect 553912 245624 553918 245636
rect 606478 245624 606484 245636
rect 606536 245624 606542 245676
rect 554498 244536 554504 244588
rect 554556 244576 554562 244588
rect 559558 244576 559564 244588
rect 554556 244548 559564 244576
rect 554556 244536 554562 244548
rect 559558 244536 559564 244548
rect 559616 244536 559622 244588
rect 37918 242836 37924 242888
rect 37976 242876 37982 242888
rect 41690 242876 41696 242888
rect 37976 242848 41696 242876
rect 37976 242836 37982 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 628558 241516 628564 241528
rect 553728 241488 628564 241516
rect 553728 241476 553734 241488
rect 628558 241476 628564 241488
rect 628616 241476 628622 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 671706 237804 671712 237856
rect 671764 237844 671770 237856
rect 672756 237844 672784 238102
rect 671764 237816 672784 237844
rect 671764 237804 671770 237816
rect 671890 237600 671896 237652
rect 671948 237640 671954 237652
rect 672874 237640 672902 237898
rect 671948 237612 672902 237640
rect 671948 237600 671954 237612
rect 672074 237396 672080 237448
rect 672132 237436 672138 237448
rect 672966 237436 672994 237694
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 672132 237408 672994 237436
rect 672132 237396 672138 237408
rect 671522 237260 671528 237312
rect 671580 237300 671586 237312
rect 671580 237272 673210 237300
rect 671580 237260 671586 237272
rect 672718 237124 672724 237176
rect 672776 237164 672782 237176
rect 672776 237136 673330 237164
rect 672776 237124 672782 237136
rect 673528 236904 673580 236910
rect 668946 236852 668952 236904
rect 669004 236892 669010 236904
rect 669004 236864 673440 236892
rect 669004 236852 669010 236864
rect 673528 236846 673580 236852
rect 673644 236496 673696 236502
rect 673644 236438 673696 236444
rect 673752 236360 673804 236366
rect 673752 236302 673804 236308
rect 673748 236116 673900 236144
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 671338 236036 671344 236088
rect 671396 236076 671402 236088
rect 673748 236076 673776 236116
rect 671396 236048 673776 236076
rect 671396 236036 671402 236048
rect 668670 235900 668676 235952
rect 668728 235940 668734 235952
rect 672074 235940 672080 235952
rect 668728 235912 672080 235940
rect 668728 235900 668734 235912
rect 672074 235900 672080 235912
rect 672132 235900 672138 235952
rect 672276 235912 673992 235940
rect 671154 235764 671160 235816
rect 671212 235804 671218 235816
rect 672276 235804 672304 235912
rect 671212 235776 672304 235804
rect 671212 235764 671218 235776
rect 672738 235220 672744 235272
rect 672796 235260 672802 235272
rect 674100 235260 674128 235654
rect 674190 235424 674196 235476
rect 674248 235424 674254 235476
rect 672796 235232 674128 235260
rect 672796 235220 672802 235232
rect 674324 234784 674352 235314
rect 674426 235136 674478 235142
rect 674426 235078 674478 235084
rect 673426 234756 674352 234784
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 571978 234580 571984 234592
rect 554464 234552 571984 234580
rect 554464 234540 554470 234552
rect 571978 234540 571984 234552
rect 572036 234540 572042 234592
rect 668302 234540 668308 234592
rect 668360 234580 668366 234592
rect 673426 234580 673454 234756
rect 674282 234608 674288 234660
rect 674340 234648 674346 234660
rect 674548 234648 674576 234906
rect 674340 234620 674576 234648
rect 674340 234608 674346 234620
rect 668360 234552 673454 234580
rect 668360 234540 668366 234552
rect 669774 234336 669780 234388
rect 669832 234376 669838 234388
rect 674668 234376 674696 234702
rect 669832 234348 674696 234376
rect 669832 234336 669838 234348
rect 674374 234200 674380 234252
rect 674432 234240 674438 234252
rect 674760 234240 674788 234498
rect 675846 234472 675852 234524
rect 675904 234512 675910 234524
rect 679802 234512 679808 234524
rect 675904 234484 679808 234512
rect 675904 234472 675910 234484
rect 679802 234472 679808 234484
rect 679860 234472 679866 234524
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674432 234212 674788 234240
rect 674432 234200 674438 234212
rect 674530 234104 674536 234116
rect 674408 234076 674536 234104
rect 672374 233996 672380 234048
rect 672432 234036 672438 234048
rect 674408 234036 674436 234076
rect 674530 234064 674536 234076
rect 674588 234064 674594 234116
rect 672432 234008 674436 234036
rect 672432 233996 672438 234008
rect 674990 233912 675018 234090
rect 675846 234064 675852 234116
rect 675904 234104 675910 234116
rect 679618 234104 679624 234116
rect 675904 234076 679624 234104
rect 675904 234064 675910 234076
rect 679618 234064 679624 234076
rect 679676 234064 679682 234116
rect 674972 233860 674978 233912
rect 675030 233860 675036 233912
rect 675108 233776 675136 233886
rect 675846 233792 675852 233844
rect 675904 233832 675910 233844
rect 677870 233832 677876 233844
rect 675904 233804 677876 233832
rect 675904 233792 675910 233804
rect 677870 233792 677876 233804
rect 677928 233792 677934 233844
rect 675108 233736 675116 233776
rect 675110 233724 675116 233736
rect 675168 233724 675174 233776
rect 674530 233588 674536 233640
rect 674588 233628 674594 233640
rect 675248 233628 675276 233682
rect 674588 233600 675276 233628
rect 674588 233588 674594 233600
rect 672902 233452 672908 233504
rect 672960 233492 672966 233504
rect 672960 233464 675018 233492
rect 672960 233452 672966 233464
rect 674990 233424 675018 233464
rect 675202 233424 675208 233436
rect 674990 233396 675208 233424
rect 675202 233384 675208 233396
rect 675260 233384 675266 233436
rect 670970 233316 670976 233368
rect 671028 233356 671034 233368
rect 671028 233328 673204 233356
rect 671028 233316 671034 233328
rect 673176 233288 673204 233328
rect 675358 233288 675386 233478
rect 673176 233260 675386 233288
rect 675846 233248 675852 233300
rect 675904 233288 675910 233300
rect 683390 233288 683396 233300
rect 675904 233260 683396 233288
rect 675904 233248 675910 233260
rect 683390 233248 683396 233260
rect 683448 233248 683454 233300
rect 671706 233180 671712 233232
rect 671764 233220 671770 233232
rect 672994 233220 673000 233232
rect 671764 233192 673000 233220
rect 671764 233180 671770 233192
rect 672994 233180 673000 233192
rect 673052 233180 673058 233232
rect 671154 232976 671160 233028
rect 671212 233016 671218 233028
rect 674834 233016 674840 233028
rect 671212 232988 674840 233016
rect 671212 232976 671218 232988
rect 674834 232976 674840 232988
rect 674892 232976 674898 233028
rect 670234 232840 670240 232892
rect 670292 232880 670298 232892
rect 674190 232880 674196 232892
rect 670292 232852 674196 232880
rect 670292 232840 670298 232852
rect 674190 232840 674196 232852
rect 674248 232840 674254 232892
rect 661862 232568 661868 232620
rect 661920 232608 661926 232620
rect 675478 232608 675484 232620
rect 661920 232580 675484 232608
rect 661920 232568 661926 232580
rect 675478 232568 675484 232580
rect 675536 232568 675542 232620
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 683666 232540 683672 232552
rect 675904 232512 683672 232540
rect 675904 232500 675910 232512
rect 683666 232500 683672 232512
rect 683724 232500 683730 232552
rect 664990 232160 664996 232212
rect 665048 232200 665054 232212
rect 665048 232172 675556 232200
rect 665048 232160 665054 232172
rect 673822 231956 673828 232008
rect 673880 231996 673886 232008
rect 673880 231968 675372 231996
rect 673880 231956 673886 231968
rect 674834 231752 674840 231804
rect 674892 231792 674898 231804
rect 674892 231764 675206 231792
rect 674892 231752 674898 231764
rect 675070 231532 675122 231538
rect 675846 231480 675852 231532
rect 675904 231520 675910 231532
rect 677594 231520 677600 231532
rect 675904 231492 677600 231520
rect 675904 231480 675910 231492
rect 677594 231480 677600 231492
rect 677652 231480 677658 231532
rect 675070 231474 675122 231480
rect 668118 231412 668124 231464
rect 668176 231452 668182 231464
rect 674512 231452 674518 231464
rect 668176 231424 674518 231452
rect 668176 231412 668182 231424
rect 674512 231412 674518 231424
rect 674570 231412 674576 231464
rect 674956 231328 675008 231334
rect 674956 231270 675008 231276
rect 674650 231140 674656 231192
rect 674708 231180 674714 231192
rect 674708 231152 674866 231180
rect 674708 231140 674714 231152
rect 662322 231072 662328 231124
rect 662380 231112 662386 231124
rect 673822 231112 673828 231124
rect 662380 231084 673828 231112
rect 662380 231072 662386 231084
rect 673822 231072 673828 231084
rect 673880 231072 673886 231124
rect 675846 231072 675852 231124
rect 675904 231112 675910 231124
rect 678422 231112 678428 231124
rect 675904 231084 678428 231112
rect 675904 231072 675910 231084
rect 678422 231072 678428 231084
rect 678480 231072 678486 231124
rect 674732 231056 674784 231062
rect 674732 230998 674784 231004
rect 674374 230976 674380 230988
rect 673518 230948 674380 230976
rect 124122 230732 124128 230784
rect 124180 230772 124186 230784
rect 194594 230772 194600 230784
rect 124180 230744 194600 230772
rect 124180 230732 124186 230744
rect 194594 230732 194600 230744
rect 194652 230732 194658 230784
rect 97902 230596 97908 230648
rect 97960 230636 97966 230648
rect 173986 230636 173992 230648
rect 97960 230608 173992 230636
rect 97960 230596 97966 230608
rect 173986 230596 173992 230608
rect 174044 230596 174050 230648
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 91002 230460 91008 230512
rect 91060 230500 91066 230512
rect 168834 230500 168840 230512
rect 91060 230472 168840 230500
rect 91060 230460 91066 230472
rect 168834 230460 168840 230472
rect 168892 230460 168898 230512
rect 184106 230392 184112 230444
rect 184164 230432 184170 230444
rect 189442 230432 189448 230444
rect 184164 230404 189448 230432
rect 184164 230392 184170 230404
rect 189442 230392 189448 230404
rect 189500 230392 189506 230444
rect 196066 230392 196072 230444
rect 196124 230432 196130 230444
rect 198458 230432 198464 230444
rect 196124 230404 198464 230432
rect 196124 230392 196130 230404
rect 198458 230392 198464 230404
rect 198516 230392 198522 230444
rect 207658 230392 207664 230444
rect 207716 230432 207722 230444
rect 251266 230432 251272 230444
rect 207716 230404 251272 230432
rect 207716 230392 207722 230404
rect 251266 230392 251272 230404
rect 251324 230392 251330 230444
rect 256602 230392 256608 230444
rect 256660 230432 256666 230444
rect 297634 230432 297640 230444
rect 256660 230404 297640 230432
rect 256660 230392 256666 230404
rect 297634 230392 297640 230404
rect 297692 230392 297698 230444
rect 323578 230392 323584 230444
rect 323636 230432 323642 230444
rect 324682 230432 324688 230444
rect 323636 230404 324688 230432
rect 323636 230392 323642 230404
rect 324682 230392 324688 230404
rect 324740 230392 324746 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443546 230432 443552 230444
rect 441948 230404 443552 230432
rect 441948 230392 441954 230404
rect 443546 230392 443552 230404
rect 443604 230392 443610 230444
rect 444466 230392 444472 230444
rect 444524 230432 444530 230444
rect 447594 230432 447600 230444
rect 444524 230404 447600 230432
rect 444524 230392 444530 230404
rect 447594 230392 447600 230404
rect 447652 230392 447658 230444
rect 468294 230392 468300 230444
rect 468352 230432 468358 230444
rect 469030 230432 469036 230444
rect 468352 230404 469036 230432
rect 468352 230392 468358 230404
rect 469030 230392 469036 230404
rect 469088 230392 469094 230444
rect 472158 230392 472164 230444
rect 472216 230432 472222 230444
rect 473078 230432 473084 230444
rect 472216 230404 473084 230432
rect 472216 230392 472222 230404
rect 473078 230392 473084 230404
rect 473136 230392 473142 230444
rect 542998 230432 543004 230444
rect 532528 230404 543004 230432
rect 376018 230324 376024 230376
rect 376076 230364 376082 230376
rect 380710 230364 380716 230376
rect 376076 230336 380716 230364
rect 376076 230324 376082 230336
rect 380710 230324 380716 230336
rect 380768 230324 380774 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 473446 230324 473452 230376
rect 473504 230364 473510 230376
rect 474550 230364 474556 230376
rect 473504 230336 474556 230364
rect 473504 230324 473510 230336
rect 474550 230324 474556 230336
rect 474608 230324 474614 230376
rect 477310 230324 477316 230376
rect 477368 230364 477374 230376
rect 480070 230364 480076 230376
rect 477368 230336 480076 230364
rect 477368 230324 477374 230336
rect 480070 230324 480076 230336
rect 480128 230324 480134 230376
rect 480530 230324 480536 230376
rect 480588 230364 480594 230376
rect 481542 230364 481548 230376
rect 480588 230336 481548 230364
rect 480588 230324 480594 230336
rect 481542 230324 481548 230336
rect 481600 230324 481606 230376
rect 499850 230324 499856 230376
rect 499908 230364 499914 230376
rect 501598 230364 501604 230376
rect 499908 230336 501604 230364
rect 499908 230324 499914 230336
rect 501598 230324 501604 230336
rect 501656 230324 501662 230376
rect 501782 230324 501788 230376
rect 501840 230364 501846 230376
rect 508498 230364 508504 230376
rect 501840 230336 508504 230364
rect 501840 230324 501846 230336
rect 508498 230324 508504 230336
rect 508556 230324 508562 230376
rect 509510 230324 509516 230376
rect 509568 230364 509574 230376
rect 518158 230364 518164 230376
rect 509568 230336 518164 230364
rect 509568 230324 509574 230336
rect 518158 230324 518164 230336
rect 518216 230324 518222 230376
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521470 230364 521476 230376
rect 520516 230336 521476 230364
rect 520516 230324 520522 230336
rect 521470 230324 521476 230336
rect 521528 230324 521534 230376
rect 530118 230324 530124 230376
rect 530176 230364 530182 230376
rect 531222 230364 531228 230376
rect 530176 230336 531228 230364
rect 530176 230324 530182 230336
rect 531222 230324 531228 230336
rect 531280 230324 531286 230376
rect 133782 230256 133788 230308
rect 133840 230296 133846 230308
rect 202322 230296 202328 230308
rect 133840 230268 202328 230296
rect 133840 230256 133846 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 240962 230296 240968 230308
rect 209746 230268 240968 230296
rect 126882 230120 126888 230172
rect 126940 230160 126946 230172
rect 197170 230160 197176 230172
rect 126940 230132 197176 230160
rect 126940 230120 126946 230132
rect 197170 230120 197176 230132
rect 197228 230120 197234 230172
rect 197446 230120 197452 230172
rect 197504 230160 197510 230172
rect 201034 230160 201040 230172
rect 197504 230132 201040 230160
rect 197504 230120 197510 230132
rect 201034 230120 201040 230132
rect 201092 230120 201098 230172
rect 202138 230120 202144 230172
rect 202196 230160 202202 230172
rect 209746 230160 209774 230268
rect 240962 230256 240968 230268
rect 241020 230256 241026 230308
rect 242526 230256 242532 230308
rect 242584 230296 242590 230308
rect 287330 230296 287336 230308
rect 242584 230268 287336 230296
rect 242584 230256 242590 230268
rect 287330 230256 287336 230268
rect 287388 230256 287394 230308
rect 305638 230256 305644 230308
rect 305696 230296 305702 230308
rect 334986 230296 334992 230308
rect 305696 230268 334992 230296
rect 305696 230256 305702 230268
rect 334986 230256 334992 230268
rect 335044 230256 335050 230308
rect 387334 230188 387340 230240
rect 387392 230228 387398 230240
rect 388438 230228 388444 230240
rect 387392 230200 388444 230228
rect 387392 230188 387398 230200
rect 388438 230188 388444 230200
rect 388496 230188 388502 230240
rect 413830 230188 413836 230240
rect 413888 230228 413894 230240
rect 419994 230228 420000 230240
rect 413888 230200 420000 230228
rect 413888 230188 413894 230200
rect 419994 230188 420000 230200
rect 420052 230188 420058 230240
rect 443822 230188 443828 230240
rect 443880 230228 443886 230240
rect 444650 230228 444656 230240
rect 443880 230200 444656 230228
rect 443880 230188 443886 230200
rect 444650 230188 444656 230200
rect 444708 230188 444714 230240
rect 470870 230188 470876 230240
rect 470928 230228 470934 230240
rect 471882 230228 471888 230240
rect 470928 230200 471888 230228
rect 470928 230188 470934 230200
rect 471882 230188 471888 230200
rect 471940 230188 471946 230240
rect 474090 230188 474096 230240
rect 474148 230228 474154 230240
rect 477402 230228 477408 230240
rect 474148 230200 477408 230228
rect 474148 230188 474154 230200
rect 477402 230188 477408 230200
rect 477460 230188 477466 230240
rect 530762 230188 530768 230240
rect 530820 230228 530826 230240
rect 532528 230228 532556 230404
rect 542998 230392 543004 230404
rect 543056 230392 543062 230444
rect 668854 230392 668860 230444
rect 668912 230432 668918 230444
rect 673518 230432 673546 230948
rect 674374 230936 674380 230948
rect 674432 230936 674438 230988
rect 673638 230800 673644 230852
rect 673696 230840 673702 230852
rect 673696 230812 674636 230840
rect 673696 230800 673702 230812
rect 674374 230636 674380 230648
rect 668912 230404 673546 230432
rect 674208 230608 674380 230636
rect 668912 230392 668918 230404
rect 533522 230256 533528 230308
rect 533580 230296 533586 230308
rect 541250 230296 541256 230308
rect 533580 230268 541256 230296
rect 533580 230256 533586 230268
rect 541250 230256 541256 230268
rect 541308 230256 541314 230308
rect 530820 230200 532556 230228
rect 674208 230228 674236 230608
rect 674374 230596 674380 230608
rect 674432 230596 674438 230648
rect 674518 230512 674570 230518
rect 674518 230454 674570 230460
rect 674396 230308 674448 230314
rect 674396 230250 674448 230256
rect 674208 230200 674314 230228
rect 530820 230188 530826 230200
rect 202196 230132 209774 230160
rect 202196 230120 202202 230132
rect 214374 230120 214380 230172
rect 214432 230160 214438 230172
rect 225506 230160 225512 230172
rect 214432 230132 225512 230160
rect 214432 230120 214438 230132
rect 225506 230120 225512 230132
rect 225564 230120 225570 230172
rect 230474 230120 230480 230172
rect 230532 230160 230538 230172
rect 277026 230160 277032 230172
rect 230532 230132 277032 230160
rect 230532 230120 230538 230132
rect 277026 230120 277032 230132
rect 277084 230120 277090 230172
rect 294598 230120 294604 230172
rect 294656 230160 294662 230172
rect 323394 230160 323400 230172
rect 294656 230132 323400 230160
rect 294656 230120 294662 230132
rect 323394 230120 323400 230132
rect 323452 230120 323458 230172
rect 324958 230120 324964 230172
rect 325016 230160 325022 230172
rect 350442 230160 350448 230172
rect 325016 230132 350448 230160
rect 325016 230120 325022 230132
rect 350442 230120 350448 230132
rect 350500 230120 350506 230172
rect 354858 230120 354864 230172
rect 354916 230160 354922 230172
rect 371050 230160 371056 230172
rect 354916 230132 371056 230160
rect 354916 230120 354922 230132
rect 371050 230120 371056 230132
rect 371108 230120 371114 230172
rect 503714 230120 503720 230172
rect 503772 230160 503778 230172
rect 512638 230160 512644 230172
rect 503772 230132 512644 230160
rect 503772 230120 503778 230132
rect 512638 230120 512644 230132
rect 512696 230120 512702 230172
rect 515306 230120 515312 230172
rect 515364 230160 515370 230172
rect 525150 230160 525156 230172
rect 515364 230132 525156 230160
rect 515364 230120 515370 230132
rect 525150 230120 525156 230132
rect 525208 230120 525214 230172
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 486326 230052 486332 230104
rect 486384 230092 486390 230104
rect 487062 230092 487068 230104
rect 486384 230064 487068 230092
rect 486384 230052 486390 230064
rect 487062 230052 487068 230064
rect 487120 230052 487126 230104
rect 490190 230052 490196 230104
rect 490248 230092 490254 230104
rect 490248 230064 499574 230092
rect 490248 230052 490254 230064
rect 86218 229984 86224 230036
rect 86276 230024 86282 230036
rect 155954 230024 155960 230036
rect 86276 229996 155960 230024
rect 86276 229984 86282 229996
rect 155954 229984 155960 229996
rect 156012 229984 156018 230036
rect 157058 229984 157064 230036
rect 157116 230024 157122 230036
rect 157116 229996 214604 230024
rect 157116 229984 157122 229996
rect 117222 229848 117228 229900
rect 117280 229888 117286 229900
rect 184106 229888 184112 229900
rect 117280 229860 184112 229888
rect 117280 229848 117286 229860
rect 184106 229848 184112 229860
rect 184164 229848 184170 229900
rect 184474 229848 184480 229900
rect 184532 229888 184538 229900
rect 214374 229888 214380 229900
rect 184532 229860 214380 229888
rect 184532 229848 184538 229860
rect 214374 229848 214380 229860
rect 214432 229848 214438 229900
rect 214576 229888 214604 229996
rect 225782 229984 225788 230036
rect 225840 230024 225846 230036
rect 271874 230024 271880 230036
rect 225840 229996 271880 230024
rect 225840 229984 225846 229996
rect 271874 229984 271880 229996
rect 271932 229984 271938 230036
rect 300118 229984 300124 230036
rect 300176 230024 300182 230036
rect 329834 230024 329840 230036
rect 300176 229996 329840 230024
rect 300176 229984 300182 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 337838 229984 337844 230036
rect 337896 230024 337902 230036
rect 360746 230024 360752 230036
rect 337896 229996 360752 230024
rect 337896 229984 337902 229996
rect 360746 229984 360752 229996
rect 360804 229984 360810 230036
rect 465442 229984 465448 230036
rect 465500 230024 465506 230036
rect 473722 230024 473728 230036
rect 465500 229996 473728 230024
rect 465500 229984 465506 229996
rect 473722 229984 473728 229996
rect 473780 229984 473786 230036
rect 484394 229916 484400 229968
rect 484452 229956 484458 229968
rect 496814 229956 496820 229968
rect 484452 229928 496820 229956
rect 484452 229916 484458 229928
rect 496814 229916 496820 229928
rect 496872 229916 496878 229968
rect 220354 229888 220360 229900
rect 214576 229860 220360 229888
rect 220354 229848 220360 229860
rect 220412 229848 220418 229900
rect 224034 229848 224040 229900
rect 224092 229888 224098 229900
rect 266722 229888 266728 229900
rect 224092 229860 266728 229888
rect 224092 229848 224098 229860
rect 266722 229848 266728 229860
rect 266780 229848 266786 229900
rect 283558 229848 283564 229900
rect 283616 229888 283622 229900
rect 318242 229888 318248 229900
rect 283616 229860 318248 229888
rect 283616 229848 283622 229860
rect 318242 229848 318248 229860
rect 318300 229848 318306 229900
rect 318426 229848 318432 229900
rect 318484 229888 318490 229900
rect 345290 229888 345296 229900
rect 318484 229860 345296 229888
rect 318484 229848 318490 229860
rect 345290 229848 345296 229860
rect 345348 229848 345354 229900
rect 361206 229848 361212 229900
rect 361264 229888 361270 229900
rect 378778 229888 378784 229900
rect 361264 229860 378784 229888
rect 361264 229848 361270 229860
rect 378778 229848 378784 229860
rect 378836 229848 378842 229900
rect 389910 229848 389916 229900
rect 389968 229888 389974 229900
rect 399386 229888 399392 229900
rect 389968 229860 399392 229888
rect 389968 229848 389974 229860
rect 399386 229848 399392 229860
rect 399444 229848 399450 229900
rect 410794 229848 410800 229900
rect 410852 229888 410858 229900
rect 417418 229888 417424 229900
rect 410852 229860 417424 229888
rect 410852 229848 410858 229860
rect 417418 229848 417424 229860
rect 417476 229848 417482 229900
rect 499546 229888 499574 230064
rect 505646 229984 505652 230036
rect 505704 230024 505710 230036
rect 505704 229996 510660 230024
rect 505704 229984 505710 229996
rect 505738 229888 505744 229900
rect 499546 229860 505744 229888
rect 505738 229848 505744 229860
rect 505796 229848 505802 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 510632 229820 510660 229996
rect 528830 229984 528836 230036
rect 528888 230024 528894 230036
rect 533522 230024 533528 230036
rect 528888 229996 533528 230024
rect 528888 229984 528894 229996
rect 533522 229984 533528 229996
rect 533580 229984 533586 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 552198 230024 552204 230036
rect 534684 229996 552204 230024
rect 534684 229984 534690 229996
rect 552198 229984 552204 229996
rect 552256 229984 552262 230036
rect 556798 229984 556804 230036
rect 556856 230024 556862 230036
rect 571334 230024 571340 230036
rect 556856 229996 571340 230024
rect 556856 229984 556862 229996
rect 571334 229984 571340 229996
rect 571392 229984 571398 230036
rect 675846 229984 675852 230036
rect 675904 230024 675910 230036
rect 677410 230024 677416 230036
rect 675904 229996 677416 230024
rect 675904 229984 675910 229996
rect 677410 229984 677416 229996
rect 677468 229984 677474 230036
rect 674172 229968 674224 229974
rect 510798 229916 510804 229968
rect 510856 229956 510862 229968
rect 511810 229956 511816 229968
rect 510856 229928 511816 229956
rect 510856 229916 510862 229928
rect 511810 229916 511816 229928
rect 511868 229916 511874 229968
rect 673914 229916 673920 229968
rect 673972 229916 673978 229968
rect 519170 229848 519176 229900
rect 519228 229888 519234 229900
rect 529198 229888 529204 229900
rect 519228 229860 529204 229888
rect 519228 229848 519234 229860
rect 529198 229848 529204 229860
rect 529256 229848 529262 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 556982 229888 556988 229900
rect 536616 229860 556988 229888
rect 536616 229848 536622 229860
rect 556982 229848 556988 229860
rect 557040 229848 557046 229900
rect 515398 229820 515404 229832
rect 510632 229792 515404 229820
rect 515398 229780 515404 229792
rect 515456 229780 515462 229832
rect 673932 229820 673960 229916
rect 674172 229910 674224 229916
rect 675846 229848 675852 229900
rect 675904 229888 675910 229900
rect 676766 229888 676772 229900
rect 675904 229860 676772 229888
rect 675904 229848 675910 229860
rect 676766 229848 676772 229860
rect 676824 229848 676830 229900
rect 673932 229792 674084 229820
rect 110322 229712 110328 229764
rect 110380 229752 110386 229764
rect 184290 229752 184296 229764
rect 110380 229724 184296 229752
rect 110380 229712 110386 229724
rect 184290 229712 184296 229724
rect 184348 229712 184354 229764
rect 185578 229712 185584 229764
rect 185636 229752 185642 229764
rect 207474 229752 207480 229764
rect 185636 229724 207480 229752
rect 185636 229712 185642 229724
rect 207474 229712 207480 229724
rect 207532 229712 207538 229764
rect 210418 229712 210424 229764
rect 210476 229752 210482 229764
rect 261570 229752 261576 229764
rect 210476 229724 261576 229752
rect 210476 229712 210482 229724
rect 261570 229712 261576 229724
rect 261628 229712 261634 229764
rect 270126 229712 270132 229764
rect 270184 229752 270190 229764
rect 307938 229752 307944 229764
rect 270184 229724 307944 229752
rect 270184 229712 270190 229724
rect 307938 229712 307944 229724
rect 307996 229712 308002 229764
rect 340138 229752 340144 229764
rect 316006 229724 340144 229752
rect 95234 229576 95240 229628
rect 95292 229616 95298 229628
rect 161106 229616 161112 229628
rect 95292 229588 161112 229616
rect 95292 229576 95298 229588
rect 161106 229576 161112 229588
rect 161164 229576 161170 229628
rect 161290 229576 161296 229628
rect 161348 229616 161354 229628
rect 175090 229616 175096 229628
rect 161348 229588 175096 229616
rect 161348 229576 161354 229588
rect 175090 229576 175096 229588
rect 175148 229576 175154 229628
rect 175274 229576 175280 229628
rect 175332 229616 175338 229628
rect 217778 229616 217784 229628
rect 175332 229588 217784 229616
rect 175332 229576 175338 229588
rect 217778 229576 217784 229588
rect 217836 229576 217842 229628
rect 251726 229576 251732 229628
rect 251784 229616 251790 229628
rect 292482 229616 292488 229628
rect 251784 229588 292488 229616
rect 251784 229576 251790 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 311894 229576 311900 229628
rect 311952 229616 311958 229628
rect 316006 229616 316034 229724
rect 340138 229712 340144 229724
rect 340196 229712 340202 229764
rect 345658 229712 345664 229764
rect 345716 229752 345722 229764
rect 355594 229752 355600 229764
rect 345716 229724 355600 229752
rect 345716 229712 345722 229724
rect 355594 229712 355600 229724
rect 355652 229712 355658 229764
rect 357066 229712 357072 229764
rect 357124 229752 357130 229764
rect 376202 229752 376208 229764
rect 357124 229724 376208 229752
rect 357124 229712 357130 229724
rect 376202 229712 376208 229724
rect 376260 229712 376266 229764
rect 380710 229712 380716 229764
rect 380768 229752 380774 229764
rect 394234 229752 394240 229764
rect 380768 229724 394240 229752
rect 380768 229712 380774 229724
rect 394234 229712 394240 229724
rect 394292 229712 394298 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 489914 229752 489920 229764
rect 479300 229724 489920 229752
rect 479300 229712 479306 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 494330 229712 494336 229764
rect 494388 229752 494394 229764
rect 509878 229752 509884 229764
rect 494388 229724 509884 229752
rect 494388 229712 494394 229724
rect 509878 229712 509884 229724
rect 509936 229712 509942 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534902 229752 534908 229764
rect 523092 229724 534908 229752
rect 523092 229712 523098 229724
rect 534902 229712 534908 229724
rect 534960 229712 534966 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 565630 229752 565636 229764
rect 538548 229724 565636 229752
rect 538548 229712 538554 229724
rect 565630 229712 565636 229724
rect 565688 229712 565694 229764
rect 311952 229588 316034 229616
rect 311952 229576 311958 229588
rect 526898 229576 526904 229628
rect 526956 229616 526962 229628
rect 534718 229616 534724 229628
rect 526956 229588 534724 229616
rect 526956 229576 526962 229588
rect 534718 229576 534724 229588
rect 534776 229576 534782 229628
rect 673948 229560 674000 229566
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 452194 229548 452200 229560
rect 449032 229520 452200 229548
rect 449032 229508 449038 229520
rect 452194 229508 452200 229520
rect 452252 229508 452258 229560
rect 673948 229502 674000 229508
rect 673828 229492 673880 229498
rect 94498 229440 94504 229492
rect 94556 229480 94562 229492
rect 145650 229480 145656 229492
rect 94556 229452 145656 229480
rect 94556 229440 94562 229452
rect 145650 229440 145656 229452
rect 145708 229440 145714 229492
rect 146202 229440 146208 229492
rect 146260 229480 146266 229492
rect 210050 229480 210056 229492
rect 146260 229452 210056 229480
rect 146260 229440 146266 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 215202 229480 215208 229492
rect 212460 229452 215208 229480
rect 137278 229304 137284 229356
rect 137336 229344 137342 229356
rect 143718 229344 143724 229356
rect 137336 229316 143724 229344
rect 137336 229304 137342 229316
rect 143718 229304 143724 229316
rect 143776 229304 143782 229356
rect 144178 229304 144184 229356
rect 144236 229344 144242 229356
rect 148870 229344 148876 229356
rect 144236 229316 148876 229344
rect 144236 229304 144242 229316
rect 148870 229304 148876 229316
rect 148928 229304 148934 229356
rect 150066 229304 150072 229356
rect 150124 229344 150130 229356
rect 212460 229344 212488 229452
rect 215202 229440 215208 229452
rect 215260 229440 215266 229492
rect 217318 229440 217324 229492
rect 217376 229480 217382 229492
rect 224034 229480 224040 229492
rect 217376 229452 224040 229480
rect 217376 229440 217382 229452
rect 224034 229440 224040 229452
rect 224092 229440 224098 229492
rect 256418 229480 256424 229492
rect 229066 229452 256424 229480
rect 150124 229316 212488 229344
rect 150124 229304 150130 229316
rect 213086 229304 213092 229356
rect 213144 229344 213150 229356
rect 229066 229344 229094 229452
rect 256418 229440 256424 229452
rect 256476 229440 256482 229492
rect 276658 229440 276664 229492
rect 276716 229480 276722 229492
rect 302786 229480 302792 229492
rect 276716 229452 302792 229480
rect 276716 229440 276722 229452
rect 302786 229440 302792 229452
rect 302844 229440 302850 229492
rect 673828 229434 673880 229440
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 453022 229412 453028 229424
rect 450964 229384 453028 229412
rect 450964 229372 450970 229384
rect 453022 229372 453028 229384
rect 453080 229372 453086 229424
rect 453482 229372 453488 229424
rect 453540 229412 453546 229424
rect 455782 229412 455788 229424
rect 453540 229384 455788 229412
rect 453540 229372 453546 229384
rect 455782 229372 455788 229384
rect 455840 229372 455846 229424
rect 213144 229316 229094 229344
rect 213144 229304 213150 229316
rect 261478 229304 261484 229356
rect 261536 229344 261542 229356
rect 282178 229344 282184 229356
rect 261536 229316 282184 229344
rect 261536 229304 261542 229316
rect 282178 229304 282184 229316
rect 282236 229304 282242 229356
rect 288710 229304 288716 229356
rect 288768 229344 288774 229356
rect 313090 229344 313096 229356
rect 288768 229316 313096 229344
rect 288768 229304 288774 229316
rect 313090 229304 313096 229316
rect 313148 229304 313154 229356
rect 517422 229304 517428 229356
rect 517480 229344 517486 229356
rect 520274 229344 520280 229356
rect 517480 229316 520280 229344
rect 517480 229304 517486 229316
rect 520274 229304 520280 229316
rect 520332 229304 520338 229356
rect 448330 229236 448336 229288
rect 448388 229276 448394 229288
rect 449802 229276 449808 229288
rect 448388 229248 449808 229276
rect 448388 229236 448394 229248
rect 449802 229236 449808 229248
rect 449860 229236 449866 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 452838 229236 452844 229288
rect 452896 229276 452902 229288
rect 454678 229276 454684 229288
rect 452896 229248 454684 229276
rect 452896 229236 452902 229248
rect 454678 229236 454684 229248
rect 454736 229236 454742 229288
rect 497918 229236 497924 229288
rect 497976 229276 497982 229288
rect 500218 229276 500224 229288
rect 497976 229248 500224 229276
rect 497976 229236 497982 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 521102 229236 521108 229288
rect 521160 229276 521166 229288
rect 526438 229276 526444 229288
rect 521160 229248 526444 229276
rect 521160 229236 521166 229248
rect 526438 229236 526444 229248
rect 526496 229236 526502 229288
rect 106918 229168 106924 229220
rect 106976 229208 106982 229220
rect 166258 229208 166264 229220
rect 106976 229180 166264 229208
rect 106976 229168 106982 229180
rect 166258 229168 166264 229180
rect 166316 229168 166322 229220
rect 167638 229168 167644 229220
rect 167696 229208 167702 229220
rect 174906 229208 174912 229220
rect 167696 229180 174912 229208
rect 167696 229168 167702 229180
rect 174906 229168 174912 229180
rect 174964 229168 174970 229220
rect 175090 229168 175096 229220
rect 175148 229208 175154 229220
rect 185578 229208 185584 229220
rect 175148 229180 185584 229208
rect 175148 229168 175154 229180
rect 185578 229168 185584 229180
rect 185636 229168 185642 229220
rect 189718 229168 189724 229220
rect 189776 229208 189782 229220
rect 235810 229208 235816 229220
rect 189776 229180 235816 229208
rect 189776 229168 189782 229180
rect 235810 229168 235816 229180
rect 235868 229168 235874 229220
rect 513374 229168 513380 229220
rect 513432 229208 513438 229220
rect 519538 229208 519544 229220
rect 513432 229180 519544 229208
rect 513432 229168 513438 229180
rect 519538 229168 519544 229180
rect 519596 229168 519602 229220
rect 673736 229152 673788 229158
rect 419626 229100 419632 229152
rect 419684 229140 419690 229152
rect 421926 229140 421932 229152
rect 419684 229112 421932 229140
rect 419684 229100 419690 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 446398 229100 446404 229152
rect 446456 229140 446462 229152
rect 448514 229140 448520 229152
rect 446456 229112 448520 229140
rect 446456 229100 446462 229112
rect 448514 229100 448520 229112
rect 448572 229100 448578 229152
rect 449618 229100 449624 229152
rect 449676 229140 449682 229152
rect 450722 229140 450728 229152
rect 449676 229112 450728 229140
rect 449676 229100 449682 229112
rect 450722 229100 450728 229112
rect 450780 229100 450786 229152
rect 451550 229100 451556 229152
rect 451608 229140 451614 229152
rect 453298 229140 453304 229152
rect 451608 229112 453304 229140
rect 451608 229100 451614 229112
rect 453298 229100 453304 229112
rect 453356 229100 453362 229152
rect 454126 229100 454132 229152
rect 454184 229140 454190 229152
rect 455322 229140 455328 229152
rect 454184 229112 455328 229140
rect 454184 229100 454190 229112
rect 455322 229100 455328 229112
rect 455380 229100 455386 229152
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 673454 229140 673460 229152
rect 672644 229112 673460 229140
rect 119982 229032 119988 229084
rect 120040 229072 120046 229084
rect 190086 229072 190092 229084
rect 120040 229044 190092 229072
rect 120040 229032 120046 229044
rect 190086 229032 190092 229044
rect 190144 229032 190150 229084
rect 193122 229032 193128 229084
rect 193180 229072 193186 229084
rect 246758 229072 246764 229084
rect 193180 229044 246764 229072
rect 193180 229032 193186 229044
rect 246758 229032 246764 229044
rect 246816 229032 246822 229084
rect 257706 229032 257712 229084
rect 257764 229072 257770 229084
rect 299566 229072 299572 229084
rect 257764 229044 299572 229072
rect 257764 229032 257770 229044
rect 299566 229032 299572 229044
rect 299624 229032 299630 229084
rect 308766 229032 308772 229084
rect 308824 229072 308830 229084
rect 336274 229072 336280 229084
rect 308824 229044 336280 229072
rect 308824 229032 308830 229044
rect 336274 229032 336280 229044
rect 336332 229032 336338 229084
rect 523310 229072 523316 229084
rect 509206 229044 523316 229072
rect 508222 228964 508228 229016
rect 508280 229004 508286 229016
rect 509206 229004 509234 229044
rect 523310 229032 523316 229044
rect 523368 229032 523374 229084
rect 508280 228976 509234 229004
rect 508280 228964 508286 228976
rect 100662 228896 100668 228948
rect 100720 228936 100726 228948
rect 174630 228936 174636 228948
rect 100720 228908 174636 228936
rect 100720 228896 100726 228908
rect 174630 228896 174636 228908
rect 174688 228896 174694 228948
rect 176378 228896 176384 228948
rect 176436 228936 176442 228948
rect 233878 228936 233884 228948
rect 176436 228908 233884 228936
rect 176436 228896 176442 228908
rect 233878 228896 233884 228908
rect 233936 228896 233942 228948
rect 234522 228896 234528 228948
rect 234580 228936 234586 228948
rect 278314 228936 278320 228948
rect 234580 228908 278320 228936
rect 234580 228896 234586 228908
rect 278314 228896 278320 228908
rect 278372 228896 278378 228948
rect 288066 228896 288072 228948
rect 288124 228936 288130 228948
rect 322750 228936 322756 228948
rect 288124 228908 322756 228936
rect 288124 228896 288130 228908
rect 322750 228896 322756 228908
rect 322808 228896 322814 228948
rect 327718 228896 327724 228948
rect 327776 228936 327782 228948
rect 337562 228936 337568 228948
rect 327776 228908 337568 228936
rect 327776 228896 327782 228908
rect 337562 228896 337568 228908
rect 337620 228896 337626 228948
rect 350166 228896 350172 228948
rect 350224 228936 350230 228948
rect 369118 228936 369124 228948
rect 350224 228908 369124 228936
rect 350224 228896 350230 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 517882 228896 517888 228948
rect 517940 228936 517946 228948
rect 540790 228936 540796 228948
rect 517940 228908 540796 228936
rect 517940 228896 517946 228908
rect 540790 228896 540796 228908
rect 540848 228896 540854 228948
rect 106182 228760 106188 228812
rect 106240 228800 106246 228812
rect 179782 228800 179788 228812
rect 106240 228772 179788 228800
rect 106240 228760 106246 228772
rect 179782 228760 179788 228772
rect 179840 228760 179846 228812
rect 183462 228760 183468 228812
rect 183520 228800 183526 228812
rect 239030 228800 239036 228812
rect 183520 228772 239036 228800
rect 183520 228760 183526 228772
rect 239030 228760 239036 228772
rect 239088 228760 239094 228812
rect 246298 228760 246304 228812
rect 246356 228800 246362 228812
rect 289262 228800 289268 228812
rect 246356 228772 289268 228800
rect 246356 228760 246362 228772
rect 289262 228760 289268 228772
rect 289320 228760 289326 228812
rect 304902 228760 304908 228812
rect 304960 228800 304966 228812
rect 333698 228800 333704 228812
rect 304960 228772 333704 228800
rect 304960 228760 304966 228772
rect 333698 228760 333704 228772
rect 333756 228760 333762 228812
rect 335262 228760 335268 228812
rect 335320 228800 335326 228812
rect 356882 228800 356888 228812
rect 335320 228772 356888 228800
rect 335320 228760 335326 228772
rect 356882 228760 356888 228772
rect 356940 228760 356946 228812
rect 373810 228760 373816 228812
rect 373868 228800 373874 228812
rect 387150 228800 387156 228812
rect 373868 228772 387156 228800
rect 373868 228760 373874 228772
rect 387150 228760 387156 228772
rect 387208 228760 387214 228812
rect 485038 228760 485044 228812
rect 485096 228800 485102 228812
rect 498746 228800 498752 228812
rect 485096 228772 498752 228800
rect 485096 228760 485102 228772
rect 498746 228760 498752 228772
rect 498804 228760 498810 228812
rect 526254 228760 526260 228812
rect 526312 228800 526318 228812
rect 550634 228800 550640 228812
rect 526312 228772 550640 228800
rect 526312 228760 526318 228772
rect 550634 228760 550640 228772
rect 550692 228760 550698 228812
rect 93762 228624 93768 228676
rect 93820 228664 93826 228676
rect 169478 228664 169484 228676
rect 93820 228636 169484 228664
rect 93820 228624 93826 228636
rect 169478 228624 169484 228636
rect 169536 228624 169542 228676
rect 169938 228624 169944 228676
rect 169996 228664 170002 228676
rect 228726 228664 228732 228676
rect 169996 228636 228732 228664
rect 169996 228624 170002 228636
rect 228726 228624 228732 228636
rect 228784 228624 228790 228676
rect 235810 228624 235816 228676
rect 235868 228664 235874 228676
rect 280246 228664 280252 228676
rect 235868 228636 280252 228664
rect 235868 228624 235874 228636
rect 280246 228624 280252 228636
rect 280304 228624 280310 228676
rect 285582 228624 285588 228676
rect 285640 228664 285646 228676
rect 318886 228664 318892 228676
rect 285640 228636 318892 228664
rect 285640 228624 285646 228636
rect 318886 228624 318892 228636
rect 318944 228624 318950 228676
rect 336550 228624 336556 228676
rect 336608 228664 336614 228676
rect 358814 228664 358820 228676
rect 336608 228636 358820 228664
rect 336608 228624 336614 228636
rect 358814 228624 358820 228636
rect 358872 228624 358878 228676
rect 371050 228624 371056 228676
rect 371108 228664 371114 228676
rect 385218 228664 385224 228676
rect 371108 228636 385224 228664
rect 371108 228624 371114 228636
rect 385218 228624 385224 228636
rect 385276 228624 385282 228676
rect 404170 228624 404176 228676
rect 404228 228664 404234 228676
rect 410978 228664 410984 228676
rect 404228 228636 410984 228664
rect 404228 228624 404234 228636
rect 410978 228624 410984 228636
rect 411036 228624 411042 228676
rect 486878 228624 486884 228676
rect 486936 228664 486942 228676
rect 500954 228664 500960 228676
rect 486936 228636 500960 228664
rect 486936 228624 486942 228636
rect 500954 228624 500960 228636
rect 501012 228624 501018 228676
rect 506290 228624 506296 228676
rect 506348 228664 506354 228676
rect 526622 228664 526628 228676
rect 506348 228636 526628 228664
rect 506348 228624 506354 228636
rect 526622 228624 526628 228636
rect 526680 228624 526686 228676
rect 531406 228624 531412 228676
rect 531464 228664 531470 228676
rect 558270 228664 558276 228676
rect 531464 228636 558276 228664
rect 531464 228624 531470 228636
rect 558270 228624 558276 228636
rect 558328 228624 558334 228676
rect 64138 228488 64144 228540
rect 64196 228528 64202 228540
rect 143074 228528 143080 228540
rect 64196 228500 143080 228528
rect 64196 228488 64202 228500
rect 143074 228488 143080 228500
rect 143132 228488 143138 228540
rect 153102 228488 153108 228540
rect 153160 228528 153166 228540
rect 215846 228528 215852 228540
rect 153160 228500 215852 228528
rect 153160 228488 153166 228500
rect 215846 228488 215852 228500
rect 215904 228488 215910 228540
rect 222010 228488 222016 228540
rect 222068 228528 222074 228540
rect 269942 228528 269948 228540
rect 222068 228500 269948 228528
rect 222068 228488 222074 228500
rect 269942 228488 269948 228500
rect 270000 228488 270006 228540
rect 274082 228488 274088 228540
rect 274140 228528 274146 228540
rect 309226 228528 309232 228540
rect 274140 228500 309232 228528
rect 274140 228488 274146 228500
rect 309226 228488 309232 228500
rect 309284 228488 309290 228540
rect 326890 228488 326896 228540
rect 326948 228528 326954 228540
rect 351086 228528 351092 228540
rect 326948 228500 351092 228528
rect 326948 228488 326954 228500
rect 351086 228488 351092 228500
rect 351144 228488 351150 228540
rect 360102 228488 360108 228540
rect 360160 228528 360166 228540
rect 376846 228528 376852 228540
rect 360160 228500 376852 228528
rect 360160 228488 360166 228500
rect 376846 228488 376852 228500
rect 376904 228488 376910 228540
rect 377766 228488 377772 228540
rect 377824 228528 377830 228540
rect 390370 228528 390376 228540
rect 377824 228500 390376 228528
rect 377824 228488 377830 228500
rect 390370 228488 390376 228500
rect 390428 228488 390434 228540
rect 400214 228488 400220 228540
rect 400272 228528 400278 228540
rect 407758 228528 407764 228540
rect 400272 228500 407764 228528
rect 400272 228488 400278 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 410978 228488 410984 228540
rect 411036 228528 411042 228540
rect 416130 228528 416136 228540
rect 411036 228500 416136 228528
rect 411036 228488 411042 228500
rect 416130 228488 416136 228500
rect 416188 228488 416194 228540
rect 480070 228488 480076 228540
rect 480128 228528 480134 228540
rect 489178 228528 489184 228540
rect 480128 228500 489184 228528
rect 480128 228488 480134 228500
rect 489178 228488 489184 228500
rect 489236 228488 489242 228540
rect 495342 228488 495348 228540
rect 495400 228528 495406 228540
rect 510614 228528 510620 228540
rect 495400 228500 510620 228528
rect 495400 228488 495406 228500
rect 510614 228488 510620 228500
rect 510672 228488 510678 228540
rect 511442 228488 511448 228540
rect 511500 228528 511506 228540
rect 531958 228528 531964 228540
rect 511500 228500 531964 228528
rect 511500 228488 511506 228500
rect 531958 228488 531964 228500
rect 532016 228488 532022 228540
rect 537846 228488 537852 228540
rect 537904 228528 537910 228540
rect 566090 228528 566096 228540
rect 537904 228500 566096 228528
rect 537904 228488 537910 228500
rect 566090 228488 566096 228500
rect 566148 228488 566154 228540
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 141142 228392 141148 228404
rect 57296 228364 141148 228392
rect 57296 228352 57302 228364
rect 141142 228352 141148 228364
rect 141200 228352 141206 228404
rect 145926 228352 145932 228404
rect 145984 228392 145990 228404
rect 210694 228392 210700 228404
rect 145984 228364 210700 228392
rect 145984 228352 145990 228364
rect 210694 228352 210700 228364
rect 210752 228352 210758 228404
rect 215202 228352 215208 228404
rect 215260 228392 215266 228404
rect 266078 228392 266084 228404
rect 215260 228364 266084 228392
rect 215260 228352 215266 228364
rect 266078 228352 266084 228364
rect 266136 228352 266142 228404
rect 271782 228352 271788 228404
rect 271840 228392 271846 228404
rect 308582 228392 308588 228404
rect 271840 228364 308588 228392
rect 271840 228352 271846 228364
rect 308582 228352 308588 228364
rect 308640 228352 308646 228404
rect 312998 228352 313004 228404
rect 313056 228392 313062 228404
rect 340782 228392 340788 228404
rect 313056 228364 340788 228392
rect 313056 228352 313062 228364
rect 340782 228352 340788 228364
rect 340840 228352 340846 228404
rect 362678 228392 362684 228404
rect 344986 228364 362684 228392
rect 126698 228216 126704 228268
rect 126756 228256 126762 228268
rect 195238 228256 195244 228268
rect 126756 228228 195244 228256
rect 126756 228216 126762 228228
rect 195238 228216 195244 228228
rect 195296 228216 195302 228268
rect 205358 228216 205364 228268
rect 205416 228256 205422 228268
rect 257062 228256 257068 228268
rect 205416 228228 257068 228256
rect 205416 228216 205422 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 265618 228216 265624 228268
rect 265676 228256 265682 228268
rect 274450 228256 274456 228268
rect 265676 228228 274456 228256
rect 265676 228216 265682 228228
rect 274450 228216 274456 228228
rect 274508 228216 274514 228268
rect 309686 228216 309692 228268
rect 309744 228256 309750 228268
rect 327258 228256 327264 228268
rect 309744 228228 327264 228256
rect 309744 228216 309750 228228
rect 327258 228216 327264 228228
rect 327316 228216 327322 228268
rect 340138 228216 340144 228268
rect 340196 228256 340202 228268
rect 344986 228256 345014 228364
rect 362678 228352 362684 228364
rect 362736 228352 362742 228404
rect 362862 228352 362868 228404
rect 362920 228392 362926 228404
rect 379422 228392 379428 228404
rect 362920 228364 379428 228392
rect 362920 228352 362926 228364
rect 379422 228352 379428 228364
rect 379480 228352 379486 228404
rect 393590 228392 393596 228404
rect 383626 228364 393596 228392
rect 340196 228228 345014 228256
rect 340196 228216 340202 228228
rect 379238 228216 379244 228268
rect 379296 228256 379302 228268
rect 383626 228256 383654 228364
rect 393590 228352 393596 228364
rect 393648 228352 393654 228404
rect 409782 228352 409788 228404
rect 409840 228392 409846 228404
rect 415486 228392 415492 228404
rect 409840 228364 415492 228392
rect 409840 228352 409846 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 470226 228352 470232 228404
rect 470284 228392 470290 228404
rect 479702 228392 479708 228404
rect 470284 228364 479708 228392
rect 470284 228352 470290 228364
rect 479702 228352 479708 228364
rect 479760 228352 479766 228404
rect 481818 228352 481824 228404
rect 481876 228392 481882 228404
rect 494698 228392 494704 228404
rect 481876 228364 494704 228392
rect 481876 228352 481882 228364
rect 494698 228352 494704 228364
rect 494756 228352 494762 228404
rect 497274 228352 497280 228404
rect 497332 228392 497338 228404
rect 514294 228392 514300 228404
rect 497332 228364 514300 228392
rect 497332 228352 497338 228364
rect 514294 228352 514300 228364
rect 514352 228352 514358 228404
rect 521746 228352 521752 228404
rect 521804 228392 521810 228404
rect 545758 228392 545764 228404
rect 521804 228364 545764 228392
rect 521804 228352 521810 228364
rect 545758 228352 545764 228364
rect 545816 228352 545822 228404
rect 554038 228352 554044 228404
rect 554096 228392 554102 228404
rect 632698 228392 632704 228404
rect 554096 228364 632704 228392
rect 554096 228352 554102 228364
rect 632698 228352 632704 228364
rect 632756 228352 632762 228404
rect 672644 228392 672672 229112
rect 673454 229100 673460 229112
rect 673512 229100 673518 229152
rect 673736 229094 673788 229100
rect 672810 228964 672816 229016
rect 672868 229004 672874 229016
rect 672868 228976 672994 229004
rect 672868 228964 672874 228976
rect 672966 228664 672994 228976
rect 673598 228948 673650 228954
rect 673598 228890 673650 228896
rect 673506 228744 673558 228750
rect 673506 228686 673558 228692
rect 672966 228636 673414 228664
rect 672810 228488 672816 228540
rect 672868 228528 672874 228540
rect 672868 228500 673302 228528
rect 672868 228488 672874 228500
rect 672810 228392 672816 228404
rect 672644 228364 672816 228392
rect 672810 228352 672816 228364
rect 672868 228352 672874 228404
rect 379296 228228 383654 228256
rect 379296 228216 379302 228228
rect 390094 228216 390100 228268
rect 390152 228256 390158 228268
rect 400030 228256 400036 228268
rect 390152 228228 400036 228256
rect 390152 228216 390158 228228
rect 400030 228216 400036 228228
rect 400088 228216 400094 228268
rect 409046 228256 409052 228268
rect 402946 228228 409052 228256
rect 133506 228080 133512 228132
rect 133564 228120 133570 228132
rect 200390 228120 200396 228132
rect 133564 228092 200396 228120
rect 133564 228080 133570 228092
rect 200390 228080 200396 228092
rect 200448 228080 200454 228132
rect 211062 228080 211068 228132
rect 211120 228120 211126 228132
rect 260282 228120 260288 228132
rect 211120 228092 260288 228120
rect 211120 228080 211126 228092
rect 260282 228080 260288 228092
rect 260340 228080 260346 228132
rect 398650 228080 398656 228132
rect 398708 228120 398714 228132
rect 402946 228120 402974 228228
rect 409046 228216 409052 228228
rect 409104 228216 409110 228268
rect 523310 228216 523316 228268
rect 523368 228256 523374 228268
rect 527726 228256 527732 228268
rect 523368 228228 527732 228256
rect 523368 228216 523374 228228
rect 527726 228216 527732 228228
rect 527784 228216 527790 228268
rect 669406 228216 669412 228268
rect 669464 228256 669470 228268
rect 669464 228228 673190 228256
rect 669464 228216 669470 228228
rect 398708 228092 402974 228120
rect 398708 228080 398714 228092
rect 672350 228012 672356 228064
rect 672408 228052 672414 228064
rect 672408 228024 673072 228052
rect 672408 228012 672414 228024
rect 139302 227944 139308 227996
rect 139360 227984 139366 227996
rect 205542 227984 205548 227996
rect 139360 227956 205548 227984
rect 139360 227944 139366 227956
rect 205542 227944 205548 227956
rect 205600 227944 205606 227996
rect 252370 227944 252376 227996
rect 252428 227984 252434 227996
rect 293126 227984 293132 227996
rect 252428 227956 293132 227984
rect 252428 227944 252434 227956
rect 293126 227944 293132 227956
rect 293184 227944 293190 227996
rect 393958 227876 393964 227928
rect 394016 227916 394022 227928
rect 401318 227916 401324 227928
rect 394016 227888 401324 227916
rect 394016 227876 394022 227888
rect 401318 227876 401324 227888
rect 401376 227876 401382 227928
rect 402238 227876 402244 227928
rect 402296 227916 402302 227928
rect 402296 227888 402974 227916
rect 402296 227876 402302 227888
rect 143442 227808 143448 227860
rect 143500 227848 143506 227860
rect 146202 227848 146208 227860
rect 143500 227820 146208 227848
rect 143500 227808 143506 227820
rect 146202 227808 146208 227820
rect 146260 227808 146266 227860
rect 169570 227808 169576 227860
rect 169628 227848 169634 227860
rect 169938 227848 169944 227860
rect 169628 227820 169944 227848
rect 169628 227808 169634 227820
rect 169938 227808 169944 227820
rect 169996 227808 170002 227860
rect 196710 227808 196716 227860
rect 196768 227848 196774 227860
rect 230658 227848 230664 227860
rect 196768 227820 230664 227848
rect 196768 227808 196774 227820
rect 230658 227808 230664 227820
rect 230716 227808 230722 227860
rect 280706 227808 280712 227860
rect 280764 227848 280770 227860
rect 284754 227848 284760 227860
rect 280764 227820 284760 227848
rect 280764 227808 280770 227820
rect 284754 227808 284760 227820
rect 284812 227808 284818 227860
rect 297358 227808 297364 227860
rect 297416 227848 297422 227860
rect 305362 227848 305368 227860
rect 297416 227820 305368 227848
rect 297416 227808 297422 227820
rect 305362 227808 305368 227820
rect 305420 227808 305426 227860
rect 396626 227740 396632 227792
rect 396684 227780 396690 227792
rect 397454 227780 397460 227792
rect 396684 227752 397460 227780
rect 396684 227740 396690 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 400766 227740 400772 227792
rect 400824 227780 400830 227792
rect 402606 227780 402612 227792
rect 400824 227752 402612 227780
rect 400824 227740 400830 227752
rect 402606 227740 402612 227752
rect 402664 227740 402670 227792
rect 402946 227780 402974 227888
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 672810 227808 672816 227860
rect 672868 227848 672874 227860
rect 672868 227820 672980 227848
rect 672868 227808 672874 227820
rect 403250 227780 403256 227792
rect 402946 227752 403256 227780
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416682 227740 416688 227792
rect 416740 227780 416746 227792
rect 420638 227780 420644 227792
rect 416740 227752 420644 227780
rect 416740 227740 416746 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 474734 227740 474740 227792
rect 474792 227780 474798 227792
rect 482922 227780 482928 227792
rect 474792 227752 482928 227780
rect 474792 227740 474798 227752
rect 482922 227740 482928 227752
rect 482980 227740 482986 227792
rect 659470 227740 659476 227792
rect 659528 227780 659534 227792
rect 665174 227780 665180 227792
rect 659528 227752 665180 227780
rect 659528 227740 659534 227752
rect 665174 227740 665180 227752
rect 665232 227740 665238 227792
rect 116946 227672 116952 227724
rect 117004 227712 117010 227724
rect 187510 227712 187516 227724
rect 117004 227684 187516 227712
rect 117004 227672 117010 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 200022 227672 200028 227724
rect 200080 227712 200086 227724
rect 251910 227712 251916 227724
rect 200080 227684 251916 227712
rect 200080 227672 200086 227684
rect 251910 227672 251916 227684
rect 251968 227672 251974 227724
rect 263410 227672 263416 227724
rect 263468 227712 263474 227724
rect 301498 227712 301504 227724
rect 263468 227684 301504 227712
rect 263468 227672 263474 227684
rect 301498 227672 301504 227684
rect 301556 227672 301562 227724
rect 110138 227536 110144 227588
rect 110196 227576 110202 227588
rect 182358 227576 182364 227588
rect 110196 227548 182364 227576
rect 110196 227536 110202 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 182818 227536 182824 227588
rect 182876 227576 182882 227588
rect 236454 227576 236460 227588
rect 182876 227548 236460 227576
rect 182876 227536 182882 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 241974 227536 241980 227588
rect 242032 227576 242038 227588
rect 285398 227576 285404 227588
rect 242032 227548 285404 227576
rect 242032 227536 242038 227548
rect 285398 227536 285404 227548
rect 285456 227536 285462 227588
rect 293770 227536 293776 227588
rect 293828 227576 293834 227588
rect 325326 227576 325332 227588
rect 293828 227548 325332 227576
rect 293828 227536 293834 227548
rect 325326 227536 325332 227548
rect 325384 227536 325390 227588
rect 515398 227536 515404 227588
rect 515456 227576 515462 227588
rect 524966 227576 524972 227588
rect 515456 227548 524972 227576
rect 515456 227536 515462 227548
rect 524966 227536 524972 227548
rect 525024 227536 525030 227588
rect 526438 227536 526444 227588
rect 526496 227576 526502 227588
rect 544378 227576 544384 227588
rect 526496 227548 544384 227576
rect 526496 227536 526502 227548
rect 544378 227536 544384 227548
rect 544436 227536 544442 227588
rect 560938 227536 560944 227588
rect 560996 227576 561002 227588
rect 568114 227576 568120 227588
rect 560996 227548 568120 227576
rect 560996 227536 561002 227548
rect 568114 227536 568120 227548
rect 568172 227536 568178 227588
rect 672816 227520 672868 227526
rect 672816 227462 672868 227468
rect 103422 227400 103428 227452
rect 103480 227440 103486 227452
rect 177206 227440 177212 227452
rect 103480 227412 177212 227440
rect 103480 227400 103486 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 185578 227440 185584 227452
rect 180766 227412 185584 227440
rect 81342 227264 81348 227316
rect 81400 227304 81406 227316
rect 95234 227304 95240 227316
rect 81400 227276 95240 227304
rect 81400 227264 81406 227276
rect 95234 227264 95240 227276
rect 95292 227264 95298 227316
rect 96246 227264 96252 227316
rect 96304 227304 96310 227316
rect 172054 227304 172060 227316
rect 96304 227276 172060 227304
rect 96304 227264 96310 227276
rect 172054 227264 172060 227276
rect 172112 227264 172118 227316
rect 173158 227264 173164 227316
rect 173216 227304 173222 227316
rect 180766 227304 180794 227412
rect 185578 227400 185584 227412
rect 185636 227400 185642 227452
rect 188982 227400 188988 227452
rect 189040 227440 189046 227452
rect 244182 227440 244188 227452
rect 189040 227412 244188 227440
rect 189040 227400 189046 227412
rect 244182 227400 244188 227412
rect 244240 227400 244246 227452
rect 251082 227400 251088 227452
rect 251140 227440 251146 227452
rect 294414 227440 294420 227452
rect 251140 227412 294420 227440
rect 251140 227400 251146 227412
rect 294414 227400 294420 227412
rect 294472 227400 294478 227452
rect 302142 227400 302148 227452
rect 302200 227440 302206 227452
rect 331122 227440 331128 227452
rect 302200 227412 331128 227440
rect 302200 227400 302206 227412
rect 331122 227400 331128 227412
rect 331180 227400 331186 227452
rect 333882 227400 333888 227452
rect 333940 227440 333946 227452
rect 356238 227440 356244 227452
rect 333940 227412 356244 227440
rect 333940 227400 333946 227412
rect 356238 227400 356244 227412
rect 356296 227400 356302 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 671724 227412 672750 227440
rect 173216 227276 180794 227304
rect 173216 227264 173222 227276
rect 184934 227264 184940 227316
rect 184992 227304 184998 227316
rect 192662 227304 192668 227316
rect 184992 227276 192668 227304
rect 184992 227264 184998 227276
rect 192662 227264 192668 227276
rect 192720 227264 192726 227316
rect 198642 227264 198648 227316
rect 198700 227304 198706 227316
rect 253198 227304 253204 227316
rect 198700 227276 253204 227304
rect 198700 227264 198706 227276
rect 253198 227264 253204 227276
rect 253256 227264 253262 227316
rect 259362 227264 259368 227316
rect 259420 227304 259426 227316
rect 298278 227304 298284 227316
rect 259420 227276 298284 227304
rect 259420 227264 259426 227276
rect 298278 227264 298284 227276
rect 298336 227264 298342 227316
rect 308950 227264 308956 227316
rect 309008 227304 309014 227316
rect 339494 227304 339500 227316
rect 309008 227276 339500 227304
rect 309008 227264 309014 227276
rect 339494 227264 339500 227276
rect 339552 227264 339558 227316
rect 351086 227264 351092 227316
rect 351144 227304 351150 227316
rect 363322 227304 363328 227316
rect 351144 227276 363328 227304
rect 351144 227264 351150 227276
rect 363322 227264 363328 227276
rect 363380 227264 363386 227316
rect 363506 227264 363512 227316
rect 363564 227304 363570 227316
rect 368474 227304 368480 227316
rect 363564 227276 368480 227304
rect 363564 227264 363570 227276
rect 368474 227264 368480 227276
rect 368532 227264 368538 227316
rect 385678 227264 385684 227316
rect 385736 227304 385742 227316
rect 391658 227304 391664 227316
rect 385736 227276 391664 227304
rect 385736 227264 385742 227276
rect 391658 227264 391664 227276
rect 391716 227264 391722 227316
rect 477402 227264 477408 227316
rect 477460 227304 477466 227316
rect 485038 227304 485044 227316
rect 477460 227276 485044 227304
rect 477460 227264 477466 227276
rect 485038 227264 485044 227276
rect 485096 227264 485102 227316
rect 490834 227264 490840 227316
rect 490892 227304 490898 227316
rect 505462 227304 505468 227316
rect 490892 227276 505468 227304
rect 490892 227264 490898 227276
rect 505462 227264 505468 227276
rect 505520 227264 505526 227316
rect 506934 227264 506940 227316
rect 506992 227304 506998 227316
rect 526346 227304 526352 227316
rect 506992 227276 526352 227304
rect 506992 227264 506998 227276
rect 526346 227264 526352 227276
rect 526404 227264 526410 227316
rect 528186 227264 528192 227316
rect 528244 227304 528250 227316
rect 554038 227304 554044 227316
rect 528244 227276 554044 227304
rect 528244 227264 528250 227276
rect 554038 227264 554044 227276
rect 554096 227264 554102 227316
rect 68278 227128 68284 227180
rect 68336 227168 68342 227180
rect 146386 227168 146392 227180
rect 68336 227140 146392 227168
rect 68336 227128 68342 227140
rect 146386 227128 146392 227140
rect 146444 227128 146450 227180
rect 152918 227128 152924 227180
rect 152976 227168 152982 227180
rect 213362 227168 213368 227180
rect 152976 227140 213368 227168
rect 152976 227128 152982 227140
rect 213362 227128 213368 227140
rect 213420 227128 213426 227180
rect 224770 227128 224776 227180
rect 224828 227168 224834 227180
rect 273806 227168 273812 227180
rect 224828 227140 273812 227168
rect 224828 227128 224834 227140
rect 273806 227128 273812 227140
rect 273864 227128 273870 227180
rect 274266 227128 274272 227180
rect 274324 227168 274330 227180
rect 312446 227168 312452 227180
rect 274324 227140 312452 227168
rect 274324 227128 274330 227140
rect 312446 227128 312452 227140
rect 312504 227128 312510 227180
rect 319806 227128 319812 227180
rect 319864 227168 319870 227180
rect 345842 227168 345848 227180
rect 319864 227140 345848 227168
rect 319864 227128 319870 227140
rect 345842 227128 345848 227140
rect 345900 227128 345906 227180
rect 346118 227128 346124 227180
rect 346176 227168 346182 227180
rect 366542 227168 366548 227180
rect 346176 227140 366548 227168
rect 346176 227128 346182 227140
rect 366542 227128 366548 227140
rect 366600 227128 366606 227180
rect 369486 227128 369492 227180
rect 369544 227168 369550 227180
rect 384574 227168 384580 227180
rect 369544 227140 384580 227168
rect 369544 227128 369550 227140
rect 384574 227128 384580 227140
rect 384632 227128 384638 227180
rect 391566 227128 391572 227180
rect 391624 227168 391630 227180
rect 400582 227168 400588 227180
rect 391624 227140 400588 227168
rect 391624 227128 391630 227140
rect 400582 227128 400588 227140
rect 400640 227128 400646 227180
rect 401502 227128 401508 227180
rect 401560 227168 401566 227180
rect 408402 227168 408408 227180
rect 401560 227140 408408 227168
rect 401560 227128 401566 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 483750 227128 483756 227180
rect 483808 227168 483814 227180
rect 497550 227168 497556 227180
rect 483808 227140 497556 227168
rect 483808 227128 483814 227140
rect 497550 227128 497556 227140
rect 497608 227128 497614 227180
rect 498562 227128 498568 227180
rect 498620 227168 498626 227180
rect 515766 227168 515772 227180
rect 498620 227140 515772 227168
rect 498620 227128 498626 227140
rect 515766 227128 515772 227140
rect 515824 227128 515830 227180
rect 525610 227128 525616 227180
rect 525668 227168 525674 227180
rect 550818 227168 550824 227180
rect 525668 227140 550824 227168
rect 525668 227128 525674 227140
rect 550818 227128 550824 227140
rect 550876 227128 550882 227180
rect 671724 227100 671752 227412
rect 671890 227196 671896 227248
rect 671948 227236 671954 227248
rect 671948 227208 672630 227236
rect 671948 227196 671954 227208
rect 671724 227072 671860 227100
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142430 227032 142436 227044
rect 56560 227004 142436 227032
rect 56560 226992 56566 227004
rect 142430 226992 142436 227004
rect 142488 226992 142494 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 208118 227032 208124 227044
rect 143316 227004 208124 227032
rect 143316 226992 143322 227004
rect 208118 226992 208124 227004
rect 208176 226992 208182 227044
rect 226150 227032 226156 227044
rect 209746 227004 226156 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 184934 226896 184940 226908
rect 122800 226868 184940 226896
rect 122800 226856 122806 226868
rect 184934 226856 184940 226868
rect 184992 226856 184998 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 209746 226896 209774 227004
rect 226150 226992 226156 227004
rect 226208 226992 226214 227044
rect 228726 226992 228732 227044
rect 228784 227032 228790 227044
rect 275094 227032 275100 227044
rect 228784 227004 275100 227032
rect 228784 226992 228790 227004
rect 275094 226992 275100 227004
rect 275152 226992 275158 227044
rect 284846 226992 284852 227044
rect 284904 227032 284910 227044
rect 320174 227032 320180 227044
rect 284904 227004 320180 227032
rect 284904 226992 284910 227004
rect 320174 226992 320180 227004
rect 320232 226992 320238 227044
rect 325510 226992 325516 227044
rect 325568 227032 325574 227044
rect 349154 227032 349160 227044
rect 325568 227004 349160 227032
rect 325568 226992 325574 227004
rect 349154 226992 349160 227004
rect 349212 226992 349218 227044
rect 357250 226992 357256 227044
rect 357308 227032 357314 227044
rect 374270 227032 374276 227044
rect 357308 227004 374276 227032
rect 357308 226992 357314 227004
rect 374270 226992 374276 227004
rect 374328 226992 374334 227044
rect 376662 226992 376668 227044
rect 376720 227032 376726 227044
rect 389726 227032 389732 227044
rect 376720 227004 389732 227032
rect 376720 226992 376726 227004
rect 389726 226992 389732 227004
rect 389784 226992 389790 227044
rect 395798 226992 395804 227044
rect 395856 227032 395862 227044
rect 406470 227032 406476 227044
rect 395856 227004 406476 227032
rect 395856 226992 395862 227004
rect 406470 226992 406476 227004
rect 406528 226992 406534 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 491478 226992 491484 227044
rect 491536 227032 491542 227044
rect 506842 227032 506848 227044
rect 491536 227004 506848 227032
rect 491536 226992 491542 227004
rect 506842 226992 506848 227004
rect 506900 226992 506906 227044
rect 512086 226992 512092 227044
rect 512144 227032 512150 227044
rect 533430 227032 533436 227044
rect 512144 227004 533436 227032
rect 512144 226992 512150 227004
rect 533430 226992 533436 227004
rect 533488 226992 533494 227044
rect 535270 226992 535276 227044
rect 535328 227032 535334 227044
rect 562778 227032 562784 227044
rect 535328 227004 562784 227032
rect 535328 226992 535334 227004
rect 562778 226992 562784 227004
rect 562836 226992 562842 227044
rect 471514 226924 471520 226976
rect 471572 226964 471578 226976
rect 479518 226964 479524 226976
rect 471572 226936 479524 226964
rect 471572 226924 471578 226936
rect 479518 226924 479524 226936
rect 479576 226924 479582 226976
rect 671338 226924 671344 226976
rect 671396 226964 671402 226976
rect 671706 226964 671712 226976
rect 671396 226936 671712 226964
rect 671396 226924 671402 226936
rect 671706 226924 671712 226936
rect 671764 226924 671770 226976
rect 185636 226868 209774 226896
rect 185636 226856 185642 226868
rect 212166 226856 212172 226908
rect 212224 226896 212230 226908
rect 262214 226896 262220 226908
rect 212224 226868 262220 226896
rect 212224 226856 212230 226868
rect 262214 226856 262220 226868
rect 262272 226856 262278 226908
rect 275646 226856 275652 226908
rect 275704 226896 275710 226908
rect 311158 226896 311164 226908
rect 275704 226868 311164 226896
rect 275704 226856 275710 226868
rect 311158 226856 311164 226868
rect 311216 226856 311222 226908
rect 384942 226856 384948 226908
rect 385000 226896 385006 226908
rect 395522 226896 395528 226908
rect 385000 226868 395528 226896
rect 385000 226856 385006 226868
rect 395522 226856 395528 226868
rect 395580 226856 395586 226908
rect 419442 226856 419448 226908
rect 419500 226896 419506 226908
rect 424502 226896 424508 226908
rect 419500 226868 424508 226896
rect 419500 226856 419506 226868
rect 424502 226856 424508 226868
rect 424560 226856 424566 226908
rect 479886 226856 479892 226908
rect 479944 226896 479950 226908
rect 491938 226896 491944 226908
rect 479944 226868 491944 226896
rect 479944 226856 479950 226868
rect 491938 226856 491944 226868
rect 491996 226856 492002 226908
rect 671706 226788 671712 226840
rect 671764 226828 671770 226840
rect 671832 226828 671860 227072
rect 672092 227004 672520 227032
rect 672092 226840 672120 227004
rect 671764 226800 671860 226828
rect 671764 226788 671770 226800
rect 672074 226788 672080 226840
rect 672132 226788 672138 226840
rect 129366 226720 129372 226772
rect 129424 226760 129430 226772
rect 197814 226760 197820 226772
rect 129424 226732 197820 226760
rect 129424 226720 129430 226732
rect 197814 226720 197820 226732
rect 197872 226720 197878 226772
rect 224586 226720 224592 226772
rect 224644 226760 224650 226772
rect 270586 226760 270592 226772
rect 224644 226732 270592 226760
rect 224644 226720 224650 226732
rect 270586 226720 270592 226732
rect 270644 226720 270650 226772
rect 672374 226652 672380 226704
rect 672432 226652 672438 226704
rect 150250 226584 150256 226636
rect 150308 226624 150314 226636
rect 152918 226624 152924 226636
rect 150308 226596 152924 226624
rect 150308 226584 150314 226596
rect 152918 226584 152924 226596
rect 152976 226584 152982 226636
rect 160002 226584 160008 226636
rect 160060 226624 160066 226636
rect 220998 226624 221004 226636
rect 160060 226596 221004 226624
rect 160060 226584 160066 226596
rect 220998 226584 221004 226596
rect 221056 226584 221062 226636
rect 671936 226584 671942 226636
rect 671994 226624 672000 226636
rect 671994 226596 672290 226624
rect 671994 226584 672000 226596
rect 177206 226448 177212 226500
rect 177264 226488 177270 226500
rect 231302 226488 231308 226500
rect 177264 226460 231308 226488
rect 177264 226448 177270 226460
rect 231302 226448 231308 226460
rect 231360 226448 231366 226500
rect 465902 226448 465908 226500
rect 465960 226488 465966 226500
rect 469858 226488 469864 226500
rect 465960 226460 469864 226488
rect 465960 226448 465966 226460
rect 469858 226448 469864 226460
rect 469916 226448 469922 226500
rect 671814 226448 671820 226500
rect 671872 226488 671878 226500
rect 671872 226460 672182 226488
rect 671872 226448 671878 226460
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 411622 226352 411628 226364
rect 407816 226324 411628 226352
rect 407816 226312 407822 226324
rect 411622 226312 411628 226324
rect 411680 226312 411686 226364
rect 135162 226244 135168 226296
rect 135220 226284 135226 226296
rect 204254 226284 204260 226296
rect 135220 226256 204260 226284
rect 135220 226244 135226 226256
rect 204254 226244 204260 226256
rect 204312 226244 204318 226296
rect 205542 226244 205548 226296
rect 205600 226284 205606 226296
rect 205600 226256 209774 226284
rect 205600 226244 205606 226256
rect 99282 226108 99288 226160
rect 99340 226148 99346 226160
rect 175918 226148 175924 226160
rect 99340 226120 175924 226148
rect 99340 226108 99346 226120
rect 175918 226108 175924 226120
rect 175976 226108 175982 226160
rect 202690 226108 202696 226160
rect 202748 226148 202754 226160
rect 206738 226148 206744 226160
rect 202748 226120 206744 226148
rect 202748 226108 202754 226120
rect 206738 226108 206744 226120
rect 206796 226108 206802 226160
rect 209746 226148 209774 226256
rect 219342 226244 219348 226296
rect 219400 226284 219406 226296
rect 267366 226284 267372 226296
rect 219400 226256 267372 226284
rect 219400 226244 219406 226256
rect 267366 226244 267372 226256
rect 267424 226244 267430 226296
rect 303246 226244 303252 226296
rect 303304 226284 303310 226296
rect 333054 226284 333060 226296
rect 303304 226256 333060 226284
rect 303304 226244 303310 226256
rect 333054 226244 333060 226256
rect 333112 226244 333118 226296
rect 672034 226160 672086 226166
rect 258350 226148 258356 226160
rect 209746 226120 258356 226148
rect 258350 226108 258356 226120
rect 258408 226108 258414 226160
rect 286686 226108 286692 226160
rect 286744 226148 286750 226160
rect 319530 226148 319536 226160
rect 286744 226120 319536 226148
rect 286744 226108 286750 226120
rect 319530 226108 319536 226120
rect 319588 226108 319594 226160
rect 350350 226108 350356 226160
rect 350408 226148 350414 226160
rect 354858 226148 354864 226160
rect 350408 226120 354864 226148
rect 350408 226108 350414 226120
rect 354858 226108 354864 226120
rect 354916 226108 354922 226160
rect 501138 226108 501144 226160
rect 501196 226148 501202 226160
rect 519262 226148 519268 226160
rect 501196 226120 519268 226148
rect 501196 226108 501202 226120
rect 519262 226108 519268 226120
rect 519320 226108 519326 226160
rect 529934 226108 529940 226160
rect 529992 226148 529998 226160
rect 549898 226148 549904 226160
rect 529992 226120 549904 226148
rect 529992 226108 529998 226120
rect 549898 226108 549904 226120
rect 549956 226108 549962 226160
rect 672034 226102 672086 226108
rect 84102 225972 84108 226024
rect 84160 226012 84166 226024
rect 161750 226012 161756 226024
rect 84160 225984 161756 226012
rect 84160 225972 84166 225984
rect 161750 225972 161756 225984
rect 161808 225972 161814 226024
rect 186038 225972 186044 226024
rect 186096 226012 186102 226024
rect 241606 226012 241612 226024
rect 186096 225984 241612 226012
rect 186096 225972 186102 225984
rect 241606 225972 241612 225984
rect 241664 225972 241670 226024
rect 245286 225972 245292 226024
rect 245344 226012 245350 226024
rect 287606 226012 287612 226024
rect 245344 225984 287612 226012
rect 245344 225972 245350 225984
rect 287606 225972 287612 225984
rect 287664 225972 287670 226024
rect 296622 225972 296628 226024
rect 296680 226012 296686 226024
rect 329190 226012 329196 226024
rect 296680 225984 329196 226012
rect 296680 225972 296686 225984
rect 329190 225972 329196 225984
rect 329248 225972 329254 226024
rect 330386 225972 330392 226024
rect 330444 226012 330450 226024
rect 351914 226012 351920 226024
rect 330444 225984 351920 226012
rect 330444 225972 330450 225984
rect 351914 225972 351920 225984
rect 351972 225972 351978 226024
rect 352558 225972 352564 226024
rect 352616 226012 352622 226024
rect 358170 226012 358176 226024
rect 352616 225984 358176 226012
rect 352616 225972 352622 225984
rect 358170 225972 358176 225984
rect 358228 225972 358234 226024
rect 515950 225972 515956 226024
rect 516008 226012 516014 226024
rect 538950 226012 538956 226024
rect 516008 225984 538956 226012
rect 516008 225972 516014 225984
rect 538950 225972 538956 225984
rect 539008 225972 539014 226024
rect 671942 225956 671994 225962
rect 671942 225898 671994 225904
rect 70302 225836 70308 225888
rect 70360 225876 70366 225888
rect 151446 225876 151452 225888
rect 70360 225848 151452 225876
rect 70360 225836 70366 225848
rect 151446 225836 151452 225848
rect 151504 225836 151510 225888
rect 158346 225836 158352 225888
rect 158404 225876 158410 225888
rect 222286 225876 222292 225888
rect 158404 225848 222292 225876
rect 158404 225836 158410 225848
rect 222286 225836 222292 225848
rect 222344 225836 222350 225888
rect 239398 225836 239404 225888
rect 239456 225876 239462 225888
rect 284110 225876 284116 225888
rect 239456 225848 284116 225876
rect 239456 225836 239462 225848
rect 284110 225836 284116 225848
rect 284168 225836 284174 225888
rect 288250 225836 288256 225888
rect 288308 225876 288314 225888
rect 321462 225876 321468 225888
rect 288308 225848 321468 225876
rect 288308 225836 288314 225848
rect 321462 225836 321468 225848
rect 321520 225836 321526 225888
rect 324222 225836 324228 225888
rect 324280 225876 324286 225888
rect 348510 225876 348516 225888
rect 324280 225848 348516 225876
rect 324280 225836 324286 225848
rect 348510 225836 348516 225848
rect 348568 225836 348574 225888
rect 355318 225836 355324 225888
rect 355376 225876 355382 225888
rect 372338 225876 372344 225888
rect 355376 225848 372344 225876
rect 355376 225836 355382 225848
rect 372338 225836 372344 225848
rect 372396 225836 372402 225888
rect 495986 225836 495992 225888
rect 496044 225876 496050 225888
rect 512454 225876 512460 225888
rect 496044 225848 512460 225876
rect 496044 225836 496050 225848
rect 512454 225836 512460 225848
rect 512512 225836 512518 225888
rect 524322 225836 524328 225888
rect 524380 225876 524386 225888
rect 547874 225876 547880 225888
rect 524380 225848 547880 225876
rect 524380 225836 524386 225848
rect 547874 225836 547880 225848
rect 547932 225836 547938 225888
rect 555418 225836 555424 225888
rect 555476 225876 555482 225888
rect 570782 225876 570788 225888
rect 555476 225848 570788 225876
rect 555476 225836 555482 225848
rect 570782 225836 570788 225848
rect 570840 225836 570846 225888
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 671820 225752 671872 225758
rect 59998 225700 60004 225752
rect 60056 225740 60062 225752
rect 141786 225740 141792 225752
rect 60056 225712 141792 225740
rect 60056 225700 60062 225712
rect 141786 225700 141792 225712
rect 141844 225700 141850 225752
rect 141970 225700 141976 225752
rect 142028 225740 142034 225752
rect 209406 225740 209412 225752
rect 142028 225712 209412 225740
rect 142028 225700 142034 225712
rect 209406 225700 209412 225712
rect 209464 225700 209470 225752
rect 209590 225700 209596 225752
rect 209648 225740 209654 225752
rect 259638 225740 259644 225752
rect 209648 225712 259644 225740
rect 209648 225700 209654 225712
rect 259638 225700 259644 225712
rect 259696 225700 259702 225752
rect 264882 225700 264888 225752
rect 264940 225740 264946 225752
rect 304718 225740 304724 225752
rect 264940 225712 304724 225740
rect 264940 225700 264946 225712
rect 304718 225700 304724 225712
rect 304776 225700 304782 225752
rect 319990 225700 319996 225752
rect 320048 225740 320054 225752
rect 347222 225740 347228 225752
rect 320048 225712 347228 225740
rect 320048 225700 320054 225712
rect 347222 225700 347228 225712
rect 347280 225700 347286 225752
rect 349062 225700 349068 225752
rect 349120 225740 349126 225752
rect 367186 225740 367192 225752
rect 349120 225712 367192 225740
rect 349120 225700 349126 225712
rect 367186 225700 367192 225712
rect 367244 225700 367250 225752
rect 375282 225700 375288 225752
rect 375340 225740 375346 225752
rect 387794 225740 387800 225752
rect 375340 225712 387800 225740
rect 375340 225700 375346 225712
rect 387794 225700 387800 225712
rect 387852 225700 387858 225752
rect 388438 225700 388444 225752
rect 388496 225740 388502 225752
rect 396442 225740 396448 225752
rect 388496 225712 396448 225740
rect 388496 225700 388502 225712
rect 396442 225700 396448 225712
rect 396500 225700 396506 225752
rect 476022 225700 476028 225752
rect 476080 225740 476086 225752
rect 483566 225740 483572 225752
rect 476080 225712 483572 225740
rect 476080 225700 476086 225712
rect 483566 225700 483572 225712
rect 483624 225700 483630 225752
rect 489546 225700 489552 225752
rect 489604 225740 489610 225752
rect 504174 225740 504180 225752
rect 489604 225712 504180 225740
rect 489604 225700 489610 225712
rect 504174 225700 504180 225712
rect 504232 225700 504238 225752
rect 510154 225700 510160 225752
rect 510212 225740 510218 225752
rect 530854 225740 530860 225752
rect 510212 225712 530860 225740
rect 510212 225700 510218 225712
rect 530854 225700 530860 225712
rect 530912 225700 530918 225752
rect 533982 225700 533988 225752
rect 534040 225740 534046 225752
rect 561490 225740 561496 225752
rect 534040 225712 561496 225740
rect 534040 225700 534046 225712
rect 561490 225700 561496 225712
rect 561548 225700 561554 225752
rect 671820 225694 671872 225700
rect 667934 225632 667940 225684
rect 667992 225672 667998 225684
rect 667992 225644 671738 225672
rect 667992 225632 667998 225644
rect 62022 225564 62028 225616
rect 62080 225604 62086 225616
rect 144362 225604 144368 225616
rect 62080 225576 144368 225604
rect 62080 225564 62086 225576
rect 144362 225564 144368 225576
rect 144420 225564 144426 225616
rect 155862 225564 155868 225616
rect 155920 225604 155926 225616
rect 219710 225604 219716 225616
rect 155920 225576 219716 225604
rect 155920 225564 155926 225576
rect 219710 225564 219716 225576
rect 219768 225564 219774 225616
rect 220446 225564 220452 225616
rect 220504 225604 220510 225616
rect 268010 225604 268016 225616
rect 220504 225576 268016 225604
rect 220504 225564 220510 225576
rect 268010 225564 268016 225576
rect 268068 225564 268074 225616
rect 269022 225564 269028 225616
rect 269080 225604 269086 225616
rect 306006 225604 306012 225616
rect 269080 225576 306012 225604
rect 269080 225564 269086 225576
rect 306006 225564 306012 225576
rect 306064 225564 306070 225616
rect 306190 225564 306196 225616
rect 306248 225604 306254 225616
rect 336918 225604 336924 225616
rect 306248 225576 336924 225604
rect 306248 225564 306254 225576
rect 336918 225564 336924 225576
rect 336976 225564 336982 225616
rect 340690 225564 340696 225616
rect 340748 225604 340754 225616
rect 361482 225604 361488 225616
rect 340748 225576 361488 225604
rect 340748 225564 340754 225576
rect 361482 225564 361488 225576
rect 361540 225564 361546 225616
rect 365530 225564 365536 225616
rect 365588 225604 365594 225616
rect 379790 225604 379796 225616
rect 365588 225576 379796 225604
rect 365588 225564 365594 225576
rect 379790 225564 379796 225576
rect 379848 225564 379854 225616
rect 380066 225564 380072 225616
rect 380124 225604 380130 225616
rect 391014 225604 391020 225616
rect 380124 225576 391020 225604
rect 380124 225564 380130 225576
rect 391014 225564 391020 225576
rect 391072 225564 391078 225616
rect 391750 225564 391756 225616
rect 391808 225604 391814 225616
rect 403526 225604 403532 225616
rect 391808 225576 403532 225604
rect 391808 225564 391814 225576
rect 403526 225564 403532 225576
rect 403584 225564 403590 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 477034 225604 477040 225616
rect 467708 225576 477040 225604
rect 467708 225564 467714 225576
rect 477034 225564 477040 225576
rect 477092 225564 477098 225616
rect 481174 225564 481180 225616
rect 481232 225604 481238 225616
rect 493686 225604 493692 225616
rect 481232 225576 493692 225604
rect 481232 225564 481238 225576
rect 493686 225564 493692 225576
rect 493744 225564 493750 225616
rect 508866 225564 508872 225616
rect 508924 225604 508930 225616
rect 529198 225604 529204 225616
rect 508924 225576 529204 225604
rect 508924 225564 508930 225576
rect 529198 225564 529204 225576
rect 529256 225564 529262 225616
rect 529474 225564 529480 225616
rect 529532 225604 529538 225616
rect 555878 225604 555884 225616
rect 529532 225576 555884 225604
rect 529532 225564 529538 225576
rect 555878 225564 555884 225576
rect 555936 225564 555942 225616
rect 132402 225428 132408 225480
rect 132460 225468 132466 225480
rect 201678 225468 201684 225480
rect 132460 225440 201684 225468
rect 132460 225428 132466 225440
rect 201678 225428 201684 225440
rect 201736 225428 201742 225480
rect 206186 225428 206192 225480
rect 206244 225468 206250 225480
rect 206244 225440 206600 225468
rect 206244 225428 206250 225440
rect 139118 225292 139124 225344
rect 139176 225332 139182 225344
rect 206370 225332 206376 225344
rect 139176 225304 206376 225332
rect 139176 225292 139182 225304
rect 206370 225292 206376 225304
rect 206428 225292 206434 225344
rect 206572 225332 206600 225440
rect 206738 225428 206744 225480
rect 206796 225468 206802 225480
rect 254486 225468 254492 225480
rect 206796 225440 254492 225468
rect 206796 225428 206802 225440
rect 254486 225428 254492 225440
rect 254544 225428 254550 225480
rect 255222 225428 255228 225480
rect 255280 225468 255286 225480
rect 296990 225468 296996 225480
rect 255280 225440 296996 225468
rect 255280 225428 255286 225440
rect 296990 225428 296996 225440
rect 297048 225428 297054 225480
rect 492766 225428 492772 225480
rect 492824 225468 492830 225480
rect 508682 225468 508688 225480
rect 492824 225440 508688 225468
rect 492824 225428 492830 225440
rect 508682 225428 508688 225440
rect 508740 225428 508746 225480
rect 671596 225344 671648 225350
rect 228082 225332 228088 225344
rect 206572 225304 228088 225332
rect 228082 225292 228088 225304
rect 228140 225292 228146 225344
rect 255038 225292 255044 225344
rect 255096 225332 255102 225344
rect 295702 225332 295708 225344
rect 255096 225304 295708 225332
rect 255096 225292 255102 225304
rect 295702 225292 295708 225304
rect 295760 225292 295766 225344
rect 671596 225286 671648 225292
rect 155678 225156 155684 225208
rect 155736 225196 155742 225208
rect 218422 225196 218428 225208
rect 155736 225168 218428 225196
rect 155736 225156 155742 225168
rect 218422 225156 218428 225168
rect 218480 225156 218486 225208
rect 225598 225156 225604 225208
rect 225656 225196 225662 225208
rect 246114 225196 246120 225208
rect 225656 225168 246120 225196
rect 225656 225156 225662 225168
rect 246114 225156 246120 225168
rect 246172 225156 246178 225208
rect 671482 225140 671534 225146
rect 671482 225082 671534 225088
rect 166258 225020 166264 225072
rect 166316 225060 166322 225072
rect 186866 225060 186872 225072
rect 166316 225032 186872 225060
rect 166316 225020 166322 225032
rect 186866 225020 186872 225032
rect 186924 225020 186930 225072
rect 195606 225020 195612 225072
rect 195664 225060 195670 225072
rect 249334 225060 249340 225072
rect 195664 225032 249340 225060
rect 195664 225020 195670 225032
rect 249334 225020 249340 225032
rect 249392 225020 249398 225072
rect 404354 225020 404360 225072
rect 404412 225060 404418 225072
rect 412266 225060 412272 225072
rect 404412 225032 412272 225060
rect 404412 225020 404418 225032
rect 412266 225020 412272 225032
rect 412324 225020 412330 225072
rect 463142 225020 463148 225072
rect 463200 225060 463206 225072
rect 467466 225060 467472 225072
rect 463200 225032 467472 225060
rect 463200 225020 463206 225032
rect 467466 225020 467472 225032
rect 467524 225020 467530 225072
rect 669406 225020 669412 225072
rect 669464 225060 669470 225072
rect 669464 225032 671398 225060
rect 669464 225020 669470 225032
rect 260006 224952 260012 225004
rect 260064 224992 260070 225004
rect 264146 224992 264152 225004
rect 260064 224964 264152 224992
rect 260064 224952 260070 224964
rect 264146 224952 264152 224964
rect 264204 224952 264210 225004
rect 367646 224952 367652 225004
rect 367704 224992 367710 225004
rect 373626 224992 373632 225004
rect 367704 224964 373632 224992
rect 367704 224952 367710 224964
rect 373626 224952 373632 224964
rect 373684 224952 373690 225004
rect 118602 224884 118608 224936
rect 118660 224924 118666 224936
rect 185578 224924 185584 224936
rect 118660 224896 185584 224924
rect 118660 224884 118666 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 191466 224884 191472 224936
rect 191524 224924 191530 224936
rect 248046 224924 248052 224936
rect 191524 224896 248052 224924
rect 191524 224884 191530 224896
rect 248046 224884 248052 224896
rect 248104 224884 248110 224936
rect 266262 224884 266268 224936
rect 266320 224924 266326 224936
rect 303430 224924 303436 224936
rect 266320 224896 303436 224924
rect 266320 224884 266326 224896
rect 303430 224884 303436 224896
rect 303488 224884 303494 224936
rect 321462 224884 321468 224936
rect 321520 224924 321526 224936
rect 346578 224924 346584 224936
rect 321520 224896 346584 224924
rect 321520 224884 321526 224896
rect 346578 224884 346584 224896
rect 346636 224884 346642 224936
rect 426434 224884 426440 224936
rect 426492 224924 426498 224936
rect 426986 224924 426992 224936
rect 426492 224896 426992 224924
rect 426492 224884 426498 224896
rect 426986 224884 426992 224896
rect 427044 224884 427050 224936
rect 460566 224884 460572 224936
rect 460624 224924 460630 224936
rect 463142 224924 463148 224936
rect 460624 224896 463148 224924
rect 460624 224884 460630 224896
rect 463142 224884 463148 224896
rect 463200 224884 463206 224936
rect 669406 224816 669412 224868
rect 669464 224856 669470 224868
rect 669464 224828 671278 224856
rect 669464 224816 669470 224828
rect 112806 224748 112812 224800
rect 112864 224788 112870 224800
rect 185854 224788 185860 224800
rect 112864 224760 185860 224788
rect 112864 224748 112870 224760
rect 185854 224748 185860 224760
rect 185912 224748 185918 224800
rect 242894 224788 242900 224800
rect 186056 224760 242900 224788
rect 105998 224612 106004 224664
rect 106056 224652 106062 224664
rect 181070 224652 181076 224664
rect 106056 224624 181076 224652
rect 106056 224612 106062 224624
rect 181070 224612 181076 224624
rect 181128 224612 181134 224664
rect 181990 224612 181996 224664
rect 182048 224652 182054 224664
rect 185210 224652 185216 224664
rect 182048 224624 185216 224652
rect 182048 224612 182054 224624
rect 185210 224612 185216 224624
rect 185268 224612 185274 224664
rect 185394 224612 185400 224664
rect 185452 224652 185458 224664
rect 186056 224652 186084 224760
rect 242894 224748 242900 224760
rect 242952 224748 242958 224800
rect 271598 224748 271604 224800
rect 271656 224788 271662 224800
rect 309870 224788 309876 224800
rect 271656 224760 309876 224788
rect 271656 224748 271662 224760
rect 309870 224748 309876 224760
rect 309928 224748 309934 224800
rect 313182 224748 313188 224800
rect 313240 224788 313246 224800
rect 342070 224788 342076 224800
rect 313240 224760 342076 224788
rect 313240 224748 313246 224760
rect 342070 224748 342076 224760
rect 342128 224748 342134 224800
rect 365898 224788 365904 224800
rect 354646 224760 365904 224788
rect 185452 224624 186084 224652
rect 185452 224612 185458 224624
rect 186222 224612 186228 224664
rect 186280 224652 186286 224664
rect 240318 224652 240324 224664
rect 186280 224624 240324 224652
rect 186280 224612 186286 224624
rect 240318 224612 240324 224624
rect 240376 224612 240382 224664
rect 249610 224612 249616 224664
rect 249668 224652 249674 224664
rect 290550 224652 290556 224664
rect 249668 224624 290556 224652
rect 249668 224612 249674 224624
rect 290550 224612 290556 224624
rect 290608 224612 290614 224664
rect 294966 224612 294972 224664
rect 295024 224652 295030 224664
rect 325970 224652 325976 224664
rect 295024 224624 325976 224652
rect 295024 224612 295030 224624
rect 325970 224612 325976 224624
rect 326028 224612 326034 224664
rect 347038 224612 347044 224664
rect 347096 224652 347102 224664
rect 354646 224652 354674 224760
rect 365898 224748 365904 224760
rect 365956 224748 365962 224800
rect 670970 224680 670976 224732
rect 671028 224720 671034 224732
rect 671028 224692 671186 224720
rect 671028 224680 671034 224692
rect 363966 224652 363972 224664
rect 347096 224624 354674 224652
rect 359292 224624 363972 224652
rect 347096 224612 347102 224624
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 172330 224476 172336 224528
rect 172388 224516 172394 224528
rect 232590 224516 232596 224528
rect 172388 224488 232596 224516
rect 172388 224476 172394 224488
rect 232590 224476 232596 224488
rect 232648 224476 232654 224528
rect 233142 224476 233148 224528
rect 233200 224516 233206 224528
rect 277670 224516 277676 224528
rect 233200 224488 277676 224516
rect 233200 224476 233206 224488
rect 277670 224476 277676 224488
rect 277728 224476 277734 224528
rect 282454 224476 282460 224528
rect 282512 224516 282518 224528
rect 316310 224516 316316 224528
rect 282512 224488 316316 224516
rect 282512 224476 282518 224488
rect 316310 224476 316316 224488
rect 316368 224476 316374 224528
rect 317138 224476 317144 224528
rect 317196 224516 317202 224528
rect 342990 224516 342996 224528
rect 317196 224488 342996 224516
rect 317196 224476 317202 224488
rect 342990 224476 342996 224488
rect 343048 224476 343054 224528
rect 343450 224476 343456 224528
rect 343508 224516 343514 224528
rect 359292 224516 359320 224624
rect 363966 224612 363972 224624
rect 364024 224612 364030 224664
rect 499206 224612 499212 224664
rect 499264 224652 499270 224664
rect 516778 224652 516784 224664
rect 499264 224624 516784 224652
rect 499264 224612 499270 224624
rect 516778 224612 516784 224624
rect 516836 224612 516842 224664
rect 518526 224612 518532 224664
rect 518584 224652 518590 224664
rect 541618 224652 541624 224664
rect 518584 224624 541624 224652
rect 518584 224612 518590 224624
rect 541618 224612 541624 224624
rect 541676 224612 541682 224664
rect 343508 224488 359320 224516
rect 343508 224476 343514 224488
rect 363782 224476 363788 224528
rect 363840 224516 363846 224528
rect 378134 224516 378140 224528
rect 363840 224488 378140 224516
rect 363840 224476 363846 224488
rect 378134 224476 378140 224488
rect 378192 224476 378198 224528
rect 387702 224476 387708 224528
rect 387760 224516 387766 224528
rect 398098 224516 398104 224528
rect 387760 224488 398104 224516
rect 387760 224476 387766 224488
rect 398098 224476 398104 224488
rect 398156 224476 398162 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 505002 224476 505008 224528
rect 505060 224516 505066 224528
rect 523034 224516 523040 224528
rect 505060 224488 523040 224516
rect 505060 224476 505066 224488
rect 523034 224476 523040 224488
rect 523092 224476 523098 224528
rect 523678 224476 523684 224528
rect 523736 224516 523742 224528
rect 548334 224516 548340 224528
rect 523736 224488 548340 224516
rect 523736 224476 523742 224488
rect 548334 224476 548340 224488
rect 548392 224476 548398 224528
rect 666830 224408 666836 224460
rect 666888 224448 666894 224460
rect 666888 224420 671048 224448
rect 666888 224408 666894 224420
rect 76558 224340 76564 224392
rect 76616 224380 76622 224392
rect 157886 224380 157892 224392
rect 76616 224352 157892 224380
rect 76616 224340 76622 224352
rect 157886 224340 157892 224352
rect 157944 224340 157950 224392
rect 165522 224340 165528 224392
rect 165580 224380 165586 224392
rect 227438 224380 227444 224392
rect 165580 224352 227444 224380
rect 165580 224340 165586 224352
rect 227438 224340 227444 224352
rect 227496 224340 227502 224392
rect 241146 224340 241152 224392
rect 241204 224380 241210 224392
rect 286502 224380 286508 224392
rect 241204 224352 286508 224380
rect 241204 224340 241210 224352
rect 286502 224340 286508 224352
rect 286560 224340 286566 224392
rect 291010 224340 291016 224392
rect 291068 224380 291074 224392
rect 324038 224380 324044 224392
rect 291068 224352 324044 224380
rect 291068 224340 291074 224352
rect 324038 224340 324044 224352
rect 324096 224340 324102 224392
rect 341978 224340 341984 224392
rect 342036 224380 342042 224392
rect 365254 224380 365260 224392
rect 342036 224352 365260 224380
rect 342036 224340 342042 224352
rect 365254 224340 365260 224352
rect 365312 224340 365318 224392
rect 368382 224340 368388 224392
rect 368440 224380 368446 224392
rect 382550 224380 382556 224392
rect 368440 224352 382556 224380
rect 368440 224340 368446 224352
rect 382550 224340 382556 224352
rect 382608 224340 382614 224392
rect 382918 224340 382924 224392
rect 382976 224380 382982 224392
rect 396166 224380 396172 224392
rect 382976 224352 396172 224380
rect 382976 224340 382982 224352
rect 396166 224340 396172 224352
rect 396224 224340 396230 224392
rect 436370 224340 436376 224392
rect 436428 224380 436434 224392
rect 436830 224380 436836 224392
rect 436428 224352 436836 224380
rect 436428 224340 436434 224352
rect 436830 224340 436836 224352
rect 436888 224340 436894 224392
rect 462498 224340 462504 224392
rect 462556 224380 462562 224392
rect 469306 224380 469312 224392
rect 462556 224352 469312 224380
rect 462556 224340 462562 224352
rect 469306 224340 469312 224352
rect 469364 224340 469370 224392
rect 478598 224340 478604 224392
rect 478656 224380 478662 224392
rect 490282 224380 490288 224392
rect 478656 224352 490288 224380
rect 478656 224340 478662 224352
rect 490282 224340 490288 224352
rect 490340 224340 490346 224392
rect 492122 224340 492128 224392
rect 492180 224380 492186 224392
rect 507762 224380 507768 224392
rect 492180 224352 507768 224380
rect 492180 224340 492186 224352
rect 507762 224340 507768 224352
rect 507820 224340 507826 224392
rect 514662 224340 514668 224392
rect 514720 224380 514726 224392
rect 535638 224380 535644 224392
rect 514720 224352 535644 224380
rect 514720 224340 514726 224352
rect 535638 224340 535644 224352
rect 535696 224340 535702 224392
rect 536006 224340 536012 224392
rect 536064 224380 536070 224392
rect 563974 224380 563980 224392
rect 536064 224352 563980 224380
rect 536064 224340 536070 224352
rect 563974 224340 563980 224352
rect 564032 224340 564038 224392
rect 565630 224272 565636 224324
rect 565688 224312 565694 224324
rect 568574 224312 568580 224324
rect 565688 224284 568580 224312
rect 565688 224272 565694 224284
rect 568574 224272 568580 224284
rect 568632 224272 568638 224324
rect 63402 224204 63408 224256
rect 63460 224244 63466 224256
rect 147582 224244 147588 224256
rect 63460 224216 147588 224244
rect 63460 224204 63466 224216
rect 147582 224204 147588 224216
rect 147640 224204 147646 224256
rect 151722 224204 151728 224256
rect 151780 224244 151786 224256
rect 217134 224244 217140 224256
rect 151780 224216 217140 224244
rect 151780 224204 151786 224216
rect 217134 224204 217140 224216
rect 217192 224204 217198 224256
rect 223482 224204 223488 224256
rect 223540 224244 223546 224256
rect 225782 224244 225788 224256
rect 223540 224216 225788 224244
rect 223540 224204 223546 224216
rect 225782 224204 225788 224216
rect 225840 224204 225846 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 281442 224204 281448 224256
rect 281500 224244 281506 224256
rect 317598 224244 317604 224256
rect 281500 224216 317604 224244
rect 281500 224204 281506 224216
rect 317598 224204 317604 224216
rect 317656 224204 317662 224256
rect 322290 224204 322296 224256
rect 322348 224244 322354 224256
rect 349798 224244 349804 224256
rect 322348 224216 349804 224244
rect 322348 224204 322354 224216
rect 349798 224204 349804 224216
rect 349856 224204 349862 224256
rect 351730 224204 351736 224256
rect 351788 224244 351794 224256
rect 369762 224244 369768 224256
rect 351788 224216 369768 224244
rect 351788 224204 351794 224216
rect 369762 224204 369768 224216
rect 369820 224204 369826 224256
rect 372430 224204 372436 224256
rect 372488 224244 372494 224256
rect 387334 224244 387340 224256
rect 372488 224216 387340 224244
rect 372488 224204 372494 224216
rect 387334 224204 387340 224216
rect 387392 224204 387398 224256
rect 394510 224204 394516 224256
rect 394568 224244 394574 224256
rect 404538 224244 404544 224256
rect 394568 224216 404544 224244
rect 394568 224204 394574 224216
rect 404538 224204 404544 224216
rect 404596 224204 404602 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 420822 224204 420828 224256
rect 420880 224244 420886 224256
rect 425146 224244 425152 224256
rect 420880 224216 425152 224244
rect 420880 224204 420886 224216
rect 425146 224204 425152 224216
rect 425204 224204 425210 224256
rect 436278 224204 436284 224256
rect 436336 224244 436342 224256
rect 437014 224244 437020 224256
rect 436336 224216 437020 224244
rect 436336 224204 436342 224216
rect 437014 224204 437020 224216
rect 437072 224204 437078 224256
rect 469582 224204 469588 224256
rect 469640 224244 469646 224256
rect 477586 224244 477592 224256
rect 469640 224216 477592 224244
rect 469640 224204 469646 224216
rect 477586 224204 477592 224216
rect 477644 224204 477650 224256
rect 488902 224204 488908 224256
rect 488960 224244 488966 224256
rect 502978 224244 502984 224256
rect 488960 224216 502984 224244
rect 488960 224204 488966 224216
rect 502978 224204 502984 224216
rect 503036 224204 503042 224256
rect 504358 224204 504364 224256
rect 504416 224244 504422 224256
rect 523494 224244 523500 224256
rect 504416 224216 523500 224244
rect 504416 224204 504422 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 533706 224204 533712 224256
rect 533764 224244 533770 224256
rect 561306 224244 561312 224256
rect 533764 224216 561312 224244
rect 533764 224204 533770 224216
rect 561306 224204 561312 224216
rect 561364 224204 561370 224256
rect 670930 224188 670982 224194
rect 563698 224136 563704 224188
rect 563756 224176 563762 224188
rect 568942 224176 568948 224188
rect 563756 224148 568948 224176
rect 563756 224136 563762 224148
rect 568942 224136 568948 224148
rect 569000 224136 569006 224188
rect 606294 224136 606300 224188
rect 606352 224176 606358 224188
rect 606352 224148 611354 224176
rect 606352 224136 606358 224148
rect 115842 224068 115848 224120
rect 115900 224108 115906 224120
rect 188798 224108 188804 224120
rect 115900 224080 188804 224108
rect 115900 224068 115906 224080
rect 188798 224068 188804 224080
rect 188856 224068 188862 224120
rect 189902 224068 189908 224120
rect 189960 224108 189966 224120
rect 212626 224108 212632 224120
rect 189960 224080 212632 224108
rect 189960 224068 189966 224080
rect 212626 224068 212632 224080
rect 212684 224068 212690 224120
rect 216582 224068 216588 224120
rect 216640 224108 216646 224120
rect 264422 224108 264428 224120
rect 216640 224080 264428 224108
rect 216640 224068 216646 224080
rect 264422 224068 264428 224080
rect 264480 224068 264486 224120
rect 275830 224068 275836 224120
rect 275888 224108 275894 224120
rect 288710 224108 288716 224120
rect 275888 224080 288716 224108
rect 275888 224068 275894 224080
rect 288710 224068 288716 224080
rect 288768 224068 288774 224120
rect 415026 224000 415032 224052
rect 415084 224040 415090 224052
rect 419626 224040 419632 224052
rect 415084 224012 419632 224040
rect 415084 224000 415090 224012
rect 419626 224000 419632 224012
rect 419684 224000 419690 224052
rect 489914 224000 489920 224052
rect 489972 224040 489978 224052
rect 491110 224040 491116 224052
rect 489972 224012 491116 224040
rect 489972 224000 489978 224012
rect 491110 224000 491116 224012
rect 491168 224000 491174 224052
rect 535638 224000 535644 224052
rect 535696 224040 535702 224052
rect 536650 224040 536656 224052
rect 535696 224012 536656 224040
rect 535696 224000 535702 224012
rect 536650 224000 536656 224012
rect 536708 224000 536714 224052
rect 567838 224000 567844 224052
rect 567896 224040 567902 224052
rect 611326 224040 611354 224148
rect 670930 224130 670982 224136
rect 616874 224040 616880 224052
rect 567896 224012 606616 224040
rect 611326 224012 616880 224040
rect 567896 224000 567902 224012
rect 122558 223932 122564 223984
rect 122616 223972 122622 223984
rect 193950 223972 193956 223984
rect 122616 223944 193956 223972
rect 122616 223932 122622 223944
rect 193950 223932 193956 223944
rect 194008 223932 194014 223984
rect 200758 223932 200764 223984
rect 200816 223972 200822 223984
rect 222930 223972 222936 223984
rect 200816 223944 222936 223972
rect 200816 223932 200822 223944
rect 222930 223932 222936 223944
rect 222988 223932 222994 223984
rect 226150 223932 226156 223984
rect 226208 223972 226214 223984
rect 272518 223972 272524 223984
rect 226208 223944 272524 223972
rect 226208 223932 226214 223944
rect 272518 223932 272524 223944
rect 272576 223932 272582 223984
rect 289078 223864 289084 223916
rect 289136 223904 289142 223916
rect 294782 223904 294788 223916
rect 289136 223876 294788 223904
rect 289136 223864 289142 223876
rect 294782 223864 294788 223876
rect 294840 223864 294846 223916
rect 512454 223864 512460 223916
rect 512512 223904 512518 223916
rect 606294 223904 606300 223916
rect 512512 223876 606300 223904
rect 512512 223864 512518 223876
rect 606294 223864 606300 223876
rect 606352 223864 606358 223916
rect 606588 223904 606616 224012
rect 616874 224000 616880 224012
rect 616932 224000 616938 224052
rect 630950 223904 630956 223916
rect 606588 223876 630956 223904
rect 630950 223864 630956 223876
rect 631008 223864 631014 223916
rect 139946 223796 139952 223848
rect 140004 223836 140010 223848
rect 171410 223836 171416 223848
rect 140004 223808 171416 223836
rect 140004 223796 140010 223808
rect 171410 223796 171416 223808
rect 171468 223796 171474 223848
rect 174906 223796 174912 223848
rect 174964 223836 174970 223848
rect 235166 223836 235172 223848
rect 174964 223808 235172 223836
rect 174964 223796 174970 223808
rect 235166 223796 235172 223808
rect 235224 223796 235230 223848
rect 496814 223728 496820 223780
rect 496872 223768 496878 223780
rect 497366 223768 497372 223780
rect 496872 223740 497372 223768
rect 496872 223728 496878 223740
rect 497366 223728 497372 223740
rect 497424 223768 497430 223780
rect 567838 223768 567844 223780
rect 497424 223740 567844 223768
rect 497424 223728 497430 223740
rect 567838 223728 567844 223740
rect 567896 223728 567902 223780
rect 568574 223728 568580 223780
rect 568632 223768 568638 223780
rect 627914 223768 627920 223780
rect 568632 223740 627920 223768
rect 568632 223728 568638 223740
rect 627914 223728 627920 223740
rect 627972 223728 627978 223780
rect 185578 223660 185584 223712
rect 185636 223700 185642 223712
rect 191006 223700 191012 223712
rect 185636 223672 191012 223700
rect 185636 223660 185642 223672
rect 191006 223660 191012 223672
rect 191064 223660 191070 223712
rect 227622 223660 227628 223712
rect 227680 223700 227686 223712
rect 273162 223700 273168 223712
rect 227680 223672 273168 223700
rect 227680 223660 227686 223672
rect 273162 223660 273168 223672
rect 273220 223660 273226 223712
rect 491110 223592 491116 223644
rect 491168 223632 491174 223644
rect 629846 223632 629852 223644
rect 491168 223604 629852 223632
rect 491168 223592 491174 223604
rect 629846 223592 629852 223604
rect 629904 223592 629910 223644
rect 654962 223592 654968 223644
rect 655020 223632 655026 223644
rect 655606 223632 655612 223644
rect 655020 223604 655612 223632
rect 655020 223592 655026 223604
rect 655606 223592 655612 223604
rect 655664 223592 655670 223644
rect 87966 223524 87972 223576
rect 88024 223564 88030 223576
rect 164970 223564 164976 223576
rect 88024 223536 164976 223564
rect 88024 223524 88030 223536
rect 164970 223524 164976 223536
rect 165028 223524 165034 223576
rect 166442 223524 166448 223576
rect 166500 223564 166506 223576
rect 192018 223564 192024 223576
rect 166500 223536 192024 223564
rect 166500 223524 166506 223536
rect 192018 223524 192024 223536
rect 192076 223524 192082 223576
rect 194502 223524 194508 223576
rect 194560 223564 194566 223576
rect 247402 223564 247408 223576
rect 194560 223536 247408 223564
rect 194560 223524 194566 223536
rect 247402 223524 247408 223536
rect 247460 223524 247466 223576
rect 253566 223524 253572 223576
rect 253624 223564 253630 223576
rect 293494 223564 293500 223576
rect 253624 223536 293500 223564
rect 253624 223524 253630 223536
rect 293494 223524 293500 223536
rect 293552 223524 293558 223576
rect 307018 223524 307024 223576
rect 307076 223564 307082 223576
rect 315666 223564 315672 223576
rect 307076 223536 315672 223564
rect 307076 223524 307082 223536
rect 315666 223524 315672 223536
rect 315724 223524 315730 223576
rect 416498 223524 416504 223576
rect 416556 223564 416562 223576
rect 422202 223564 422208 223576
rect 416556 223536 422208 223564
rect 416556 223524 416562 223536
rect 422202 223524 422208 223536
rect 422260 223524 422266 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 102042 223388 102048 223440
rect 102100 223428 102106 223440
rect 178494 223428 178500 223440
rect 102100 223400 178500 223428
rect 102100 223388 102106 223400
rect 178494 223388 178500 223400
rect 178552 223388 178558 223440
rect 197262 223388 197268 223440
rect 197320 223428 197326 223440
rect 249978 223428 249984 223440
rect 197320 223400 249984 223428
rect 197320 223388 197326 223400
rect 249978 223388 249984 223400
rect 250036 223388 250042 223440
rect 267550 223388 267556 223440
rect 267608 223428 267614 223440
rect 307294 223428 307300 223440
rect 267608 223400 307300 223428
rect 267608 223388 267614 223400
rect 307294 223388 307300 223400
rect 307352 223388 307358 223440
rect 322842 223388 322848 223440
rect 322900 223428 322906 223440
rect 332410 223428 332416 223440
rect 322900 223400 332416 223428
rect 322900 223388 322906 223400
rect 332410 223388 332416 223400
rect 332468 223388 332474 223440
rect 520274 223388 520280 223440
rect 520332 223428 520338 223440
rect 539962 223428 539968 223440
rect 520332 223400 539968 223428
rect 520332 223388 520338 223400
rect 539962 223388 539968 223400
rect 540020 223388 540026 223440
rect 78582 223252 78588 223304
rect 78640 223292 78646 223304
rect 157242 223292 157248 223304
rect 78640 223264 157248 223292
rect 78640 223252 78646 223264
rect 157242 223252 157248 223264
rect 157300 223252 157306 223304
rect 159358 223252 159364 223304
rect 159416 223292 159422 223304
rect 181714 223292 181720 223304
rect 159416 223264 181720 223292
rect 159416 223252 159422 223264
rect 181714 223252 181720 223264
rect 181772 223252 181778 223304
rect 191650 223252 191656 223304
rect 191708 223292 191714 223304
rect 244826 223292 244832 223304
rect 191708 223264 244832 223292
rect 191708 223252 191714 223264
rect 244826 223252 244832 223264
rect 244884 223252 244890 223304
rect 261846 223252 261852 223304
rect 261904 223292 261910 223304
rect 300854 223292 300860 223304
rect 261904 223264 300860 223292
rect 261904 223252 261910 223264
rect 300854 223252 300860 223264
rect 300912 223252 300918 223304
rect 315850 223252 315856 223304
rect 315908 223292 315914 223304
rect 341426 223292 341432 223304
rect 315908 223264 341432 223292
rect 315908 223252 315914 223264
rect 341426 223252 341432 223264
rect 341484 223252 341490 223304
rect 342162 223252 342168 223304
rect 342220 223292 342226 223304
rect 362034 223292 362040 223304
rect 342220 223264 362040 223292
rect 342220 223252 342226 223264
rect 362034 223252 362040 223264
rect 362092 223252 362098 223304
rect 366726 223252 366732 223304
rect 366784 223292 366790 223304
rect 381998 223292 382004 223304
rect 366784 223264 382004 223292
rect 366784 223252 366790 223264
rect 381998 223252 382004 223264
rect 382056 223252 382062 223304
rect 406746 223252 406752 223304
rect 406804 223292 406810 223304
rect 414842 223292 414848 223304
rect 406804 223264 414848 223292
rect 406804 223252 406810 223264
rect 414842 223252 414848 223264
rect 414900 223252 414906 223304
rect 513098 223252 513104 223304
rect 513156 223292 513162 223304
rect 534534 223292 534540 223304
rect 513156 223264 534540 223292
rect 513156 223252 513162 223264
rect 534534 223252 534540 223264
rect 534592 223252 534598 223304
rect 541250 223252 541256 223304
rect 541308 223292 541314 223304
rect 554866 223292 554872 223304
rect 541308 223264 554872 223292
rect 541308 223252 541314 223264
rect 554866 223252 554872 223264
rect 554924 223252 554930 223304
rect 81158 223116 81164 223168
rect 81216 223156 81222 223168
rect 159818 223156 159824 223168
rect 81216 223128 159824 223156
rect 81216 223116 81222 223128
rect 159818 223116 159824 223128
rect 159876 223116 159882 223168
rect 168282 223116 168288 223168
rect 168340 223156 168346 223168
rect 226794 223156 226800 223168
rect 168340 223128 226800 223156
rect 168340 223116 168346 223128
rect 226794 223116 226800 223128
rect 226852 223116 226858 223168
rect 248230 223116 248236 223168
rect 248288 223156 248294 223168
rect 291838 223156 291844 223168
rect 248288 223128 291844 223156
rect 248288 223116 248294 223128
rect 291838 223116 291844 223128
rect 291896 223116 291902 223168
rect 300762 223116 300768 223168
rect 300820 223156 300826 223168
rect 330110 223156 330116 223168
rect 300820 223128 330116 223156
rect 300820 223116 300826 223128
rect 330110 223116 330116 223128
rect 330168 223116 330174 223168
rect 336366 223116 336372 223168
rect 336424 223156 336430 223168
rect 359734 223156 359740 223168
rect 336424 223128 359740 223156
rect 336424 223116 336430 223128
rect 359734 223116 359740 223128
rect 359792 223116 359798 223168
rect 366910 223116 366916 223168
rect 366968 223156 366974 223168
rect 383930 223156 383936 223168
rect 366968 223128 383936 223156
rect 366968 223116 366974 223128
rect 383930 223116 383936 223128
rect 383988 223116 383994 223168
rect 477954 223116 477960 223168
rect 478012 223156 478018 223168
rect 489454 223156 489460 223168
rect 478012 223128 489460 223156
rect 478012 223116 478018 223128
rect 489454 223116 489460 223128
rect 489512 223116 489518 223168
rect 496630 223116 496636 223168
rect 496688 223156 496694 223168
rect 513558 223156 513564 223168
rect 496688 223128 513564 223156
rect 496688 223116 496694 223128
rect 513558 223116 513564 223128
rect 513616 223116 513622 223168
rect 519814 223116 519820 223168
rect 519872 223156 519878 223168
rect 542354 223156 542360 223168
rect 519872 223128 542360 223156
rect 519872 223116 519878 223128
rect 542354 223116 542360 223128
rect 542412 223116 542418 223168
rect 552198 223116 552204 223168
rect 552256 223156 552262 223168
rect 561674 223156 561680 223168
rect 552256 223128 561680 223156
rect 552256 223116 552262 223128
rect 561674 223116 561680 223128
rect 561732 223116 561738 223168
rect 75822 222980 75828 223032
rect 75880 223020 75886 223032
rect 154666 223020 154672 223032
rect 75880 222992 154672 223020
rect 75880 222980 75886 222992
rect 154666 222980 154672 222992
rect 154724 222980 154730 223032
rect 164050 222980 164056 223032
rect 164108 223020 164114 223032
rect 224218 223020 224224 223032
rect 164108 222992 224224 223020
rect 164108 222980 164114 222992
rect 224218 222980 224224 222992
rect 224276 222980 224282 223032
rect 238662 222980 238668 223032
rect 238720 223020 238726 223032
rect 282822 223020 282828 223032
rect 238720 222992 282828 223020
rect 238720 222980 238726 222992
rect 282822 222980 282828 222992
rect 282880 222980 282886 223032
rect 292482 222980 292488 223032
rect 292540 223020 292546 223032
rect 326614 223020 326620 223032
rect 292540 222992 326620 223020
rect 292540 222980 292546 222992
rect 326614 222980 326620 222992
rect 326672 222980 326678 223032
rect 329742 222980 329748 223032
rect 329800 223020 329806 223032
rect 353662 223020 353668 223032
rect 329800 222992 353668 223020
rect 329800 222980 329806 222992
rect 353662 222980 353668 222992
rect 353720 222980 353726 223032
rect 355962 222980 355968 223032
rect 356020 223020 356026 223032
rect 375558 223020 375564 223032
rect 356020 222992 375564 223020
rect 356020 222980 356026 222992
rect 375558 222980 375564 222992
rect 375616 222980 375622 223032
rect 382090 222980 382096 223032
rect 382148 223020 382154 223032
rect 392946 223020 392952 223032
rect 382148 222992 392952 223020
rect 382148 222980 382154 222992
rect 392946 222980 392952 222992
rect 393004 222980 393010 223032
rect 483106 222980 483112 223032
rect 483164 223020 483170 223032
rect 496078 223020 496084 223032
rect 483164 222992 496084 223020
rect 483164 222980 483170 222992
rect 496078 222980 496084 222992
rect 496136 222980 496142 223032
rect 502426 222980 502432 223032
rect 502484 223020 502490 223032
rect 521010 223020 521016 223032
rect 502484 222992 521016 223020
rect 502484 222980 502490 222992
rect 521010 222980 521016 222992
rect 521068 222980 521074 223032
rect 527542 222980 527548 223032
rect 527600 223020 527606 223032
rect 553302 223020 553308 223032
rect 527600 222992 553308 223020
rect 527600 222980 527606 222992
rect 553302 222980 553308 222992
rect 553360 222980 553366 223032
rect 68922 222844 68928 222896
rect 68980 222884 68986 222896
rect 149514 222884 149520 222896
rect 68980 222856 149520 222884
rect 68980 222844 68986 222856
rect 149514 222844 149520 222856
rect 149572 222844 149578 222896
rect 154206 222844 154212 222896
rect 154264 222884 154270 222896
rect 216214 222884 216220 222896
rect 154264 222856 216220 222884
rect 154264 222844 154270 222856
rect 216214 222844 216220 222856
rect 216272 222844 216278 222896
rect 217870 222844 217876 222896
rect 217928 222884 217934 222896
rect 268654 222884 268660 222896
rect 217928 222856 268660 222884
rect 217928 222844 217934 222856
rect 268654 222844 268660 222856
rect 268712 222844 268718 222896
rect 278406 222844 278412 222896
rect 278464 222884 278470 222896
rect 313734 222884 313740 222896
rect 278464 222856 313740 222884
rect 278464 222844 278470 222856
rect 313734 222844 313740 222856
rect 313792 222844 313798 222896
rect 315666 222844 315672 222896
rect 315724 222884 315730 222896
rect 344646 222884 344652 222896
rect 315724 222856 344652 222884
rect 315724 222844 315730 222856
rect 344646 222844 344652 222856
rect 344704 222844 344710 222896
rect 346302 222844 346308 222896
rect 346360 222884 346366 222896
rect 367462 222884 367468 222896
rect 346360 222856 367468 222884
rect 346360 222844 346366 222856
rect 367462 222844 367468 222856
rect 367520 222844 367526 222896
rect 386322 222844 386328 222896
rect 386380 222884 386386 222896
rect 398282 222884 398288 222896
rect 386380 222856 398288 222884
rect 386380 222844 386386 222856
rect 398282 222844 398288 222856
rect 398340 222844 398346 222896
rect 398466 222844 398472 222896
rect 398524 222884 398530 222896
rect 405826 222884 405832 222896
rect 398524 222856 405832 222884
rect 398524 222844 398530 222856
rect 405826 222844 405832 222856
rect 405884 222844 405890 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467282 222844 467288 222896
rect 467340 222884 467346 222896
rect 475378 222884 475384 222896
rect 467340 222856 475384 222884
rect 467340 222844 467346 222856
rect 475378 222844 475384 222856
rect 475436 222844 475442 222896
rect 476666 222844 476672 222896
rect 476724 222884 476730 222896
rect 487798 222884 487804 222896
rect 476724 222856 487804 222884
rect 476724 222844 476730 222856
rect 487798 222844 487804 222856
rect 487856 222844 487862 222896
rect 488258 222844 488264 222896
rect 488316 222884 488322 222896
rect 503162 222884 503168 222896
rect 488316 222856 503168 222884
rect 488316 222844 488322 222856
rect 503162 222844 503168 222856
rect 503220 222844 503226 222896
rect 507578 222844 507584 222896
rect 507636 222884 507642 222896
rect 527542 222884 527548 222896
rect 507636 222856 527548 222884
rect 507636 222844 507642 222856
rect 527542 222844 527548 222856
rect 527600 222844 527606 222896
rect 532418 222844 532424 222896
rect 532476 222884 532482 222896
rect 559006 222884 559012 222896
rect 532476 222856 559012 222884
rect 532476 222844 532482 222856
rect 559006 222844 559012 222856
rect 559064 222844 559070 222896
rect 559558 222844 559564 222896
rect 559616 222884 559622 222896
rect 633710 222884 633716 222896
rect 559616 222856 633716 222884
rect 559616 222844 559622 222856
rect 633710 222844 633716 222856
rect 633768 222844 633774 222896
rect 131022 222708 131028 222760
rect 131080 222748 131086 222760
rect 196066 222748 196072 222760
rect 131080 222720 196072 222748
rect 131080 222708 131086 222720
rect 196066 222708 196072 222720
rect 196124 222708 196130 222760
rect 208026 222708 208032 222760
rect 208084 222748 208090 222760
rect 260926 222748 260932 222760
rect 208084 222720 260932 222748
rect 208084 222708 208090 222720
rect 260926 222708 260932 222720
rect 260984 222708 260990 222760
rect 290826 222708 290832 222760
rect 290884 222748 290890 222760
rect 321830 222748 321836 222760
rect 290884 222720 321836 222748
rect 290884 222708 290890 222720
rect 321830 222708 321836 222720
rect 321888 222708 321894 222760
rect 503346 222708 503352 222760
rect 503404 222748 503410 222760
rect 521838 222748 521844 222760
rect 503404 222720 521844 222748
rect 503404 222708 503410 222720
rect 521838 222708 521844 222720
rect 521896 222708 521902 222760
rect 558638 222708 558644 222760
rect 558696 222748 558702 222760
rect 568758 222748 568764 222760
rect 558696 222720 568764 222748
rect 558696 222708 558702 222720
rect 568758 222708 568764 222720
rect 568816 222708 568822 222760
rect 146110 222572 146116 222624
rect 146168 222612 146174 222624
rect 211982 222612 211988 222624
rect 146168 222584 211988 222612
rect 146168 222572 146174 222584
rect 211982 222572 211988 222584
rect 212040 222572 212046 222624
rect 213822 222572 213828 222624
rect 213880 222612 213886 222624
rect 262858 222612 262864 222624
rect 213880 222584 262864 222612
rect 213880 222572 213886 222584
rect 262858 222572 262864 222584
rect 262916 222572 262922 222624
rect 561674 222572 561680 222624
rect 561732 222612 561738 222624
rect 562134 222612 562140 222624
rect 561732 222584 562140 222612
rect 561732 222572 561738 222584
rect 562134 222572 562140 222584
rect 562192 222612 562198 222624
rect 563146 222612 563152 222624
rect 562192 222584 563152 222612
rect 562192 222572 562198 222584
rect 563146 222572 563152 222584
rect 563204 222572 563210 222624
rect 565446 222572 565452 222624
rect 565504 222612 565510 222624
rect 567102 222612 567108 222624
rect 565504 222584 567108 222612
rect 565504 222572 565510 222584
rect 567102 222572 567108 222584
rect 567160 222572 567166 222624
rect 567654 222572 567660 222624
rect 567712 222612 567718 222624
rect 571610 222612 571616 222624
rect 567712 222584 571616 222612
rect 567712 222572 567718 222584
rect 571610 222572 571616 222584
rect 571668 222572 571674 222624
rect 134978 222436 134984 222488
rect 135036 222476 135042 222488
rect 197446 222476 197452 222488
rect 135036 222448 197452 222476
rect 135036 222436 135042 222448
rect 197446 222436 197452 222448
rect 197504 222436 197510 222488
rect 203886 222436 203892 222488
rect 203944 222476 203950 222488
rect 254854 222476 254860 222488
rect 203944 222448 254860 222476
rect 203944 222436 203950 222448
rect 254854 222436 254860 222448
rect 254912 222436 254918 222488
rect 482922 222436 482928 222488
rect 482980 222476 482986 222488
rect 593966 222476 593972 222488
rect 482980 222448 593972 222476
rect 482980 222436 482986 222448
rect 593966 222436 593972 222448
rect 594024 222436 594030 222488
rect 244090 222300 244096 222352
rect 244148 222340 244154 222352
rect 286042 222340 286048 222352
rect 244148 222312 286048 222340
rect 244148 222300 244154 222312
rect 286042 222300 286048 222312
rect 286100 222300 286106 222352
rect 556062 222300 556068 222352
rect 556120 222340 556126 222352
rect 557350 222340 557356 222352
rect 556120 222312 557356 222340
rect 556120 222300 556126 222312
rect 557350 222300 557356 222312
rect 557408 222340 557414 222352
rect 626534 222340 626540 222352
rect 557408 222312 626540 222340
rect 557408 222300 557414 222312
rect 626534 222300 626540 222312
rect 626592 222300 626598 222352
rect 553366 222244 553532 222272
rect 550818 222164 550824 222216
rect 550876 222204 550882 222216
rect 553366 222204 553394 222244
rect 550876 222176 553394 222204
rect 550876 222164 550882 222176
rect 111150 222096 111156 222148
rect 111208 222136 111214 222148
rect 182542 222136 182548 222148
rect 111208 222108 182548 222136
rect 111208 222096 111214 222108
rect 182542 222096 182548 222108
rect 182600 222096 182606 222148
rect 184014 222096 184020 222148
rect 184072 222136 184078 222148
rect 239214 222136 239220 222148
rect 184072 222108 239220 222136
rect 184072 222096 184078 222108
rect 239214 222096 239220 222108
rect 239272 222096 239278 222148
rect 282638 222096 282644 222148
rect 282696 222136 282702 222148
rect 283558 222136 283564 222148
rect 282696 222108 283564 222136
rect 282696 222096 282702 222108
rect 283558 222096 283564 222108
rect 283616 222096 283622 222148
rect 283742 222096 283748 222148
rect 283800 222136 283806 222148
rect 314838 222136 314844 222148
rect 283800 222108 314844 222136
rect 283800 222096 283806 222108
rect 314838 222096 314844 222108
rect 314896 222096 314902 222148
rect 386874 222096 386880 222148
rect 386932 222136 386938 222148
rect 389910 222136 389916 222148
rect 386932 222108 389916 222136
rect 386932 222096 386938 222108
rect 389910 222096 389916 222108
rect 389968 222096 389974 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468662 222136 468668 222148
rect 462188 222108 468668 222136
rect 462188 222096 462194 222108
rect 468662 222096 468668 222108
rect 468720 222096 468726 222148
rect 553504 222136 553532 222244
rect 563146 222164 563152 222216
rect 563204 222204 563210 222216
rect 628190 222204 628196 222216
rect 563204 222176 628196 222204
rect 563204 222164 563210 222176
rect 628190 222164 628196 222176
rect 628248 222164 628254 222216
rect 558362 222136 558368 222148
rect 553504 222108 558368 222136
rect 558362 222096 558368 222108
rect 558420 222096 558426 222148
rect 560754 222096 560760 222148
rect 560812 222136 560818 222148
rect 561306 222136 561312 222148
rect 560812 222108 561312 222136
rect 560812 222096 560818 222108
rect 561306 222096 561312 222108
rect 561364 222136 561370 222148
rect 563008 222136 563014 222148
rect 561364 222108 563014 222136
rect 561364 222096 561370 222108
rect 563008 222096 563014 222108
rect 563066 222096 563072 222148
rect 542998 222028 543004 222080
rect 543056 222068 543062 222080
rect 543056 222040 553394 222068
rect 543056 222028 543062 222040
rect 104526 221960 104532 222012
rect 104584 222000 104590 222012
rect 177390 222000 177396 222012
rect 104584 221972 177396 222000
rect 104584 221960 104590 221972
rect 177390 221960 177396 221972
rect 177448 221960 177454 222012
rect 194778 221960 194784 222012
rect 194836 222000 194842 222012
rect 250162 222000 250168 222012
rect 194836 221972 250168 222000
rect 194836 221960 194842 221972
rect 250162 221960 250168 221972
rect 250220 221960 250226 222012
rect 258074 221960 258080 222012
rect 258132 222000 258138 222012
rect 269206 222000 269212 222012
rect 258132 221972 269212 222000
rect 258132 221960 258138 221972
rect 269206 221960 269212 221972
rect 269264 221960 269270 222012
rect 270034 221960 270040 222012
rect 270092 222000 270098 222012
rect 306558 222000 306564 222012
rect 270092 221972 306564 222000
rect 270092 221960 270098 221972
rect 306558 221960 306564 221972
rect 306616 221960 306622 222012
rect 330570 221960 330576 222012
rect 330628 222000 330634 222012
rect 345658 222000 345664 222012
rect 330628 221972 345664 222000
rect 330628 221960 330634 221972
rect 345658 221960 345664 221972
rect 345716 221960 345722 222012
rect 553366 222000 553394 222040
rect 556062 222000 556068 222012
rect 553366 221972 556068 222000
rect 556062 221960 556068 221972
rect 556120 221960 556126 222012
rect 556246 221960 556252 222012
rect 556304 222000 556310 222012
rect 559558 222000 559564 222012
rect 556304 221972 559564 222000
rect 556304 221960 556310 221972
rect 559558 221960 559564 221972
rect 559616 221960 559622 222012
rect 562318 221960 562324 222012
rect 562376 222000 562382 222012
rect 571426 222000 571432 222012
rect 562376 221972 571432 222000
rect 562376 221960 562382 221972
rect 571426 221960 571432 221972
rect 571484 221960 571490 222012
rect 571610 221960 571616 222012
rect 571668 222000 571674 222012
rect 577682 222000 577688 222012
rect 571668 221972 577688 222000
rect 571668 221960 571674 221972
rect 577682 221960 577688 221972
rect 577740 221960 577746 222012
rect 596266 221960 596272 222012
rect 596324 222000 596330 222012
rect 597002 222000 597008 222012
rect 596324 221972 597008 222000
rect 596324 221960 596330 221972
rect 597002 221960 597008 221972
rect 597060 221960 597066 222012
rect 101214 221824 101220 221876
rect 101272 221864 101278 221876
rect 175458 221864 175464 221876
rect 101272 221836 175464 221864
rect 101272 221824 101278 221836
rect 175458 221824 175464 221836
rect 175516 221824 175522 221876
rect 189166 221824 189172 221876
rect 189224 221864 189230 221876
rect 245010 221864 245016 221876
rect 189224 221836 245016 221864
rect 189224 221824 189230 221836
rect 245010 221824 245016 221836
rect 245068 221824 245074 221876
rect 252554 221824 252560 221876
rect 252612 221864 252618 221876
rect 258626 221864 258632 221876
rect 252612 221836 258632 221864
rect 252612 221824 252618 221836
rect 258626 221824 258632 221836
rect 258684 221824 258690 221876
rect 266814 221824 266820 221876
rect 266872 221864 266878 221876
rect 297174 221864 297180 221876
rect 266872 221836 297180 221864
rect 266872 221824 266878 221836
rect 297174 221824 297180 221836
rect 297232 221824 297238 221876
rect 298554 221864 298560 221876
rect 297652 221836 298560 221864
rect 60642 221688 60648 221740
rect 60700 221728 60706 221740
rect 94406 221728 94412 221740
rect 60700 221700 94412 221728
rect 60700 221688 60706 221700
rect 94406 221688 94412 221700
rect 94464 221688 94470 221740
rect 94590 221688 94596 221740
rect 94648 221728 94654 221740
rect 169754 221728 169760 221740
rect 94648 221700 169760 221728
rect 94648 221688 94654 221700
rect 169754 221688 169760 221700
rect 169812 221688 169818 221740
rect 177390 221688 177396 221740
rect 177448 221728 177454 221740
rect 234154 221728 234160 221740
rect 177448 221700 234160 221728
rect 177448 221688 177454 221700
rect 234154 221688 234160 221700
rect 234212 221688 234218 221740
rect 247126 221688 247132 221740
rect 247184 221728 247190 221740
rect 253382 221728 253388 221740
rect 247184 221700 253388 221728
rect 247184 221688 247190 221700
rect 253382 221688 253388 221700
rect 253440 221688 253446 221740
rect 260190 221688 260196 221740
rect 260248 221728 260254 221740
rect 297652 221728 297680 221836
rect 298554 221824 298560 221836
rect 298612 221824 298618 221876
rect 306558 221824 306564 221876
rect 306616 221864 306622 221876
rect 335446 221864 335452 221876
rect 306616 221836 335452 221864
rect 306616 221824 306622 221836
rect 335446 221824 335452 221836
rect 335504 221824 335510 221876
rect 344646 221824 344652 221876
rect 344704 221864 344710 221876
rect 364518 221864 364524 221876
rect 344704 221836 364524 221864
rect 344704 221824 344710 221836
rect 364518 221824 364524 221836
rect 364576 221824 364582 221876
rect 512638 221824 512644 221876
rect 512696 221864 512702 221876
rect 522574 221864 522580 221876
rect 512696 221836 522580 221864
rect 512696 221824 512702 221836
rect 522574 221824 522580 221836
rect 522632 221824 522638 221876
rect 525150 221824 525156 221876
rect 525208 221864 525214 221876
rect 537478 221864 537484 221876
rect 525208 221836 537484 221864
rect 525208 221824 525214 221836
rect 537478 221824 537484 221836
rect 537536 221824 537542 221876
rect 547138 221824 547144 221876
rect 547196 221864 547202 221876
rect 559834 221864 559840 221876
rect 547196 221836 559840 221864
rect 547196 221824 547202 221836
rect 559834 221824 559840 221836
rect 559892 221824 559898 221876
rect 562778 221824 562784 221876
rect 562836 221864 562842 221876
rect 610526 221864 610532 221876
rect 562836 221836 610532 221864
rect 562836 221824 562842 221836
rect 610526 221824 610532 221836
rect 610584 221824 610590 221876
rect 260248 221700 297680 221728
rect 260248 221688 260254 221700
rect 298278 221688 298284 221740
rect 298336 221728 298342 221740
rect 328546 221728 328552 221740
rect 298336 221700 328552 221728
rect 298336 221688 298342 221700
rect 328546 221688 328552 221700
rect 328604 221688 328610 221740
rect 331398 221688 331404 221740
rect 331456 221728 331462 221740
rect 353846 221728 353852 221740
rect 331456 221700 353852 221728
rect 331456 221688 331462 221700
rect 353846 221688 353852 221700
rect 353904 221688 353910 221740
rect 362034 221688 362040 221740
rect 362092 221728 362098 221740
rect 376018 221728 376024 221740
rect 362092 221700 376024 221728
rect 362092 221688 362098 221700
rect 376018 221688 376024 221700
rect 376076 221688 376082 221740
rect 382734 221728 382740 221740
rect 378428 221700 382740 221728
rect 73890 221552 73896 221604
rect 73948 221592 73954 221604
rect 86218 221592 86224 221604
rect 73948 221564 86224 221592
rect 73948 221552 73954 221564
rect 86218 221552 86224 221564
rect 86276 221552 86282 221604
rect 91278 221552 91284 221604
rect 91336 221592 91342 221604
rect 167086 221592 167092 221604
rect 91336 221564 167092 221592
rect 91336 221552 91342 221564
rect 167086 221552 167092 221564
rect 167144 221552 167150 221604
rect 178218 221552 178224 221604
rect 178276 221592 178282 221604
rect 237374 221592 237380 221604
rect 178276 221564 237380 221592
rect 178276 221552 178282 221564
rect 237374 221552 237380 221564
rect 237432 221552 237438 221604
rect 238846 221552 238852 221604
rect 238904 221592 238910 221604
rect 248598 221592 248604 221604
rect 238904 221564 248604 221592
rect 238904 221552 238910 221564
rect 248598 221552 248604 221564
rect 248656 221552 248662 221604
rect 250254 221552 250260 221604
rect 250312 221592 250318 221604
rect 291378 221592 291384 221604
rect 250312 221564 291384 221592
rect 250312 221552 250318 221564
rect 291378 221552 291384 221564
rect 291436 221552 291442 221604
rect 327534 221592 327540 221604
rect 296686 221564 327540 221592
rect 84654 221416 84660 221468
rect 84712 221456 84718 221468
rect 161474 221456 161480 221468
rect 84712 221428 161480 221456
rect 84712 221416 84718 221428
rect 161474 221416 161480 221428
rect 161532 221416 161538 221468
rect 161658 221416 161664 221468
rect 161716 221456 161722 221468
rect 224402 221456 224408 221468
rect 161716 221428 224408 221456
rect 161716 221416 161722 221428
rect 224402 221416 224408 221428
rect 224460 221416 224466 221468
rect 234338 221416 234344 221468
rect 234396 221456 234402 221468
rect 234396 221428 277394 221456
rect 234396 221416 234402 221428
rect 121086 221280 121092 221332
rect 121144 221320 121150 221332
rect 190638 221320 190644 221332
rect 121144 221292 190644 221320
rect 121144 221280 121150 221292
rect 190638 221280 190644 221292
rect 190696 221280 190702 221332
rect 201402 221280 201408 221332
rect 201460 221320 201466 221332
rect 255406 221320 255412 221332
rect 201460 221292 255412 221320
rect 201460 221280 201466 221292
rect 255406 221280 255412 221292
rect 255464 221280 255470 221332
rect 277366 221320 277394 221428
rect 277578 221416 277584 221468
rect 277636 221456 277642 221468
rect 283742 221456 283748 221468
rect 277636 221428 283748 221456
rect 277636 221416 277642 221428
rect 283742 221416 283748 221428
rect 283800 221416 283806 221468
rect 284018 221416 284024 221468
rect 284076 221456 284082 221468
rect 289906 221456 289912 221468
rect 284076 221428 289912 221456
rect 284076 221416 284082 221428
rect 289906 221416 289912 221428
rect 289964 221416 289970 221468
rect 296438 221416 296444 221468
rect 296496 221456 296502 221468
rect 296686 221456 296714 221564
rect 327534 221552 327540 221564
rect 327592 221552 327598 221604
rect 328086 221552 328092 221604
rect 328144 221592 328150 221604
rect 351270 221592 351276 221604
rect 328144 221564 351276 221592
rect 328144 221552 328150 221564
rect 351270 221552 351276 221564
rect 351328 221552 351334 221604
rect 353294 221552 353300 221604
rect 353352 221592 353358 221604
rect 369946 221592 369952 221604
rect 353352 221564 369952 221592
rect 353352 221552 353358 221564
rect 369946 221552 369952 221564
rect 370004 221552 370010 221604
rect 370498 221552 370504 221604
rect 370556 221592 370562 221604
rect 378428 221592 378456 221700
rect 382734 221688 382740 221700
rect 382792 221688 382798 221740
rect 475746 221688 475752 221740
rect 475804 221728 475810 221740
rect 486142 221728 486148 221740
rect 475804 221700 486148 221728
rect 475804 221688 475810 221700
rect 486142 221688 486148 221700
rect 486200 221688 486206 221740
rect 487062 221688 487068 221740
rect 487120 221728 487126 221740
rect 500034 221728 500040 221740
rect 487120 221700 500040 221728
rect 487120 221688 487126 221700
rect 500034 221688 500040 221700
rect 500092 221688 500098 221740
rect 501598 221688 501604 221740
rect 501656 221728 501662 221740
rect 517698 221728 517704 221740
rect 501656 221700 517704 221728
rect 501656 221688 501662 221700
rect 517698 221688 517704 221700
rect 517756 221688 517762 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 546586 221728 546592 221740
rect 522908 221700 546592 221728
rect 522908 221688 522914 221700
rect 546586 221688 546592 221700
rect 546644 221688 546650 221740
rect 548334 221688 548340 221740
rect 548392 221728 548398 221740
rect 553026 221728 553032 221740
rect 548392 221700 553032 221728
rect 548392 221688 548398 221700
rect 553026 221688 553032 221700
rect 553084 221688 553090 221740
rect 553302 221688 553308 221740
rect 553360 221728 553366 221740
rect 608594 221728 608600 221740
rect 553360 221700 608600 221728
rect 553360 221688 553366 221700
rect 608594 221688 608600 221700
rect 608652 221688 608658 221740
rect 370556 221564 378456 221592
rect 370556 221552 370562 221564
rect 382734 221552 382740 221604
rect 382792 221592 382798 221604
rect 394878 221592 394884 221604
rect 382792 221564 394884 221592
rect 382792 221552 382798 221564
rect 394878 221552 394884 221564
rect 394936 221552 394942 221604
rect 396810 221552 396816 221604
rect 396868 221592 396874 221604
rect 407298 221592 407304 221604
rect 396868 221564 407304 221592
rect 396868 221552 396874 221564
rect 407298 221552 407304 221564
rect 407356 221552 407362 221604
rect 469030 221552 469036 221604
rect 469088 221592 469094 221604
rect 474550 221592 474556 221604
rect 469088 221564 474556 221592
rect 469088 221552 469094 221564
rect 474550 221552 474556 221564
rect 474608 221552 474614 221604
rect 485498 221552 485504 221604
rect 485556 221592 485562 221604
rect 499390 221592 499396 221604
rect 485556 221564 499396 221592
rect 485556 221552 485562 221564
rect 499390 221552 499396 221564
rect 499448 221552 499454 221604
rect 500218 221552 500224 221604
rect 500276 221592 500282 221604
rect 517514 221592 517520 221604
rect 500276 221564 517520 221592
rect 500276 221552 500282 221564
rect 517514 221552 517520 221564
rect 517572 221552 517578 221604
rect 518158 221552 518164 221604
rect 518216 221592 518222 221604
rect 530026 221592 530032 221604
rect 518216 221564 530032 221592
rect 518216 221552 518222 221564
rect 530026 221552 530032 221564
rect 530084 221552 530090 221604
rect 531222 221552 531228 221604
rect 531280 221592 531286 221604
rect 556522 221592 556528 221604
rect 531280 221564 556528 221592
rect 531280 221552 531286 221564
rect 556522 221552 556528 221564
rect 556580 221552 556586 221604
rect 556982 221552 556988 221604
rect 557040 221592 557046 221604
rect 564894 221592 564900 221604
rect 557040 221564 564900 221592
rect 557040 221552 557046 221564
rect 564894 221552 564900 221564
rect 564952 221592 564958 221604
rect 567654 221592 567660 221604
rect 564952 221564 567660 221592
rect 564952 221552 564958 221564
rect 567654 221552 567660 221564
rect 567712 221552 567718 221604
rect 567838 221552 567844 221604
rect 567896 221592 567902 221604
rect 596266 221592 596272 221604
rect 567896 221564 596272 221592
rect 567896 221552 567902 221564
rect 596266 221552 596272 221564
rect 596324 221552 596330 221604
rect 596450 221552 596456 221604
rect 596508 221592 596514 221604
rect 607306 221592 607312 221604
rect 596508 221564 607312 221592
rect 596508 221552 596514 221564
rect 607306 221552 607312 221564
rect 607364 221552 607370 221604
rect 296496 221428 296714 221456
rect 296496 221416 296502 221428
rect 297174 221416 297180 221468
rect 297232 221456 297238 221468
rect 297232 221428 300164 221456
rect 297232 221416 297238 221428
rect 281718 221320 281724 221332
rect 277366 221292 281724 221320
rect 281718 221280 281724 221292
rect 281776 221280 281782 221332
rect 292298 221280 292304 221332
rect 292356 221320 292362 221332
rect 299934 221320 299940 221332
rect 292356 221292 299940 221320
rect 292356 221280 292362 221292
rect 299934 221280 299940 221292
rect 299992 221280 299998 221332
rect 300136 221320 300164 221428
rect 302418 221416 302424 221468
rect 302476 221456 302482 221468
rect 334066 221456 334072 221468
rect 302476 221428 334072 221456
rect 302476 221416 302482 221428
rect 334066 221416 334072 221428
rect 334124 221416 334130 221468
rect 334986 221416 334992 221468
rect 335044 221456 335050 221468
rect 357526 221456 357532 221468
rect 335044 221428 357532 221456
rect 335044 221416 335050 221428
rect 357526 221416 357532 221428
rect 357584 221416 357590 221468
rect 357894 221416 357900 221468
rect 357952 221456 357958 221468
rect 374546 221456 374552 221468
rect 357952 221428 374552 221456
rect 357952 221416 357958 221428
rect 374546 221416 374552 221428
rect 374604 221416 374610 221468
rect 375466 221416 375472 221468
rect 375524 221456 375530 221468
rect 386506 221456 386512 221468
rect 375524 221428 386512 221456
rect 375524 221416 375530 221428
rect 386506 221416 386512 221428
rect 386564 221416 386570 221468
rect 390278 221416 390284 221468
rect 390336 221456 390342 221468
rect 401686 221456 401692 221468
rect 390336 221428 401692 221456
rect 390336 221416 390342 221428
rect 401686 221416 401692 221428
rect 401744 221416 401750 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 473078 221416 473084 221468
rect 473136 221456 473142 221468
rect 481174 221456 481180 221468
rect 473136 221428 481180 221456
rect 473136 221416 473142 221428
rect 481174 221416 481180 221428
rect 481232 221416 481238 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538766 221456 538772 221468
rect 483808 221428 538772 221456
rect 483808 221416 483814 221428
rect 538766 221416 538772 221428
rect 538824 221416 538830 221468
rect 540882 221416 540888 221468
rect 540940 221456 540946 221468
rect 605466 221456 605472 221468
rect 540940 221428 605472 221456
rect 540940 221416 540946 221428
rect 605466 221416 605472 221428
rect 605524 221416 605530 221468
rect 606478 221416 606484 221468
rect 606536 221456 606542 221468
rect 633434 221456 633440 221468
rect 606536 221428 633440 221456
rect 606536 221416 606542 221428
rect 633434 221416 633440 221428
rect 633492 221416 633498 221468
rect 303798 221320 303804 221332
rect 300136 221292 303804 221320
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 534902 221280 534908 221332
rect 534960 221320 534966 221332
rect 546770 221320 546776 221332
rect 534960 221292 546776 221320
rect 534960 221280 534966 221292
rect 546770 221280 546776 221292
rect 546828 221280 546834 221332
rect 547708 221292 552704 221320
rect 148410 221144 148416 221196
rect 148468 221184 148474 221196
rect 214098 221184 214104 221196
rect 148468 221156 214104 221184
rect 148468 221144 148474 221156
rect 214098 221144 214104 221156
rect 214156 221144 214162 221196
rect 214282 221144 214288 221196
rect 214340 221184 214346 221196
rect 263134 221184 263140 221196
rect 214340 221156 263140 221184
rect 214340 221144 214346 221156
rect 263134 221144 263140 221156
rect 263192 221144 263198 221196
rect 373994 221144 374000 221196
rect 374052 221184 374058 221196
rect 381078 221184 381084 221196
rect 374052 221156 381084 221184
rect 374052 221144 374058 221156
rect 381078 221144 381084 221156
rect 381136 221144 381142 221196
rect 542354 221144 542360 221196
rect 542412 221184 542418 221196
rect 543274 221184 543280 221196
rect 542412 221156 543280 221184
rect 542412 221144 542418 221156
rect 543274 221144 543280 221156
rect 543332 221184 543338 221196
rect 547708 221184 547736 221292
rect 543332 221156 547736 221184
rect 543332 221144 543338 221156
rect 552676 221116 552704 221292
rect 552842 221212 552848 221264
rect 552900 221252 552906 221264
rect 558178 221252 558184 221264
rect 552900 221224 558184 221252
rect 552900 221212 552906 221224
rect 558178 221212 558184 221224
rect 558236 221212 558242 221264
rect 558362 221212 558368 221264
rect 558420 221252 558426 221264
rect 596450 221252 596456 221264
rect 558420 221224 596456 221252
rect 558420 221212 558426 221224
rect 596450 221212 596456 221224
rect 596508 221212 596514 221264
rect 596634 221212 596640 221264
rect 596692 221252 596698 221264
rect 607490 221252 607496 221264
rect 596692 221224 607496 221252
rect 596692 221212 596698 221224
rect 607490 221212 607496 221224
rect 607548 221212 607554 221264
rect 552676 221088 596864 221116
rect 140958 221008 140964 221060
rect 141016 221048 141022 221060
rect 205818 221048 205824 221060
rect 141016 221020 205824 221048
rect 141016 221008 141022 221020
rect 205818 221008 205824 221020
rect 205876 221008 205882 221060
rect 222562 221008 222568 221060
rect 222620 221048 222626 221060
rect 270862 221048 270868 221060
rect 222620 221020 270868 221048
rect 222620 221008 222626 221020
rect 270862 221008 270868 221020
rect 270920 221008 270926 221060
rect 545758 221008 545764 221060
rect 545816 221048 545822 221060
rect 545816 221020 547874 221048
rect 545816 221008 545822 221020
rect 547846 220980 547874 221020
rect 552842 220980 552848 220992
rect 547846 220952 552848 220980
rect 552842 220940 552848 220952
rect 552900 220940 552906 220992
rect 553026 220940 553032 220992
rect 553084 220980 553090 220992
rect 596634 220980 596640 220992
rect 553084 220952 596640 220980
rect 553084 220940 553090 220952
rect 596634 220940 596640 220952
rect 596692 220940 596698 220992
rect 596836 220980 596864 221088
rect 597002 221076 597008 221128
rect 597060 221116 597066 221128
rect 606938 221116 606944 221128
rect 597060 221088 606944 221116
rect 597060 221076 597066 221088
rect 606938 221076 606944 221088
rect 606996 221076 607002 221128
rect 606202 220980 606208 220992
rect 596836 220952 606208 220980
rect 606202 220940 606208 220952
rect 606260 220940 606266 220992
rect 172606 220872 172612 220924
rect 172664 220912 172670 220924
rect 199470 220912 199476 220924
rect 172664 220884 199476 220912
rect 172664 220872 172670 220884
rect 199470 220872 199476 220884
rect 199528 220872 199534 220924
rect 227898 220872 227904 220924
rect 227956 220912 227962 220924
rect 276106 220912 276112 220924
rect 227956 220884 276112 220912
rect 227956 220872 227962 220884
rect 276106 220872 276112 220884
rect 276164 220872 276170 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423858 220844 423864 220856
rect 420696 220816 423864 220844
rect 420696 220804 420702 220816
rect 423858 220804 423864 220816
rect 423916 220804 423922 220856
rect 456702 220804 456708 220856
rect 456760 220844 456766 220856
rect 462130 220844 462136 220856
rect 456760 220816 462136 220844
rect 456760 220804 456766 220816
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 558178 220804 558184 220856
rect 558236 220844 558242 220856
rect 567838 220844 567844 220856
rect 558236 220816 567844 220844
rect 558236 220804 558242 220816
rect 567838 220804 567844 220816
rect 567896 220804 567902 220856
rect 577682 220804 577688 220856
rect 577740 220844 577746 220856
rect 628374 220844 628380 220856
rect 577740 220816 628380 220844
rect 577740 220804 577746 220816
rect 628374 220804 628380 220816
rect 628432 220804 628438 220856
rect 107838 220736 107844 220788
rect 107896 220776 107902 220788
rect 179966 220776 179972 220788
rect 107896 220748 179972 220776
rect 107896 220736 107902 220748
rect 179966 220736 179972 220748
rect 180024 220736 180030 220788
rect 187326 220736 187332 220788
rect 187384 220776 187390 220788
rect 241790 220776 241796 220788
rect 187384 220748 241796 220776
rect 187384 220736 187390 220748
rect 241790 220736 241796 220748
rect 241848 220736 241854 220788
rect 261018 220736 261024 220788
rect 261076 220776 261082 220788
rect 301682 220776 301688 220788
rect 261076 220748 301688 220776
rect 261076 220736 261082 220748
rect 301682 220736 301688 220748
rect 301740 220736 301746 220788
rect 313826 220736 313832 220788
rect 313884 220776 313890 220788
rect 320358 220776 320364 220788
rect 313884 220748 320364 220776
rect 313884 220736 313890 220748
rect 320358 220736 320364 220748
rect 320416 220736 320422 220788
rect 339218 220736 339224 220788
rect 339276 220776 339282 220788
rect 342438 220776 342444 220788
rect 339276 220748 342444 220776
rect 339276 220736 339282 220748
rect 342438 220736 342444 220748
rect 342496 220736 342502 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418338 220776 418344 220788
rect 414256 220748 418344 220776
rect 414256 220736 414262 220748
rect 418338 220736 418344 220748
rect 418396 220736 418402 220788
rect 465718 220736 465724 220788
rect 465776 220776 465782 220788
rect 469582 220776 469588 220788
rect 465776 220748 469588 220776
rect 465776 220736 465782 220748
rect 469582 220736 469588 220748
rect 469640 220736 469646 220788
rect 471882 220736 471888 220788
rect 471940 220776 471946 220788
rect 477862 220776 477868 220788
rect 471940 220748 477868 220776
rect 471940 220736 471946 220748
rect 477862 220736 477868 220748
rect 477920 220736 477926 220788
rect 552474 220736 552480 220788
rect 552532 220776 552538 220788
rect 552532 220748 553394 220776
rect 552532 220736 552538 220748
rect 455322 220668 455328 220720
rect 455380 220708 455386 220720
rect 458818 220708 458824 220720
rect 455380 220680 458824 220708
rect 455380 220668 455386 220680
rect 458818 220668 458824 220680
rect 458876 220668 458882 220720
rect 553366 220708 553394 220748
rect 568022 220736 568028 220788
rect 568080 220776 568086 220788
rect 577314 220776 577320 220788
rect 568080 220748 577320 220776
rect 568080 220736 568086 220748
rect 577314 220736 577320 220748
rect 577372 220736 577378 220788
rect 563054 220708 563060 220720
rect 553366 220680 563060 220708
rect 563054 220668 563060 220680
rect 563112 220668 563118 220720
rect 563256 220680 567056 220708
rect 66438 220600 66444 220652
rect 66496 220640 66502 220652
rect 144086 220640 144092 220652
rect 66496 220612 144092 220640
rect 66496 220600 66502 220612
rect 144086 220600 144092 220612
rect 144144 220600 144150 220652
rect 144270 220600 144276 220652
rect 144328 220640 144334 220652
rect 208578 220640 208584 220652
rect 144328 220612 208584 220640
rect 144328 220600 144334 220612
rect 208578 220600 208584 220612
rect 208636 220600 208642 220652
rect 216306 220600 216312 220652
rect 216364 220640 216370 220652
rect 217318 220640 217324 220652
rect 216364 220612 217324 220640
rect 216364 220600 216370 220612
rect 217318 220600 217324 220612
rect 217376 220600 217382 220652
rect 217502 220600 217508 220652
rect 217560 220640 217566 220652
rect 265066 220640 265072 220652
rect 217560 220612 265072 220640
rect 217560 220600 217566 220612
rect 265066 220600 265072 220612
rect 265124 220600 265130 220652
rect 280062 220600 280068 220652
rect 280120 220640 280126 220652
rect 314010 220640 314016 220652
rect 280120 220612 314016 220640
rect 280120 220600 280126 220612
rect 314010 220600 314016 220612
rect 314068 220600 314074 220652
rect 318150 220600 318156 220652
rect 318208 220640 318214 220652
rect 343818 220640 343824 220652
rect 318208 220612 343824 220640
rect 318208 220600 318214 220612
rect 343818 220600 343824 220612
rect 343876 220600 343882 220652
rect 508498 220600 508504 220652
rect 508556 220640 508562 220652
rect 520182 220640 520188 220652
rect 508556 220612 520188 220640
rect 508556 220600 508562 220612
rect 520182 220600 520188 220612
rect 520240 220600 520246 220652
rect 521470 220600 521476 220652
rect 521528 220640 521534 220652
rect 544102 220640 544108 220652
rect 521528 220612 544108 220640
rect 521528 220600 521534 220612
rect 544102 220600 544108 220612
rect 544160 220600 544166 220652
rect 553670 220532 553676 220584
rect 553728 220572 553734 220584
rect 553728 220544 560294 220572
rect 553728 220532 553734 220544
rect 86310 220464 86316 220516
rect 86368 220504 86374 220516
rect 164326 220504 164332 220516
rect 86368 220476 164332 220504
rect 86368 220464 86374 220476
rect 164326 220464 164332 220476
rect 164384 220464 164390 220516
rect 180702 220464 180708 220516
rect 180760 220504 180766 220516
rect 180760 220476 232544 220504
rect 180760 220464 180766 220476
rect 76374 220328 76380 220380
rect 76432 220368 76438 220380
rect 156138 220368 156144 220380
rect 76432 220340 156144 220368
rect 76432 220328 76438 220340
rect 156138 220328 156144 220340
rect 156196 220328 156202 220380
rect 170766 220328 170772 220380
rect 170824 220368 170830 220380
rect 229094 220368 229100 220380
rect 170824 220340 229100 220368
rect 170824 220328 170830 220340
rect 229094 220328 229100 220340
rect 229152 220328 229158 220380
rect 232516 220368 232544 220476
rect 232682 220464 232688 220516
rect 232740 220504 232746 220516
rect 238018 220504 238024 220516
rect 232740 220476 238024 220504
rect 232740 220464 232746 220476
rect 238018 220464 238024 220476
rect 238076 220464 238082 220516
rect 240318 220464 240324 220516
rect 240376 220504 240382 220516
rect 283098 220504 283104 220516
rect 240376 220476 283104 220504
rect 240376 220464 240382 220476
rect 283098 220464 283104 220476
rect 283156 220464 283162 220516
rect 283374 220464 283380 220516
rect 283432 220504 283438 220516
rect 316586 220504 316592 220516
rect 283432 220476 316592 220504
rect 283432 220464 283438 220476
rect 316586 220464 316592 220476
rect 316644 220464 316650 220516
rect 328914 220464 328920 220516
rect 328972 220504 328978 220516
rect 354674 220504 354680 220516
rect 328972 220476 354680 220504
rect 328972 220464 328978 220476
rect 354674 220464 354680 220476
rect 354732 220464 354738 220516
rect 385402 220504 385408 220516
rect 373966 220476 385408 220504
rect 232516 220340 233648 220368
rect 79686 220192 79692 220244
rect 79744 220232 79750 220244
rect 158898 220232 158904 220244
rect 79744 220204 158904 220232
rect 79744 220192 79750 220204
rect 158898 220192 158904 220204
rect 158956 220192 158962 220244
rect 161934 220192 161940 220244
rect 161992 220232 161998 220244
rect 161992 220204 219434 220232
rect 161992 220192 161998 220204
rect 73062 220056 73068 220108
rect 73120 220096 73126 220108
rect 153746 220096 153752 220108
rect 73120 220068 153752 220096
rect 73120 220056 73126 220068
rect 153746 220056 153752 220068
rect 153804 220056 153810 220108
rect 157518 220056 157524 220108
rect 157576 220096 157582 220108
rect 218698 220096 218704 220108
rect 157576 220068 218704 220096
rect 157576 220056 157582 220068
rect 218698 220056 218704 220068
rect 218756 220056 218762 220108
rect 219406 220096 219434 220204
rect 220814 220192 220820 220244
rect 220872 220232 220878 220244
rect 233418 220232 233424 220244
rect 220872 220204 233424 220232
rect 220872 220192 220878 220204
rect 233418 220192 233424 220204
rect 233476 220192 233482 220244
rect 233620 220232 233648 220340
rect 235626 220328 235632 220380
rect 235684 220368 235690 220380
rect 243078 220368 243084 220380
rect 235684 220340 243084 220368
rect 235684 220328 235690 220340
rect 243078 220328 243084 220340
rect 243136 220328 243142 220380
rect 246942 220328 246948 220380
rect 247000 220368 247006 220380
rect 288526 220368 288532 220380
rect 247000 220340 288532 220368
rect 247000 220328 247006 220340
rect 288526 220328 288532 220340
rect 288584 220328 288590 220380
rect 309870 220328 309876 220380
rect 309928 220368 309934 220380
rect 338114 220368 338120 220380
rect 309928 220340 338120 220368
rect 309928 220328 309934 220340
rect 338114 220328 338120 220340
rect 338172 220328 338178 220380
rect 343634 220328 343640 220380
rect 343692 220368 343698 220380
rect 347866 220368 347872 220380
rect 343692 220340 347872 220368
rect 343692 220328 343698 220340
rect 347866 220328 347872 220340
rect 347924 220328 347930 220380
rect 352926 220328 352932 220380
rect 352984 220368 352990 220380
rect 371418 220368 371424 220380
rect 352984 220340 371424 220368
rect 352984 220328 352990 220340
rect 371418 220328 371424 220340
rect 371476 220328 371482 220380
rect 372246 220328 372252 220380
rect 372304 220368 372310 220380
rect 373966 220368 373994 220476
rect 385402 220464 385408 220476
rect 385460 220464 385466 220516
rect 488074 220464 488080 220516
rect 488132 220504 488138 220516
rect 501874 220504 501880 220516
rect 488132 220476 501880 220504
rect 488132 220464 488138 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 519538 220464 519544 220516
rect 519596 220504 519602 220516
rect 534350 220504 534356 220516
rect 519596 220476 534356 220504
rect 519596 220464 519602 220476
rect 534350 220464 534356 220476
rect 534408 220464 534414 220516
rect 534718 220464 534724 220516
rect 534776 220504 534782 220516
rect 552474 220504 552480 220516
rect 534776 220476 552480 220504
rect 534776 220464 534782 220476
rect 552474 220464 552480 220476
rect 552532 220464 552538 220516
rect 560266 220504 560294 220544
rect 563256 220504 563284 220680
rect 567028 220640 567056 220680
rect 572070 220640 572076 220652
rect 567028 220612 572076 220640
rect 572070 220600 572076 220612
rect 572128 220600 572134 220652
rect 605282 220600 605288 220652
rect 605340 220640 605346 220652
rect 608962 220640 608968 220652
rect 605340 220612 608968 220640
rect 605340 220600 605346 220612
rect 608962 220600 608968 220612
rect 609020 220600 609026 220652
rect 560266 220476 563284 220504
rect 563422 220464 563428 220516
rect 563480 220504 563486 220516
rect 565446 220504 565452 220516
rect 563480 220476 565452 220504
rect 563480 220464 563486 220476
rect 565446 220464 565452 220476
rect 565504 220464 565510 220516
rect 565630 220464 565636 220516
rect 565688 220504 565694 220516
rect 566366 220504 566372 220516
rect 565688 220476 566372 220504
rect 565688 220464 565694 220476
rect 566366 220464 566372 220476
rect 566424 220464 566430 220516
rect 566826 220464 566832 220516
rect 566884 220504 566890 220516
rect 606478 220504 606484 220516
rect 566884 220476 606484 220504
rect 566884 220464 566890 220476
rect 606478 220464 606484 220476
rect 606536 220464 606542 220516
rect 558380 220408 558960 220436
rect 372304 220340 373994 220368
rect 372304 220328 372310 220340
rect 493962 220328 493968 220380
rect 494020 220368 494026 220380
rect 494020 220340 499574 220368
rect 494020 220328 494026 220340
rect 236638 220232 236644 220244
rect 233620 220204 236644 220232
rect 236638 220192 236644 220204
rect 236696 220192 236702 220244
rect 237006 220192 237012 220244
rect 237064 220232 237070 220244
rect 280430 220232 280436 220244
rect 237064 220204 280436 220232
rect 237064 220192 237070 220204
rect 280430 220192 280436 220204
rect 280488 220192 280494 220244
rect 299106 220192 299112 220244
rect 299164 220232 299170 220244
rect 331214 220232 331220 220244
rect 299164 220204 331220 220232
rect 299164 220192 299170 220204
rect 331214 220192 331220 220204
rect 331272 220192 331278 220244
rect 338022 220192 338028 220244
rect 338080 220232 338086 220244
rect 358998 220232 359004 220244
rect 338080 220204 359004 220232
rect 338080 220192 338086 220204
rect 358998 220192 359004 220204
rect 359056 220192 359062 220244
rect 361114 220192 361120 220244
rect 361172 220232 361178 220244
rect 377030 220232 377036 220244
rect 361172 220204 377036 220232
rect 361172 220192 361178 220204
rect 377030 220192 377036 220204
rect 377088 220192 377094 220244
rect 378042 220192 378048 220244
rect 378100 220232 378106 220244
rect 388622 220232 388628 220244
rect 378100 220204 388628 220232
rect 378100 220192 378106 220204
rect 388622 220192 388628 220204
rect 388680 220192 388686 220244
rect 432230 220192 432236 220244
rect 432288 220232 432294 220244
rect 434806 220232 434812 220244
rect 432288 220204 434812 220232
rect 432288 220192 432294 220204
rect 434806 220192 434812 220204
rect 434864 220192 434870 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 468846 220192 468852 220244
rect 468904 220232 468910 220244
rect 476206 220232 476212 220244
rect 468904 220204 476212 220232
rect 468904 220192 468910 220204
rect 476206 220192 476212 220204
rect 476264 220192 476270 220244
rect 481542 220192 481548 220244
rect 481600 220232 481606 220244
rect 492766 220232 492772 220244
rect 481600 220204 492772 220232
rect 481600 220192 481606 220204
rect 492766 220192 492772 220204
rect 492824 220192 492830 220244
rect 495158 220192 495164 220244
rect 495216 220232 495222 220244
rect 499546 220232 499574 220340
rect 500402 220328 500408 220380
rect 500460 220368 500466 220380
rect 515122 220368 515128 220380
rect 500460 220340 515128 220368
rect 500460 220328 500466 220340
rect 515122 220328 515128 220340
rect 515180 220328 515186 220380
rect 517146 220328 517152 220380
rect 517204 220368 517210 220380
rect 539226 220368 539232 220380
rect 517204 220340 539232 220368
rect 517204 220328 517210 220340
rect 539226 220328 539232 220340
rect 539284 220328 539290 220380
rect 553118 220328 553124 220380
rect 553176 220368 553182 220380
rect 554222 220368 554228 220380
rect 553176 220340 554228 220368
rect 553176 220328 553182 220340
rect 554222 220328 554228 220340
rect 554280 220328 554286 220380
rect 555418 220328 555424 220380
rect 555476 220368 555482 220380
rect 558380 220368 558408 220408
rect 555476 220340 558408 220368
rect 558932 220368 558960 220408
rect 566550 220368 566556 220380
rect 558932 220340 566556 220368
rect 555476 220328 555482 220340
rect 566550 220328 566556 220340
rect 566608 220328 566614 220380
rect 606294 220368 606300 220380
rect 567764 220340 606300 220368
rect 509326 220232 509332 220244
rect 495216 220204 495572 220232
rect 499546 220204 509332 220232
rect 495216 220192 495222 220204
rect 427906 220124 427912 220176
rect 427964 220164 427970 220176
rect 428734 220164 428740 220176
rect 427964 220136 428740 220164
rect 427964 220124 427970 220136
rect 428734 220124 428740 220136
rect 428792 220124 428798 220176
rect 221274 220096 221280 220108
rect 219406 220068 221280 220096
rect 221274 220056 221280 220068
rect 221332 220056 221338 220108
rect 230198 220056 230204 220108
rect 230256 220096 230262 220108
rect 275278 220096 275284 220108
rect 230256 220068 275284 220096
rect 230256 220056 230262 220068
rect 275278 220056 275284 220068
rect 275336 220056 275342 220108
rect 276842 220056 276848 220108
rect 276900 220096 276906 220108
rect 311342 220096 311348 220108
rect 276900 220068 311348 220096
rect 276900 220056 276906 220068
rect 311342 220056 311348 220068
rect 311400 220056 311406 220108
rect 311526 220056 311532 220108
rect 311584 220096 311590 220108
rect 338390 220096 338396 220108
rect 311584 220068 338396 220096
rect 311584 220056 311590 220068
rect 338390 220056 338396 220068
rect 338448 220056 338454 220108
rect 342714 220056 342720 220108
rect 342772 220096 342778 220108
rect 352374 220096 352380 220108
rect 342772 220068 352380 220096
rect 342772 220056 342778 220068
rect 352374 220056 352380 220068
rect 352432 220056 352438 220108
rect 354398 220056 354404 220108
rect 354456 220096 354462 220108
rect 372798 220096 372804 220108
rect 354456 220068 372804 220096
rect 354456 220056 354462 220068
rect 372798 220056 372804 220068
rect 372856 220056 372862 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 473262 220056 473268 220108
rect 473320 220096 473326 220108
rect 482002 220096 482008 220108
rect 473320 220068 482008 220096
rect 473320 220056 473326 220068
rect 482002 220056 482008 220068
rect 482060 220056 482066 220108
rect 482738 220056 482744 220108
rect 482796 220096 482802 220108
rect 495250 220096 495256 220108
rect 482796 220068 495256 220096
rect 482796 220056 482802 220068
rect 495250 220056 495256 220068
rect 495308 220056 495314 220108
rect 495544 220096 495572 220204
rect 509326 220192 509332 220204
rect 509384 220192 509390 220244
rect 536926 220192 536932 220244
rect 536984 220232 536990 220244
rect 558822 220232 558828 220244
rect 536984 220204 558828 220232
rect 536984 220192 536990 220204
rect 558822 220192 558828 220204
rect 558880 220192 558886 220244
rect 559374 220192 559380 220244
rect 559432 220232 559438 220244
rect 567764 220232 567792 220340
rect 606294 220328 606300 220340
rect 606352 220328 606358 220380
rect 559432 220204 567792 220232
rect 572686 220204 615494 220232
rect 559432 220192 559438 220204
rect 572686 220164 572714 220204
rect 567856 220136 572714 220164
rect 510982 220096 510988 220108
rect 495544 220068 510988 220096
rect 510982 220056 510988 220068
rect 511040 220056 511046 220108
rect 511810 220056 511816 220108
rect 511868 220096 511874 220108
rect 531682 220096 531688 220108
rect 511868 220068 531688 220096
rect 511868 220056 511874 220068
rect 531682 220056 531688 220068
rect 531740 220056 531746 220108
rect 534350 220056 534356 220108
rect 534408 220096 534414 220108
rect 534994 220096 535000 220108
rect 534408 220068 535000 220096
rect 534408 220056 534414 220068
rect 534994 220056 535000 220068
rect 535052 220096 535058 220108
rect 567856 220096 567884 220136
rect 535052 220068 558270 220096
rect 535052 220056 535058 220068
rect 558242 220028 558270 220068
rect 558840 220068 567884 220096
rect 558242 220000 558408 220028
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 185026 219960 185032 219972
rect 114520 219932 185032 219960
rect 114520 219920 114526 219932
rect 185026 219920 185032 219932
rect 185084 219920 185090 219972
rect 200574 219920 200580 219972
rect 200632 219960 200638 219972
rect 252738 219960 252744 219972
rect 200632 219932 252744 219960
rect 200632 219920 200638 219932
rect 252738 219920 252744 219932
rect 252796 219920 252802 219972
rect 256878 219920 256884 219972
rect 256936 219960 256942 219972
rect 295978 219960 295984 219972
rect 256936 219932 295984 219960
rect 256936 219920 256942 219932
rect 295978 219920 295984 219932
rect 296036 219920 296042 219972
rect 556246 219960 556252 219972
rect 547846 219932 556252 219960
rect 529014 219852 529020 219904
rect 529072 219892 529078 219904
rect 542538 219892 542544 219904
rect 529072 219864 542544 219892
rect 529072 219852 529078 219864
rect 542538 219852 542544 219864
rect 542596 219892 542602 219904
rect 547846 219892 547874 219932
rect 556246 219920 556252 219932
rect 556304 219920 556310 219972
rect 558380 219960 558408 220000
rect 558840 219960 558868 220068
rect 577314 220056 577320 220108
rect 577372 220096 577378 220108
rect 611354 220096 611360 220108
rect 577372 220068 611360 220096
rect 577372 220056 577378 220068
rect 611354 220056 611360 220068
rect 611412 220056 611418 220108
rect 615466 220096 615494 220204
rect 621106 220096 621112 220108
rect 615466 220068 621112 220096
rect 621106 220056 621112 220068
rect 621164 220056 621170 220108
rect 636470 220056 636476 220108
rect 636528 220096 636534 220108
rect 653398 220096 653404 220108
rect 636528 220068 653404 220096
rect 636528 220056 636534 220068
rect 653398 220056 653404 220068
rect 653456 220056 653462 220108
rect 676490 220056 676496 220108
rect 676548 220096 676554 220108
rect 677042 220096 677048 220108
rect 676548 220068 677048 220096
rect 676548 220056 676554 220068
rect 677042 220056 677048 220068
rect 677100 220056 677106 220108
rect 568298 219988 568304 220040
rect 568356 220028 568362 220040
rect 574462 220028 574468 220040
rect 568356 220000 574468 220028
rect 568356 219988 568362 220000
rect 574462 219988 574468 220000
rect 574520 219988 574526 220040
rect 558380 219932 558868 219960
rect 559558 219920 559564 219972
rect 559616 219960 559622 219972
rect 559616 219932 563054 219960
rect 559616 219920 559622 219932
rect 542596 219864 547874 219892
rect 563026 219892 563054 219932
rect 622486 219892 622492 219904
rect 563026 219864 622492 219892
rect 542596 219852 542602 219864
rect 622486 219852 622492 219864
rect 622544 219852 622550 219904
rect 127710 219784 127716 219836
rect 127768 219824 127774 219836
rect 195422 219824 195428 219836
rect 127768 219796 195428 219824
rect 127768 219784 127774 219796
rect 195422 219784 195428 219796
rect 195480 219784 195486 219836
rect 207198 219784 207204 219836
rect 207256 219824 207262 219836
rect 257246 219824 257252 219836
rect 207256 219796 257252 219824
rect 207256 219784 207262 219796
rect 257246 219784 257252 219796
rect 257304 219784 257310 219836
rect 288434 219784 288440 219836
rect 288492 219824 288498 219836
rect 310698 219824 310704 219836
rect 288492 219796 310704 219824
rect 288492 219784 288498 219796
rect 310698 219784 310704 219796
rect 310756 219784 310762 219836
rect 555786 219784 555792 219836
rect 555844 219824 555850 219836
rect 558454 219824 558460 219836
rect 555844 219796 558460 219824
rect 555844 219784 555850 219796
rect 558454 219784 558460 219796
rect 558512 219784 558518 219836
rect 558822 219784 558828 219836
rect 558880 219824 558886 219836
rect 558880 219796 562916 219824
rect 558880 219784 558886 219796
rect 546770 219716 546776 219768
rect 546828 219756 546834 219768
rect 547414 219756 547420 219768
rect 546828 219728 547420 219756
rect 546828 219716 546834 219728
rect 547414 219716 547420 219728
rect 547472 219756 547478 219768
rect 555418 219756 555424 219768
rect 547472 219728 555424 219756
rect 547472 219716 547478 219728
rect 555418 219716 555424 219728
rect 555476 219716 555482 219768
rect 562888 219756 562916 219796
rect 563422 219756 563428 219768
rect 562888 219728 563428 219756
rect 563422 219716 563428 219728
rect 563480 219716 563486 219768
rect 564342 219716 564348 219768
rect 564400 219756 564406 219768
rect 568574 219756 568580 219768
rect 564400 219728 568580 219756
rect 564400 219716 564406 219728
rect 568574 219716 568580 219728
rect 568632 219716 568638 219768
rect 568758 219716 568764 219768
rect 568816 219756 568822 219768
rect 605650 219756 605656 219768
rect 568816 219728 605656 219756
rect 568816 219716 568822 219728
rect 605650 219716 605656 219728
rect 605708 219716 605714 219768
rect 606478 219716 606484 219768
rect 606536 219756 606542 219768
rect 624326 219756 624332 219768
rect 606536 219728 624332 219756
rect 606536 219716 606542 219728
rect 624326 219716 624332 219728
rect 624384 219716 624390 219768
rect 137646 219648 137652 219700
rect 137704 219688 137710 219700
rect 203150 219688 203156 219700
rect 137704 219660 203156 219688
rect 137704 219648 137710 219660
rect 203150 219648 203156 219660
rect 203208 219648 203214 219700
rect 236178 219648 236184 219700
rect 236236 219688 236242 219700
rect 261478 219688 261484 219700
rect 236236 219660 261484 219688
rect 236236 219648 236242 219660
rect 261478 219648 261484 219660
rect 261536 219648 261542 219700
rect 558822 219648 558828 219700
rect 558880 219688 558886 219700
rect 559374 219688 559380 219700
rect 558880 219660 559380 219688
rect 558880 219648 558886 219660
rect 559374 219648 559380 219660
rect 559432 219648 559438 219700
rect 563790 219648 563796 219700
rect 563848 219688 563854 219700
rect 563848 219660 564112 219688
rect 563848 219648 563854 219660
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 539962 219580 539968 219632
rect 540020 219620 540026 219632
rect 558362 219620 558368 219632
rect 540020 219592 558368 219620
rect 540020 219580 540026 219592
rect 558362 219580 558368 219592
rect 558420 219580 558426 219632
rect 563514 219620 563520 219632
rect 560128 219592 563520 219620
rect 179414 219512 179420 219564
rect 179472 219552 179478 219564
rect 231946 219552 231952 219564
rect 179472 219524 231952 219552
rect 179472 219512 179478 219524
rect 231946 219512 231952 219524
rect 232004 219512 232010 219564
rect 270770 219512 270776 219564
rect 270828 219552 270834 219564
rect 279234 219552 279240 219564
rect 270828 219524 279240 219552
rect 270828 219512 270834 219524
rect 279234 219512 279240 219524
rect 279292 219512 279298 219564
rect 432046 219552 432052 219564
rect 431926 219524 432052 219552
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 70578 219376 70584 219428
rect 70636 219416 70642 219428
rect 149054 219416 149060 219428
rect 70636 219388 149060 219416
rect 70636 219376 70642 219388
rect 149054 219376 149060 219388
rect 149112 219376 149118 219428
rect 149238 219376 149244 219428
rect 149296 219416 149302 219428
rect 150250 219416 150256 219428
rect 149296 219388 150256 219416
rect 149296 219376 149302 219388
rect 150250 219376 150256 219388
rect 150308 219376 150314 219428
rect 152550 219376 152556 219428
rect 152608 219416 152614 219428
rect 153102 219416 153108 219428
rect 152608 219388 153108 219416
rect 152608 219376 152614 219388
rect 153102 219376 153108 219388
rect 153160 219376 153166 219428
rect 155034 219376 155040 219428
rect 155092 219416 155098 219428
rect 155954 219416 155960 219428
rect 155092 219388 155960 219416
rect 155092 219376 155098 219388
rect 155954 219376 155960 219388
rect 156012 219376 156018 219428
rect 156138 219376 156144 219428
rect 156196 219416 156202 219428
rect 162854 219416 162860 219428
rect 156196 219388 162860 219416
rect 156196 219376 156202 219388
rect 162854 219376 162860 219388
rect 162912 219376 162918 219428
rect 165798 219376 165804 219428
rect 165856 219416 165862 219428
rect 173158 219416 173164 219428
rect 165856 219388 173164 219416
rect 165856 219376 165862 219388
rect 173158 219376 173164 219388
rect 173216 219376 173222 219428
rect 179046 219376 179052 219428
rect 179104 219416 179110 219428
rect 182818 219416 182824 219428
rect 179104 219388 182824 219416
rect 179104 219376 179110 219388
rect 182818 219376 182824 219388
rect 182876 219376 182882 219428
rect 183186 219376 183192 219428
rect 183244 219416 183250 219428
rect 199286 219416 199292 219428
rect 183244 219388 199292 219416
rect 183244 219376 183250 219388
rect 199286 219376 199292 219388
rect 199344 219376 199350 219428
rect 199746 219376 199752 219428
rect 199804 219416 199810 219428
rect 203058 219416 203064 219428
rect 199804 219388 203064 219416
rect 199804 219376 199810 219388
rect 203058 219376 203064 219388
rect 203116 219376 203122 219428
rect 204714 219376 204720 219428
rect 204772 219416 204778 219428
rect 205634 219416 205640 219428
rect 204772 219388 205640 219416
rect 204772 219376 204778 219388
rect 205634 219376 205640 219388
rect 205692 219376 205698 219428
rect 209682 219376 209688 219428
rect 209740 219416 209746 219428
rect 210326 219416 210332 219428
rect 209740 219388 210332 219416
rect 209740 219376 209746 219388
rect 210326 219376 210332 219388
rect 210384 219376 210390 219428
rect 212810 219376 212816 219428
rect 212868 219416 212874 219428
rect 252554 219416 252560 219428
rect 212868 219388 252560 219416
rect 212868 219376 212874 219388
rect 252554 219376 252560 219388
rect 252612 219376 252618 219428
rect 254394 219376 254400 219428
rect 254452 219416 254458 219428
rect 255314 219416 255320 219428
rect 254452 219388 255320 219416
rect 254452 219376 254458 219388
rect 255314 219376 255320 219388
rect 255372 219376 255378 219428
rect 272426 219376 272432 219428
rect 272484 219416 272490 219428
rect 297358 219416 297364 219428
rect 272484 219388 297364 219416
rect 272484 219376 272490 219388
rect 297358 219376 297364 219388
rect 297416 219376 297422 219428
rect 312354 219376 312360 219428
rect 312412 219416 312418 219428
rect 313274 219416 313280 219428
rect 312412 219388 313280 219416
rect 312412 219376 312418 219388
rect 313274 219376 313280 219388
rect 313332 219376 313338 219428
rect 323118 219376 323124 219428
rect 323176 219416 323182 219428
rect 324222 219416 324228 219428
rect 323176 219388 324228 219416
rect 323176 219376 323182 219388
rect 324222 219376 324228 219388
rect 324280 219376 324286 219428
rect 324774 219376 324780 219428
rect 324832 219416 324838 219428
rect 325510 219416 325516 219428
rect 324832 219388 325516 219416
rect 324832 219376 324838 219388
rect 325510 219376 325516 219388
rect 325568 219376 325574 219428
rect 326430 219376 326436 219428
rect 326488 219416 326494 219428
rect 326890 219416 326896 219428
rect 326488 219388 326896 219416
rect 326488 219376 326494 219388
rect 326890 219376 326896 219388
rect 326948 219376 326954 219428
rect 327718 219416 327724 219428
rect 327092 219388 327724 219416
rect 63954 219240 63960 219292
rect 64012 219280 64018 219292
rect 65518 219280 65524 219292
rect 64012 219252 65524 219280
rect 64012 219240 64018 219252
rect 65518 219240 65524 219252
rect 65576 219240 65582 219292
rect 113634 219240 113640 219292
rect 113692 219280 113698 219292
rect 166258 219280 166264 219292
rect 113692 219252 166264 219280
rect 113692 219240 113698 219252
rect 166258 219240 166264 219252
rect 166316 219240 166322 219292
rect 192938 219240 192944 219292
rect 192996 219280 193002 219292
rect 233878 219280 233884 219292
rect 192996 219252 233884 219280
rect 192996 219240 193002 219252
rect 233878 219240 233884 219252
rect 233936 219240 233942 219292
rect 237834 219240 237840 219292
rect 237892 219280 237898 219292
rect 239398 219280 239404 219292
rect 237892 219252 239404 219280
rect 237892 219240 237898 219252
rect 239398 219240 239404 219252
rect 239456 219240 239462 219292
rect 252738 219240 252744 219292
rect 252796 219280 252802 219292
rect 252796 219252 258074 219280
rect 252796 219240 252802 219252
rect 87138 219104 87144 219156
rect 87196 219144 87202 219156
rect 106918 219144 106924 219156
rect 87196 219116 106924 219144
rect 87196 219104 87202 219116
rect 106918 219104 106924 219116
rect 106976 219104 106982 219156
rect 107102 219104 107108 219156
rect 107160 219144 107166 219156
rect 159358 219144 159364 219156
rect 107160 219116 159364 219144
rect 107160 219104 107166 219116
rect 159358 219104 159364 219116
rect 159416 219104 159422 219156
rect 163314 219104 163320 219156
rect 163372 219144 163378 219156
rect 163372 219116 169110 219144
rect 163372 219104 163378 219116
rect 59814 218968 59820 219020
rect 59872 219008 59878 219020
rect 137278 219008 137284 219020
rect 59872 218980 137284 219008
rect 59872 218968 59878 218980
rect 137278 218968 137284 218980
rect 137336 218968 137342 219020
rect 143718 218968 143724 219020
rect 143776 219008 143782 219020
rect 160738 219008 160744 219020
rect 143776 218980 160744 219008
rect 143776 218968 143782 218980
rect 160738 218968 160744 218980
rect 160796 218968 160802 219020
rect 162486 218968 162492 219020
rect 162544 219008 162550 219020
rect 168926 219008 168932 219020
rect 162544 218980 168932 219008
rect 162544 218968 162550 218980
rect 168926 218968 168932 218980
rect 168984 218968 168990 219020
rect 169082 219008 169110 219116
rect 169938 219104 169944 219156
rect 169996 219144 170002 219156
rect 196618 219144 196624 219156
rect 169996 219116 196624 219144
rect 169996 219104 170002 219116
rect 196618 219104 196624 219116
rect 196676 219104 196682 219156
rect 203058 219104 203064 219156
rect 203116 219144 203122 219156
rect 247126 219144 247132 219156
rect 203116 219116 247132 219144
rect 203116 219104 203122 219116
rect 247126 219104 247132 219116
rect 247184 219104 247190 219156
rect 258046 219144 258074 219252
rect 259178 219240 259184 219292
rect 259236 219280 259242 219292
rect 292298 219280 292304 219292
rect 259236 219252 292304 219280
rect 259236 219240 259242 219252
rect 292298 219240 292304 219252
rect 292356 219240 292362 219292
rect 307386 219240 307392 219292
rect 307444 219280 307450 219292
rect 307444 219252 323808 219280
rect 307444 219240 307450 219252
rect 258046 219116 287054 219144
rect 184198 219008 184204 219020
rect 169082 218980 184204 219008
rect 184198 218968 184204 218980
rect 184256 218968 184262 219020
rect 186498 218968 186504 219020
rect 186556 219008 186562 219020
rect 235626 219008 235632 219020
rect 186556 218980 235632 219008
rect 186556 218968 186562 218980
rect 235626 218968 235632 218980
rect 235684 218968 235690 219020
rect 246114 218968 246120 219020
rect 246172 219008 246178 219020
rect 284018 219008 284024 219020
rect 246172 218980 284024 219008
rect 246172 218968 246178 218980
rect 284018 218968 284024 218980
rect 284076 218968 284082 219020
rect 287026 219008 287054 219116
rect 300578 219104 300584 219156
rect 300636 219144 300642 219156
rect 322842 219144 322848 219156
rect 300636 219116 322848 219144
rect 300636 219104 300642 219116
rect 322842 219104 322848 219116
rect 322900 219104 322906 219156
rect 323780 219144 323808 219252
rect 323946 219240 323952 219292
rect 324004 219280 324010 219292
rect 324958 219280 324964 219292
rect 324004 219252 324964 219280
rect 324004 219240 324010 219252
rect 324958 219240 324964 219252
rect 325016 219240 325022 219292
rect 327092 219280 327120 219388
rect 327718 219376 327724 219388
rect 327776 219376 327782 219428
rect 341334 219376 341340 219428
rect 341392 219416 341398 219428
rect 342254 219416 342260 219428
rect 341392 219388 342260 219416
rect 341392 219376 341398 219388
rect 342254 219376 342260 219388
rect 342312 219376 342318 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 354582 219376 354588 219428
rect 354640 219416 354646 219428
rect 355318 219416 355324 219428
rect 354640 219388 355324 219416
rect 354640 219376 354646 219388
rect 355318 219376 355324 219388
rect 355376 219376 355382 219428
rect 373626 219376 373632 219428
rect 373684 219416 373690 219428
rect 378042 219416 378048 219428
rect 373684 219388 378048 219416
rect 373684 219376 373690 219388
rect 378042 219376 378048 219388
rect 378100 219376 378106 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 403434 219376 403440 219428
rect 403492 219416 403498 219428
rect 404354 219416 404360 219428
rect 403492 219388 404360 219416
rect 403492 219376 403498 219388
rect 404354 219376 404360 219388
rect 404412 219376 404418 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 431926 219484 431954 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 558638 219512 558644 219564
rect 558696 219552 558702 219564
rect 560128 219552 560156 219592
rect 563514 219580 563520 219592
rect 563572 219580 563578 219632
rect 564084 219620 564112 219660
rect 676214 219648 676220 219700
rect 676272 219688 676278 219700
rect 678422 219688 678428 219700
rect 676272 219660 678428 219688
rect 676272 219648 676278 219660
rect 678422 219648 678428 219660
rect 678480 219648 678486 219700
rect 605282 219620 605288 219632
rect 564084 219592 605288 219620
rect 605282 219580 605288 219592
rect 605340 219580 605346 219632
rect 606294 219580 606300 219632
rect 606352 219620 606358 219632
rect 622670 219620 622676 219632
rect 606352 219592 622676 219620
rect 606352 219580 606358 219592
rect 622670 219580 622676 219592
rect 622728 219580 622734 219632
rect 558696 219524 560156 219552
rect 558696 219512 558702 219524
rect 563008 219484 563014 219496
rect 429212 219456 431954 219484
rect 560266 219456 563014 219484
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219456
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 438210 219376 438216 219428
rect 438268 219416 438274 219428
rect 438854 219416 438860 219428
rect 438268 219388 438860 219416
rect 438268 219376 438274 219388
rect 438854 219376 438860 219388
rect 438912 219376 438918 219428
rect 439866 219376 439872 219428
rect 439924 219416 439930 219428
rect 440326 219416 440332 219428
rect 439924 219388 440332 219416
rect 439924 219376 439930 219388
rect 440326 219376 440332 219388
rect 440384 219376 440390 219428
rect 527726 219376 527732 219428
rect 527784 219416 527790 219428
rect 528278 219416 528284 219428
rect 527784 219388 528284 219416
rect 527784 219376 527790 219388
rect 528278 219376 528284 219388
rect 528336 219376 528342 219428
rect 548150 219376 548156 219428
rect 548208 219416 548214 219428
rect 552658 219416 552664 219428
rect 548208 219388 552664 219416
rect 548208 219376 548214 219388
rect 552658 219376 552664 219388
rect 552716 219376 552722 219428
rect 560266 219416 560294 219456
rect 563008 219444 563014 219456
rect 563066 219444 563072 219496
rect 563698 219484 563704 219496
rect 563164 219456 563704 219484
rect 554516 219388 560294 219416
rect 553854 219348 553860 219360
rect 552860 219320 553860 219348
rect 325160 219252 327120 219280
rect 325160 219144 325188 219252
rect 327258 219240 327264 219292
rect 327316 219280 327322 219292
rect 342714 219280 342720 219292
rect 327316 219252 342720 219280
rect 327316 219240 327322 219252
rect 342714 219240 342720 219252
rect 342772 219240 342778 219292
rect 358722 219240 358728 219292
rect 358780 219280 358786 219292
rect 363782 219280 363788 219292
rect 358780 219252 363788 219280
rect 358780 219240 358786 219252
rect 363782 219240 363788 219252
rect 363840 219240 363846 219292
rect 479702 219240 479708 219292
rect 479760 219280 479766 219292
rect 480346 219280 480352 219292
rect 479760 219252 480352 219280
rect 479760 219240 479766 219252
rect 480346 219240 480352 219252
rect 480404 219240 480410 219292
rect 533706 219240 533712 219292
rect 533764 219280 533770 219292
rect 534442 219280 534448 219292
rect 533764 219252 534448 219280
rect 533764 219240 533770 219252
rect 534442 219240 534448 219252
rect 534500 219240 534506 219292
rect 547874 219240 547880 219292
rect 547932 219280 547938 219292
rect 549070 219280 549076 219292
rect 547932 219252 549076 219280
rect 547932 219240 547938 219252
rect 549070 219240 549076 219252
rect 549128 219240 549134 219292
rect 549898 219240 549904 219292
rect 549956 219280 549962 219292
rect 552860 219280 552888 219320
rect 553854 219308 553860 219320
rect 553912 219308 553918 219360
rect 549956 219252 552888 219280
rect 549956 219240 549962 219252
rect 323780 219116 325188 219144
rect 325602 219104 325608 219156
rect 325660 219144 325666 219156
rect 330386 219144 330392 219156
rect 325660 219116 330392 219144
rect 325660 219104 325666 219116
rect 330386 219104 330392 219116
rect 330444 219104 330450 219156
rect 363690 219104 363696 219156
rect 363748 219144 363754 219156
rect 373994 219144 374000 219156
rect 363748 219116 374000 219144
rect 363748 219104 363754 219116
rect 373994 219104 374000 219116
rect 374052 219104 374058 219156
rect 419166 219104 419172 219156
rect 419224 219144 419230 219156
rect 422662 219144 422668 219156
rect 419224 219116 422668 219144
rect 419224 219104 419230 219116
rect 422662 219104 422668 219116
rect 422720 219104 422726 219156
rect 466086 219104 466092 219156
rect 466144 219144 466150 219156
rect 472894 219144 472900 219156
rect 466144 219116 472900 219144
rect 466144 219104 466150 219116
rect 472894 219104 472900 219116
rect 472952 219104 472958 219156
rect 531958 219104 531964 219156
rect 532016 219144 532022 219156
rect 532510 219144 532516 219156
rect 532016 219116 532516 219144
rect 532016 219104 532022 219116
rect 532510 219104 532516 219116
rect 532568 219144 532574 219156
rect 534258 219144 534264 219156
rect 532568 219116 534264 219144
rect 532568 219104 532574 219116
rect 534258 219104 534264 219116
rect 534316 219104 534322 219156
rect 537478 219104 537484 219156
rect 537536 219144 537542 219156
rect 539686 219144 539692 219156
rect 537536 219116 539692 219144
rect 537536 219104 537542 219116
rect 539686 219104 539692 219116
rect 539744 219104 539750 219156
rect 544378 219104 544384 219156
rect 544436 219144 544442 219156
rect 545022 219144 545028 219156
rect 544436 219116 545028 219144
rect 544436 219104 544442 219116
rect 545022 219104 545028 219116
rect 545080 219144 545086 219156
rect 548150 219144 548156 219156
rect 545080 219116 548156 219144
rect 545080 219104 545086 219116
rect 548150 219104 548156 219116
rect 548208 219104 548214 219156
rect 554516 219144 554544 219388
rect 563164 219280 563192 219456
rect 563698 219444 563704 219456
rect 563756 219444 563762 219496
rect 564158 219444 564164 219496
rect 564216 219484 564222 219496
rect 625154 219484 625160 219496
rect 564216 219456 625160 219484
rect 564216 219444 564222 219456
rect 625154 219444 625160 219456
rect 625212 219444 625218 219496
rect 605650 219308 605656 219360
rect 605708 219348 605714 219360
rect 608778 219348 608784 219360
rect 605708 219320 608784 219348
rect 605708 219308 605714 219320
rect 608778 219308 608784 219320
rect 608836 219308 608842 219360
rect 548352 219116 554544 219144
rect 554700 219252 563192 219280
rect 289078 219008 289084 219020
rect 287026 218980 289084 219008
rect 289078 218968 289084 218980
rect 289136 218968 289142 219020
rect 294138 218968 294144 219020
rect 294196 219008 294202 219020
rect 309686 219008 309692 219020
rect 294196 218980 309692 219008
rect 294196 218968 294202 218980
rect 309686 218968 309692 218980
rect 309744 218968 309750 219020
rect 314010 218968 314016 219020
rect 314068 219008 314074 219020
rect 339218 219008 339224 219020
rect 314068 218980 339224 219008
rect 314068 218968 314074 218980
rect 339218 218968 339224 218980
rect 339276 218968 339282 219020
rect 340506 218968 340512 219020
rect 340564 219008 340570 219020
rect 351086 219008 351092 219020
rect 340564 218980 351092 219008
rect 340564 218968 340570 218980
rect 351086 218968 351092 218980
rect 351144 218968 351150 219020
rect 370314 218968 370320 219020
rect 370372 219008 370378 219020
rect 375466 219008 375472 219020
rect 370372 218980 375472 219008
rect 370372 218968 370378 218980
rect 375466 218968 375472 218980
rect 375524 218968 375530 219020
rect 383562 218968 383568 219020
rect 383620 219008 383626 219020
rect 388438 219008 388444 219020
rect 383620 218980 388444 219008
rect 383620 218968 383626 218980
rect 388438 218968 388444 218980
rect 388496 218968 388502 219020
rect 505094 218968 505100 219020
rect 505152 219008 505158 219020
rect 505152 218980 514754 219008
rect 505152 218968 505158 218980
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 156138 218872 156144 218884
rect 83884 218844 156144 218872
rect 83884 218832 83890 218844
rect 156138 218832 156144 218844
rect 156196 218832 156202 218884
rect 167638 218872 167644 218884
rect 161446 218844 167644 218872
rect 92934 218696 92940 218748
rect 92992 218736 92998 218748
rect 93762 218736 93768 218748
rect 92992 218708 93768 218736
rect 92992 218696 92998 218708
rect 93762 218696 93768 218708
rect 93820 218696 93826 218748
rect 100386 218696 100392 218748
rect 100444 218736 100450 218748
rect 146938 218736 146944 218748
rect 100444 218708 146944 218736
rect 100444 218696 100450 218708
rect 146938 218696 146944 218708
rect 146996 218696 147002 218748
rect 149054 218696 149060 218748
rect 149112 218736 149118 218748
rect 153194 218736 153200 218748
rect 149112 218708 153200 218736
rect 149112 218696 149118 218708
rect 153194 218696 153200 218708
rect 153252 218696 153258 218748
rect 153378 218696 153384 218748
rect 153436 218736 153442 218748
rect 161446 218736 161474 218844
rect 167638 218832 167644 218844
rect 167696 218832 167702 218884
rect 173250 218832 173256 218884
rect 173308 218872 173314 218884
rect 210878 218872 210884 218884
rect 173308 218844 210884 218872
rect 173308 218832 173314 218844
rect 210878 218832 210884 218844
rect 210936 218832 210942 218884
rect 232866 218832 232872 218884
rect 232924 218872 232930 218884
rect 270770 218872 270776 218884
rect 232924 218844 270776 218872
rect 232924 218832 232930 218844
rect 270770 218832 270776 218844
rect 270828 218832 270834 218884
rect 285858 218832 285864 218884
rect 285916 218872 285922 218884
rect 313826 218872 313832 218884
rect 285916 218844 313832 218872
rect 285916 218832 285922 218844
rect 313826 218832 313832 218844
rect 313884 218832 313890 218884
rect 343634 218872 343640 218884
rect 331186 218844 343640 218872
rect 153436 218708 161474 218736
rect 153436 218696 153442 218708
rect 166626 218696 166632 218748
rect 166684 218736 166690 218748
rect 169754 218736 169760 218748
rect 166684 218708 169760 218736
rect 166684 218696 166690 218708
rect 169754 218696 169760 218708
rect 169812 218696 169818 218748
rect 171410 218696 171416 218748
rect 171468 218736 171474 218748
rect 175918 218736 175924 218748
rect 171468 218708 175924 218736
rect 171468 218696 171474 218708
rect 175918 218696 175924 218708
rect 175976 218696 175982 218748
rect 176286 218696 176292 218748
rect 176344 218736 176350 218748
rect 189718 218736 189724 218748
rect 176344 218708 189724 218736
rect 176344 218696 176350 218708
rect 189718 218696 189724 218708
rect 189776 218696 189782 218748
rect 232682 218736 232688 218748
rect 190426 218708 232688 218736
rect 63126 218628 63132 218680
rect 63184 218668 63190 218680
rect 68278 218668 68284 218680
rect 63184 218640 68284 218668
rect 63184 218628 63190 218640
rect 68278 218628 68284 218640
rect 68336 218628 68342 218680
rect 93762 218560 93768 218612
rect 93820 218600 93826 218612
rect 139946 218600 139952 218612
rect 93820 218572 139952 218600
rect 93820 218560 93826 218572
rect 139946 218560 139952 218572
rect 140004 218560 140010 218612
rect 140130 218560 140136 218612
rect 140188 218600 140194 218612
rect 143718 218600 143724 218612
rect 140188 218572 143724 218600
rect 140188 218560 140194 218572
rect 143718 218560 143724 218572
rect 143776 218560 143782 218612
rect 146754 218560 146760 218612
rect 146812 218600 146818 218612
rect 189902 218600 189908 218612
rect 146812 218572 189908 218600
rect 146812 218560 146818 218572
rect 189902 218560 189908 218572
rect 189960 218560 189966 218612
rect 166442 218464 166448 218476
rect 122806 218436 166448 218464
rect 68738 218288 68744 218340
rect 68796 218328 68802 218340
rect 72418 218328 72424 218340
rect 68796 218300 72424 218328
rect 68796 218288 68802 218300
rect 72418 218288 72424 218300
rect 72476 218288 72482 218340
rect 120258 218288 120264 218340
rect 120316 218328 120322 218340
rect 122806 218328 122834 218436
rect 166442 218424 166448 218436
rect 166500 218424 166506 218476
rect 168098 218424 168104 218476
rect 168156 218464 168162 218476
rect 171042 218464 171048 218476
rect 168156 218436 171048 218464
rect 168156 218424 168162 218436
rect 171042 218424 171048 218436
rect 171100 218424 171106 218476
rect 172146 218424 172152 218476
rect 172204 218464 172210 218476
rect 177206 218464 177212 218476
rect 172204 218436 177212 218464
rect 172204 218424 172210 218436
rect 177206 218424 177212 218436
rect 177264 218424 177270 218476
rect 179874 218424 179880 218476
rect 179932 218464 179938 218476
rect 190426 218464 190454 218708
rect 232682 218696 232688 218708
rect 232740 218696 232746 218748
rect 233878 218696 233884 218748
rect 233936 218736 233942 218748
rect 238846 218736 238852 218748
rect 233936 218708 238852 218736
rect 233936 218696 233942 218708
rect 238846 218696 238852 218708
rect 238904 218696 238910 218748
rect 239490 218696 239496 218748
rect 239548 218736 239554 218748
rect 280706 218736 280712 218748
rect 239548 218708 280712 218736
rect 239548 218696 239554 218708
rect 280706 218696 280712 218708
rect 280764 218696 280770 218748
rect 291654 218696 291660 218748
rect 291712 218736 291718 218748
rect 323578 218736 323584 218748
rect 291712 218708 323584 218736
rect 291712 218696 291718 218708
rect 323578 218696 323584 218708
rect 323636 218696 323642 218748
rect 198918 218560 198924 218612
rect 198976 218600 198982 218612
rect 200022 218600 200028 218612
rect 198976 218572 200028 218600
rect 198976 218560 198982 218572
rect 200022 218560 200028 218572
rect 200080 218560 200086 218612
rect 201862 218560 201868 218612
rect 201920 218600 201926 218612
rect 206186 218600 206192 218612
rect 201920 218572 206192 218600
rect 201920 218560 201926 218572
rect 206186 218560 206192 218572
rect 206244 218560 206250 218612
rect 206370 218560 206376 218612
rect 206428 218600 206434 218612
rect 212810 218600 212816 218612
rect 206428 218572 212816 218600
rect 206428 218560 206434 218572
rect 212810 218560 212816 218572
rect 212868 218560 212874 218612
rect 212994 218560 213000 218612
rect 213052 218600 213058 218612
rect 260006 218600 260012 218612
rect 213052 218572 260012 218600
rect 213052 218560 213058 218572
rect 260006 218560 260012 218572
rect 260064 218560 260070 218612
rect 262674 218560 262680 218612
rect 262732 218600 262738 218612
rect 276566 218600 276572 218612
rect 262732 218572 276572 218600
rect 262732 218560 262738 218572
rect 276566 218560 276572 218572
rect 276624 218560 276630 218612
rect 279234 218560 279240 218612
rect 279292 218600 279298 218612
rect 307018 218600 307024 218612
rect 279292 218572 307024 218600
rect 279292 218560 279298 218572
rect 307018 218560 307024 218572
rect 307076 218560 307082 218612
rect 320634 218560 320640 218612
rect 320692 218600 320698 218612
rect 331186 218600 331214 218844
rect 343634 218832 343640 218844
rect 343692 218832 343698 218884
rect 347130 218832 347136 218884
rect 347188 218872 347194 218884
rect 363506 218872 363512 218884
rect 347188 218844 363512 218872
rect 347188 218832 347194 218844
rect 363506 218832 363512 218844
rect 363564 218832 363570 218884
rect 392670 218832 392676 218884
rect 392728 218872 392734 218884
rect 400766 218872 400772 218884
rect 392728 218844 400772 218872
rect 392728 218832 392734 218844
rect 400766 218832 400772 218844
rect 400824 218832 400830 218884
rect 401778 218832 401784 218884
rect 401836 218872 401842 218884
rect 407758 218872 407764 218884
rect 401836 218844 407764 218872
rect 401836 218832 401842 218844
rect 407758 218832 407764 218844
rect 407816 218832 407822 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 499574 218832 499580 218884
rect 499632 218872 499638 218884
rect 505278 218872 505284 218884
rect 499632 218844 505284 218872
rect 499632 218832 499638 218844
rect 505278 218832 505284 218844
rect 505336 218832 505342 218884
rect 514726 218804 514754 218980
rect 534074 218968 534080 219020
rect 534132 219008 534138 219020
rect 548352 219008 548380 219116
rect 534132 218980 548380 219008
rect 534132 218968 534138 218980
rect 548702 218968 548708 219020
rect 548760 219008 548766 219020
rect 554700 219008 554728 219252
rect 563422 219240 563428 219292
rect 563480 219280 563486 219292
rect 572438 219280 572444 219292
rect 563480 219252 572444 219280
rect 563480 219240 563486 219252
rect 572438 219240 572444 219252
rect 572496 219240 572502 219292
rect 572622 219240 572628 219292
rect 572680 219280 572686 219292
rect 575658 219280 575664 219292
rect 572680 219252 575664 219280
rect 572680 219240 572686 219252
rect 575658 219240 575664 219252
rect 575716 219240 575722 219292
rect 591390 219172 591396 219224
rect 591448 219212 591454 219224
rect 594150 219212 594156 219224
rect 591448 219184 594156 219212
rect 591448 219172 591454 219184
rect 594150 219172 594156 219184
rect 594208 219172 594214 219224
rect 554866 219104 554872 219156
rect 554924 219144 554930 219156
rect 554924 219116 556476 219144
rect 554924 219104 554930 219116
rect 548760 218980 554728 219008
rect 556448 219008 556476 219116
rect 556890 219104 556896 219156
rect 556948 219144 556954 219156
rect 587342 219144 587348 219156
rect 556948 219116 587348 219144
rect 556948 219104 556954 219116
rect 587342 219104 587348 219116
rect 587400 219104 587406 219156
rect 566734 219008 566740 219020
rect 556448 218980 566740 219008
rect 548760 218968 548766 218980
rect 566734 218968 566740 218980
rect 566792 218968 566798 219020
rect 572254 219008 572260 219020
rect 566936 218980 572260 219008
rect 518894 218900 518900 218952
rect 518952 218940 518958 218952
rect 519446 218940 519452 218952
rect 518952 218912 519452 218940
rect 518952 218900 518958 218912
rect 519446 218900 519452 218912
rect 519504 218900 519510 218952
rect 524782 218900 524788 218952
rect 524840 218940 524846 218952
rect 528462 218940 528468 218952
rect 524840 218912 528468 218940
rect 524840 218900 524846 218912
rect 528462 218900 528468 218912
rect 528520 218900 528526 218952
rect 534442 218832 534448 218884
rect 534500 218872 534506 218884
rect 553670 218872 553676 218884
rect 534500 218844 553676 218872
rect 534500 218832 534506 218844
rect 553670 218832 553676 218844
rect 553728 218832 553734 218884
rect 553854 218832 553860 218884
rect 553912 218872 553918 218884
rect 558178 218872 558184 218884
rect 553912 218844 558184 218872
rect 553912 218832 553918 218844
rect 558178 218832 558184 218844
rect 558236 218832 558242 218884
rect 559834 218832 559840 218884
rect 559892 218872 559898 218884
rect 563008 218872 563014 218884
rect 559892 218844 563014 218872
rect 559892 218832 559898 218844
rect 563008 218832 563014 218844
rect 563066 218832 563072 218884
rect 563146 218832 563152 218884
rect 563204 218872 563210 218884
rect 566936 218872 566964 218980
rect 572254 218968 572260 218980
rect 572312 218968 572318 219020
rect 572438 218968 572444 219020
rect 572496 219008 572502 219020
rect 575842 219008 575848 219020
rect 572496 218980 575848 219008
rect 572496 218968 572502 218980
rect 575842 218968 575848 218980
rect 575900 218968 575906 219020
rect 597738 219008 597744 219020
rect 582346 218980 597744 219008
rect 563204 218844 566964 218872
rect 563204 218832 563210 218844
rect 567102 218832 567108 218884
rect 567160 218872 567166 218884
rect 582346 218872 582374 218980
rect 597738 218968 597744 218980
rect 597796 218968 597802 219020
rect 567160 218844 582374 218872
rect 567160 218832 567166 218844
rect 587158 218832 587164 218884
rect 587216 218872 587222 218884
rect 596818 218872 596824 218884
rect 587216 218844 596824 218872
rect 587216 218832 587222 218844
rect 596818 218832 596824 218844
rect 596876 218832 596882 218884
rect 519078 218804 519084 218816
rect 514726 218776 519084 218804
rect 519078 218764 519084 218776
rect 519136 218764 519142 218816
rect 524414 218764 524420 218816
rect 524472 218804 524478 218816
rect 533890 218804 533896 218816
rect 524472 218776 533896 218804
rect 524472 218764 524478 218776
rect 533890 218764 533896 218776
rect 533948 218764 533954 218816
rect 333698 218696 333704 218748
rect 333756 218736 333762 218748
rect 352558 218736 352564 218748
rect 333756 218708 352564 218736
rect 333756 218696 333762 218708
rect 352558 218696 352564 218708
rect 352616 218696 352622 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 367646 218736 367652 218748
rect 353812 218708 367652 218736
rect 353812 218696 353818 218708
rect 367646 218696 367652 218708
rect 367704 218696 367710 218748
rect 376938 218696 376944 218748
rect 376996 218736 377002 218748
rect 385678 218736 385684 218748
rect 376996 218708 385684 218736
rect 376996 218696 377002 218708
rect 385678 218696 385684 218708
rect 385736 218696 385742 218748
rect 386046 218696 386052 218748
rect 386104 218736 386110 218748
rect 396626 218736 396632 218748
rect 386104 218708 396632 218736
rect 386104 218696 386110 218708
rect 396626 218696 396632 218708
rect 396684 218696 396690 218748
rect 402606 218696 402612 218748
rect 402664 218736 402670 218748
rect 409046 218736 409052 218748
rect 402664 218708 409052 218736
rect 402664 218696 402670 218708
rect 409046 218696 409052 218708
rect 409104 218696 409110 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 482922 218696 482928 218748
rect 482980 218736 482986 218748
rect 485314 218736 485320 218748
rect 482980 218708 485320 218736
rect 482980 218696 482986 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 502794 218696 502800 218748
rect 502852 218736 502858 218748
rect 503162 218736 503168 218748
rect 502852 218708 503168 218736
rect 502852 218696 502858 218708
rect 503162 218696 503168 218708
rect 503220 218736 503226 218748
rect 503220 218708 505094 218736
rect 503220 218696 503226 218708
rect 320692 218572 331214 218600
rect 320692 218560 320698 218572
rect 388530 218560 388536 218612
rect 388588 218600 388594 218612
rect 393958 218600 393964 218612
rect 388588 218572 393964 218600
rect 388588 218560 388594 218572
rect 393958 218560 393964 218572
rect 394016 218560 394022 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 474734 218560 474740 218612
rect 474792 218600 474798 218612
rect 482830 218600 482836 218612
rect 474792 218572 482836 218600
rect 474792 218560 474798 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 505066 218600 505094 218708
rect 505278 218696 505284 218748
rect 505336 218736 505342 218748
rect 505738 218736 505744 218748
rect 505336 218708 505744 218736
rect 505336 218696 505342 218708
rect 505738 218696 505744 218708
rect 505796 218696 505802 218748
rect 534074 218696 534080 218748
rect 534132 218736 534138 218748
rect 548702 218736 548708 218748
rect 534132 218708 548708 218736
rect 534132 218696 534138 218708
rect 548702 218696 548708 218708
rect 548760 218696 548766 218748
rect 556890 218736 556896 218748
rect 550468 218708 556896 218736
rect 550468 218600 550496 218708
rect 556890 218696 556896 218708
rect 556948 218696 556954 218748
rect 618162 218736 618168 218748
rect 557092 218708 618168 218736
rect 505066 218572 550496 218600
rect 550634 218560 550640 218612
rect 550692 218600 550698 218612
rect 551554 218600 551560 218612
rect 550692 218572 551560 218600
rect 550692 218560 550698 218572
rect 551554 218560 551560 218572
rect 551612 218560 551618 218612
rect 552658 218560 552664 218612
rect 552716 218600 552722 218612
rect 557092 218600 557120 218708
rect 618162 218696 618168 218708
rect 618220 218696 618226 218748
rect 552716 218572 557120 218600
rect 552716 218560 552722 218572
rect 558178 218560 558184 218612
rect 558236 218600 558242 218612
rect 587158 218600 587164 218612
rect 558236 218572 587164 218600
rect 558236 218560 558242 218572
rect 587158 218560 587164 218572
rect 587216 218560 587222 218612
rect 587342 218560 587348 218612
rect 587400 218600 587406 218612
rect 611538 218600 611544 218612
rect 587400 218572 611544 218600
rect 587400 218560 587406 218572
rect 611538 218560 611544 218572
rect 611596 218560 611602 218612
rect 179932 218436 190454 218464
rect 179932 218424 179938 218436
rect 196434 218424 196440 218476
rect 196492 218464 196498 218476
rect 207658 218464 207664 218476
rect 196492 218436 207664 218464
rect 196492 218424 196498 218436
rect 207658 218424 207664 218436
rect 207716 218424 207722 218476
rect 210878 218424 210884 218476
rect 210936 218464 210942 218476
rect 220814 218464 220820 218476
rect 210936 218436 220820 218464
rect 210936 218424 210942 218436
rect 220814 218424 220820 218436
rect 220872 218424 220878 218476
rect 225966 218424 225972 218476
rect 226024 218464 226030 218476
rect 265618 218464 265624 218476
rect 226024 218436 265624 218464
rect 226024 218424 226030 218436
rect 265618 218424 265624 218436
rect 265676 218424 265682 218476
rect 265986 218424 265992 218476
rect 266044 218464 266050 218476
rect 272426 218464 272432 218476
rect 266044 218436 272432 218464
rect 266044 218424 266050 218436
rect 272426 218424 272432 218436
rect 272484 218424 272490 218476
rect 272610 218424 272616 218476
rect 272668 218464 272674 218476
rect 288434 218464 288440 218476
rect 272668 218436 288440 218464
rect 272668 218424 272674 218436
rect 288434 218424 288440 218436
rect 288492 218424 288498 218476
rect 500034 218424 500040 218476
rect 500092 218464 500098 218476
rect 500218 218464 500224 218476
rect 500092 218436 500224 218464
rect 500092 218424 500098 218436
rect 500218 218424 500224 218436
rect 500276 218464 500282 218476
rect 604362 218464 604368 218476
rect 500276 218436 604368 218464
rect 500276 218424 500282 218436
rect 604362 218424 604368 218436
rect 604420 218424 604426 218476
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 120316 218300 122834 218328
rect 120316 218288 120322 218300
rect 136818 218288 136824 218340
rect 136876 218328 136882 218340
rect 139486 218328 139492 218340
rect 136876 218300 139492 218328
rect 136876 218288 136882 218300
rect 139486 218288 139492 218300
rect 139544 218288 139550 218340
rect 172606 218328 172612 218340
rect 142126 218300 172612 218328
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 64138 218192 64144 218204
rect 57480 218164 64144 218192
rect 57480 218152 57486 218164
rect 64138 218152 64144 218164
rect 64196 218152 64202 218204
rect 67266 218152 67272 218204
rect 67324 218192 67330 218204
rect 71038 218192 71044 218204
rect 67324 218164 71044 218192
rect 67324 218152 67330 218164
rect 71038 218152 71044 218164
rect 71096 218152 71102 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 130194 218152 130200 218204
rect 130252 218192 130258 218204
rect 142126 218192 142154 218300
rect 172606 218288 172612 218300
rect 172664 218288 172670 218340
rect 174078 218288 174084 218340
rect 174136 218328 174142 218340
rect 179414 218328 179420 218340
rect 174136 218300 179420 218328
rect 174136 218288 174142 218300
rect 179414 218288 179420 218300
rect 179472 218288 179478 218340
rect 190638 218288 190644 218340
rect 190696 218328 190702 218340
rect 191650 218328 191656 218340
rect 190696 218300 191656 218328
rect 190696 218288 190702 218300
rect 191650 218288 191656 218300
rect 191708 218288 191714 218340
rect 192294 218288 192300 218340
rect 192352 218328 192358 218340
rect 193122 218328 193128 218340
rect 192352 218300 193128 218328
rect 192352 218288 192358 218300
rect 193122 218288 193128 218300
rect 193180 218288 193186 218340
rect 193950 218288 193956 218340
rect 194008 218328 194014 218340
rect 194502 218328 194508 218340
rect 194008 218300 194508 218328
rect 194008 218288 194014 218300
rect 194502 218288 194508 218300
rect 194560 218288 194566 218340
rect 198090 218288 198096 218340
rect 198148 218328 198154 218340
rect 198642 218328 198648 218340
rect 198148 218300 198648 218328
rect 198148 218288 198154 218300
rect 198642 218288 198648 218300
rect 198700 218288 198706 218340
rect 199286 218288 199292 218340
rect 199344 218328 199350 218340
rect 202046 218328 202052 218340
rect 199344 218300 202052 218328
rect 199344 218288 199350 218300
rect 202046 218288 202052 218300
rect 202104 218288 202110 218340
rect 203058 218288 203064 218340
rect 203116 218328 203122 218340
rect 213178 218328 213184 218340
rect 203116 218300 213184 218328
rect 203116 218288 203122 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 219618 218288 219624 218340
rect 219676 218328 219682 218340
rect 258074 218328 258080 218340
rect 219676 218300 258080 218328
rect 219676 218288 219682 218300
rect 258074 218288 258080 218300
rect 258132 218288 258138 218340
rect 365346 218288 365352 218340
rect 365404 218328 365410 218340
rect 370498 218328 370504 218340
rect 365404 218300 370504 218328
rect 365404 218288 365410 218300
rect 370498 218288 370504 218300
rect 370556 218288 370562 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429562 218328 429568 218340
rect 426676 218300 429568 218328
rect 426676 218288 426682 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 510154 218288 510160 218340
rect 510212 218328 510218 218340
rect 616138 218328 616144 218340
rect 510212 218300 616144 218328
rect 510212 218288 510218 218300
rect 616138 218288 616144 218300
rect 616196 218288 616202 218340
rect 130252 218164 142154 218192
rect 130252 218152 130258 218164
rect 142614 218152 142620 218204
rect 142672 218192 142678 218204
rect 143258 218192 143264 218204
rect 142672 218164 143264 218192
rect 142672 218152 142678 218164
rect 143258 218152 143264 218164
rect 143316 218152 143322 218204
rect 145098 218152 145104 218204
rect 145156 218192 145162 218204
rect 146110 218192 146116 218204
rect 145156 218164 146116 218192
rect 145156 218152 145162 218164
rect 146110 218152 146116 218164
rect 146168 218152 146174 218204
rect 159174 218152 159180 218204
rect 159232 218192 159238 218204
rect 160002 218192 160008 218204
rect 159232 218164 160008 218192
rect 159232 218152 159238 218164
rect 160002 218152 160008 218164
rect 160060 218152 160066 218204
rect 160830 218152 160836 218204
rect 160888 218192 160894 218204
rect 161934 218192 161940 218204
rect 160888 218164 161940 218192
rect 160888 218152 160894 218164
rect 161934 218152 161940 218164
rect 161992 218152 161998 218204
rect 164970 218152 164976 218204
rect 165028 218192 165034 218204
rect 165522 218192 165528 218204
rect 165028 218164 165528 218192
rect 165028 218152 165034 218164
rect 165522 218152 165528 218164
rect 165580 218152 165586 218204
rect 167454 218152 167460 218204
rect 167512 218192 167518 218204
rect 168282 218192 168288 218204
rect 167512 218164 168288 218192
rect 167512 218152 167518 218164
rect 168282 218152 168288 218164
rect 168340 218152 168346 218204
rect 169110 218152 169116 218204
rect 169168 218192 169174 218204
rect 169570 218192 169576 218204
rect 169168 218164 169576 218192
rect 169168 218152 169174 218164
rect 169570 218152 169576 218164
rect 169628 218152 169634 218204
rect 169754 218152 169760 218204
rect 169812 218192 169818 218204
rect 201862 218192 201868 218204
rect 169812 218164 201868 218192
rect 169812 218152 169818 218164
rect 201862 218152 201868 218164
rect 201920 218152 201926 218204
rect 202230 218152 202236 218204
rect 202288 218192 202294 218204
rect 202690 218192 202696 218204
rect 202288 218164 202696 218192
rect 202288 218152 202294 218164
rect 202690 218152 202696 218164
rect 202748 218152 202754 218204
rect 208854 218152 208860 218204
rect 208912 218192 208918 218204
rect 209498 218192 209504 218204
rect 208912 218164 209504 218192
rect 208912 218152 208918 218164
rect 209498 218152 209504 218164
rect 209556 218152 209562 218204
rect 210510 218152 210516 218204
rect 210568 218192 210574 218204
rect 211062 218192 211068 218204
rect 210568 218164 211068 218192
rect 210568 218152 210574 218164
rect 211062 218152 211068 218164
rect 211120 218152 211126 218204
rect 211338 218152 211344 218204
rect 211396 218192 211402 218204
rect 214282 218192 214288 218204
rect 211396 218164 214288 218192
rect 211396 218152 211402 218164
rect 214282 218152 214288 218164
rect 214340 218152 214346 218204
rect 214650 218152 214656 218204
rect 214708 218192 214714 218204
rect 215202 218192 215208 218204
rect 214708 218164 215208 218192
rect 214708 218152 214714 218164
rect 215202 218152 215208 218164
rect 215260 218152 215266 218204
rect 215478 218152 215484 218204
rect 215536 218192 215542 218204
rect 216582 218192 216588 218204
rect 215536 218164 216588 218192
rect 215536 218152 215542 218164
rect 216582 218152 216588 218164
rect 216640 218152 216646 218204
rect 218790 218152 218796 218204
rect 218848 218192 218854 218204
rect 219342 218192 219348 218204
rect 218848 218164 219348 218192
rect 218848 218152 218854 218164
rect 219342 218152 219348 218164
rect 219400 218152 219406 218204
rect 225598 218192 225604 218204
rect 221108 218164 225604 218192
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59998 218056 60004 218068
rect 58216 218028 60004 218056
rect 58216 218016 58222 218028
rect 59998 218016 60004 218028
rect 60056 218016 60062 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62022 218056 62028 218068
rect 61528 218028 62028 218056
rect 61528 218016 61534 218028
rect 62022 218016 62028 218028
rect 62080 218016 62086 218068
rect 62298 218016 62304 218068
rect 62356 218056 62362 218068
rect 63402 218056 63408 218068
rect 62356 218028 63408 218056
rect 62356 218016 62362 218028
rect 63402 218016 63408 218028
rect 63460 218016 63466 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66898 218056 66904 218068
rect 65668 218028 66904 218056
rect 65668 218016 65674 218028
rect 66898 218016 66904 218028
rect 66956 218016 66962 218068
rect 68094 218016 68100 218068
rect 68152 218056 68158 218068
rect 68922 218056 68928 218068
rect 68152 218028 68928 218056
rect 68152 218016 68158 218028
rect 68922 218016 68928 218028
rect 68980 218016 68986 218068
rect 69750 218016 69756 218068
rect 69808 218056 69814 218068
rect 70302 218056 70308 218068
rect 69808 218028 70308 218056
rect 69808 218016 69814 218028
rect 70302 218016 70308 218028
rect 70360 218016 70366 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 80514 218016 80520 218068
rect 80572 218056 80578 218068
rect 81434 218056 81440 218068
rect 80572 218028 81440 218056
rect 80572 218016 80578 218028
rect 81434 218016 81440 218028
rect 81492 218016 81498 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 82722 218056 82728 218068
rect 82228 218028 82728 218056
rect 82228 218016 82234 218028
rect 82722 218016 82728 218028
rect 82780 218016 82786 218068
rect 82998 218016 83004 218068
rect 83056 218056 83062 218068
rect 84102 218056 84108 218068
rect 83056 218028 84108 218056
rect 83056 218016 83062 218028
rect 84102 218016 84108 218028
rect 84160 218016 84166 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 90450 218016 90456 218068
rect 90508 218056 90514 218068
rect 91002 218056 91008 218068
rect 90508 218028 91008 218056
rect 90508 218016 90514 218028
rect 91002 218016 91008 218028
rect 91060 218016 91066 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 111978 218016 111984 218068
rect 112036 218056 112042 218068
rect 112806 218056 112812 218068
rect 112036 218028 112812 218056
rect 112036 218016 112042 218028
rect 112806 218016 112812 218028
rect 112864 218016 112870 218068
rect 115290 218016 115296 218068
rect 115348 218056 115354 218068
rect 115842 218056 115848 218068
rect 115348 218028 115848 218056
rect 115348 218016 115354 218028
rect 115842 218016 115848 218028
rect 115900 218016 115906 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 116946 218056 116952 218068
rect 116176 218028 116952 218056
rect 116176 218016 116182 218028
rect 116946 218016 116952 218028
rect 117004 218016 117010 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 123570 218016 123576 218068
rect 123628 218056 123634 218068
rect 124122 218056 124128 218068
rect 123628 218028 124128 218056
rect 123628 218016 123634 218028
rect 124122 218016 124128 218028
rect 124180 218016 124186 218068
rect 126054 218016 126060 218068
rect 126112 218056 126118 218068
rect 126698 218056 126704 218068
rect 126112 218028 126704 218056
rect 126112 218016 126118 218028
rect 126698 218016 126704 218028
rect 126756 218016 126762 218068
rect 131850 218016 131856 218068
rect 131908 218056 131914 218068
rect 132402 218056 132408 218068
rect 131908 218028 132408 218056
rect 131908 218016 131914 218028
rect 132402 218016 132408 218028
rect 132460 218016 132466 218068
rect 132678 218016 132684 218068
rect 132736 218056 132742 218068
rect 133506 218056 133512 218068
rect 132736 218028 133512 218056
rect 132736 218016 132742 218028
rect 133506 218016 133512 218028
rect 133564 218016 133570 218068
rect 134334 218016 134340 218068
rect 134392 218056 134398 218068
rect 134978 218056 134984 218068
rect 134392 218028 134984 218056
rect 134392 218016 134398 218028
rect 134978 218016 134984 218028
rect 135036 218016 135042 218068
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 136542 218056 136548 218068
rect 136048 218028 136548 218056
rect 136048 218016 136054 218028
rect 136542 218016 136548 218028
rect 136600 218016 136606 218068
rect 138474 218016 138480 218068
rect 138532 218056 138538 218068
rect 139118 218056 139124 218068
rect 138532 218028 139124 218056
rect 138532 218016 138538 218028
rect 139118 218016 139124 218028
rect 139176 218016 139182 218068
rect 139486 218016 139492 218068
rect 139544 218056 139550 218068
rect 171410 218056 171416 218068
rect 139544 218028 171416 218056
rect 139544 218016 139550 218028
rect 171410 218016 171416 218028
rect 171468 218016 171474 218068
rect 171594 218016 171600 218068
rect 171652 218056 171658 218068
rect 172330 218056 172336 218068
rect 171652 218028 172336 218056
rect 171652 218016 171658 218028
rect 172330 218016 172336 218028
rect 172388 218016 172394 218068
rect 175734 218016 175740 218068
rect 175792 218056 175798 218068
rect 176470 218056 176476 218068
rect 175792 218028 176476 218056
rect 175792 218016 175798 218028
rect 176470 218016 176476 218028
rect 176528 218016 176534 218068
rect 181530 218016 181536 218068
rect 181588 218056 181594 218068
rect 181990 218056 181996 218068
rect 181588 218028 181996 218056
rect 181588 218016 181594 218028
rect 181990 218016 181996 218028
rect 182048 218016 182054 218068
rect 182358 218016 182364 218068
rect 182416 218056 182422 218068
rect 183462 218056 183468 218068
rect 182416 218028 183468 218056
rect 182416 218016 182422 218028
rect 183462 218016 183468 218028
rect 183520 218016 183526 218068
rect 184842 218016 184848 218068
rect 184900 218056 184906 218068
rect 185486 218056 185492 218068
rect 184900 218028 185492 218056
rect 184900 218016 184906 218028
rect 185486 218016 185492 218028
rect 185544 218016 185550 218068
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 188154 218016 188160 218068
rect 188212 218056 188218 218068
rect 189166 218056 189172 218068
rect 188212 218028 189172 218056
rect 188212 218016 188218 218028
rect 189166 218016 189172 218028
rect 189224 218016 189230 218068
rect 189810 218016 189816 218068
rect 189868 218056 189874 218068
rect 221108 218056 221136 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251726 218192 251732 218204
rect 249484 218164 251732 218192
rect 249484 218152 249490 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 289170 218152 289176 218204
rect 289228 218192 289234 218204
rect 294598 218192 294604 218204
rect 289228 218164 294604 218192
rect 289228 218152 289234 218164
rect 294598 218152 294604 218164
rect 294656 218152 294662 218204
rect 297450 218152 297456 218204
rect 297508 218192 297514 218204
rect 300118 218192 300124 218204
rect 297508 218164 300124 218192
rect 297508 218152 297514 218164
rect 300118 218152 300124 218164
rect 300176 218152 300182 218204
rect 304074 218152 304080 218204
rect 304132 218192 304138 218204
rect 305638 218192 305644 218204
rect 304132 218164 305644 218192
rect 304132 218152 304138 218164
rect 305638 218152 305644 218164
rect 305696 218152 305702 218204
rect 332226 218152 332232 218204
rect 332284 218192 332290 218204
rect 334986 218192 334992 218204
rect 332284 218164 334992 218192
rect 332284 218152 332290 218164
rect 334986 218152 334992 218164
rect 335044 218152 335050 218204
rect 338850 218152 338856 218204
rect 338908 218192 338914 218204
rect 340138 218192 340144 218204
rect 338908 218164 340144 218192
rect 338908 218152 338914 218164
rect 340138 218152 340144 218164
rect 340196 218152 340202 218204
rect 348786 218152 348792 218204
rect 348844 218192 348850 218204
rect 353294 218192 353300 218204
rect 348844 218164 353300 218192
rect 348844 218152 348850 218164
rect 353294 218152 353300 218164
rect 353352 218152 353358 218204
rect 368658 218152 368664 218204
rect 368716 218192 368722 218204
rect 372246 218192 372252 218204
rect 368716 218164 372252 218192
rect 368716 218152 368722 218164
rect 372246 218152 372252 218164
rect 372304 218152 372310 218204
rect 375098 218152 375104 218204
rect 375156 218192 375162 218204
rect 380066 218192 380072 218204
rect 375156 218164 380072 218192
rect 375156 218152 375162 218164
rect 380066 218152 380072 218164
rect 380124 218152 380130 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 394326 218152 394332 218204
rect 394384 218192 394390 218204
rect 402238 218192 402244 218204
rect 394384 218164 402244 218192
rect 394384 218152 394390 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 428458 218192 428464 218204
rect 425848 218164 428464 218192
rect 425848 218152 425854 218164
rect 428458 218152 428464 218164
rect 428516 218152 428522 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 435726 218152 435732 218204
rect 435784 218192 435790 218204
rect 436830 218192 436836 218204
rect 435784 218164 436836 218192
rect 435784 218152 435790 218164
rect 436830 218152 436836 218164
rect 436888 218152 436894 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 498654 218152 498660 218204
rect 498712 218192 498718 218204
rect 503622 218192 503628 218204
rect 498712 218164 503628 218192
rect 498712 218152 498718 218164
rect 503622 218152 503628 218164
rect 503680 218152 503686 218204
rect 505278 218152 505284 218204
rect 505336 218192 505342 218204
rect 605742 218192 605748 218204
rect 505336 218164 605748 218192
rect 505336 218152 505342 218164
rect 605742 218152 605748 218164
rect 605800 218152 605806 218204
rect 648246 218152 648252 218204
rect 648304 218192 648310 218204
rect 654778 218192 654784 218204
rect 648304 218164 654784 218192
rect 648304 218152 648310 218164
rect 654778 218152 654784 218164
rect 654836 218152 654842 218204
rect 189868 218028 221136 218056
rect 189868 218016 189874 218028
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 222562 218056 222568 218068
rect 221332 218028 222568 218056
rect 221332 218016 221338 218028
rect 222562 218016 222568 218028
rect 222620 218016 222626 218068
rect 222930 218016 222936 218068
rect 222988 218056 222994 218068
rect 223482 218056 223488 218068
rect 222988 218028 223488 218056
rect 222988 218016 222994 218028
rect 223482 218016 223488 218028
rect 223540 218016 223546 218068
rect 223758 218016 223764 218068
rect 223816 218056 223822 218068
rect 224586 218056 224592 218068
rect 223816 218028 224592 218056
rect 223816 218016 223822 218028
rect 224586 218016 224592 218028
rect 224644 218016 224650 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 227070 218016 227076 218068
rect 227128 218056 227134 218068
rect 227622 218056 227628 218068
rect 227128 218028 227628 218056
rect 227128 218016 227134 218028
rect 227622 218016 227628 218028
rect 227680 218016 227686 218068
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 230474 218056 230480 218068
rect 229612 218028 230480 218056
rect 229612 218016 229618 218028
rect 230474 218016 230480 218028
rect 230532 218016 230538 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 233694 218016 233700 218068
rect 233752 218056 233758 218068
rect 234614 218056 234620 218068
rect 233752 218028 234620 218056
rect 233752 218016 233758 218028
rect 234614 218016 234620 218028
rect 234672 218016 234678 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 246298 218056 246304 218068
rect 244516 218028 246304 218056
rect 244516 218016 244522 218028
rect 246298 218016 246304 218028
rect 246356 218016 246362 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249610 218056 249616 218068
rect 248656 218028 249616 218056
rect 248656 218016 248662 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252370 218056 252376 218068
rect 251968 218028 252376 218056
rect 251968 218016 251974 218028
rect 252370 218016 252376 218028
rect 252428 218016 252434 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259362 218056 259368 218068
rect 258592 218028 259368 218056
rect 258592 218016 258598 218028
rect 259362 218016 259368 218028
rect 259420 218016 259426 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264882 218056 264888 218068
rect 264388 218028 264888 218056
rect 264388 218016 264394 218028
rect 264882 218016 264888 218028
rect 264940 218016 264946 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 269022 218056 269028 218068
rect 268528 218028 269028 218056
rect 268528 218016 268534 218028
rect 269022 218016 269028 218028
rect 269080 218016 269086 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270218 218056 270224 218068
rect 269356 218028 270224 218056
rect 269356 218016 269362 218028
rect 270218 218016 270224 218028
rect 270276 218016 270282 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 271598 218056 271604 218068
rect 271012 218028 271604 218056
rect 271012 218016 271018 218028
rect 271598 218016 271604 218028
rect 271656 218016 271662 218068
rect 273438 218016 273444 218068
rect 273496 218056 273502 218068
rect 274082 218056 274088 218068
rect 273496 218028 274088 218056
rect 273496 218016 273502 218028
rect 274082 218016 274088 218028
rect 274140 218016 274146 218068
rect 275094 218016 275100 218068
rect 275152 218056 275158 218068
rect 275646 218056 275652 218068
rect 275152 218028 275652 218056
rect 275152 218016 275158 218028
rect 275646 218016 275652 218028
rect 275704 218016 275710 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282454 218056 282460 218068
rect 281776 218028 282460 218056
rect 281776 218016 281782 218028
rect 282454 218016 282460 218028
rect 282512 218016 282518 218068
rect 284202 218016 284208 218068
rect 284260 218056 284266 218068
rect 284846 218056 284852 218068
rect 284260 218028 284852 218056
rect 284260 218016 284266 218028
rect 284846 218016 284852 218028
rect 284904 218016 284910 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288066 218056 288072 218068
rect 287572 218028 288072 218056
rect 287572 218016 287578 218028
rect 288066 218016 288072 218028
rect 288124 218016 288130 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 290826 218056 290832 218068
rect 290056 218028 290832 218056
rect 290056 218016 290062 218028
rect 290826 218016 290832 218028
rect 290884 218016 290890 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 295794 218016 295800 218068
rect 295852 218056 295858 218068
rect 296714 218056 296720 218068
rect 295852 218028 296720 218056
rect 295852 218016 295858 218028
rect 296714 218016 296720 218028
rect 296772 218016 296778 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300762 218056 300768 218068
rect 299992 218028 300768 218056
rect 299992 218016 299998 218028
rect 300762 218016 300768 218028
rect 300820 218016 300826 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308766 218056 308772 218068
rect 308272 218028 308772 218056
rect 308272 218016 308278 218028
rect 308766 218016 308772 218028
rect 308824 218016 308830 218068
rect 310698 218016 310704 218068
rect 310756 218056 310762 218068
rect 311802 218056 311808 218068
rect 310756 218028 311808 218056
rect 310756 218016 310762 218028
rect 311802 218016 311808 218028
rect 311860 218016 311866 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315850 218056 315856 218068
rect 314896 218028 315856 218056
rect 314896 218016 314902 218028
rect 315850 218016 315856 218028
rect 315908 218016 315914 218068
rect 316494 218016 316500 218068
rect 316552 218056 316558 218068
rect 317138 218056 317144 218068
rect 316552 218028 317144 218056
rect 316552 218016 316558 218028
rect 317138 218016 317144 218028
rect 317196 218016 317202 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319990 218056 319996 218068
rect 319036 218028 319996 218056
rect 319036 218016 319042 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335262 218056 335268 218068
rect 334768 218028 335268 218056
rect 334768 218016 334774 218028
rect 335262 218016 335268 218028
rect 335320 218016 335326 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 336366 218056 336372 218068
rect 335596 218028 336372 218056
rect 335596 218016 335602 218028
rect 336366 218016 336372 218028
rect 336424 218016 336430 218068
rect 337194 218016 337200 218068
rect 337252 218056 337258 218068
rect 337838 218056 337844 218068
rect 337252 218028 337844 218056
rect 337252 218016 337258 218028
rect 337838 218016 337844 218028
rect 337896 218016 337902 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 342990 218016 342996 218068
rect 343048 218056 343054 218068
rect 343450 218056 343456 218068
rect 343048 218028 343456 218056
rect 343048 218016 343054 218028
rect 343450 218016 343456 218028
rect 343508 218016 343514 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 346394 218056 346400 218068
rect 345532 218028 346400 218056
rect 345532 218016 345538 218028
rect 346394 218016 346400 218028
rect 346452 218016 346458 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 351270 218016 351276 218068
rect 351328 218056 351334 218068
rect 351730 218056 351736 218068
rect 351328 218028 351736 218056
rect 351328 218016 351334 218028
rect 351730 218016 351736 218028
rect 351788 218016 351794 218068
rect 352098 218016 352104 218068
rect 352156 218056 352162 218068
rect 354398 218056 354404 218068
rect 352156 218028 354404 218056
rect 352156 218016 352162 218028
rect 354398 218016 354404 218028
rect 354456 218016 354462 218068
rect 355410 218016 355416 218068
rect 355468 218056 355474 218068
rect 355962 218056 355968 218068
rect 355468 218028 355968 218056
rect 355468 218016 355474 218028
rect 355962 218016 355968 218028
rect 356020 218016 356026 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357250 218056 357256 218068
rect 356296 218028 357256 218056
rect 356296 218016 356302 218028
rect 357250 218016 357256 218028
rect 357308 218016 357314 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361298 218056 361304 218068
rect 360436 218028 361304 218056
rect 360436 218016 360442 218028
rect 361298 218016 361304 218028
rect 361356 218016 361362 218068
rect 364518 218016 364524 218068
rect 364576 218056 364582 218068
rect 365530 218056 365536 218068
rect 364576 218028 365536 218056
rect 364576 218016 364582 218028
rect 365530 218016 365536 218028
rect 365588 218016 365594 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366726 218056 366732 218068
rect 366232 218028 366732 218056
rect 366232 218016 366238 218028
rect 366726 218016 366732 218028
rect 366784 218016 366790 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372430 218056 372436 218068
rect 372028 218028 372436 218056
rect 372028 218016 372034 218028
rect 372430 218016 372436 218028
rect 372488 218016 372494 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373810 218056 373816 218068
rect 372856 218028 373816 218056
rect 372856 218016 372862 218028
rect 373810 218016 373816 218028
rect 373868 218016 373874 218068
rect 374454 218016 374460 218068
rect 374512 218056 374518 218068
rect 375282 218056 375288 218068
rect 374512 218028 375288 218056
rect 374512 218016 374518 218028
rect 375282 218016 375288 218028
rect 375340 218016 375346 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 380250 218016 380256 218068
rect 380308 218056 380314 218068
rect 380710 218056 380716 218068
rect 380308 218028 380716 218056
rect 380308 218016 380314 218028
rect 380710 218016 380716 218028
rect 380768 218016 380774 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 384390 218016 384396 218068
rect 384448 218056 384454 218068
rect 384942 218056 384948 218068
rect 384448 218028 384948 218056
rect 384448 218016 384454 218028
rect 384942 218016 384948 218028
rect 385000 218016 385006 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386322 218056 386328 218068
rect 385276 218028 386328 218056
rect 385276 218016 385282 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390094 218056 390100 218068
rect 389416 218028 390100 218056
rect 389416 218016 389422 218028
rect 390094 218016 390100 218028
rect 390152 218016 390158 218068
rect 391014 218016 391020 218068
rect 391072 218056 391078 218068
rect 391566 218056 391572 218068
rect 391072 218028 391572 218056
rect 391072 218016 391078 218028
rect 391566 218016 391572 218028
rect 391624 218016 391630 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 398466 218056 398472 218068
rect 397696 218028 398472 218056
rect 397696 218016 397702 218028
rect 398466 218016 398472 218028
rect 398524 218016 398530 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 401502 218056 401508 218068
rect 401008 218028 401508 218056
rect 401008 218016 401014 218028
rect 401502 218016 401508 218028
rect 401560 218016 401566 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 418338 218016 418344 218068
rect 418396 218056 418402 218068
rect 419442 218056 419448 218068
rect 418396 218028 419448 218056
rect 418396 218016 418402 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434898 218016 434904 218068
rect 434956 218056 434962 218068
rect 436278 218056 436284 218068
rect 434956 218028 436284 218056
rect 434956 218016 434962 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436462 218016 436468 218068
rect 436520 218056 436526 218068
rect 437750 218056 437756 218068
rect 436520 218028 437756 218056
rect 436520 218016 436526 218028
rect 437750 218016 437756 218028
rect 437808 218016 437814 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 483566 218016 483572 218068
rect 483624 218056 483630 218068
rect 486970 218056 486976 218068
rect 483624 218028 486976 218056
rect 483624 218016 483630 218028
rect 486970 218016 486976 218028
rect 487028 218056 487034 218068
rect 519446 218056 519452 218068
rect 487028 218028 519452 218056
rect 487028 218016 487034 218028
rect 519446 218016 519452 218028
rect 519504 218016 519510 218068
rect 520182 218016 520188 218068
rect 520240 218056 520246 218068
rect 524782 218056 524788 218068
rect 520240 218028 524788 218056
rect 520240 218016 520246 218028
rect 524782 218016 524788 218028
rect 524840 218016 524846 218068
rect 539686 218016 539692 218068
rect 539744 218056 539750 218068
rect 563008 218056 563014 218068
rect 539744 218028 563014 218056
rect 539744 218016 539750 218028
rect 563008 218016 563014 218028
rect 563066 218016 563072 218068
rect 573174 218016 573180 218068
rect 573232 218056 573238 218068
rect 582282 218056 582288 218068
rect 573232 218028 582288 218056
rect 573232 218016 573238 218028
rect 582282 218016 582288 218028
rect 582340 218016 582346 218068
rect 655422 218016 655428 218068
rect 655480 218056 655486 218068
rect 656158 218056 656164 218068
rect 655480 218028 656164 218056
rect 655480 218016 655486 218028
rect 656158 218016 656164 218028
rect 656216 218016 656222 218068
rect 534074 217988 534080 218000
rect 525628 217960 534080 217988
rect 518894 217880 518900 217932
rect 518952 217920 518958 217932
rect 524598 217920 524604 217932
rect 518952 217892 524604 217920
rect 518952 217880 518958 217892
rect 524598 217880 524604 217892
rect 524656 217880 524662 217932
rect 514938 217744 514944 217796
rect 514996 217784 515002 217796
rect 518710 217784 518716 217796
rect 514996 217756 518716 217784
rect 514996 217744 515002 217756
rect 518710 217744 518716 217756
rect 518768 217744 518774 217796
rect 518894 217744 518900 217796
rect 518952 217784 518958 217796
rect 525628 217784 525656 217960
rect 534074 217948 534080 217960
rect 534132 217948 534138 218000
rect 538398 217948 538404 218000
rect 538456 217988 538462 218000
rect 538950 217988 538956 218000
rect 538456 217960 538956 217988
rect 538456 217948 538462 217960
rect 538950 217948 538956 217960
rect 539008 217988 539014 218000
rect 539502 217988 539508 218000
rect 539008 217960 539508 217988
rect 539008 217948 539014 217960
rect 539502 217948 539508 217960
rect 539560 217948 539566 218000
rect 563146 217948 563152 218000
rect 563204 217988 563210 218000
rect 568298 217988 568304 218000
rect 563204 217960 568304 217988
rect 563204 217948 563210 217960
rect 568298 217948 568304 217960
rect 568356 217948 568362 218000
rect 568666 217948 568672 218000
rect 568724 217988 568730 218000
rect 572162 217988 572168 218000
rect 568724 217960 572168 217988
rect 568724 217948 568730 217960
rect 572162 217948 572168 217960
rect 572220 217948 572226 218000
rect 572300 217948 572306 218000
rect 572358 217988 572364 218000
rect 572358 217960 572944 217988
rect 572358 217948 572364 217960
rect 572916 217920 572944 217960
rect 572916 217892 573036 217920
rect 525978 217812 525984 217864
rect 526036 217852 526042 217864
rect 526714 217852 526720 217864
rect 526036 217824 526720 217852
rect 526036 217812 526042 217824
rect 526714 217812 526720 217824
rect 526772 217812 526778 217864
rect 534166 217812 534172 217864
rect 534224 217852 534230 217864
rect 563238 217852 563244 217864
rect 534224 217824 563244 217852
rect 534224 217812 534230 217824
rect 563238 217812 563244 217824
rect 563296 217812 563302 217864
rect 563422 217812 563428 217864
rect 563480 217852 563486 217864
rect 567562 217852 567568 217864
rect 563480 217824 567568 217852
rect 563480 217812 563486 217824
rect 567562 217812 567568 217824
rect 567620 217812 567626 217864
rect 572714 217852 572720 217864
rect 567948 217824 572720 217852
rect 567948 217784 567976 217824
rect 572714 217812 572720 217824
rect 572772 217812 572778 217864
rect 573008 217852 573036 217892
rect 610066 217852 610072 217864
rect 573008 217824 610072 217852
rect 610066 217812 610072 217824
rect 610124 217812 610130 217864
rect 518952 217756 525656 217784
rect 567764 217756 567976 217784
rect 518952 217744 518958 217756
rect 528278 217676 528284 217728
rect 528336 217716 528342 217728
rect 539042 217716 539048 217728
rect 528336 217688 539048 217716
rect 528336 217676 528342 217688
rect 539042 217676 539048 217688
rect 539100 217676 539106 217728
rect 539502 217676 539508 217728
rect 539560 217716 539566 217728
rect 567764 217716 567792 217756
rect 539560 217688 567792 217716
rect 539560 217676 539566 217688
rect 568114 217676 568120 217728
rect 568172 217716 568178 217728
rect 572070 217716 572076 217728
rect 568172 217688 572076 217716
rect 568172 217676 568178 217688
rect 572070 217676 572076 217688
rect 572128 217676 572134 217728
rect 572254 217676 572260 217728
rect 572312 217716 572318 217728
rect 572714 217716 572720 217728
rect 572312 217688 572720 217716
rect 572312 217676 572318 217688
rect 572714 217676 572720 217688
rect 572772 217676 572778 217728
rect 573082 217676 573088 217728
rect 573140 217716 573146 217728
rect 577314 217716 577320 217728
rect 573140 217688 577320 217716
rect 573140 217676 573146 217688
rect 577314 217676 577320 217688
rect 577372 217676 577378 217728
rect 582098 217676 582104 217728
rect 582156 217716 582162 217728
rect 586882 217716 586888 217728
rect 582156 217688 586888 217716
rect 582156 217676 582162 217688
rect 586882 217676 586888 217688
rect 586940 217676 586946 217728
rect 592034 217676 592040 217728
rect 592092 217716 592098 217728
rect 594978 217716 594984 217728
rect 592092 217688 594984 217716
rect 592092 217676 592098 217688
rect 594978 217676 594984 217688
rect 595036 217676 595042 217728
rect 605742 217676 605748 217728
rect 605800 217716 605806 217728
rect 615034 217716 615040 217728
rect 605800 217688 615040 217716
rect 605800 217676 605806 217688
rect 615034 217676 615040 217688
rect 615092 217676 615098 217728
rect 517698 217608 517704 217660
rect 517756 217648 517762 217660
rect 517756 217620 519308 217648
rect 517756 217608 517762 217620
rect 518342 217472 518348 217524
rect 518400 217512 518406 217524
rect 519078 217512 519084 217524
rect 518400 217484 519084 217512
rect 518400 217472 518406 217484
rect 519078 217472 519084 217484
rect 519136 217472 519142 217524
rect 519280 217512 519308 217620
rect 526714 217540 526720 217592
rect 526772 217580 526778 217592
rect 526772 217552 596864 217580
rect 526772 217540 526778 217552
rect 519280 217484 524414 217512
rect 128538 217404 128544 217456
rect 128596 217444 128602 217456
rect 199102 217444 199108 217456
rect 128596 217416 199108 217444
rect 128596 217404 128602 217416
rect 199102 217404 199108 217416
rect 199160 217404 199166 217456
rect 524386 217444 524414 217484
rect 534166 217444 534172 217456
rect 524386 217416 534172 217444
rect 534166 217404 534172 217416
rect 534224 217404 534230 217456
rect 596634 217444 596640 217456
rect 538876 217416 596640 217444
rect 535914 217336 535920 217388
rect 535972 217376 535978 217388
rect 538674 217376 538680 217388
rect 535972 217348 538680 217376
rect 535972 217336 535978 217348
rect 538674 217336 538680 217348
rect 538732 217336 538738 217388
rect 178402 217308 178408 217320
rect 113146 217280 178408 217308
rect 103652 217200 103658 217252
rect 103710 217240 103716 217252
rect 113146 217240 113174 217280
rect 178402 217268 178408 217280
rect 178460 217268 178466 217320
rect 103710 217212 113174 217240
rect 103710 217200 103716 217212
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 477586 217200 477592 217252
rect 477644 217240 477650 217252
rect 478736 217240 478742 217252
rect 477644 217212 478742 217240
rect 477644 217200 477650 217212
rect 478736 217200 478742 217212
rect 478794 217200 478800 217252
rect 510614 217200 510620 217252
rect 510672 217240 510678 217252
rect 511856 217240 511862 217252
rect 510672 217212 511862 217240
rect 510672 217200 510678 217212
rect 511856 217200 511862 217212
rect 511914 217200 511920 217252
rect 523034 217200 523040 217252
rect 523092 217240 523098 217252
rect 524276 217240 524282 217252
rect 523092 217212 524282 217240
rect 523092 217200 523098 217212
rect 524276 217200 524282 217212
rect 524334 217200 524340 217252
rect 533338 217200 533344 217252
rect 533396 217240 533402 217252
rect 538876 217240 538904 217416
rect 596634 217404 596640 217416
rect 596692 217404 596698 217456
rect 596836 217444 596864 217552
rect 602062 217540 602068 217592
rect 602120 217580 602126 217592
rect 613378 217580 613384 217592
rect 602120 217552 613384 217580
rect 602120 217540 602126 217552
rect 613378 217540 613384 217552
rect 613436 217540 613442 217592
rect 602338 217444 602344 217456
rect 596836 217416 602344 217444
rect 602338 217404 602344 217416
rect 602396 217404 602402 217456
rect 604362 217404 604368 217456
rect 604420 217444 604426 217456
rect 614114 217444 614120 217456
rect 604420 217416 614120 217444
rect 604420 217404 604426 217416
rect 614114 217404 614120 217416
rect 614172 217404 614178 217456
rect 539042 217268 539048 217320
rect 539100 217308 539106 217320
rect 603074 217308 603080 217320
rect 539100 217280 603080 217308
rect 539100 217268 539106 217280
rect 603074 217268 603080 217280
rect 603132 217268 603138 217320
rect 612734 217268 612740 217320
rect 612792 217308 612798 217320
rect 629386 217308 629392 217320
rect 612792 217280 629392 217308
rect 612792 217268 612798 217280
rect 629386 217268 629392 217280
rect 629444 217268 629450 217320
rect 533396 217212 538904 217240
rect 533396 217200 533402 217212
rect 539042 217132 539048 217184
rect 539100 217172 539106 217184
rect 604546 217172 604552 217184
rect 539100 217144 604552 217172
rect 539100 217132 539106 217144
rect 604546 217132 604552 217144
rect 604604 217132 604610 217184
rect 523448 217064 523454 217116
rect 523506 217104 523512 217116
rect 523506 217064 523540 217104
rect 523512 217036 523540 217064
rect 575474 217036 575480 217048
rect 523512 217008 575480 217036
rect 575474 216996 575480 217008
rect 575532 216996 575538 217048
rect 577314 216996 577320 217048
rect 577372 217036 577378 217048
rect 605098 217036 605104 217048
rect 577372 217008 605104 217036
rect 577372 216996 577378 217008
rect 605098 216996 605104 217008
rect 605156 216996 605162 217048
rect 582374 216860 582380 216912
rect 582432 216900 582438 216912
rect 592034 216900 592040 216912
rect 582432 216872 592040 216900
rect 582432 216860 582438 216872
rect 592034 216860 592040 216872
rect 592092 216860 592098 216912
rect 596634 216860 596640 216912
rect 596692 216900 596698 216912
rect 603994 216900 604000 216912
rect 596692 216872 604000 216900
rect 596692 216860 596698 216872
rect 603994 216860 604000 216872
rect 604052 216860 604058 216912
rect 618162 216656 618168 216708
rect 618220 216696 618226 216708
rect 623866 216696 623872 216708
rect 618220 216668 623872 216696
rect 618220 216656 618226 216668
rect 623866 216656 623872 216668
rect 623924 216656 623930 216708
rect 597738 216044 597744 216096
rect 597796 216084 597802 216096
rect 626074 216084 626080 216096
rect 597796 216056 626080 216084
rect 597796 216044 597802 216056
rect 626074 216044 626080 216056
rect 626132 216044 626138 216096
rect 596818 215908 596824 215960
rect 596876 215948 596882 215960
rect 625246 215948 625252 215960
rect 596876 215920 625252 215948
rect 596876 215908 596882 215920
rect 625246 215908 625252 215920
rect 625304 215908 625310 215960
rect 577038 215840 577044 215892
rect 577096 215880 577102 215892
rect 582558 215880 582564 215892
rect 577096 215852 582564 215880
rect 577096 215840 577102 215852
rect 582558 215840 582564 215852
rect 582616 215840 582622 215892
rect 594610 215568 594616 215620
rect 594668 215608 594674 215620
rect 598474 215608 598480 215620
rect 594668 215580 598480 215608
rect 594668 215568 594674 215580
rect 598474 215568 598480 215580
rect 598532 215568 598538 215620
rect 596174 215296 596180 215348
rect 596232 215336 596238 215348
rect 596818 215336 596824 215348
rect 596232 215308 596824 215336
rect 596232 215296 596238 215308
rect 596818 215296 596824 215308
rect 596876 215296 596882 215348
rect 611538 215296 611544 215348
rect 611596 215336 611602 215348
rect 614482 215336 614488 215348
rect 611596 215308 614488 215336
rect 611596 215296 611602 215308
rect 614482 215296 614488 215308
rect 614540 215296 614546 215348
rect 676030 215092 676036 215144
rect 676088 215132 676094 215144
rect 677594 215132 677600 215144
rect 676088 215104 677600 215132
rect 676088 215092 676094 215104
rect 677594 215092 677600 215104
rect 677652 215092 677658 215144
rect 575842 214956 575848 215008
rect 575900 214996 575906 215008
rect 612274 214996 612280 215008
rect 575900 214968 612280 214996
rect 575900 214956 575906 214968
rect 612274 214956 612280 214968
rect 612332 214956 612338 215008
rect 574462 214820 574468 214872
rect 574520 214860 574526 214872
rect 612826 214860 612832 214872
rect 574520 214832 612832 214860
rect 574520 214820 574526 214832
rect 612826 214820 612832 214832
rect 612884 214820 612890 214872
rect 675846 214820 675852 214872
rect 675904 214860 675910 214872
rect 677318 214860 677324 214872
rect 675904 214832 677324 214860
rect 675904 214820 675910 214832
rect 677318 214820 677324 214832
rect 677376 214820 677382 214872
rect 575658 214684 575664 214736
rect 575716 214724 575722 214736
rect 622302 214724 622308 214736
rect 575716 214696 622308 214724
rect 575716 214684 575722 214696
rect 622302 214684 622308 214696
rect 622360 214684 622366 214736
rect 628558 214684 628564 214736
rect 628616 214724 628622 214736
rect 632882 214724 632888 214736
rect 628616 214696 632888 214724
rect 628616 214684 628622 214696
rect 632882 214684 632888 214696
rect 632940 214684 632946 214736
rect 652846 214684 652852 214736
rect 652904 214724 652910 214736
rect 661678 214724 661684 214736
rect 652904 214696 661684 214724
rect 652904 214684 652910 214696
rect 661678 214684 661684 214696
rect 661736 214684 661742 214736
rect 574094 214548 574100 214600
rect 574152 214588 574158 214600
rect 574152 214560 605834 214588
rect 574152 214548 574158 214560
rect 605806 214452 605834 214560
rect 607306 214548 607312 214600
rect 607364 214588 607370 214600
rect 607858 214588 607864 214600
rect 607364 214560 607864 214588
rect 607364 214548 607370 214560
rect 607858 214548 607864 214560
rect 607916 214548 607922 214600
rect 608778 214548 608784 214600
rect 608836 214588 608842 214600
rect 609514 214588 609520 214600
rect 608836 214560 609520 214588
rect 608836 214548 608842 214560
rect 609514 214548 609520 214560
rect 609572 214548 609578 214600
rect 621106 214548 621112 214600
rect 621164 214588 621170 214600
rect 621658 214588 621664 214600
rect 621164 214560 621664 214588
rect 621164 214548 621170 214560
rect 621658 214548 621664 214560
rect 621716 214548 621722 214600
rect 622486 214548 622492 214600
rect 622544 214588 622550 214600
rect 623314 214588 623320 214600
rect 622544 214560 623320 214588
rect 622544 214548 622550 214560
rect 623314 214548 623320 214560
rect 623372 214548 623378 214600
rect 627914 214548 627920 214600
rect 627972 214588 627978 214600
rect 628834 214588 628840 214600
rect 627972 214560 628840 214588
rect 627972 214548 627978 214560
rect 628834 214548 628840 214560
rect 628892 214548 628898 214600
rect 636286 214548 636292 214600
rect 636344 214588 636350 214600
rect 639598 214588 639604 214600
rect 636344 214560 639604 214588
rect 636344 214548 636350 214560
rect 639598 214548 639604 214560
rect 639656 214548 639662 214600
rect 648430 214548 648436 214600
rect 648488 214588 648494 214600
rect 658918 214588 658924 214600
rect 648488 214560 658924 214588
rect 648488 214548 648494 214560
rect 658918 214548 658924 214560
rect 658976 214548 658982 214600
rect 627178 214452 627184 214464
rect 605806 214424 627184 214452
rect 627178 214412 627184 214424
rect 627236 214412 627242 214464
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 41690 213976 41696 213988
rect 35860 213948 41696 213976
rect 35860 213936 35866 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 627730 213936 627736 213988
rect 627788 213976 627794 213988
rect 631594 213976 631600 213988
rect 627788 213948 631600 213976
rect 627788 213936 627794 213948
rect 631594 213936 631600 213948
rect 631652 213936 631658 213988
rect 637574 213868 637580 213920
rect 637632 213908 637638 213920
rect 638218 213908 638224 213920
rect 637632 213880 638224 213908
rect 637632 213868 637638 213880
rect 638218 213868 638224 213880
rect 638276 213868 638282 213920
rect 645486 213868 645492 213920
rect 645544 213908 645550 213920
rect 646130 213908 646136 213920
rect 645544 213880 646136 213908
rect 645544 213868 645550 213880
rect 646130 213868 646136 213880
rect 646188 213868 646194 213920
rect 648614 213868 648620 213920
rect 648672 213908 648678 213920
rect 649258 213908 649264 213920
rect 648672 213880 649264 213908
rect 648672 213868 648678 213880
rect 649258 213868 649264 213880
rect 649316 213868 649322 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 638034 213732 638040 213784
rect 638092 213772 638098 213784
rect 641162 213772 641168 213784
rect 638092 213744 641168 213772
rect 638092 213732 638098 213744
rect 641162 213732 641168 213744
rect 641220 213732 641226 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 663058 213772 663064 213784
rect 661000 213744 663064 213772
rect 661000 213732 661006 213744
rect 663058 213732 663064 213744
rect 663116 213732 663122 213784
rect 641622 213596 641628 213648
rect 641680 213636 641686 213648
rect 650638 213636 650644 213648
rect 641680 213608 650644 213636
rect 641680 213596 641686 213608
rect 650638 213596 650644 213608
rect 650696 213596 650702 213648
rect 651834 213596 651840 213648
rect 651892 213636 651898 213648
rect 657538 213636 657544 213648
rect 651892 213608 657544 213636
rect 651892 213596 651898 213608
rect 657538 213596 657544 213608
rect 657596 213596 657602 213648
rect 676030 213596 676036 213648
rect 676088 213636 676094 213648
rect 676950 213636 676956 213648
rect 676088 213608 676956 213636
rect 676088 213596 676094 213608
rect 676950 213596 676956 213608
rect 677008 213596 677014 213648
rect 635550 213460 635556 213512
rect 635608 213500 635614 213512
rect 652386 213500 652392 213512
rect 635608 213472 652392 213500
rect 635608 213460 635614 213472
rect 652386 213460 652392 213472
rect 652444 213460 652450 213512
rect 663150 213460 663156 213512
rect 663208 213500 663214 213512
rect 665818 213500 665824 213512
rect 663208 213472 665824 213500
rect 663208 213460 663214 213472
rect 665818 213460 665824 213472
rect 665876 213460 665882 213512
rect 575474 213324 575480 213376
rect 575532 213364 575538 213376
rect 601786 213364 601792 213376
rect 575532 213336 601792 213364
rect 575532 213324 575538 213336
rect 601786 213324 601792 213336
rect 601844 213324 601850 213376
rect 640242 213324 640248 213376
rect 640300 213364 640306 213376
rect 660758 213364 660764 213376
rect 640300 213336 660764 213364
rect 640300 213324 640306 213336
rect 660758 213324 660764 213336
rect 660816 213324 660822 213376
rect 574278 213188 574284 213240
rect 574336 213228 574342 213240
rect 615586 213228 615592 213240
rect 574336 213200 615592 213228
rect 574336 213188 574342 213200
rect 615586 213188 615592 213200
rect 615644 213188 615650 213240
rect 642174 213188 642180 213240
rect 642232 213228 642238 213240
rect 642232 213200 644474 213228
rect 642232 213188 642238 213200
rect 644446 213160 644474 213200
rect 664162 213160 664168 213172
rect 644446 213132 664168 213160
rect 664162 213120 664168 213132
rect 664220 213120 664226 213172
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 632698 212712 632704 212764
rect 632756 212752 632762 212764
rect 634354 212752 634360 212764
rect 632756 212724 634360 212752
rect 632756 212712 632762 212724
rect 634354 212712 634360 212724
rect 634412 212712 634418 212764
rect 658734 212712 658740 212764
rect 658792 212752 658798 212764
rect 659470 212752 659476 212764
rect 658792 212724 659476 212752
rect 658792 212712 658798 212724
rect 659470 212712 659476 212724
rect 659528 212712 659534 212764
rect 600314 212372 600320 212424
rect 600372 212412 600378 212424
rect 601234 212412 601240 212424
rect 600372 212384 601240 212412
rect 600372 212372 600378 212384
rect 601234 212372 601240 212384
rect 601292 212372 601298 212424
rect 35618 211284 35624 211336
rect 35676 211324 35682 211336
rect 41690 211324 41696 211336
rect 35676 211296 41696 211324
rect 35676 211284 35682 211296
rect 41690 211284 41696 211296
rect 41748 211284 41754 211336
rect 578234 211284 578240 211336
rect 578292 211324 578298 211336
rect 580442 211324 580448 211336
rect 578292 211296 580448 211324
rect 578292 211284 578298 211296
rect 580442 211284 580448 211296
rect 580500 211284 580506 211336
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 41690 211188 41696 211200
rect 35860 211160 41696 211188
rect 35860 211148 35866 211160
rect 41690 211148 41696 211160
rect 41748 211148 41754 211200
rect 600498 211012 600504 211064
rect 600556 211052 600562 211064
rect 600866 211052 600872 211064
rect 600556 211024 600872 211052
rect 600556 211012 600562 211024
rect 600866 211012 600872 211024
rect 600924 211012 600930 211064
rect 619634 211012 619640 211064
rect 619692 211052 619698 211064
rect 620002 211052 620008 211064
rect 619692 211024 620008 211052
rect 619692 211012 619698 211024
rect 620002 211012 620008 211024
rect 620060 211012 620066 211064
rect 35802 209788 35808 209840
rect 35860 209828 35866 209840
rect 41322 209828 41328 209840
rect 35860 209800 41328 209828
rect 35860 209788 35866 209800
rect 41322 209788 41328 209800
rect 41380 209788 41386 209840
rect 579246 209788 579252 209840
rect 579304 209828 579310 209840
rect 581730 209828 581736 209840
rect 579304 209800 581736 209828
rect 579304 209788 579310 209800
rect 581730 209788 581736 209800
rect 581788 209788 581794 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 581546 208564 581552 208616
rect 581604 208604 581610 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652018 209516 652024 209568
rect 652076 209516 652082 209568
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 666830 209556 666836 209568
rect 652260 209528 666836 209556
rect 652260 209516 652266 209528
rect 666830 209516 666836 209528
rect 666888 209516 666894 209568
rect 652036 209420 652064 209516
rect 652036 209392 654134 209420
rect 654106 209080 654134 209392
rect 666646 209080 666652 209092
rect 654106 209052 666652 209080
rect 666646 209040 666652 209052
rect 666704 209040 666710 209092
rect 581604 208576 625154 208604
rect 581604 208564 581610 208576
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 580442 207612 580448 207664
rect 580500 207652 580506 207664
rect 589458 207652 589464 207664
rect 580500 207624 589464 207652
rect 580500 207612 580506 207624
rect 589458 207612 589464 207624
rect 589516 207612 589522 207664
rect 581730 206252 581736 206304
rect 581788 206292 581794 206304
rect 589642 206292 589648 206304
rect 581788 206264 589648 206292
rect 581788 206252 581794 206264
rect 589642 206252 589648 206264
rect 589700 206252 589706 206304
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 667934 199180 667940 199232
rect 667992 199220 667998 199232
rect 670786 199220 670792 199232
rect 667992 199192 670792 199220
rect 667992 199180 667998 199192
rect 670786 199180 670792 199192
rect 670844 199180 670850 199232
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 667934 194284 667940 194336
rect 667992 194324 667998 194336
rect 670786 194324 670792 194336
rect 667992 194296 670792 194324
rect 667992 194284 667998 194296
rect 670786 194284 670792 194296
rect 670844 194284 670850 194336
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 667934 189388 667940 189440
rect 667992 189428 667998 189440
rect 670786 189428 670792 189440
rect 667992 189400 670792 189428
rect 667992 189388 667998 189400
rect 670786 189388 670792 189400
rect 670844 189388 670850 189440
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 669222 184492 669228 184544
rect 669280 184532 669286 184544
rect 669774 184532 669780 184544
rect 669280 184504 669780 184532
rect 669280 184492 669286 184504
rect 669774 184492 669780 184504
rect 669832 184492 669838 184544
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 667934 174700 667940 174752
rect 667992 174740 667998 174752
rect 670234 174740 670240 174752
rect 667992 174712 670240 174740
rect 667992 174700 667998 174712
rect 670234 174700 670240 174712
rect 670292 174700 670298 174752
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 667934 169668 667940 169720
rect 667992 169708 667998 169720
rect 670050 169708 670056 169720
rect 667992 169680 670056 169708
rect 667992 169668 667998 169680
rect 670050 169668 670056 169680
rect 670108 169668 670114 169720
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 675846 162528 675852 162580
rect 675904 162568 675910 162580
rect 680998 162568 681004 162580
rect 675904 162540 681004 162568
rect 675904 162528 675910 162540
rect 680998 162528 681004 162540
rect 681056 162528 681062 162580
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580442 151784 580448 151836
rect 580500 151824 580506 151836
rect 589458 151824 589464 151836
rect 580500 151796 589464 151824
rect 580500 151784 580506 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 668302 150220 668308 150272
rect 668360 150260 668366 150272
rect 670786 150260 670792 150272
rect 668360 150232 670792 150260
rect 668360 150220 668366 150232
rect 670786 150220 670792 150232
rect 670844 150220 670850 150272
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 579246 145256 579252 145308
rect 579304 145296 579310 145308
rect 585134 145296 585140 145308
rect 579304 145268 585140 145296
rect 579304 145256 579310 145268
rect 585134 145256 585140 145268
rect 585192 145256 585198 145308
rect 585962 144916 585968 144968
rect 586020 144956 586026 144968
rect 589458 144956 589464 144968
rect 586020 144928 589464 144956
rect 586020 144916 586026 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579522 144644 579528 144696
rect 579580 144684 579586 144696
rect 584398 144684 584404 144696
rect 579580 144656 584404 144684
rect 579580 144644 579586 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 584582 143556 584588 143608
rect 584640 143596 584646 143608
rect 589458 143596 589464 143608
rect 584640 143568 589464 143596
rect 584640 143556 584646 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 583018 140768 583024 140820
rect 583076 140808 583082 140820
rect 589458 140808 589464 140820
rect 583076 140780 589464 140808
rect 583076 140768 583082 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580442 140740 580448 140752
rect 578660 140712 580448 140740
rect 578660 140700 578666 140712
rect 580442 140700 580448 140712
rect 580500 140700 580506 140752
rect 580258 139408 580264 139460
rect 580316 139448 580322 139460
rect 589458 139448 589464 139460
rect 580316 139420 589464 139448
rect 580316 139408 580322 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579062 136824 579068 136876
rect 579120 136864 579126 136876
rect 585962 136864 585968 136876
rect 579120 136836 585968 136864
rect 579120 136824 579126 136836
rect 585962 136824 585968 136836
rect 586020 136824 586026 136876
rect 585778 136620 585784 136672
rect 585836 136660 585842 136672
rect 589458 136660 589464 136672
rect 585836 136632 589464 136660
rect 585836 136620 585842 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 584398 135260 584404 135312
rect 584456 135300 584462 135312
rect 589458 135300 589464 135312
rect 584456 135272 589464 135300
rect 584456 135260 584462 135272
rect 589458 135260 589464 135272
rect 589516 135260 589522 135312
rect 579522 135124 579528 135176
rect 579580 135164 579586 135176
rect 588538 135164 588544 135176
rect 579580 135136 588544 135164
rect 579580 135124 579586 135136
rect 588538 135124 588544 135136
rect 588596 135124 588602 135176
rect 580626 131724 580632 131776
rect 580684 131764 580690 131776
rect 590286 131764 590292 131776
rect 580684 131736 590292 131764
rect 580684 131724 580690 131736
rect 590286 131724 590292 131736
rect 590344 131724 590350 131776
rect 578878 131248 578884 131300
rect 578936 131288 578942 131300
rect 589458 131288 589464 131300
rect 578936 131260 589464 131288
rect 578936 131248 578942 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 579062 131112 579068 131164
rect 579120 131152 579126 131164
rect 584582 131152 584588 131164
rect 579120 131124 584588 131152
rect 579120 131112 579126 131124
rect 584582 131112 584588 131124
rect 584640 131112 584646 131164
rect 579154 128256 579160 128308
rect 579212 128296 579218 128308
rect 587158 128296 587164 128308
rect 579212 128268 587164 128296
rect 579212 128256 579218 128268
rect 587158 128256 587164 128268
rect 587216 128256 587222 128308
rect 587618 127168 587624 127220
rect 587676 127208 587682 127220
rect 589458 127208 589464 127220
rect 587676 127180 589464 127208
rect 587676 127168 587682 127180
rect 589458 127168 589464 127180
rect 589516 127168 589522 127220
rect 579062 126216 579068 126268
rect 579120 126256 579126 126268
rect 587618 126256 587624 126268
rect 579120 126228 587624 126256
rect 579120 126216 579126 126228
rect 587618 126216 587624 126228
rect 587676 126216 587682 126268
rect 579522 125332 579528 125384
rect 579580 125372 579586 125384
rect 583018 125372 583024 125384
rect 579580 125344 583024 125372
rect 579580 125332 579586 125344
rect 583018 125332 583024 125344
rect 583076 125332 583082 125384
rect 583202 124856 583208 124908
rect 583260 124896 583266 124908
rect 589642 124896 589648 124908
rect 583260 124868 589648 124896
rect 583260 124856 583266 124868
rect 589642 124856 589648 124868
rect 589700 124856 589706 124908
rect 578326 124108 578332 124160
rect 578384 124148 578390 124160
rect 580258 124148 580264 124160
rect 578384 124120 580264 124148
rect 578384 124108 578390 124120
rect 580258 124108 580264 124120
rect 580316 124108 580322 124160
rect 580442 122816 580448 122868
rect 580500 122856 580506 122868
rect 589458 122856 589464 122868
rect 580500 122828 589464 122856
rect 580500 122816 580506 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 581822 122068 581828 122120
rect 581880 122108 581886 122120
rect 590102 122108 590108 122120
rect 581880 122080 590108 122108
rect 581880 122068 581886 122080
rect 590102 122068 590108 122080
rect 590160 122068 590166 122120
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 579522 121388 579528 121440
rect 579580 121428 579586 121440
rect 585778 121428 585784 121440
rect 579580 121400 585784 121428
rect 579580 121388 579586 121400
rect 585778 121388 585784 121400
rect 585836 121388 585842 121440
rect 667934 120096 667940 120148
rect 667992 120136 667998 120148
rect 670142 120136 670148 120148
rect 667992 120108 670148 120136
rect 667992 120096 667998 120108
rect 670142 120096 670148 120108
rect 670200 120096 670206 120148
rect 584582 118668 584588 118720
rect 584640 118708 584646 118720
rect 589458 118708 589464 118720
rect 584640 118680 589464 118708
rect 584640 118668 584646 118680
rect 589458 118668 589464 118680
rect 589516 118668 589522 118720
rect 578694 118532 578700 118584
rect 578752 118572 578758 118584
rect 584398 118572 584404 118584
rect 578752 118544 584404 118572
rect 578752 118532 578758 118544
rect 584398 118532 584404 118544
rect 584456 118532 584462 118584
rect 668026 118532 668032 118584
rect 668084 118572 668090 118584
rect 670326 118572 670332 118584
rect 668084 118544 670332 118572
rect 668084 118532 668090 118544
rect 670326 118532 670332 118544
rect 670384 118532 670390 118584
rect 585962 117308 585968 117360
rect 586020 117348 586026 117360
rect 589458 117348 589464 117360
rect 586020 117320 589464 117348
rect 586020 117308 586026 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 678238 117280 678244 117292
rect 675904 117252 678244 117280
rect 675904 117240 675910 117252
rect 678238 117240 678244 117252
rect 678296 117240 678302 117292
rect 578694 117172 578700 117224
rect 578752 117212 578758 117224
rect 580626 117212 580632 117224
rect 578752 117184 580632 117212
rect 578752 117172 578758 117184
rect 580626 117172 580632 117184
rect 580684 117172 580690 117224
rect 585778 115948 585784 116000
rect 585836 115988 585842 116000
rect 589458 115988 589464 116000
rect 585836 115960 589464 115988
rect 585836 115948 585842 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 584398 113160 584404 113212
rect 584456 113200 584462 113212
rect 589458 113200 589464 113212
rect 584456 113172 589464 113200
rect 584456 113160 584462 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579154 113024 579160 113076
rect 579212 113064 579218 113076
rect 588722 113064 588728 113076
rect 579212 113036 588728 113064
rect 579212 113024 579218 113036
rect 588722 113024 588728 113036
rect 588780 113024 588786 113076
rect 588538 111800 588544 111852
rect 588596 111840 588602 111852
rect 590378 111840 590384 111852
rect 588596 111812 590384 111840
rect 588596 111800 588602 111812
rect 590378 111800 590384 111812
rect 590436 111800 590442 111852
rect 581638 111052 581644 111104
rect 581696 111092 581702 111104
rect 589918 111092 589924 111104
rect 581696 111064 589924 111092
rect 581696 111052 581702 111064
rect 589918 111052 589924 111064
rect 589976 111052 589982 111104
rect 583018 109692 583024 109744
rect 583076 109732 583082 109744
rect 589366 109732 589372 109744
rect 583076 109704 589372 109732
rect 583076 109692 583082 109704
rect 589366 109692 589372 109704
rect 589424 109692 589430 109744
rect 578878 108944 578884 108996
rect 578936 108984 578942 108996
rect 581822 108984 581828 108996
rect 578936 108956 581828 108984
rect 578936 108944 578942 108956
rect 581822 108944 581828 108956
rect 581880 108944 581886 108996
rect 581270 107652 581276 107704
rect 581328 107692 581334 107704
rect 589458 107692 589464 107704
rect 581328 107664 589464 107692
rect 581328 107652 581334 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 666554 106088 666560 106140
rect 666612 106128 666618 106140
rect 666830 106128 666836 106140
rect 666612 106100 666836 106128
rect 666612 106088 666618 106100
rect 666830 106088 666836 106100
rect 666888 106128 666894 106140
rect 670694 106128 670700 106140
rect 666888 106100 670700 106128
rect 666888 106088 666894 106100
rect 670694 106088 670700 106100
rect 670752 106088 670758 106140
rect 579338 105136 579344 105188
rect 579396 105176 579402 105188
rect 581270 105176 581276 105188
rect 579396 105148 581276 105176
rect 579396 105136 579402 105148
rect 581270 105136 581276 105148
rect 581328 105136 581334 105188
rect 581822 104864 581828 104916
rect 581880 104904 581886 104916
rect 589458 104904 589464 104916
rect 581880 104876 589464 104904
rect 581880 104864 581886 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 580258 104116 580264 104168
rect 580316 104156 580322 104168
rect 589642 104156 589648 104168
rect 580316 104128 589648 104156
rect 580316 104116 580322 104128
rect 589642 104116 589648 104128
rect 589700 104116 589706 104168
rect 578326 103300 578332 103352
rect 578384 103340 578390 103352
rect 583202 103340 583208 103352
rect 578384 103312 583208 103340
rect 578384 103300 578390 103312
rect 583202 103300 583208 103312
rect 583260 103300 583266 103352
rect 578510 102076 578516 102128
rect 578568 102116 578574 102128
rect 580442 102116 580448 102128
rect 578568 102088 580448 102116
rect 578568 102076 578574 102088
rect 580442 102076 580448 102088
rect 580500 102076 580506 102128
rect 587158 100716 587164 100768
rect 587216 100756 587222 100768
rect 590286 100756 590292 100768
rect 587216 100728 590292 100756
rect 587216 100716 587222 100728
rect 590286 100716 590292 100728
rect 590344 100716 590350 100768
rect 624786 100104 624792 100156
rect 624844 100144 624850 100156
rect 668394 100144 668400 100156
rect 624844 100116 668400 100144
rect 624844 100104 624850 100116
rect 668394 100104 668400 100116
rect 668452 100104 668458 100156
rect 580442 99968 580448 100020
rect 580500 100008 580506 100020
rect 590102 100008 590108 100020
rect 580500 99980 590108 100008
rect 580500 99968 580506 99980
rect 590102 99968 590108 99980
rect 590160 99968 590166 100020
rect 594058 99968 594064 100020
rect 594116 100008 594122 100020
rect 667934 100008 667940 100020
rect 594116 99980 667940 100008
rect 594116 99968 594122 99980
rect 667934 99968 667940 99980
rect 667992 99968 667998 100020
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 579154 99220 579160 99272
rect 579212 99260 579218 99272
rect 581638 99260 581644 99272
rect 579212 99232 581644 99260
rect 579212 99220 579218 99232
rect 581638 99220 581644 99232
rect 581696 99220 581702 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 627546 98880 627552 98932
rect 627604 98920 627610 98932
rect 640702 98920 640708 98932
rect 627604 98892 640708 98920
rect 627604 98880 627610 98892
rect 640702 98880 640708 98892
rect 640760 98880 640766 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98744 647148 98796
rect 647200 98784 647206 98796
rect 661954 98784 661960 98796
rect 647200 98756 661960 98784
rect 647200 98744 647206 98756
rect 661954 98744 661960 98756
rect 662012 98744 662018 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 631410 98200 631416 98252
rect 631468 98240 631474 98252
rect 631468 98212 634814 98240
rect 631468 98200 631474 98212
rect 634786 98172 634814 98212
rect 642174 98172 642180 98184
rect 634786 98144 642180 98172
rect 642174 98132 642180 98144
rect 642232 98132 642238 98184
rect 631980 98076 632192 98104
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 632164 98036 632192 98076
rect 645118 98036 645124 98048
rect 632164 98008 645124 98036
rect 645118 97996 645124 98008
rect 645176 97996 645182 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 653950 97928 653956 97980
rect 654008 97968 654014 97980
rect 655054 97968 655060 97980
rect 654008 97940 655060 97968
rect 654008 97928 654014 97940
rect 655054 97928 655060 97940
rect 655112 97928 655118 97980
rect 628282 97792 628288 97844
rect 628340 97832 628346 97844
rect 631410 97832 631416 97844
rect 628340 97804 631416 97832
rect 628340 97792 628346 97804
rect 631410 97792 631416 97804
rect 631468 97792 631474 97844
rect 631594 97792 631600 97844
rect 631652 97832 631658 97844
rect 637758 97832 637764 97844
rect 631652 97804 637764 97832
rect 631652 97792 631658 97804
rect 637758 97792 637764 97804
rect 637816 97792 637822 97844
rect 644290 97792 644296 97844
rect 644348 97832 644354 97844
rect 658826 97832 658832 97844
rect 644348 97804 658832 97832
rect 644348 97792 644354 97804
rect 658826 97792 658832 97804
rect 658884 97792 658890 97844
rect 591298 97656 591304 97708
rect 591356 97696 591362 97708
rect 598198 97696 598204 97708
rect 591356 97668 598204 97696
rect 591356 97656 591362 97668
rect 598198 97656 598204 97668
rect 598256 97656 598262 97708
rect 620186 97656 620192 97708
rect 620244 97696 620250 97708
rect 625982 97696 625988 97708
rect 620244 97668 625988 97696
rect 620244 97656 620250 97668
rect 625982 97656 625988 97668
rect 626040 97656 626046 97708
rect 626810 97656 626816 97708
rect 626868 97696 626874 97708
rect 639230 97696 639236 97708
rect 626868 97668 639236 97696
rect 626868 97656 626874 97668
rect 639230 97656 639236 97668
rect 639288 97656 639294 97708
rect 643002 97656 643008 97708
rect 643060 97696 643066 97708
rect 657998 97696 658004 97708
rect 643060 97668 658004 97696
rect 643060 97656 643066 97668
rect 657998 97656 658004 97668
rect 658056 97656 658062 97708
rect 658182 97656 658188 97708
rect 658240 97696 658246 97708
rect 663058 97696 663064 97708
rect 658240 97668 663064 97696
rect 658240 97656 658246 97668
rect 663058 97656 663064 97668
rect 663116 97656 663122 97708
rect 626166 97520 626172 97572
rect 626224 97560 626230 97572
rect 631594 97560 631600 97572
rect 626224 97532 631600 97560
rect 626224 97520 626230 97532
rect 631594 97520 631600 97532
rect 631652 97520 631658 97572
rect 631962 97520 631968 97572
rect 632020 97560 632026 97572
rect 648614 97560 648620 97572
rect 632020 97532 648620 97560
rect 632020 97520 632026 97532
rect 648614 97520 648620 97532
rect 648672 97520 648678 97572
rect 650362 97520 650368 97572
rect 650420 97560 650426 97572
rect 658274 97560 658280 97572
rect 650420 97532 658280 97560
rect 650420 97520 650426 97532
rect 658274 97520 658280 97532
rect 658332 97520 658338 97572
rect 659194 97520 659200 97572
rect 659252 97560 659258 97572
rect 663886 97560 663892 97572
rect 659252 97532 663892 97560
rect 659252 97520 659258 97532
rect 663886 97520 663892 97532
rect 663944 97520 663950 97572
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 620278 97424 620284 97436
rect 612700 97396 620284 97424
rect 612700 97384 612706 97396
rect 620278 97384 620284 97396
rect 620336 97384 620342 97436
rect 623130 97384 623136 97436
rect 623188 97424 623194 97436
rect 632054 97424 632060 97436
rect 623188 97396 632060 97424
rect 623188 97384 623194 97396
rect 632054 97384 632060 97396
rect 632112 97384 632118 97436
rect 632698 97384 632704 97436
rect 632756 97424 632762 97436
rect 650270 97424 650276 97436
rect 632756 97396 650276 97424
rect 632756 97384 632762 97396
rect 650270 97384 650276 97396
rect 650328 97384 650334 97436
rect 651834 97384 651840 97436
rect 651892 97424 651898 97436
rect 659562 97424 659568 97436
rect 651892 97396 659568 97424
rect 651892 97384 651898 97396
rect 659562 97384 659568 97396
rect 659620 97384 659626 97436
rect 659930 97384 659936 97436
rect 659988 97424 659994 97436
rect 665358 97424 665364 97436
rect 659988 97396 665364 97424
rect 659988 97384 659994 97396
rect 665358 97384 665364 97396
rect 665416 97384 665422 97436
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 613378 97288 613384 97300
rect 605524 97260 613384 97288
rect 605524 97248 605530 97260
rect 613378 97248 613384 97260
rect 613436 97248 613442 97300
rect 621658 97248 621664 97300
rect 621716 97288 621722 97300
rect 629294 97288 629300 97300
rect 621716 97260 629300 97288
rect 621716 97248 621722 97260
rect 629294 97248 629300 97260
rect 629352 97248 629358 97300
rect 633250 97248 633256 97300
rect 633308 97288 633314 97300
rect 650546 97288 650552 97300
rect 633308 97260 650552 97288
rect 633308 97248 633314 97260
rect 650546 97248 650552 97260
rect 650604 97248 650610 97300
rect 656802 97180 656808 97232
rect 656860 97220 656866 97232
rect 661402 97220 661408 97232
rect 656860 97192 661408 97220
rect 656860 97180 656866 97192
rect 661402 97180 661408 97192
rect 661460 97180 661466 97232
rect 634722 97112 634728 97164
rect 634780 97152 634786 97164
rect 649074 97152 649080 97164
rect 634780 97124 649080 97152
rect 634780 97112 634786 97124
rect 649074 97112 649080 97124
rect 649132 97112 649138 97164
rect 657998 97044 658004 97096
rect 658056 97084 658062 97096
rect 660114 97084 660120 97096
rect 658056 97056 660120 97084
rect 658056 97044 658062 97056
rect 660114 97044 660120 97056
rect 660172 97044 660178 97096
rect 624602 96976 624608 97028
rect 624660 97016 624666 97028
rect 634998 97016 635004 97028
rect 624660 96988 635004 97016
rect 624660 96976 624666 96988
rect 634998 96976 635004 96988
rect 635056 96976 635062 97028
rect 638586 96976 638592 97028
rect 638644 97016 638650 97028
rect 647786 97016 647792 97028
rect 638644 96988 647792 97016
rect 638644 96976 638650 96988
rect 647786 96976 647792 96988
rect 647844 96976 647850 97028
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 610618 96908 610624 96960
rect 610676 96948 610682 96960
rect 611078 96948 611084 96960
rect 610676 96920 611084 96948
rect 610676 96908 610682 96920
rect 611078 96908 611084 96920
rect 611136 96908 611142 96960
rect 614022 96908 614028 96960
rect 614080 96948 614086 96960
rect 614758 96948 614764 96960
rect 614080 96920 614764 96948
rect 614080 96908 614086 96920
rect 614758 96908 614764 96920
rect 614816 96908 614822 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 660666 96908 660672 96960
rect 660724 96948 660730 96960
rect 663242 96948 663248 96960
rect 660724 96920 663248 96948
rect 660724 96908 660730 96920
rect 663242 96908 663248 96920
rect 663300 96908 663306 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 634170 96840 634176 96892
rect 634228 96880 634234 96892
rect 647970 96880 647976 96892
rect 634228 96852 647976 96880
rect 634228 96840 634234 96852
rect 647970 96840 647976 96852
rect 648028 96840 648034 96892
rect 613562 96772 613568 96824
rect 613620 96812 613626 96824
rect 614022 96812 614028 96824
rect 613620 96784 614028 96812
rect 613620 96772 613626 96784
rect 614022 96772 614028 96784
rect 614080 96772 614086 96824
rect 655238 96772 655244 96824
rect 655296 96812 655302 96824
rect 662506 96812 662512 96824
rect 655296 96784 662512 96812
rect 655296 96772 655302 96784
rect 662506 96772 662512 96784
rect 662564 96772 662570 96824
rect 639046 96568 639052 96620
rect 639104 96608 639110 96620
rect 640334 96608 640340 96620
rect 639104 96580 640340 96608
rect 639104 96568 639110 96580
rect 640334 96568 640340 96580
rect 640392 96568 640398 96620
rect 640518 96568 640524 96620
rect 640576 96608 640582 96620
rect 648430 96608 648436 96620
rect 640576 96580 648436 96608
rect 640576 96568 640582 96580
rect 648430 96568 648436 96580
rect 648488 96568 648494 96620
rect 653306 96568 653312 96620
rect 653364 96608 653370 96620
rect 665174 96608 665180 96620
rect 653364 96580 665180 96608
rect 653364 96568 653370 96580
rect 665174 96568 665180 96580
rect 665232 96568 665238 96620
rect 640058 96432 640064 96484
rect 640116 96472 640122 96484
rect 652018 96472 652024 96484
rect 640116 96444 652024 96472
rect 640116 96432 640122 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 652570 96432 652576 96484
rect 652628 96472 652634 96484
rect 664162 96472 664168 96484
rect 652628 96444 664168 96472
rect 652628 96432 652634 96444
rect 664162 96432 664168 96444
rect 664220 96432 664226 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 647142 96336 647148 96348
rect 631284 96308 647148 96336
rect 631284 96296 631290 96308
rect 647142 96296 647148 96308
rect 647200 96296 647206 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664346 96336 664352 96348
rect 648948 96308 664352 96336
rect 648948 96296 648954 96308
rect 664346 96296 664352 96308
rect 664404 96296 664410 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 663702 96064 663708 96076
rect 641588 96036 663708 96064
rect 641588 96024 641594 96036
rect 663702 96024 663708 96036
rect 663760 96024 663766 96076
rect 577498 95888 577504 95940
rect 577556 95928 577562 95940
rect 600406 95928 600412 95940
rect 577556 95900 600412 95928
rect 577556 95888 577562 95900
rect 600406 95888 600412 95900
rect 600464 95888 600470 95940
rect 609146 95888 609152 95940
rect 609204 95928 609210 95940
rect 621658 95928 621664 95940
rect 609204 95900 621664 95928
rect 609204 95888 609210 95900
rect 621658 95888 621664 95900
rect 621716 95888 621722 95940
rect 644842 95888 644848 95940
rect 644900 95928 644906 95940
rect 648062 95928 648068 95940
rect 644900 95900 648068 95928
rect 644900 95888 644906 95900
rect 648062 95888 648068 95900
rect 648120 95888 648126 95940
rect 648430 95888 648436 95940
rect 648488 95928 648494 95940
rect 664530 95928 664536 95940
rect 648488 95900 664536 95928
rect 648488 95888 648494 95900
rect 664530 95888 664536 95900
rect 664588 95888 664594 95940
rect 645762 95752 645768 95804
rect 645820 95792 645826 95804
rect 652202 95792 652208 95804
rect 645820 95764 652208 95792
rect 645820 95752 645826 95764
rect 652202 95752 652208 95764
rect 652260 95752 652266 95804
rect 656158 95792 656164 95804
rect 654106 95764 656164 95792
rect 646406 95616 646412 95668
rect 646464 95656 646470 95668
rect 653398 95656 653404 95668
rect 646464 95628 653404 95656
rect 646464 95616 646470 95628
rect 653398 95616 653404 95628
rect 653456 95616 653462 95668
rect 640334 95412 640340 95464
rect 640392 95412 640398 95464
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 643520 95424 647924 95452
rect 643520 95412 643526 95424
rect 640352 95316 640380 95412
rect 640352 95288 647464 95316
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 579522 95004 579528 95056
rect 579580 95044 579586 95056
rect 584582 95044 584588 95056
rect 579580 95016 584588 95044
rect 579580 95004 579586 95016
rect 584582 95004 584588 95016
rect 584640 95004 584646 95056
rect 647436 95044 647464 95288
rect 647896 95192 647924 95424
rect 648154 95344 648160 95396
rect 648212 95384 648218 95396
rect 654106 95384 654134 95764
rect 656158 95752 656164 95764
rect 656216 95752 656222 95804
rect 648212 95356 654134 95384
rect 648212 95344 648218 95356
rect 647878 95140 647884 95192
rect 647936 95140 647942 95192
rect 648062 95140 648068 95192
rect 648120 95180 648126 95192
rect 649994 95180 650000 95192
rect 648120 95152 650000 95180
rect 648120 95140 648126 95152
rect 649994 95140 650000 95152
rect 650052 95140 650058 95192
rect 648798 95044 648804 95056
rect 647436 95016 648804 95044
rect 648798 95004 648804 95016
rect 648856 95004 648862 95056
rect 607674 94596 607680 94648
rect 607732 94636 607738 94648
rect 620922 94636 620928 94648
rect 607732 94608 620928 94636
rect 607732 94596 607738 94608
rect 620922 94596 620928 94608
rect 620980 94596 620986 94648
rect 606938 94460 606944 94512
rect 606996 94500 607002 94512
rect 623038 94500 623044 94512
rect 606996 94472 623044 94500
rect 606996 94460 607002 94472
rect 623038 94460 623044 94472
rect 623096 94460 623102 94512
rect 648430 93848 648436 93900
rect 648488 93888 648494 93900
rect 654778 93888 654784 93900
rect 648488 93860 654784 93888
rect 648488 93848 648494 93860
rect 654778 93848 654784 93860
rect 654836 93848 654842 93900
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 651282 93508 651288 93560
rect 651340 93548 651346 93560
rect 655422 93548 655428 93560
rect 651340 93520 655428 93548
rect 651340 93508 651346 93520
rect 655422 93508 655428 93520
rect 655480 93508 655486 93560
rect 579154 93372 579160 93424
rect 579212 93412 579218 93424
rect 585962 93412 585968 93424
rect 579212 93384 585968 93412
rect 579212 93372 579218 93384
rect 585962 93372 585968 93384
rect 586020 93372 586026 93424
rect 611078 93100 611084 93152
rect 611136 93140 611142 93152
rect 618530 93140 618536 93152
rect 611136 93112 618536 93140
rect 611136 93100 611142 93112
rect 618530 93100 618536 93112
rect 618588 93100 618594 93152
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 616598 91740 616604 91792
rect 616656 91780 616662 91792
rect 626258 91780 626264 91792
rect 616656 91752 626264 91780
rect 616656 91740 616662 91752
rect 626258 91740 626264 91752
rect 626316 91740 626322 91792
rect 578510 91672 578516 91724
rect 578568 91712 578574 91724
rect 585778 91712 585784 91724
rect 578568 91684 585784 91712
rect 578568 91672 578574 91684
rect 585778 91672 585784 91684
rect 585836 91672 585842 91724
rect 647694 91672 647700 91724
rect 647752 91712 647758 91724
rect 654686 91712 654692 91724
rect 647752 91684 654692 91712
rect 647752 91672 647758 91684
rect 654686 91672 654692 91684
rect 654744 91672 654750 91724
rect 618162 91128 618168 91180
rect 618220 91168 618226 91180
rect 618220 91140 618392 91168
rect 618220 91128 618226 91140
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 618162 91032 618168 91044
rect 611320 91004 618168 91032
rect 611320 90992 611326 91004
rect 618162 90992 618168 91004
rect 618220 90992 618226 91044
rect 618364 91032 618392 91140
rect 626442 91032 626448 91044
rect 618364 91004 626448 91032
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 648798 90652 648804 90704
rect 648856 90692 648862 90704
rect 655422 90692 655428 90704
rect 648856 90664 655428 90692
rect 648856 90652 648862 90664
rect 655422 90652 655428 90664
rect 655480 90652 655486 90704
rect 620922 89632 620928 89684
rect 620980 89672 620986 89684
rect 626442 89672 626448 89684
rect 620980 89644 626448 89672
rect 620980 89632 620986 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 581638 88952 581644 89004
rect 581696 88992 581702 89004
rect 601694 88992 601700 89004
rect 581696 88964 601700 88992
rect 581696 88952 581702 88964
rect 601694 88952 601700 88964
rect 601752 88952 601758 89004
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 578510 88272 578516 88324
rect 578568 88312 578574 88324
rect 588538 88312 588544 88324
rect 578568 88284 588544 88312
rect 578568 88272 578574 88284
rect 588538 88272 588544 88284
rect 588596 88272 588602 88324
rect 618162 88272 618168 88324
rect 618220 88312 618226 88324
rect 625614 88312 625620 88324
rect 618220 88284 625620 88312
rect 618220 88272 618226 88284
rect 625614 88272 625620 88284
rect 625672 88272 625678 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 623038 88136 623044 88188
rect 623096 88176 623102 88188
rect 626442 88176 626448 88188
rect 623096 88148 626448 88176
rect 623096 88136 623102 88148
rect 626442 88136 626448 88148
rect 626500 88136 626506 88188
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 659562 86912 659568 86964
rect 659620 86952 659626 86964
rect 663242 86952 663248 86964
rect 659620 86924 663248 86952
rect 659620 86912 659626 86924
rect 663242 86912 663248 86924
rect 663300 86912 663306 86964
rect 652202 86844 652208 86896
rect 652260 86884 652266 86896
rect 657722 86884 657728 86896
rect 652260 86856 657728 86884
rect 652260 86844 652266 86856
rect 657722 86844 657728 86856
rect 657780 86844 657786 86896
rect 647878 86708 647884 86760
rect 647936 86748 647942 86760
rect 661402 86748 661408 86760
rect 647936 86720 661408 86748
rect 647936 86708 647942 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 652018 86572 652024 86624
rect 652076 86612 652082 86624
rect 660114 86612 660120 86624
rect 652076 86584 660120 86612
rect 652076 86572 652082 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 656158 86436 656164 86488
rect 656216 86476 656222 86488
rect 660666 86476 660672 86488
rect 656216 86448 660672 86476
rect 656216 86436 656222 86448
rect 660666 86436 660672 86448
rect 660724 86436 660730 86488
rect 618530 86300 618536 86352
rect 618588 86340 618594 86352
rect 626442 86340 626448 86352
rect 618588 86312 626448 86340
rect 618588 86300 618594 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 654870 86300 654876 86352
rect 654928 86340 654934 86352
rect 662506 86340 662512 86352
rect 654928 86312 662512 86340
rect 654928 86300 654934 86312
rect 662506 86300 662512 86312
rect 662564 86300 662570 86352
rect 653398 86164 653404 86216
rect 653456 86204 653462 86216
rect 657170 86204 657176 86216
rect 653456 86176 657176 86204
rect 653456 86164 653462 86176
rect 657170 86164 657176 86176
rect 657228 86164 657234 86216
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 579062 85416 579068 85468
rect 579120 85456 579126 85468
rect 581822 85456 581828 85468
rect 579120 85428 581828 85456
rect 579120 85416 579126 85428
rect 581822 85416 581828 85428
rect 581880 85416 581886 85468
rect 621658 85348 621664 85400
rect 621716 85388 621722 85400
rect 625246 85388 625252 85400
rect 621716 85360 625252 85388
rect 621716 85348 621722 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 626442 84164 626448 84176
rect 608560 84136 626448 84164
rect 608560 84124 608566 84136
rect 626442 84124 626448 84136
rect 626500 84124 626506 84176
rect 579522 83988 579528 84040
rect 579580 84028 579586 84040
rect 583018 84028 583024 84040
rect 579580 84000 583024 84028
rect 579580 83988 579586 84000
rect 583018 83988 583024 84000
rect 583076 83988 583082 84040
rect 578510 82560 578516 82612
rect 578568 82600 578574 82612
rect 584398 82600 584404 82612
rect 578568 82572 584404 82600
rect 578568 82560 578574 82572
rect 584398 82560 584404 82572
rect 584456 82560 584462 82612
rect 628742 80928 628748 80980
rect 628800 80968 628806 80980
rect 642450 80968 642456 80980
rect 628800 80940 642456 80968
rect 628800 80928 628806 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 615402 80792 615408 80844
rect 615460 80832 615466 80844
rect 646130 80832 646136 80844
rect 615460 80804 646136 80832
rect 615460 80792 615466 80804
rect 646130 80792 646136 80804
rect 646188 80792 646194 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 612642 79432 612648 79484
rect 612700 79472 612706 79484
rect 645946 79472 645952 79484
rect 612700 79444 645952 79472
rect 612700 79432 612706 79444
rect 645946 79432 645952 79444
rect 646004 79432 646010 79484
rect 584398 79296 584404 79348
rect 584456 79336 584462 79348
rect 589918 79336 589924 79348
rect 584456 79308 589924 79336
rect 584456 79296 584462 79308
rect 589918 79296 589924 79308
rect 589976 79296 589982 79348
rect 614758 79296 614764 79348
rect 614816 79336 614822 79348
rect 648706 79336 648712 79348
rect 614816 79308 648712 79336
rect 614816 79296 614822 79308
rect 648706 79296 648712 79308
rect 648764 79296 648770 79348
rect 578510 78412 578516 78464
rect 578568 78452 578574 78464
rect 580258 78452 580264 78464
rect 578568 78424 580264 78452
rect 578568 78412 578574 78424
rect 580258 78412 580264 78424
rect 580316 78412 580322 78464
rect 633434 78208 633440 78260
rect 633492 78248 633498 78260
rect 645302 78248 645308 78260
rect 633492 78220 645308 78248
rect 633492 78208 633498 78220
rect 645302 78208 645308 78220
rect 645360 78208 645366 78260
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 643094 78112 643100 78124
rect 631100 78084 643100 78112
rect 631100 78072 631106 78084
rect 643094 78072 643100 78084
rect 643152 78072 643158 78124
rect 614022 77936 614028 77988
rect 614080 77976 614086 77988
rect 647234 77976 647240 77988
rect 614080 77948 647240 77976
rect 614080 77936 614086 77948
rect 647234 77936 647240 77948
rect 647292 77936 647298 77988
rect 628466 77392 628472 77444
rect 628524 77432 628530 77444
rect 632790 77432 632796 77444
rect 628524 77404 632796 77432
rect 628524 77392 628530 77404
rect 632790 77392 632796 77404
rect 632848 77392 632854 77444
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 616782 76644 616788 76696
rect 616840 76684 616846 76696
rect 646498 76684 646504 76696
rect 616840 76656 646504 76684
rect 616840 76644 616846 76656
rect 646498 76644 646504 76656
rect 646556 76644 646562 76696
rect 579338 76508 579344 76560
rect 579396 76548 579402 76560
rect 666554 76548 666560 76560
rect 579396 76520 666560 76548
rect 579396 76508 579402 76520
rect 666554 76508 666560 76520
rect 666612 76508 666618 76560
rect 621658 75896 621664 75948
rect 621716 75936 621722 75948
rect 628466 75936 628472 75948
rect 621716 75908 628472 75936
rect 621716 75896 621722 75908
rect 628466 75896 628472 75908
rect 628524 75896 628530 75948
rect 620278 75420 620284 75472
rect 620336 75460 620342 75472
rect 648890 75460 648896 75472
rect 620336 75432 648896 75460
rect 620336 75420 620342 75432
rect 648890 75420 648896 75432
rect 648948 75420 648954 75472
rect 607122 75284 607128 75336
rect 607180 75324 607186 75336
rect 646314 75324 646320 75336
rect 607180 75296 646320 75324
rect 607180 75284 607186 75296
rect 646314 75284 646320 75296
rect 646372 75284 646378 75336
rect 613378 75148 613384 75200
rect 613436 75188 613442 75200
rect 662598 75188 662604 75200
rect 613436 75160 662604 75188
rect 613436 75148 613442 75160
rect 662598 75148 662604 75160
rect 662656 75148 662662 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 587158 73148 587164 73160
rect 579580 73120 587164 73148
rect 579580 73108 579586 73120
rect 587158 73108 587164 73120
rect 587216 73108 587222 73160
rect 578510 71544 578516 71596
rect 578568 71584 578574 71596
rect 584398 71584 584404 71596
rect 578568 71556 584404 71584
rect 578568 71544 578574 71556
rect 584398 71544 584404 71556
rect 584456 71544 584462 71596
rect 584398 68280 584404 68332
rect 584456 68320 584462 68332
rect 604454 68320 604460 68332
rect 584456 68292 604460 68320
rect 584456 68280 584462 68292
rect 604454 68280 604460 68292
rect 604512 68280 604518 68332
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 623038 66280 623044 66292
rect 579580 66252 623044 66280
rect 579580 66240 579586 66252
rect 623038 66240 623044 66252
rect 623096 66240 623102 66292
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 594058 64852 594064 64864
rect 579580 64824 594064 64852
rect 579580 64812 579586 64824
rect 594058 64812 594064 64824
rect 594116 64812 594122 64864
rect 579522 62024 579528 62076
rect 579580 62064 579586 62076
rect 611998 62064 612004 62076
rect 579580 62036 612004 62064
rect 579580 62024 579586 62036
rect 611998 62024 612004 62036
rect 612056 62024 612062 62076
rect 579522 60664 579528 60716
rect 579580 60704 579586 60716
rect 624418 60704 624424 60716
rect 579580 60676 624424 60704
rect 579580 60664 579586 60676
rect 624418 60664 624424 60676
rect 624476 60664 624482 60716
rect 579062 58760 579068 58812
rect 579120 58800 579126 58812
rect 597554 58800 597560 58812
rect 579120 58772 597560 58800
rect 579120 58760 579126 58772
rect 597554 58760 597560 58772
rect 597612 58760 597618 58812
rect 577682 58624 577688 58676
rect 577740 58664 577746 58676
rect 603074 58664 603080 58676
rect 577740 58636 603080 58664
rect 577740 58624 577746 58636
rect 603074 58624 603080 58636
rect 603132 58624 603138 58676
rect 574922 57332 574928 57384
rect 574980 57372 574986 57384
rect 600498 57372 600504 57384
rect 574980 57344 600504 57372
rect 574980 57332 574986 57344
rect 600498 57332 600504 57344
rect 600556 57332 600562 57384
rect 575474 57196 575480 57248
rect 575532 57236 575538 57248
rect 601878 57236 601884 57248
rect 575532 57208 601884 57236
rect 575532 57196 575538 57208
rect 601878 57196 601884 57208
rect 601936 57196 601942 57248
rect 578510 56516 578516 56568
rect 578568 56556 578574 56568
rect 621658 56556 621664 56568
rect 578568 56528 621664 56556
rect 578568 56516 578574 56528
rect 621658 56516 621664 56528
rect 621716 56516 621722 56568
rect 574738 55972 574744 56024
rect 574796 56012 574802 56024
rect 598934 56012 598940 56024
rect 574796 55984 598940 56012
rect 574796 55972 574802 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574554 55836 574560 55888
rect 574612 55876 574618 55888
rect 599118 55876 599124 55888
rect 574612 55848 599124 55876
rect 574612 55836 574618 55848
rect 599118 55836 599124 55848
rect 599176 55836 599182 55888
rect 577498 55196 577504 55208
rect 462838 55168 577504 55196
rect 462838 54856 462866 55168
rect 577498 55156 577504 55168
rect 577556 55156 577562 55208
rect 591298 55060 591304 55072
rect 462332 54828 462866 54856
rect 462976 55032 591304 55060
rect 462130 53592 462136 53644
rect 462188 53632 462194 53644
rect 462332 53632 462360 54828
rect 462976 54516 463004 55032
rect 591298 55020 591304 55032
rect 591356 55020 591362 55072
rect 596450 54924 596456 54936
rect 462884 54488 463004 54516
rect 464080 54896 596456 54924
rect 462884 54380 462912 54488
rect 462884 54352 463004 54380
rect 462188 53604 462360 53632
rect 462976 53632 463004 54352
rect 464080 53644 464108 54896
rect 596450 54884 596456 54896
rect 596508 54884 596514 54936
rect 596266 54788 596272 54800
rect 465000 54760 596272 54788
rect 465000 53644 465028 54760
rect 596266 54748 596272 54760
rect 596324 54748 596330 54800
rect 625982 54652 625988 54664
rect 467760 54624 625988 54652
rect 463326 53632 463332 53644
rect 462976 53604 463332 53632
rect 462188 53592 462194 53604
rect 463326 53592 463332 53604
rect 463384 53592 463390 53644
rect 464062 53592 464068 53644
rect 464120 53592 464126 53644
rect 464982 53592 464988 53644
rect 465040 53592 465046 53644
rect 465902 53592 465908 53644
rect 465960 53632 465966 53644
rect 467760 53632 467788 54624
rect 625982 54612 625988 54624
rect 626040 54612 626046 54664
rect 625798 54516 625804 54528
rect 467944 54488 625804 54516
rect 467944 53644 467972 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 580442 54380 580448 54392
rect 468588 54352 580448 54380
rect 468588 53644 468616 54352
rect 580442 54340 580448 54352
rect 580500 54340 580506 54392
rect 579062 54244 579068 54256
rect 468772 54216 579068 54244
rect 468772 53644 468800 54216
rect 579062 54204 579068 54216
rect 579120 54204 579126 54256
rect 574554 54108 574560 54120
rect 473326 54080 574560 54108
rect 473326 53972 473354 54080
rect 574554 54068 574560 54080
rect 574612 54068 574618 54120
rect 574922 53972 574928 53984
rect 468956 53944 473354 53972
rect 480226 53944 574928 53972
rect 465960 53604 467788 53632
rect 465960 53592 465966 53604
rect 467926 53592 467932 53644
rect 467984 53592 467990 53644
rect 468570 53592 468576 53644
rect 468628 53592 468634 53644
rect 468754 53592 468760 53644
rect 468812 53592 468818 53644
rect 461302 53456 461308 53508
rect 461360 53496 461366 53508
rect 468956 53496 468984 53944
rect 480226 53904 480254 53944
rect 574922 53932 574928 53944
rect 574980 53932 574986 53984
rect 476086 53876 480254 53904
rect 476086 53836 476114 53876
rect 461360 53468 468984 53496
rect 469140 53808 476114 53836
rect 461360 53456 461366 53468
rect 49142 53320 49148 53372
rect 49200 53360 49206 53372
rect 129182 53360 129188 53372
rect 49200 53332 129188 53360
rect 49200 53320 49206 53332
rect 129182 53320 129188 53332
rect 129240 53320 129246 53372
rect 463142 53320 463148 53372
rect 463200 53360 463206 53372
rect 469140 53360 469168 53808
rect 463200 53332 469168 53360
rect 463200 53320 463206 53332
rect 50338 53184 50344 53236
rect 50396 53224 50402 53236
rect 130378 53224 130384 53236
rect 50396 53196 130384 53224
rect 50396 53184 50402 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 465442 53116 465448 53168
rect 465500 53156 465506 53168
rect 468570 53156 468576 53168
rect 465500 53128 468576 53156
rect 465500 53116 465506 53128
rect 468570 53116 468576 53128
rect 468628 53116 468634 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 128998 53088 129004 53100
rect 46256 53060 129004 53088
rect 46256 53048 46262 53060
rect 128998 53048 129004 53060
rect 129056 53048 129062 53100
rect 467926 52952 467932 52964
rect 462286 52924 467932 52952
rect 460060 52776 460066 52828
rect 460118 52816 460124 52828
rect 462286 52816 462314 52924
rect 467926 52912 467932 52924
rect 467984 52912 467990 52964
rect 460118 52788 462314 52816
rect 460118 52776 460124 52788
rect 464200 52776 464206 52828
rect 464258 52816 464264 52828
rect 468754 52816 468760 52828
rect 464258 52788 468760 52816
rect 464258 52776 464264 52788
rect 468754 52776 468760 52788
rect 468812 52776 468818 52828
rect 48958 51960 48964 52012
rect 49016 52000 49022 52012
rect 129550 52000 129556 52012
rect 49016 51972 129556 52000
rect 49016 51960 49022 51972
rect 129550 51960 129556 51972
rect 129608 51960 129614 52012
rect 47578 51824 47584 51876
rect 47636 51864 47642 51876
rect 129366 51864 129372 51876
rect 47636 51836 129372 51864
rect 47636 51824 47642 51836
rect 129366 51824 129372 51836
rect 129424 51824 129430 51876
rect 46382 51688 46388 51740
rect 46440 51728 46446 51740
rect 130562 51728 130568 51740
rect 46440 51700 130568 51728
rect 46440 51688 46446 51700
rect 130562 51688 130568 51700
rect 130620 51688 130626 51740
rect 145374 51688 145380 51740
rect 145432 51728 145438 51740
rect 306006 51728 306012 51740
rect 145432 51700 306012 51728
rect 145432 51688 145438 51700
rect 306006 51688 306012 51700
rect 306064 51688 306070 51740
rect 50522 50464 50528 50516
rect 50580 50504 50586 50516
rect 128722 50504 128728 50516
rect 50580 50476 128728 50504
rect 50580 50464 50586 50476
rect 128722 50464 128728 50476
rect 128780 50464 128786 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 128538 50368 128544 50380
rect 45520 50340 128544 50368
rect 45520 50328 45526 50340
rect 128538 50328 128544 50340
rect 128596 50328 128602 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 128906 49144 128912 49156
rect 51776 49116 128912 49144
rect 51776 49104 51782 49116
rect 128906 49104 128912 49116
rect 128964 49104 128970 49156
rect 47762 48968 47768 49020
rect 47820 49008 47826 49020
rect 131022 49008 131028 49020
rect 47820 48980 131028 49008
rect 47820 48968 47826 48980
rect 131022 48968 131028 48980
rect 131080 48968 131086 49020
rect 128906 47812 128912 47864
rect 128964 47852 128970 47864
rect 131574 47852 131580 47864
rect 128964 47824 131580 47852
rect 128964 47812 128970 47824
rect 131574 47812 131580 47824
rect 131632 47812 131638 47864
rect 128722 47676 128728 47728
rect 128780 47716 128786 47728
rect 132034 47716 132040 47728
rect 128780 47688 132040 47716
rect 128780 47676 128786 47688
rect 132034 47676 132040 47688
rect 132092 47676 132098 47728
rect 623038 46452 623044 46504
rect 623096 46492 623102 46504
rect 661586 46492 661592 46504
rect 623096 46464 661592 46492
rect 623096 46452 623102 46464
rect 661586 46452 661592 46464
rect 661644 46452 661650 46504
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 129608 45036 131160 45064
rect 129608 45024 129614 45036
rect 129366 44752 129372 44804
rect 129424 44792 129430 44804
rect 131408 44792 131436 44978
rect 131592 44804 131620 44894
rect 129424 44764 131436 44792
rect 129424 44752 129430 44764
rect 131574 44752 131580 44804
rect 131632 44752 131638 44804
rect 129182 44616 129188 44668
rect 129240 44656 129246 44668
rect 131776 44656 131804 44810
rect 131960 44724 131988 44726
rect 129240 44628 131804 44656
rect 131868 44696 131988 44724
rect 129240 44616 129246 44628
rect 131868 44572 131896 44696
rect 130396 44544 131896 44572
rect 132052 44628 132158 44656
rect 128998 44480 129004 44532
rect 129056 44520 129062 44532
rect 130396 44520 130424 44544
rect 132052 44532 132080 44628
rect 129056 44492 130424 44520
rect 129056 44480 129062 44492
rect 132034 44480 132040 44532
rect 132092 44480 132098 44532
rect 132420 44464 132448 44558
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 130562 44276 130568 44328
rect 130620 44316 130626 44328
rect 132604 44316 132632 44474
rect 130620 44288 132632 44316
rect 130620 44276 130626 44288
rect 128538 44140 128544 44192
rect 128596 44180 128602 44192
rect 132218 44180 132224 44192
rect 128596 44152 132224 44180
rect 128596 44140 128602 44152
rect 132218 44140 132224 44152
rect 132276 44140 132282 44192
rect 132788 44180 132816 44362
rect 132420 44152 132816 44180
rect 130378 44004 130384 44056
rect 130436 44044 130442 44056
rect 132420 44044 132448 44152
rect 130436 44016 132448 44044
rect 130436 44004 130442 44016
rect 131022 43868 131028 43920
rect 131080 43908 131086 43920
rect 132972 43908 133000 44250
rect 131080 43880 133000 43908
rect 131080 43868 131086 43880
rect 43438 42780 43444 42832
rect 43496 42820 43502 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 439590 43596 439596 43648
rect 439648 43636 439654 43648
rect 441614 43636 441620 43648
rect 439648 43608 441620 43636
rect 439648 43596 439654 43608
rect 441614 43596 441620 43608
rect 441672 43596 441678 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43496 42792 133184 42820
rect 43496 42780 43502 42792
rect 310422 42712 310428 42764
rect 310480 42752 310486 42764
rect 431218 42752 431224 42764
rect 310480 42724 431224 42752
rect 310480 42712 310486 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 463050 42752 463056 42764
rect 456116 42724 463056 42752
rect 456116 42712 456122 42724
rect 463050 42712 463056 42724
rect 463108 42712 463114 42764
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405550 42344 405556 42356
rect 404504 42316 405556 42344
rect 404504 42304 404510 42316
rect 405550 42304 405556 42316
rect 405608 42304 405614 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 427078 42344 427084 42356
rect 420788 42316 427084 42344
rect 420788 42304 420794 42316
rect 427078 42304 427084 42316
rect 427136 42304 427142 42356
rect 662414 42173 662420 42225
rect 662472 42173 662478 42225
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 427078 41420 427084 41472
rect 427136 41460 427142 41472
rect 459186 41460 459192 41472
rect 427136 41432 459192 41460
rect 427136 41420 427142 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 428004 1006816 428056 1006868
rect 428372 1006680 428424 1006732
rect 434444 1006680 434496 1006732
rect 357716 1006612 357768 1006664
rect 371884 1006612 371936 1006664
rect 145564 1006544 145616 1006596
rect 152924 1006544 152976 1006596
rect 300124 1006544 300176 1006596
rect 308128 1006544 308180 1006596
rect 359740 1006476 359792 1006528
rect 370504 1006476 370556 1006528
rect 422668 1006476 422720 1006528
rect 426532 1006476 426584 1006528
rect 94504 1006408 94556 1006460
rect 103980 1006408 104032 1006460
rect 145748 1006408 145800 1006460
rect 152096 1006408 152148 1006460
rect 157432 1006408 157484 1006460
rect 166264 1006408 166316 1006460
rect 94688 1006272 94740 1006324
rect 101128 1006272 101180 1006324
rect 144276 1006272 144328 1006324
rect 93308 1006136 93360 1006188
rect 98276 1006136 98328 1006188
rect 107660 1006136 107712 1006188
rect 124864 1006136 124916 1006188
rect 144092 1006136 144144 1006188
rect 151268 1006136 151320 1006188
rect 158260 1006272 158312 1006324
rect 171784 1006408 171836 1006460
rect 431684 1006408 431736 1006460
rect 425336 1006340 425388 1006392
rect 204904 1006272 204956 1006324
rect 210056 1006272 210108 1006324
rect 249248 1006272 249300 1006324
rect 254124 1006272 254176 1006324
rect 298928 1006272 298980 1006324
rect 311808 1006272 311860 1006324
rect 358544 1006272 358596 1006324
rect 377404 1006272 377456 1006324
rect 431684 1006204 431736 1006256
rect 153752 1006136 153804 1006188
rect 160284 1006136 160336 1006188
rect 164884 1006136 164936 1006188
rect 166264 1006136 166316 1006188
rect 175924 1006136 175976 1006188
rect 210424 1006136 210476 1006188
rect 228364 1006136 228416 1006188
rect 247040 1006136 247092 1006188
rect 255320 1006136 255372 1006188
rect 261852 1006136 261904 1006188
rect 279424 1006136 279476 1006188
rect 299480 1006136 299532 1006188
rect 306104 1006136 306156 1006188
rect 361396 1006136 361448 1006188
rect 367008 1006136 367060 1006188
rect 402244 1006136 402296 1006188
rect 429200 1006136 429252 1006188
rect 504548 1006816 504600 1006868
rect 516968 1006816 517020 1006868
rect 556988 1006816 557040 1006868
rect 559656 1006816 559708 1006868
rect 505376 1006680 505428 1006732
rect 515404 1006680 515456 1006732
rect 554320 1006680 554372 1006732
rect 562324 1006680 562376 1006732
rect 506204 1006408 506256 1006460
rect 464988 1006272 465040 1006324
rect 555976 1006408 556028 1006460
rect 566464 1006408 566516 1006460
rect 520924 1006272 520976 1006324
rect 471244 1006136 471296 1006188
rect 508228 1006136 508280 1006188
rect 93124 1006000 93176 1006052
rect 99472 1006000 99524 1006052
rect 102784 1006000 102836 1006052
rect 104808 1006000 104860 1006052
rect 108488 1006000 108540 1006052
rect 126244 1006000 126296 1006052
rect 148876 1006000 148928 1006052
rect 150072 1006000 150124 1006052
rect 159456 1006000 159508 1006052
rect 177304 1006000 177356 1006052
rect 198372 1006000 198424 1006052
rect 201040 1006000 201092 1006052
rect 208400 1006000 208452 1006052
rect 229744 1006000 229796 1006052
rect 251088 1006000 251140 1006052
rect 252468 1006000 252520 1006052
rect 260196 1006000 260248 1006052
rect 280804 1006000 280856 1006052
rect 298744 1006000 298796 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 314660 1006000 314712 1006052
rect 319444 1006000 319496 1006052
rect 363420 1005932 363472 1005984
rect 382924 1006000 382976 1006052
rect 400864 1006000 400916 1006052
rect 425336 1006000 425388 1006052
rect 425520 1006000 425572 1006052
rect 429200 1006000 429252 1006052
rect 430856 1005932 430908 1005984
rect 469864 1006000 469916 1006052
rect 498108 1006000 498160 1006052
rect 498844 1006000 498896 1006052
rect 509056 1006000 509108 1006052
rect 557172 1006136 557224 1006188
rect 567844 1006136 567896 1006188
rect 522304 1006000 522356 1006052
rect 549168 1006000 549220 1006052
rect 550272 1006000 550324 1006052
rect 553952 1006000 554004 1006052
rect 556160 1006000 556212 1006052
rect 562324 1006000 562376 1006052
rect 573364 1006000 573416 1006052
rect 514024 1005932 514076 1005984
rect 304080 1005796 304132 1005848
rect 426348 1005728 426400 1005780
rect 440884 1005728 440936 1005780
rect 367008 1005660 367060 1005712
rect 380164 1005660 380216 1005712
rect 360568 1005524 360620 1005576
rect 378784 1005524 378836 1005576
rect 426348 1005524 426400 1005576
rect 443644 1005524 443696 1005576
rect 556160 1005524 556212 1005576
rect 570604 1005524 570656 1005576
rect 358544 1005388 358596 1005440
rect 373264 1005388 373316 1005440
rect 430028 1005388 430080 1005440
rect 431960 1005388 432012 1005440
rect 434444 1005388 434496 1005440
rect 458824 1005388 458876 1005440
rect 502156 1005388 502208 1005440
rect 518164 1005388 518216 1005440
rect 551468 1005388 551520 1005440
rect 569224 1005388 569276 1005440
rect 354864 1005252 354916 1005304
rect 374644 1005252 374696 1005304
rect 423496 1005252 423548 1005304
rect 456064 1005252 456116 1005304
rect 499672 1005252 499724 1005304
rect 516784 1005252 516836 1005304
rect 551468 1005116 551520 1005168
rect 574744 1005252 574796 1005304
rect 149888 1005048 149940 1005100
rect 152924 1005048 152976 1005100
rect 158628 1005048 158680 1005100
rect 162124 1005048 162176 1005100
rect 263048 1005048 263100 1005100
rect 268384 1005048 268436 1005100
rect 354404 1005048 354456 1005100
rect 356520 1005048 356572 1005100
rect 361396 1005048 361448 1005100
rect 364892 1005048 364944 1005100
rect 430028 1005048 430080 1005100
rect 432604 1005048 432656 1005100
rect 151084 1004912 151136 1004964
rect 153752 1004912 153804 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 313832 1004912 313884 1004964
rect 316040 1004912 316092 1004964
rect 353208 1004912 353260 1004964
rect 355692 1004912 355744 1004964
rect 422208 1004912 422260 1004964
rect 423496 1004912 423548 1004964
rect 431224 1004912 431276 1004964
rect 433524 1004912 433576 1004964
rect 507032 1004912 507084 1004964
rect 509700 1004912 509752 1004964
rect 556804 1004912 556856 1004964
rect 558920 1004912 558972 1004964
rect 149704 1004776 149756 1004828
rect 151728 1004776 151780 1004828
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 207572 1004776 207624 1004828
rect 209780 1004776 209832 1004828
rect 211252 1004776 211304 1004828
rect 215944 1004776 215996 1004828
rect 314660 1004776 314712 1004828
rect 316684 1004776 316736 1004828
rect 362592 1004776 362644 1004828
rect 365260 1004776 365312 1004828
rect 420828 1004776 420880 1004828
rect 422668 1004776 422720 1004828
rect 507860 1004776 507912 1004828
rect 510068 1004776 510120 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 151268 1004640 151320 1004692
rect 154120 1004640 154172 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 212540 1004640 212592 1004692
rect 217324 1004640 217376 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 499304 1004640 499356 1004692
rect 501328 1004640 501380 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 505376 1004572 505428 1004624
rect 510252 1004572 510304 1004624
rect 429200 1004028 429252 1004080
rect 446404 1004028 446456 1004080
rect 558920 1004028 558972 1004080
rect 571984 1004028 572036 1004080
rect 92664 1003892 92716 1003944
rect 104808 1003892 104860 1003944
rect 356888 1003892 356940 1003944
rect 375380 1003892 375432 1003944
rect 427176 1003892 427228 1003944
rect 464804 1003892 464856 1003944
rect 505008 1003892 505060 1003944
rect 517520 1003892 517572 1003944
rect 552296 1003892 552348 1003944
rect 572628 1003892 572680 1003944
rect 464988 1003280 465040 1003332
rect 472440 1003280 472492 1003332
rect 424324 1002804 424376 1002856
rect 426532 1002668 426584 1002720
rect 106832 1002600 106884 1002652
rect 109500 1002600 109552 1002652
rect 253480 1002600 253532 1002652
rect 256148 1002600 256200 1002652
rect 261024 1002600 261076 1002652
rect 264244 1002600 264296 1002652
rect 303252 1002600 303304 1002652
rect 306932 1002600 306984 1002652
rect 422208 1002532 422260 1002584
rect 427728 1002532 427780 1002584
rect 449164 1002668 449216 1002720
rect 504180 1002668 504232 1002720
rect 518900 1002668 518952 1002720
rect 464988 1002532 465040 1002584
rect 501696 1002532 501748 1002584
rect 523316 1002532 523368 1002584
rect 98644 1002464 98696 1002516
rect 101496 1002464 101548 1002516
rect 108028 1002464 108080 1002516
rect 110696 1002464 110748 1002516
rect 251916 1002464 251968 1002516
rect 255320 1002464 255372 1002516
rect 358728 1002464 358780 1002516
rect 359372 1002464 359424 1002516
rect 558828 1002464 558880 1002516
rect 562508 1002464 562560 1002516
rect 261024 1002396 261076 1002448
rect 263692 1002396 263744 1002448
rect 97264 1002328 97316 1002380
rect 100300 1002328 100352 1002380
rect 100484 1002328 100536 1002380
rect 103152 1002328 103204 1002380
rect 106832 1002328 106884 1002380
rect 109040 1002328 109092 1002380
rect 148508 1002328 148560 1002380
rect 150900 1002328 150952 1002380
rect 210884 1002328 210936 1002380
rect 213184 1002328 213236 1002380
rect 253020 1002328 253072 1002380
rect 256148 1002328 256200 1002380
rect 357348 1002328 357400 1002380
rect 359464 1002328 359516 1002380
rect 500316 1002328 500368 1002380
rect 503352 1002328 503404 1002380
rect 560852 1002328 560904 1002380
rect 565268 1002328 565320 1002380
rect 262680 1002260 262732 1002312
rect 265808 1002260 265860 1002312
rect 365076 1002260 365128 1002312
rect 367928 1002260 367980 1002312
rect 95884 1002192 95936 1002244
rect 99104 1002192 99156 1002244
rect 100024 1002192 100076 1002244
rect 101956 1002192 102008 1002244
rect 106004 1002192 106056 1002244
rect 108304 1002192 108356 1002244
rect 108856 1002192 108908 1002244
rect 111892 1002192 111944 1002244
rect 153844 1002192 153896 1002244
rect 155776 1002192 155828 1002244
rect 156604 1002192 156656 1002244
rect 158720 1002192 158772 1002244
rect 203340 1002192 203392 1002244
rect 206376 1002192 206428 1002244
rect 251456 1002192 251508 1002244
rect 254492 1002192 254544 1002244
rect 357716 1002192 357768 1002244
rect 360844 1002192 360896 1002244
rect 428372 1002192 428424 1002244
rect 431408 1002192 431460 1002244
rect 432052 1002192 432104 1002244
rect 435548 1002192 435600 1002244
rect 500500 1002192 500552 1002244
rect 502984 1002192 503036 1002244
rect 509884 1002192 509936 1002244
rect 512828 1002192 512880 1002244
rect 560024 1002192 560076 1002244
rect 562324 1002192 562376 1002244
rect 263876 1002124 263928 1002176
rect 267004 1002124 267056 1002176
rect 365904 1002124 365956 1002176
rect 369124 1002124 369176 1002176
rect 97448 1002056 97500 1002108
rect 100300 1002056 100352 1002108
rect 101588 1002056 101640 1002108
rect 103152 1002056 103204 1002108
rect 105636 1002056 105688 1002108
rect 107752 1002056 107804 1002108
rect 109684 1002056 109736 1002108
rect 112076 1002056 112128 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 195152 1002056 195204 1002108
rect 203524 1002056 203576 1002108
rect 206744 1002056 206796 1002108
rect 208400 1002056 208452 1002108
rect 210884 1002056 210936 1002108
rect 212540 1002056 212592 1002108
rect 301504 1002056 301556 1002108
rect 304908 1002056 304960 1002108
rect 360568 1002056 360620 1002108
rect 363604 1002056 363656 1002108
rect 419448 1002056 419500 1002108
rect 421472 1002056 421524 1002108
rect 427544 1002056 427596 1002108
rect 429936 1002056 429988 1002108
rect 433340 1002056 433392 1002108
rect 435364 1002056 435416 1002108
rect 503352 1002056 503404 1002108
rect 505744 1002056 505796 1002108
rect 510344 1002056 510396 1002108
rect 512644 1002056 512696 1002108
rect 552296 1002056 552348 1002108
rect 555424 1002056 555476 1002108
rect 558000 1002056 558052 1002108
rect 560668 1002056 560720 1002108
rect 560852 1002056 560904 1002108
rect 565084 1002056 565136 1002108
rect 263508 1001988 263560 1002040
rect 265624 1001988 265676 1002040
rect 365076 1001988 365128 1002040
rect 367744 1001988 367796 1002040
rect 96068 1001920 96120 1001972
rect 98276 1001920 98328 1001972
rect 98828 1001920 98880 1001972
rect 101128 1001920 101180 1001972
rect 101404 1001920 101456 1001972
rect 102324 1001920 102376 1001972
rect 106004 1001920 106056 1001972
rect 108120 1001920 108172 1001972
rect 108856 1001920 108908 1001972
rect 110512 1001920 110564 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 152464 1001920 152516 1001972
rect 154580 1001920 154632 1001972
rect 154948 1001920 155000 1001972
rect 157340 1001920 157392 1001972
rect 157800 1001920 157852 1001972
rect 160100 1001920 160152 1001972
rect 202696 1001920 202748 1001972
rect 204168 1001920 204220 1001972
rect 205548 1001920 205600 1001972
rect 206284 1001920 206336 1001972
rect 207572 1001920 207624 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 355692 1001920 355744 1001972
rect 356704 1001920 356756 1001972
rect 360200 1001920 360252 1001972
rect 362224 1001920 362276 1001972
rect 399944 1001920 399996 1001972
rect 422300 1001920 422352 1001972
rect 423404 1001920 423456 1001972
rect 424324 1001920 424376 1001972
rect 425520 1001920 425572 1001972
rect 428464 1001920 428516 1001972
rect 429200 1001920 429252 1001972
rect 431224 1001920 431276 1001972
rect 432880 1001920 432932 1001972
rect 436744 1001920 436796 1001972
rect 496728 1001920 496780 1001972
rect 498476 1001920 498528 1001972
rect 499580 1001920 499632 1001972
rect 500500 1001920 500552 1001972
rect 500960 1001920 501012 1001972
rect 502156 1001920 502208 1001972
rect 502524 1001920 502576 1001972
rect 504364 1001920 504416 1001972
rect 553308 1001920 553360 1001972
rect 555148 1001920 555200 1001972
rect 558828 1001920 558880 1001972
rect 560300 1001920 560352 1001972
rect 561680 1001920 561732 1001972
rect 563704 1001920 563756 1001972
rect 195888 1001784 195940 1001836
rect 510160 1001716 510212 1001768
rect 516692 1001716 516744 1001768
rect 446404 1001580 446456 1001632
rect 453212 1001580 453264 1001632
rect 428464 1001444 428516 1001496
rect 446404 1001444 446456 1001496
rect 359464 1001308 359516 1001360
rect 372712 1001308 372764 1001360
rect 431408 1001308 431460 1001360
rect 461860 1001308 461912 1001360
rect 93492 1001172 93544 1001224
rect 101588 1001172 101640 1001224
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 423404 1001172 423456 1001224
rect 466460 1001172 466512 1001224
rect 496728 1001172 496780 1001224
rect 522764 1001172 522816 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 98000 1000492 98052 1000544
rect 100484 1000492 100536 1000544
rect 92848 999744 92900 999796
rect 98828 999744 98880 999796
rect 504364 999744 504416 999796
rect 519820 999744 519872 999796
rect 558184 999744 558236 999796
rect 568120 999744 568172 999796
rect 518900 999200 518952 999252
rect 524052 999200 524104 999252
rect 256700 999132 256752 999184
rect 258172 999132 258224 999184
rect 440884 999064 440936 999116
rect 444288 999064 444340 999116
rect 516968 999064 517020 999116
rect 520188 999064 520240 999116
rect 370504 998792 370556 998844
rect 378048 998792 378100 998844
rect 499304 998792 499356 998844
rect 516876 998792 516928 998844
rect 517520 998792 517572 998844
rect 523684 998792 523736 998844
rect 92480 998656 92532 998708
rect 93308 998656 93360 998708
rect 196624 998656 196676 998708
rect 204352 998656 204404 998708
rect 443644 998656 443696 998708
rect 472624 998656 472676 998708
rect 499580 998656 499632 998708
rect 517520 998656 517572 998708
rect 303068 998588 303120 998640
rect 308956 998588 309008 998640
rect 200856 998520 200908 998572
rect 203892 998520 203944 998572
rect 351828 998520 351880 998572
rect 382280 998520 382332 998572
rect 427728 998520 427780 998572
rect 456064 998520 456116 998572
rect 464804 998520 464856 998572
rect 472256 998520 472308 998572
rect 500316 998520 500368 998572
rect 522948 998520 523000 998572
rect 303252 998452 303304 998504
rect 305276 998452 305328 998504
rect 92296 998384 92348 998436
rect 98000 998384 98052 998436
rect 144184 998384 144236 998436
rect 155224 998384 155276 998436
rect 195520 998384 195572 998436
rect 204168 998384 204220 998436
rect 247408 998384 247460 998436
rect 259000 998384 259052 998436
rect 354404 998384 354456 998436
rect 383568 998384 383620 998436
rect 429936 998384 429988 998436
rect 472072 998384 472124 998436
rect 500960 998384 501012 998436
rect 523868 998384 523920 998436
rect 196808 998248 196860 998300
rect 202696 998248 202748 998300
rect 247224 998248 247276 998300
rect 251088 998248 251140 998300
rect 304264 998248 304316 998300
rect 307300 998248 307352 998300
rect 371884 998248 371936 998300
rect 372988 998248 373040 998300
rect 374644 998248 374696 998300
rect 379152 998248 379204 998300
rect 456064 998248 456116 998300
rect 461124 998248 461176 998300
rect 202144 998112 202196 998164
rect 205548 998112 205600 998164
rect 249064 998112 249116 998164
rect 253664 998112 253716 998164
rect 256332 998112 256384 998164
rect 257344 998112 257396 998164
rect 304448 998112 304500 998164
rect 306932 998112 306984 998164
rect 199384 998044 199436 998096
rect 201868 998044 201920 998096
rect 555424 998044 555476 998096
rect 557172 998044 557224 998096
rect 591488 998044 591540 998096
rect 625712 998044 625764 998096
rect 202328 997976 202380 998028
rect 204720 997976 204772 998028
rect 250444 997976 250496 998028
rect 253296 997976 253348 998028
rect 302884 997976 302936 998028
rect 306104 997976 306156 998028
rect 307024 997976 307076 998028
rect 308956 997976 309008 998028
rect 550548 997976 550600 998028
rect 553124 997976 553176 998028
rect 195336 997908 195388 997960
rect 200672 997908 200724 997960
rect 254584 997908 254636 997960
rect 256516 997908 256568 997960
rect 257344 997908 257396 997960
rect 259000 997908 259052 997960
rect 259828 997908 259880 997960
rect 262312 997908 262364 997960
rect 377404 997908 377456 997960
rect 383200 997908 383252 997960
rect 591120 997908 591172 997960
rect 625528 997908 625580 997960
rect 201040 997840 201092 997892
rect 203524 997840 203576 997892
rect 247776 997840 247828 997892
rect 252468 997840 252520 997892
rect 305644 997840 305696 997892
rect 307760 997840 307812 997892
rect 308404 997840 308456 997892
rect 310612 997840 310664 997892
rect 461860 997840 461912 997892
rect 463884 997840 463936 997892
rect 196072 997772 196124 997824
rect 198372 997772 198424 997824
rect 254952 997772 255004 997824
rect 256976 997772 257028 997824
rect 258172 997772 258224 997824
rect 259460 997772 259512 997824
rect 260196 997772 260248 997824
rect 262496 997772 262548 997824
rect 378784 997772 378836 997824
rect 383384 997772 383436 997824
rect 551744 997772 551796 997824
rect 553124 997772 553176 997824
rect 591304 997772 591356 997824
rect 625344 997772 625396 997824
rect 93308 997704 93360 997756
rect 103520 997704 103572 997756
rect 109500 997704 109552 997756
rect 116308 997704 116360 997756
rect 144000 997704 144052 997756
rect 160100 997704 160152 997756
rect 162124 997704 162176 997756
rect 170312 997704 170364 997756
rect 195704 997636 195756 997688
rect 209780 997704 209832 997756
rect 246580 997704 246632 997756
rect 254768 997704 254820 997756
rect 299112 997704 299164 997756
rect 311900 997704 311952 997756
rect 365260 997704 365312 997756
rect 372528 997704 372580 997756
rect 399944 997704 399996 997756
rect 431960 997704 432012 997756
rect 432604 997704 432656 997756
rect 439872 997704 439924 997756
rect 464988 997704 465040 997756
rect 471060 997704 471112 997756
rect 488908 997704 488960 997756
rect 507860 997704 507912 997756
rect 509700 997704 509752 997756
rect 516692 997704 516744 997756
rect 540520 997636 540572 997688
rect 556988 997636 557040 997688
rect 566464 997636 566516 997688
rect 591488 997636 591540 997688
rect 108304 997568 108356 997620
rect 117228 997568 117280 997620
rect 144828 997568 144880 997620
rect 158720 997568 158772 997620
rect 360844 997568 360896 997620
rect 372344 997568 372396 997620
rect 422300 997568 422352 997620
rect 426256 997568 426308 997620
rect 431224 997568 431276 997620
rect 439688 997568 439740 997620
rect 489092 997568 489144 997620
rect 506480 997568 506532 997620
rect 509976 997568 510028 997620
rect 517060 997568 517112 997620
rect 554504 997500 554556 997552
rect 591120 997500 591172 997552
rect 540336 997364 540388 997416
rect 560300 997364 560352 997416
rect 573364 997364 573416 997416
rect 591304 997364 591356 997416
rect 200212 997228 200264 997280
rect 204904 997228 204956 997280
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 554688 997160 554740 997212
rect 568948 997160 569000 997212
rect 572628 997160 572680 997212
rect 623688 997160 623740 997212
rect 444288 997024 444340 997076
rect 470508 997024 470560 997076
rect 505744 997024 505796 997076
rect 520004 997024 520056 997076
rect 550548 997024 550600 997076
rect 620100 997024 620152 997076
rect 197360 996888 197412 996940
rect 200948 996888 201000 996940
rect 570604 996888 570656 996940
rect 590568 996888 590620 996940
rect 106924 996752 106976 996804
rect 110512 996752 110564 996804
rect 303252 996684 303304 996736
rect 304448 996684 304500 996736
rect 144828 996480 144880 996532
rect 150440 996480 150492 996532
rect 103888 996344 103940 996396
rect 144000 996344 144052 996396
rect 151268 996344 151320 996396
rect 199384 996344 199436 996396
rect 299388 996344 299440 996396
rect 360200 996344 360252 996396
rect 200948 996276 201000 996328
rect 206284 996276 206336 996328
rect 553308 996276 553360 996328
rect 93308 996208 93360 996260
rect 195704 996208 195756 996260
rect 247592 996208 247644 996260
rect 263692 996208 263744 996260
rect 618168 996208 618220 996260
rect 171784 996072 171836 996124
rect 211160 996072 211212 996124
rect 211804 996072 211856 996124
rect 262496 996072 262548 996124
rect 265808 996072 265860 996124
rect 316040 996072 316092 996124
rect 382924 996072 382976 996124
rect 433524 996072 433576 996124
rect 169392 995936 169444 995988
rect 171508 995936 171560 995988
rect 177304 995936 177356 995988
rect 212540 995936 212592 995988
rect 229744 995936 229796 995988
rect 262312 995936 262364 995988
rect 264244 995936 264296 995988
rect 299296 995936 299348 995988
rect 366364 995936 366416 995988
rect 400864 995936 400916 995988
rect 136456 995800 136508 995852
rect 143816 995800 143868 995852
rect 170680 995800 170732 995852
rect 171692 995800 171744 995852
rect 213184 995800 213236 995852
rect 261300 995800 261352 995852
rect 364892 995800 364944 995852
rect 402244 995800 402296 995852
rect 518164 995800 518216 995852
rect 524052 995800 524104 995852
rect 92664 995528 92716 995580
rect 97448 995528 97500 995580
rect 171048 995528 171100 995580
rect 246212 995528 246264 995580
rect 256332 995528 256384 995580
rect 383200 995528 383252 995580
rect 385040 995528 385092 995580
rect 415952 995528 416004 995580
rect 472624 995528 472676 995580
rect 473360 995528 473412 995580
rect 494704 995528 494756 995580
rect 511080 995528 511132 995580
rect 523684 995528 523736 995580
rect 524788 995528 524840 995580
rect 625712 995528 625764 995580
rect 626540 995528 626592 995580
rect 194876 995460 194928 995512
rect 197360 995460 197412 995512
rect 246764 995392 246816 995444
rect 253480 995392 253532 995444
rect 383476 995392 383528 995444
rect 385684 995392 385736 995444
rect 171692 995277 171744 995329
rect 189448 995324 189500 995376
rect 192944 995324 192996 995376
rect 193128 995324 193180 995376
rect 196072 995324 196124 995376
rect 228364 995324 228416 995376
rect 245292 995324 245344 995376
rect 245568 995324 245620 995376
rect 246580 995324 246632 995376
rect 292304 995324 292356 995376
rect 295984 995324 296036 995376
rect 296168 995324 296220 995376
rect 298468 995324 298520 995376
rect 396632 995324 396684 995376
rect 400128 995324 400180 995376
rect 362224 995256 362276 995308
rect 387800 995256 387852 995308
rect 171508 995165 171560 995217
rect 184802 995188 184854 995240
rect 194140 995188 194192 995240
rect 194324 995188 194376 995240
rect 195520 995188 195572 995240
rect 244234 995188 244286 995240
rect 247224 995188 247276 995240
rect 283472 995188 283524 995240
rect 300124 995188 300176 995240
rect 380900 995120 380952 995172
rect 489736 995120 489788 995172
rect 489920 995120 489972 995172
rect 172336 995052 172388 995104
rect 180616 995052 180668 995104
rect 202144 995052 202196 995104
rect 232872 995052 232924 995104
rect 257344 995052 257396 995104
rect 285956 995052 286008 995104
rect 309140 995052 309192 995104
rect 425152 995052 425204 995104
rect 484124 995052 484176 995104
rect 515404 995052 515456 995104
rect 537392 995052 537444 995104
rect 568120 995052 568172 995104
rect 629668 995052 629720 995104
rect 358728 994984 358780 995036
rect 398840 994984 398892 995036
rect 638868 994984 638920 995036
rect 640800 994984 640852 995036
rect 641720 994984 641772 995036
rect 660580 994983 660632 995035
rect 181444 994916 181496 994968
rect 200948 994916 201000 994968
rect 229008 994916 229060 994968
rect 246212 994916 246264 994968
rect 284116 994916 284168 994968
rect 308404 994916 308456 994968
rect 419448 994916 419500 994968
rect 568212 994916 568264 994968
rect 568948 994916 569000 994968
rect 78312 994780 78364 994832
rect 102784 994780 102836 994832
rect 129740 994780 129792 994832
rect 155960 994780 156012 994832
rect 170864 994829 170916 994881
rect 171232 994829 171284 994881
rect 363604 994848 363656 994900
rect 397000 994848 397052 994900
rect 640984 994848 641036 994900
rect 245292 994780 245344 994832
rect 247592 994780 247644 994832
rect 287152 994780 287204 994832
rect 296720 994780 296772 994832
rect 456248 994780 456300 994832
rect 471244 994780 471296 994832
rect 472440 994780 472492 994832
rect 475936 994780 475988 994832
rect 476120 994780 476172 994832
rect 485228 994780 485280 994832
rect 486608 994780 486660 994832
rect 489736 994780 489788 994832
rect 502984 994780 503036 994832
rect 534356 994780 534408 994832
rect 569224 994780 569276 994832
rect 635832 994780 635884 994832
rect 169392 994712 169444 994764
rect 243176 994712 243228 994764
rect 253204 994712 253256 994764
rect 259460 994712 259512 994764
rect 379152 994712 379204 994764
rect 397644 994712 397696 994764
rect 74632 994644 74684 994696
rect 81992 994644 82044 994696
rect 85488 994644 85540 994696
rect 98644 994644 98696 994696
rect 128452 994644 128504 994696
rect 153844 994644 153896 994696
rect 289544 994644 289596 994696
rect 305644 994644 305696 994696
rect 420828 994644 420880 994696
rect 590568 994644 590620 994696
rect 625344 994644 625396 994696
rect 630220 994644 630272 994696
rect 171048 994576 171100 994628
rect 287704 994576 287756 994628
rect 372712 994576 372764 994628
rect 393320 994576 393372 994628
rect 660764 994576 660816 994628
rect 74448 994508 74500 994560
rect 97264 994508 97316 994560
rect 132408 994508 132460 994560
rect 149704 994508 149756 994560
rect 170680 994440 170732 994492
rect 301320 994508 301372 994560
rect 470508 994508 470560 994560
rect 475660 994508 475712 994560
rect 475936 994508 475988 994560
rect 490104 994508 490156 994560
rect 520004 994508 520056 994560
rect 539232 994508 539284 994560
rect 567844 994508 567896 994560
rect 591304 994508 591356 994560
rect 660948 994508 661000 994560
rect 356704 994440 356756 994492
rect 393964 994440 394016 994492
rect 81348 994372 81400 994424
rect 85488 994372 85540 994424
rect 85672 994372 85724 994424
rect 100024 994372 100076 994424
rect 103888 994372 103940 994424
rect 121736 994372 121788 994424
rect 129096 994372 129148 994424
rect 151084 994372 151136 994424
rect 296812 994372 296864 994424
rect 304264 994372 304316 994424
rect 463884 994372 463936 994424
rect 191748 994304 191800 994356
rect 197360 994304 197412 994356
rect 229192 994304 229244 994356
rect 234068 994304 234120 994356
rect 73160 994236 73212 994288
rect 111892 994236 111944 994288
rect 150440 994236 150492 994288
rect 186504 994236 186556 994288
rect 139216 994168 139268 994220
rect 144552 994168 144604 994220
rect 231584 994168 231636 994220
rect 256700 994304 256752 994356
rect 287704 994304 287756 994356
rect 298836 994236 298888 994288
rect 360200 994236 360252 994288
rect 381176 994236 381228 994288
rect 426256 994236 426308 994288
rect 446128 994236 446180 994288
rect 466552 994372 466604 994424
rect 475752 994372 475804 994424
rect 476074 994372 476126 994424
rect 485228 994372 485280 994424
rect 487804 994372 487856 994424
rect 498108 994372 498160 994424
rect 538036 994372 538088 994424
rect 571984 994372 572036 994424
rect 639052 994372 639104 994424
rect 237472 994168 237524 994220
rect 254584 994168 254636 994220
rect 286508 994168 286560 994220
rect 289544 994168 289596 994220
rect 80704 994100 80756 994152
rect 85672 994100 85724 994152
rect 184940 994100 184992 994152
rect 196624 994100 196676 994152
rect 471060 994100 471112 994152
rect 476028 994100 476080 994152
rect 137560 994032 137612 994084
rect 141792 994032 141844 994084
rect 235908 994032 235960 994084
rect 253020 994032 253072 994084
rect 471244 993964 471296 994016
rect 481640 994100 481692 994152
rect 489920 994236 489972 994288
rect 524052 994236 524104 994288
rect 535552 994236 535604 994288
rect 482284 994100 482336 994152
rect 489552 994100 489604 994152
rect 574100 994032 574152 994084
rect 485964 993964 486016 994016
rect 228824 993896 228876 993948
rect 253204 993896 253256 993948
rect 574744 993896 574796 993948
rect 171232 993760 171284 993812
rect 195152 993760 195204 993812
rect 232228 993760 232280 993812
rect 237472 993760 237524 993812
rect 243176 993760 243228 993812
rect 247776 993760 247828 993812
rect 522764 993760 522816 993812
rect 660764 993760 660816 993812
rect 170864 993624 170916 993676
rect 195704 993624 195756 993676
rect 229376 993624 229428 993676
rect 238392 993624 238444 993676
rect 516508 993624 516560 993676
rect 660948 993624 661000 993676
rect 549168 993488 549220 993540
rect 639512 993488 639564 993540
rect 551744 993352 551796 993404
rect 637028 993352 637080 993404
rect 51724 993148 51776 993200
rect 107752 993148 107804 993200
rect 50344 993012 50396 993064
rect 108120 993012 108172 993064
rect 202880 993012 202932 993064
rect 213920 993012 213972 993064
rect 563704 993012 563756 993064
rect 608600 993012 608652 993064
rect 55864 992876 55916 992928
rect 146944 992876 146996 992928
rect 197360 992876 197412 992928
rect 251456 992876 251508 992928
rect 316684 992876 316736 992928
rect 364984 992876 365036 992928
rect 367928 992876 367980 992928
rect 429936 992876 429988 992928
rect 435548 992876 435600 992928
rect 494704 992876 494756 992928
rect 512828 992876 512880 992928
rect 527272 992876 527324 992928
rect 562508 992876 562560 992928
rect 660304 992876 660356 992928
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 48964 991584 49016 991636
rect 110696 991584 110748 991636
rect 138296 991584 138348 991636
rect 163136 991584 163188 991636
rect 54484 991448 54536 991500
rect 148324 991448 148376 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 318064 991448 318116 991500
rect 349160 991448 349212 991500
rect 367744 991448 367796 991500
rect 397828 991448 397880 991500
rect 435364 991448 435416 991500
rect 478972 991448 479024 991500
rect 512644 991448 512696 991500
rect 543832 991448 543884 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 164884 990836 164936 990888
rect 170772 990836 170824 990888
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 89720 990224 89772 990276
rect 112076 990224 112128 990276
rect 560944 990224 560996 990276
rect 668584 990224 668636 990276
rect 44824 990088 44876 990140
rect 109040 990088 109092 990140
rect 319444 990088 319496 990140
rect 332968 990088 333020 990140
rect 369124 990088 369176 990140
rect 414112 990088 414164 990140
rect 562324 990088 562376 990140
rect 669964 990088 670016 990140
rect 53288 988728 53340 988780
rect 95884 988728 95936 988780
rect 217324 986620 217376 986672
rect 219440 986620 219492 986672
rect 105820 986552 105872 986604
rect 106924 986552 106976 986604
rect 565084 986076 565136 986128
rect 592500 986076 592552 986128
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 436744 985940 436796 985992
rect 462780 985940 462832 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565268 985940 565320 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 667204 975672 667256 975724
rect 43444 961868 43496 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952416 36596 952468
rect 41696 952416 41748 952468
rect 37924 952212 37976 952264
rect 41696 952212 41748 952264
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 663064 948064 663116 948116
rect 46296 945956 46348 946008
rect 62120 945956 62172 946008
rect 35808 942692 35860 942744
rect 40408 942692 40460 942744
rect 35808 941332 35860 941384
rect 38476 941332 38528 941384
rect 35808 939836 35860 939888
rect 39488 939836 39540 939888
rect 39488 938136 39540 938188
rect 41696 938136 41748 938188
rect 38476 937524 38528 937576
rect 41696 937524 41748 937576
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 41328 934328 41380 934380
rect 41696 934328 41748 934380
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 663064 921816 663116 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 665824 909440 665876 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 670976 895636 671028 895688
rect 44088 892712 44140 892764
rect 42938 892202 42990 892254
rect 43076 891896 43128 891948
rect 44088 891828 44140 891880
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 651472 852116 651524 852168
rect 664444 852116 664496 852168
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 651840 841780 651892 841832
rect 669964 841780 670016 841832
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 35808 817028 35860 817080
rect 41696 817028 41748 817080
rect 35808 815600 35860 815652
rect 41604 815600 41656 815652
rect 651472 815600 651524 815652
rect 661684 815600 661736 815652
rect 35808 814240 35860 814292
rect 41420 814240 41472 814292
rect 41328 810704 41380 810756
rect 41696 810704 41748 810756
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 33048 802408 33100 802460
rect 41696 802408 41748 802460
rect 39304 801660 39356 801712
rect 41604 801660 41656 801712
rect 44824 793568 44876 793620
rect 62120 793568 62172 793620
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 652392 775548 652444 775600
rect 668400 775548 668452 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35532 768952 35584 769004
rect 39304 768952 39356 769004
rect 35348 768816 35400 768868
rect 40408 768816 40460 768868
rect 35808 768680 35860 768732
rect 40592 768680 40644 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35624 767320 35676 767372
rect 41328 767320 41380 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 35808 763240 35860 763292
rect 37924 763240 37976 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 31024 759636 31076 759688
rect 41512 759636 41564 759688
rect 35164 758276 35216 758328
rect 40592 758344 40644 758396
rect 37924 757732 37976 757784
rect 41604 757732 41656 757784
rect 675852 754264 675904 754316
rect 683120 754264 683172 754316
rect 676036 753584 676088 753636
rect 676588 753584 676640 753636
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 672908 734000 672960 734052
rect 673552 734000 673604 734052
rect 35808 730056 35860 730108
rect 41696 730056 41748 730108
rect 674104 728628 674156 728680
rect 673092 728424 673144 728476
rect 673920 728152 673972 728204
rect 674150 728084 674202 728136
rect 41328 725908 41380 725960
rect 41696 725908 41748 725960
rect 41328 724480 41380 724532
rect 41696 724480 41748 724532
rect 677324 724208 677376 724260
rect 683856 724208 683908 724260
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 36544 717340 36596 717392
rect 41420 717340 41472 717392
rect 34520 715640 34572 715692
rect 41696 715640 41748 715692
rect 33784 715504 33836 715556
rect 40316 715504 40368 715556
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 651472 709316 651524 709368
rect 664444 709316 664496 709368
rect 672540 707208 672592 707260
rect 673276 707208 673328 707260
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 651472 696940 651524 696992
rect 669964 696940 670016 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 35808 687216 35860 687268
rect 41420 687216 41472 687268
rect 35808 683340 35860 683392
rect 41512 683272 41564 683324
rect 35808 683136 35860 683188
rect 41696 683136 41748 683188
rect 651656 683136 651708 683188
rect 658924 683136 658976 683188
rect 35808 681980 35860 682032
rect 36544 681980 36596 682032
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35440 681708 35492 681760
rect 40960 681708 41012 681760
rect 35624 674092 35676 674144
rect 39672 674092 39724 674144
rect 36544 673140 36596 673192
rect 40592 673140 40644 673192
rect 32404 672732 32456 672784
rect 41696 672732 41748 672784
rect 37188 670964 37240 671016
rect 40132 670964 40184 671016
rect 651472 669332 651524 669384
rect 661684 669332 661736 669384
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651472 656888 651524 656940
rect 663064 656888 663116 656940
rect 54484 647844 54536 647896
rect 62120 647844 62172 647896
rect 35808 644444 35860 644496
rect 41696 644444 41748 644496
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639208 35860 639260
rect 40040 639208 40092 639260
rect 35348 639072 35400 639124
rect 41696 639072 41748 639124
rect 35532 638936 35584 638988
rect 36544 638936 36596 638988
rect 35808 637576 35860 637628
rect 41328 637576 41380 637628
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 33784 629892 33836 629944
rect 41696 629892 41748 629944
rect 651564 628532 651616 628584
rect 667204 628532 667256 628584
rect 48964 623772 49016 623824
rect 62120 623772 62172 623824
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 671068 616156 671120 616208
rect 671712 616156 671764 616208
rect 43628 612688 43680 612740
rect 43812 612620 43864 612672
rect 43996 612484 44048 612536
rect 43582 612280 43634 612332
rect 43720 612280 43772 612332
rect 46940 611872 46992 611924
rect 46112 611668 46164 611720
rect 45560 611464 45612 611516
rect 45744 611260 45796 611312
rect 44272 610920 44324 610972
rect 44379 610784 44431 610836
rect 44502 610716 44554 610768
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 661684 603100 661736 603152
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 41328 596028 41380 596080
rect 41604 596028 41656 596080
rect 41144 594736 41196 594788
rect 41696 594736 41748 594788
rect 40868 593240 40920 593292
rect 41604 593240 41656 593292
rect 40500 592288 40552 592340
rect 41604 592288 41656 592340
rect 675852 591336 675904 591388
rect 682384 591336 682436 591388
rect 652392 590656 652444 590708
rect 665824 590656 665876 590708
rect 33048 587120 33100 587172
rect 40132 587120 40184 587172
rect 35164 585896 35216 585948
rect 41696 585896 41748 585948
rect 31024 585760 31076 585812
rect 39396 585760 39448 585812
rect 40868 584536 40920 584588
rect 41604 584536 41656 584588
rect 50344 583720 50396 583772
rect 62120 583720 62172 583772
rect 671620 578212 671672 578264
rect 671436 577940 671488 577992
rect 651472 576852 651524 576904
rect 664444 576852 664496 576904
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 41328 557540 41380 557592
rect 41512 557540 41564 557592
rect 41328 554752 41380 554804
rect 41696 554752 41748 554804
rect 41144 552100 41196 552152
rect 41604 552100 41656 552152
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 40592 549380 40644 549432
rect 41604 549380 41656 549432
rect 41236 549244 41288 549296
rect 41696 549244 41748 549296
rect 41236 548088 41288 548140
rect 41696 548088 41748 548140
rect 31760 547816 31812 547868
rect 38292 547816 38344 547868
rect 675944 547612 675996 547664
rect 678244 547612 678296 547664
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 32404 542988 32456 543040
rect 41512 542988 41564 543040
rect 38292 542308 38344 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669964 536800 670016 536852
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 676864 520276 676916 520328
rect 683120 520276 683172 520328
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 676036 518780 676088 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 675852 503616 675904 503668
rect 679624 503616 679676 503668
rect 675852 500896 675904 500948
rect 681004 500896 681056 500948
rect 652576 494708 652628 494760
rect 663248 494708 663300 494760
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 677416 489880 677468 489932
rect 683120 489880 683172 489932
rect 651472 484440 651524 484492
rect 667204 484372 667256 484424
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 651472 470568 651524 470620
rect 665824 470568 665876 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 652392 456764 652444 456816
rect 661684 456764 661736 456816
rect 673460 456560 673512 456612
rect 673828 456016 673880 456068
rect 673736 455744 673788 455796
rect 673598 455540 673650 455592
rect 675852 455540 675904 455592
rect 677048 455540 677100 455592
rect 672264 455336 672316 455388
rect 673388 455200 673440 455252
rect 671804 454996 671856 455048
rect 673046 454860 673098 454912
rect 672908 454656 672960 454708
rect 673164 454588 673216 454640
rect 672816 454180 672868 454232
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672264 453908 672316 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 671344 430584 671396 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 41328 425008 41380 425060
rect 41696 425008 41748 425060
rect 41328 423784 41380 423836
rect 41604 423784 41656 423836
rect 41328 422288 41380 422340
rect 41604 422288 41656 422340
rect 41328 420928 41380 420980
rect 41604 420928 41656 420980
rect 651840 416780 651892 416832
rect 663064 416780 663116 416832
rect 33692 416168 33744 416220
rect 41696 416168 41748 416220
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 41144 387064 41196 387116
rect 41696 387064 41748 387116
rect 44640 385432 44692 385484
rect 45008 385432 45060 385484
rect 41328 382372 41380 382424
rect 41696 382372 41748 382424
rect 41144 382236 41196 382288
rect 41696 382236 41748 382288
rect 35808 379516 35860 379568
rect 41696 379516 41748 379568
rect 35808 375980 35860 376032
rect 39580 375980 39632 376032
rect 51724 375368 51776 375420
rect 62120 375368 62172 375420
rect 28908 371832 28960 371884
rect 41696 371832 41748 371884
rect 651840 364352 651892 364404
rect 661868 364352 661920 364404
rect 46388 362924 46440 362976
rect 62120 362924 62172 362976
rect 45008 355784 45060 355836
rect 45652 355784 45704 355836
rect 44640 355648 44692 355700
rect 44575 354832 44627 354884
rect 44575 354628 44627 354680
rect 44799 354424 44851 354476
rect 44686 354288 44738 354340
rect 45652 354016 45704 354068
rect 45928 353744 45980 353796
rect 45560 353200 45612 353252
rect 652392 350548 652444 350600
rect 667388 350548 667440 350600
rect 35808 343612 35860 343664
rect 40224 343612 40276 343664
rect 35808 339464 35860 339516
rect 36636 339464 36688 339516
rect 46204 336744 46256 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 667756 324300 667808 324352
rect 53288 322940 53340 322992
rect 62120 322940 62172 322992
rect 54484 310496 54536 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667204 310496 667256 310548
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675852 298052 675904 298104
rect 678980 298052 679032 298104
rect 676036 297916 676088 297968
rect 681004 297916 681056 297968
rect 41328 284928 41380 284980
rect 41696 284928 41748 284980
rect 37924 284724 37976 284776
rect 41696 284724 41748 284776
rect 651472 284316 651524 284368
rect 667572 284316 667624 284368
rect 464804 276768 464856 276820
rect 532792 276768 532844 276820
rect 482836 276632 482888 276684
rect 558828 276632 558880 276684
rect 103704 275952 103756 276004
rect 160744 275952 160796 276004
rect 166356 275952 166408 276004
rect 182088 275952 182140 276004
rect 188804 275952 188856 276004
rect 222844 275952 222896 276004
rect 385960 275952 386012 276004
rect 401600 275952 401652 276004
rect 432972 275952 433024 276004
rect 487896 275952 487948 276004
rect 512552 275952 512604 276004
rect 526904 275952 526956 276004
rect 527364 275952 527416 276004
rect 607312 275952 607364 276004
rect 88340 275816 88392 275868
rect 146944 275816 146996 275868
rect 149796 275816 149848 275868
rect 187884 275816 187936 275868
rect 393872 275816 393924 275868
rect 411076 275816 411128 275868
rect 411260 275816 411312 275868
rect 415768 275816 415820 275868
rect 423588 275816 423640 275868
rect 439412 275816 439464 275868
rect 443644 275816 443696 275868
rect 498568 275816 498620 275868
rect 504732 275816 504784 275868
rect 590752 275816 590804 275868
rect 260932 275748 260984 275800
rect 263508 275748 263560 275800
rect 96620 275680 96672 275732
rect 156604 275680 156656 275732
rect 174636 275680 174688 275732
rect 208676 275680 208728 275732
rect 212448 275680 212500 275732
rect 220544 275680 220596 275732
rect 232504 275680 232556 275732
rect 220728 275612 220780 275664
rect 224960 275612 225012 275664
rect 85948 275544 86000 275596
rect 150808 275544 150860 275596
rect 160468 275544 160520 275596
rect 172428 275544 172480 275596
rect 181720 275544 181772 275596
rect 218612 275544 218664 275596
rect 225420 275544 225472 275596
rect 242256 275544 242308 275596
rect 244372 275680 244424 275732
rect 247040 275680 247092 275732
rect 268016 275680 268068 275732
rect 269120 275680 269172 275732
rect 365904 275680 365956 275732
rect 369676 275680 369728 275732
rect 373080 275680 373132 275732
rect 385040 275680 385092 275732
rect 400220 275680 400272 275732
rect 418160 275680 418212 275732
rect 418344 275680 418396 275732
rect 435916 275680 435968 275732
rect 457444 275680 457496 275732
rect 516232 275680 516284 275732
rect 516692 275680 516744 275732
rect 604920 275680 604972 275732
rect 605104 275680 605156 275732
rect 616788 275680 616840 275732
rect 245660 275544 245712 275596
rect 347412 275544 347464 275596
rect 349620 275544 349672 275596
rect 352380 275544 352432 275596
rect 360200 275544 360252 275596
rect 376576 275544 376628 275596
rect 393320 275544 393372 275596
rect 395068 275544 395120 275596
rect 403992 275544 404044 275596
rect 407672 275544 407724 275596
rect 432328 275544 432380 275596
rect 438860 275544 438912 275596
rect 446496 275544 446548 275596
rect 453948 275544 454000 275596
rect 464252 275544 464304 275596
rect 464436 275544 464488 275596
rect 523408 275544 523460 275596
rect 525800 275544 525852 275596
rect 527364 275544 527416 275596
rect 532700 275544 532752 275596
rect 626172 275544 626224 275596
rect 76472 275408 76524 275460
rect 143264 275408 143316 275460
rect 148600 275408 148652 275460
rect 164148 275408 164200 275460
rect 167552 275408 167604 275460
rect 209044 275408 209096 275460
rect 218336 275408 218388 275460
rect 239404 275408 239456 275460
rect 253848 275408 253900 275460
rect 261484 275408 261536 275460
rect 349712 275408 349764 275460
rect 361396 275408 361448 275460
rect 362960 275408 363012 275460
rect 367284 275408 367336 275460
rect 367836 275408 367888 275460
rect 377956 275408 378008 275460
rect 382464 275408 382516 275460
rect 400404 275408 400456 275460
rect 403624 275408 403676 275460
rect 428832 275408 428884 275460
rect 435732 275408 435784 275460
rect 491484 275408 491536 275460
rect 494060 275408 494112 275460
rect 502064 275408 502116 275460
rect 505836 275408 505888 275460
rect 512736 275408 512788 275460
rect 525616 275408 525668 275460
rect 619088 275408 619140 275460
rect 626448 275408 626500 275460
rect 640432 275408 640484 275460
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 156880 275272 156932 275324
rect 199292 275272 199344 275324
rect 211252 275272 211304 275324
rect 232688 275272 232740 275324
rect 259736 275272 259788 275324
rect 268844 275272 268896 275324
rect 276296 275272 276348 275324
rect 284300 275272 284352 275324
rect 284576 275272 284628 275324
rect 290096 275272 290148 275324
rect 339132 275272 339184 275324
rect 353116 275272 353168 275324
rect 359464 275272 359516 275324
rect 370872 275272 370924 275324
rect 377404 275272 377456 275324
rect 396908 275272 396960 275324
rect 400404 275272 400456 275324
rect 425244 275272 425296 275324
rect 427820 275272 427872 275324
rect 443000 275272 443052 275324
rect 448244 275272 448296 275324
rect 509148 275272 509200 275324
rect 513748 275272 513800 275324
rect 533988 275272 534040 275324
rect 539508 275272 539560 275324
rect 542268 275272 542320 275324
rect 543280 275272 543332 275324
rect 645124 275272 645176 275324
rect 249064 275204 249116 275256
rect 253572 275204 253624 275256
rect 110788 275136 110840 275188
rect 164976 275136 165028 275188
rect 171048 275136 171100 275188
rect 191104 275136 191156 275188
rect 429200 275136 429252 275188
rect 480812 275136 480864 275188
rect 487160 275136 487212 275188
rect 544660 275136 544712 275188
rect 552572 275136 552624 275188
rect 560024 275136 560076 275188
rect 246764 275068 246816 275120
rect 256700 275068 256752 275120
rect 270408 275068 270460 275120
rect 276204 275068 276256 275120
rect 580264 275068 580316 275120
rect 583668 275068 583720 275120
rect 135628 275000 135680 275052
rect 167644 275000 167696 275052
rect 426256 275000 426308 275052
rect 477224 275000 477276 275052
rect 485044 275000 485096 275052
rect 494060 275000 494112 275052
rect 494428 275000 494480 275052
rect 537300 275000 537352 275052
rect 537668 275000 537720 275052
rect 538772 275000 538824 275052
rect 541992 275000 542044 275052
rect 549352 275000 549404 275052
rect 81256 274932 81308 274984
rect 86224 274932 86276 274984
rect 241980 274932 242032 274984
rect 244096 274932 244148 274984
rect 129648 274864 129700 274916
rect 136088 274864 136140 274916
rect 142712 274864 142764 274916
rect 166264 274864 166316 274916
rect 210056 274864 210108 274916
rect 212448 274864 212500 274916
rect 418528 274864 418580 274916
rect 422852 274864 422904 274916
rect 478972 274864 479024 274916
rect 482008 274864 482060 274916
rect 487804 274864 487856 274916
rect 530492 274864 530544 274916
rect 530676 274864 530728 274916
rect 541072 274864 541124 274916
rect 545120 274864 545172 274916
rect 552940 274864 552992 274916
rect 559196 274864 559248 274916
rect 567016 274864 567068 274916
rect 199476 274796 199528 274848
rect 202788 274796 202840 274848
rect 243176 274796 243228 274848
rect 249064 274796 249116 274848
rect 263232 274796 263284 274848
rect 266452 274796 266504 274848
rect 277492 274796 277544 274848
rect 283196 274796 283248 274848
rect 289268 274796 289320 274848
rect 293408 274796 293460 274848
rect 336648 274796 336700 274848
rect 343640 274796 343692 274848
rect 369860 274796 369912 274848
rect 375564 274796 375616 274848
rect 146208 274728 146260 274780
rect 149704 274728 149756 274780
rect 150992 274728 151044 274780
rect 152740 274728 152792 274780
rect 163964 274728 164016 274780
rect 170404 274728 170456 274780
rect 172244 274728 172296 274780
rect 174912 274728 174964 274780
rect 208860 274728 208912 274780
rect 210608 274728 210660 274780
rect 415308 274728 415360 274780
rect 419356 274728 419408 274780
rect 423036 274728 423088 274780
rect 424048 274728 424100 274780
rect 471888 274728 471940 274780
rect 496176 274728 496228 274780
rect 510528 274728 510580 274780
rect 519820 274728 519872 274780
rect 523684 274728 523736 274780
rect 545856 274728 545908 274780
rect 551284 274728 551336 274780
rect 574192 274728 574244 274780
rect 71780 274660 71832 274712
rect 73804 274660 73856 274712
rect 74080 274660 74132 274712
rect 77208 274660 77260 274712
rect 257344 274660 257396 274712
rect 260196 274660 260248 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 290464 274660 290516 274712
rect 294328 274660 294380 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 298744 274660 298796 274712
rect 300124 274660 300176 274712
rect 324964 274660 325016 274712
rect 327080 274660 327132 274712
rect 331404 274660 331456 274712
rect 335360 274660 335412 274712
rect 337108 274660 337160 274712
rect 338948 274660 339000 274712
rect 344284 274660 344336 274712
rect 347228 274660 347280 274712
rect 360200 274660 360252 274712
rect 363788 274660 363840 274712
rect 368756 274660 368808 274712
rect 373264 274660 373316 274712
rect 120264 274592 120316 274644
rect 175280 274592 175332 274644
rect 204720 274592 204772 274644
rect 218796 274592 218848 274644
rect 403992 274592 404044 274644
rect 438860 274592 438912 274644
rect 114284 274456 114336 274508
rect 171600 274456 171652 274508
rect 179328 274456 179380 274508
rect 213184 274456 213236 274508
rect 378784 274456 378836 274508
rect 395712 274456 395764 274508
rect 409236 274456 409288 274508
rect 453580 274660 453632 274712
rect 498476 274660 498528 274712
rect 499764 274660 499816 274712
rect 501604 274660 501656 274712
rect 505652 274660 505704 274712
rect 506480 274660 506532 274712
rect 510344 274660 510396 274712
rect 619180 274660 619232 274712
rect 623872 274660 623924 274712
rect 458824 274592 458876 274644
rect 484308 274592 484360 274644
rect 493140 274592 493192 274644
rect 494428 274592 494480 274644
rect 522396 274592 522448 274644
rect 595444 274592 595496 274644
rect 453304 274456 453356 274508
rect 478420 274456 478472 274508
rect 481364 274456 481416 274508
rect 556436 274456 556488 274508
rect 559564 274456 559616 274508
rect 587164 274456 587216 274508
rect 93032 274320 93084 274372
rect 95884 274320 95936 274372
rect 97724 274320 97776 274372
rect 158812 274320 158864 274372
rect 180524 274320 180576 274372
rect 216956 274320 217008 274372
rect 223120 274320 223172 274372
rect 247224 274320 247276 274372
rect 384948 274320 385000 274372
rect 400220 274320 400272 274372
rect 416596 274320 416648 274372
rect 453948 274320 454000 274372
rect 474372 274320 474424 274372
rect 523684 274320 523736 274372
rect 537484 274320 537536 274372
rect 613200 274320 613252 274372
rect 95424 274184 95476 274236
rect 157616 274184 157668 274236
rect 165620 274184 165672 274236
rect 205732 274184 205784 274236
rect 213644 274184 213696 274236
rect 240416 274184 240468 274236
rect 362776 274184 362828 274236
rect 386236 274184 386288 274236
rect 400128 274184 400180 274236
rect 423588 274184 423640 274236
rect 427452 274184 427504 274236
rect 479340 274184 479392 274236
rect 486976 274184 487028 274236
rect 563520 274184 563572 274236
rect 563704 274184 563756 274236
rect 612004 274184 612056 274236
rect 75276 274048 75328 274100
rect 142160 274048 142212 274100
rect 147404 274048 147456 274100
rect 193312 274048 193364 274100
rect 193496 274048 193548 274100
rect 204720 274048 204772 274100
rect 206560 274048 206612 274100
rect 234620 274048 234672 274100
rect 245660 274048 245712 274100
rect 254032 274048 254084 274100
rect 269120 274048 269172 274100
rect 278780 274048 278832 274100
rect 349896 274048 349948 274100
rect 362592 274048 362644 274100
rect 368296 274048 368348 274100
rect 394516 274048 394568 274100
rect 395344 274048 395396 274100
rect 426440 274048 426492 274100
rect 431684 274048 431736 274100
rect 485504 274048 485556 274100
rect 529848 274048 529900 274100
rect 532700 274048 532752 274100
rect 540888 274048 540940 274100
rect 626448 274048 626500 274100
rect 77668 273912 77720 273964
rect 145104 273912 145156 273964
rect 145288 273912 145340 273964
rect 130844 273776 130896 273828
rect 181444 273776 181496 273828
rect 191840 273912 191892 273964
rect 191840 273776 191892 273828
rect 224960 273912 225012 273964
rect 245752 273912 245804 273964
rect 247040 273912 247092 273964
rect 262220 273912 262272 273964
rect 263508 273912 263560 273964
rect 273536 273912 273588 273964
rect 279792 273912 279844 273964
rect 287152 273912 287204 273964
rect 333796 273912 333848 273964
rect 344468 273912 344520 273964
rect 344652 273912 344704 273964
rect 349712 273912 349764 273964
rect 224960 273776 225012 273828
rect 350356 273776 350408 273828
rect 365904 273912 365956 273964
rect 367008 273912 367060 273964
rect 376576 273912 376628 273964
rect 376576 273776 376628 273828
rect 407488 273912 407540 273964
rect 420736 273912 420788 273964
rect 470140 273912 470192 273964
rect 470416 273912 470468 273964
rect 539876 273912 539928 273964
rect 542176 273912 542228 273964
rect 642732 273912 642784 273964
rect 397276 273776 397328 273828
rect 418344 273776 418396 273828
rect 439320 273776 439372 273828
rect 471336 273776 471388 273828
rect 473084 273776 473136 273828
rect 487160 273776 487212 273828
rect 488356 273776 488408 273828
rect 559196 273776 559248 273828
rect 124956 273640 125008 273692
rect 148416 273640 148468 273692
rect 155684 273640 155736 273692
rect 198096 273640 198148 273692
rect 438124 273640 438176 273692
rect 467840 273640 467892 273692
rect 484308 273640 484360 273692
rect 552572 273640 552624 273692
rect 446404 273504 446456 273556
rect 468944 273504 468996 273556
rect 478788 273504 478840 273556
rect 545120 273504 545172 273556
rect 552664 273504 552716 273556
rect 580080 273504 580132 273556
rect 475752 273368 475804 273420
rect 541992 273368 542044 273420
rect 330484 273232 330536 273284
rect 333060 273232 333112 273284
rect 128544 273164 128596 273216
rect 181260 273164 181312 273216
rect 268844 273164 268896 273216
rect 272616 273164 272668 273216
rect 401508 273164 401560 273216
rect 427820 273164 427872 273216
rect 438768 273164 438820 273216
rect 471888 273164 471940 273216
rect 475936 273164 475988 273216
rect 548156 273164 548208 273216
rect 111984 273028 112036 273080
rect 168380 273028 168432 273080
rect 182088 273028 182140 273080
rect 207296 273028 207348 273080
rect 102508 272892 102560 272944
rect 162124 272892 162176 272944
rect 190000 272892 190052 272944
rect 217416 273028 217468 273080
rect 382004 273028 382056 273080
rect 414572 273028 414624 273080
rect 424968 273028 425020 273080
rect 474924 273028 474976 273080
rect 500868 273028 500920 273080
rect 580264 273028 580316 273080
rect 217140 272892 217192 272944
rect 242900 272892 242952 272944
rect 388812 272892 388864 272944
rect 400404 272892 400456 272944
rect 406844 272892 406896 272944
rect 450084 272892 450136 272944
rect 451096 272892 451148 272944
rect 513932 272892 513984 272944
rect 520096 272892 520148 272944
rect 610808 272892 610860 272944
rect 94228 272756 94280 272808
rect 155960 272756 156012 272808
rect 187608 272756 187660 272808
rect 220084 272756 220136 272808
rect 220544 272756 220596 272808
rect 239220 272756 239272 272808
rect 343548 272756 343600 272808
rect 359004 272756 359056 272808
rect 360844 272756 360896 272808
rect 381544 272756 381596 272808
rect 394332 272756 394384 272808
rect 407672 272756 407724 272808
rect 408132 272756 408184 272808
rect 452108 272756 452160 272808
rect 452292 272756 452344 272808
rect 515128 272756 515180 272808
rect 524052 272756 524104 272808
rect 617984 272756 618036 272808
rect 82360 272620 82412 272672
rect 148232 272620 148284 272672
rect 161572 272620 161624 272672
rect 203064 272620 203116 272672
rect 203248 272620 203300 272672
rect 233240 272620 233292 272672
rect 239588 272620 239640 272672
rect 251824 272620 251876 272672
rect 252652 272620 252704 272672
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 187700 272484 187752 272536
rect 192300 272484 192352 272536
rect 225512 272484 225564 272536
rect 228824 272484 228876 272536
rect 238024 272484 238076 272536
rect 238484 272484 238536 272536
rect 258080 272484 258132 272536
rect 347596 272620 347648 272672
rect 366088 272620 366140 272672
rect 370964 272620 371016 272672
rect 399208 272620 399260 272672
rect 412272 272620 412324 272672
rect 457168 272620 457220 272672
rect 457996 272620 458048 272672
rect 522212 272620 522264 272672
rect 526812 272620 526864 272672
rect 621480 272620 621532 272672
rect 267832 272484 267884 272536
rect 273904 272484 273956 272536
rect 283012 272484 283064 272536
rect 322756 272484 322808 272536
rect 330668 272484 330720 272536
rect 331036 272484 331088 272536
rect 342444 272484 342496 272536
rect 356704 272484 356756 272536
rect 376760 272484 376812 272536
rect 380808 272484 380860 272536
rect 411996 272484 412048 272536
rect 413836 272484 413888 272536
rect 460664 272484 460716 272536
rect 461952 272484 462004 272536
rect 529296 272484 529348 272536
rect 529480 272484 529532 272536
rect 624700 272484 624752 272536
rect 127348 272348 127400 272400
rect 179880 272348 179932 272400
rect 258540 272348 258592 272400
rect 269764 272348 269816 272400
rect 429844 272348 429896 272400
rect 447692 272348 447744 272400
rect 471612 272348 471664 272400
rect 543464 272348 543516 272400
rect 116676 272212 116728 272264
rect 166080 272212 166132 272264
rect 166264 272212 166316 272264
rect 192024 272212 192076 272264
rect 467748 272212 467800 272264
rect 536380 272212 536432 272264
rect 541624 272212 541676 272264
rect 603724 272212 603776 272264
rect 152188 272076 152240 272128
rect 189816 272076 189868 272128
rect 447784 272076 447836 272128
rect 506848 272076 506900 272128
rect 507308 272076 507360 272128
rect 565912 272076 565964 272128
rect 516048 271940 516100 271992
rect 516692 271940 516744 271992
rect 517336 271940 517388 271992
rect 525800 271940 525852 271992
rect 121368 271804 121420 271856
rect 176752 271804 176804 271856
rect 187884 271804 187936 271856
rect 196440 271804 196492 271856
rect 283196 271804 283248 271856
rect 285128 271804 285180 271856
rect 375288 271804 375340 271856
rect 395068 271804 395120 271856
rect 433156 271804 433208 271856
rect 486700 271804 486752 271856
rect 496544 271804 496596 271856
rect 578884 271804 578936 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 104900 271668 104952 271720
rect 163320 271668 163372 271720
rect 164148 271668 164200 271720
rect 194784 271668 194836 271720
rect 197084 271668 197136 271720
rect 224224 271668 224276 271720
rect 224592 271668 224644 271720
rect 247776 271668 247828 271720
rect 363604 271668 363656 271720
rect 374368 271668 374420 271720
rect 384764 271668 384816 271720
rect 415308 271668 415360 271720
rect 437204 271668 437256 271720
rect 493784 271668 493836 271720
rect 499488 271668 499540 271720
rect 582472 271668 582524 271720
rect 106004 271532 106056 271584
rect 164792 271532 164844 271584
rect 178132 271532 178184 271584
rect 184204 271532 184256 271584
rect 184480 271532 184532 271584
rect 215944 271532 215996 271584
rect 216312 271532 216364 271584
rect 242072 271532 242124 271584
rect 340604 271532 340656 271584
rect 355140 271532 355192 271584
rect 355324 271532 355376 271584
rect 368480 271532 368532 271584
rect 369492 271532 369544 271584
rect 377404 271532 377456 271584
rect 379336 271532 379388 271584
rect 393872 271532 393924 271584
rect 395528 271532 395580 271584
rect 427636 271532 427688 271584
rect 434444 271532 434496 271584
rect 490288 271532 490340 271584
rect 494704 271532 494756 271584
rect 500500 271532 500552 271584
rect 501972 271532 502024 271584
rect 585600 271532 585652 271584
rect 585784 271532 585836 271584
rect 608508 271532 608560 271584
rect 89536 271396 89588 271448
rect 152372 271396 152424 271448
rect 162768 271396 162820 271448
rect 204720 271396 204772 271448
rect 205364 271396 205416 271448
rect 234988 271396 235040 271448
rect 248420 271396 248472 271448
rect 264336 271396 264388 271448
rect 348884 271396 348936 271448
rect 362960 271396 363012 271448
rect 366364 271396 366416 271448
rect 379152 271396 379204 271448
rect 383384 271396 383436 271448
rect 416964 271396 417016 271448
rect 418988 271396 419040 271448
rect 429660 271396 429712 271448
rect 439964 271396 440016 271448
rect 497372 271396 497424 271448
rect 504916 271396 504968 271448
rect 589556 271396 589608 271448
rect 592684 271396 592736 271448
rect 622676 271396 622728 271448
rect 68192 271260 68244 271312
rect 138480 271260 138532 271312
rect 139124 271260 139176 271312
rect 141608 271260 141660 271312
rect 141792 271260 141844 271312
rect 189632 271260 189684 271312
rect 195704 271260 195756 271312
rect 227904 271260 227956 271312
rect 237288 271260 237340 271312
rect 256976 271260 257028 271312
rect 260196 271260 260248 271312
rect 270960 271260 271012 271312
rect 271512 271260 271564 271312
rect 280896 271260 280948 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 325516 271260 325568 271312
rect 334164 271260 334216 271312
rect 334624 271260 334676 271312
rect 341340 271260 341392 271312
rect 354588 271260 354640 271312
rect 369860 271260 369912 271312
rect 372528 271260 372580 271312
rect 382464 271260 382516 271312
rect 387524 271260 387576 271312
rect 421380 271260 421432 271312
rect 421564 271260 421616 271312
rect 437020 271260 437072 271312
rect 445668 271260 445720 271312
rect 455788 271260 455840 271312
rect 465724 271260 465776 271312
rect 465908 271260 465960 271312
rect 507952 271260 508004 271312
rect 509148 271260 509200 271312
rect 596640 271260 596692 271312
rect 596824 271260 596876 271312
rect 629760 271260 629812 271312
rect 72976 271124 73028 271176
rect 142344 271124 142396 271176
rect 143264 271124 143316 271176
rect 144368 271124 144420 271176
rect 154304 271124 154356 271176
rect 197912 271124 197964 271176
rect 198280 271124 198332 271176
rect 229560 271124 229612 271176
rect 231400 271124 231452 271176
rect 252744 271124 252796 271176
rect 253572 271124 253624 271176
rect 265256 271124 265308 271176
rect 269488 271124 269540 271176
rect 279240 271124 279292 271176
rect 285772 271124 285824 271176
rect 291200 271124 291252 271176
rect 328092 271124 328144 271176
rect 337752 271124 337804 271176
rect 339316 271124 339368 271176
rect 354312 271124 354364 271176
rect 362684 271124 362736 271176
rect 387156 271124 387208 271176
rect 391756 271124 391808 271176
rect 403624 271124 403676 271176
rect 404176 271124 404228 271176
rect 445300 271124 445352 271176
rect 449808 271124 449860 271176
rect 456340 271124 456392 271176
rect 504180 271124 504232 271176
rect 83556 270988 83608 271040
rect 123484 270988 123536 271040
rect 123760 270988 123812 271040
rect 177488 270988 177540 271040
rect 418068 270988 418120 271040
rect 463792 270988 463844 271040
rect 465724 270988 465776 271040
rect 511540 271124 511592 271176
rect 511908 271124 511960 271176
rect 600228 271124 600280 271176
rect 623044 271124 623096 271176
rect 643928 271124 643980 271176
rect 504548 270988 504600 271040
rect 575388 270988 575440 271040
rect 576124 270988 576176 271040
rect 594340 270988 594392 271040
rect 134432 270852 134484 270904
rect 184940 270852 184992 270904
rect 405004 270852 405056 270904
rect 434720 270852 434772 270904
rect 456064 270852 456116 270904
rect 465908 270852 465960 270904
rect 492036 270852 492088 270904
rect 571800 270852 571852 270904
rect 113180 270716 113232 270768
rect 154028 270716 154080 270768
rect 175832 270716 175884 270768
rect 206284 270716 206336 270768
rect 425704 270716 425756 270768
rect 448888 270716 448940 270768
rect 463792 270716 463844 270768
rect 466644 270716 466696 270768
rect 467104 270716 467156 270768
rect 525340 270716 525392 270768
rect 526444 270716 526496 270768
rect 576584 270716 576636 270768
rect 414480 270580 414532 270632
rect 437940 270580 437992 270632
rect 445024 270580 445076 270632
rect 494704 270580 494756 270632
rect 495348 270580 495400 270632
rect 504548 270580 504600 270632
rect 100668 270444 100720 270496
rect 119804 270444 119856 270496
rect 122748 270444 122800 270496
rect 176200 270444 176252 270496
rect 176936 270444 176988 270496
rect 214748 270444 214800 270496
rect 230388 270444 230440 270496
rect 252100 270444 252152 270496
rect 275100 270444 275152 270496
rect 276020 270444 276072 270496
rect 281448 270444 281500 270496
rect 285680 270444 285732 270496
rect 292856 270444 292908 270496
rect 293960 270444 294012 270496
rect 297916 270444 297968 270496
rect 299572 270444 299624 270496
rect 299940 270444 299992 270496
rect 300860 270444 300912 270496
rect 327080 270444 327132 270496
rect 328460 270444 328512 270496
rect 78864 270308 78916 270360
rect 132592 270308 132644 270360
rect 133788 270308 133840 270360
rect 183652 270308 183704 270360
rect 185216 270308 185268 270360
rect 186320 270308 186372 270360
rect 186504 270308 186556 270360
rect 202328 270308 202380 270360
rect 202788 270308 202840 270360
rect 205916 270308 205968 270360
rect 219532 270308 219584 270360
rect 244924 270308 244976 270360
rect 278596 270308 278648 270360
rect 286324 270308 286376 270360
rect 291660 270308 291712 270360
rect 295524 270308 295576 270360
rect 85488 270172 85540 270224
rect 149428 270172 149480 270224
rect 153292 270172 153344 270224
rect 169852 270172 169904 270224
rect 170036 270172 170088 270224
rect 210148 270172 210200 270224
rect 210608 270172 210660 270224
rect 237472 270172 237524 270224
rect 255228 270172 255280 270224
rect 269396 270172 269448 270224
rect 288256 270172 288308 270224
rect 292948 270172 293000 270224
rect 321100 270172 321152 270224
rect 327448 270172 327500 270224
rect 329380 270172 329432 270224
rect 339500 270172 339552 270224
rect 345940 270172 345992 270224
rect 360200 270444 360252 270496
rect 359188 270308 359240 270360
rect 382280 270444 382332 270496
rect 383844 270444 383896 270496
rect 391940 270444 391992 270496
rect 400588 270444 400640 270496
rect 441620 270444 441672 270496
rect 453580 270444 453632 270496
rect 516508 270444 516560 270496
rect 517796 270444 517848 270496
rect 597560 270444 597612 270496
rect 377956 270308 378008 270360
rect 387800 270308 387852 270360
rect 407212 270308 407264 270360
rect 451464 270308 451516 270360
rect 456432 270308 456484 270360
rect 520280 270308 520332 270360
rect 523132 270308 523184 270360
rect 605104 270308 605156 270360
rect 360200 270172 360252 270224
rect 383660 270172 383712 270224
rect 387708 270172 387760 270224
rect 401784 270172 401836 270224
rect 410524 270172 410576 270224
rect 455420 270172 455472 270224
rect 461400 270172 461452 270224
rect 527180 270172 527232 270224
rect 528100 270172 528152 270224
rect 619180 270172 619232 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 67548 270036 67600 270088
rect 75920 270036 75972 270088
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 158628 270036 158680 270088
rect 201040 270036 201092 270088
rect 201776 270036 201828 270088
rect 77208 269900 77260 269952
rect 143908 269900 143960 269952
rect 144092 269900 144144 269952
rect 190828 269900 190880 269952
rect 204168 269900 204220 269952
rect 205088 269900 205140 269952
rect 205916 270036 205968 270088
rect 230848 270036 230900 270088
rect 244096 270036 244148 270088
rect 260656 270036 260708 270088
rect 262036 270036 262088 270088
rect 274732 270036 274784 270088
rect 316960 270036 317012 270088
rect 321560 270036 321612 270088
rect 332232 270036 332284 270088
rect 336648 270036 336700 270088
rect 232504 269900 232556 269952
rect 233700 269900 233752 269952
rect 243912 269900 243964 269952
rect 245476 269900 245528 269952
rect 263140 269900 263192 269952
rect 266268 269900 266320 269952
rect 272892 269900 272944 269952
rect 286968 269900 287020 269952
rect 292120 269900 292172 269952
rect 323584 269900 323636 269952
rect 331220 269900 331272 269952
rect 336004 269900 336056 269952
rect 347412 270036 347464 270088
rect 349712 270036 349764 270088
rect 357440 270036 357492 270088
rect 364156 270036 364208 270088
rect 389180 270036 389232 270088
rect 389640 270036 389692 270088
rect 405740 270036 405792 270088
rect 409696 270036 409748 270088
rect 454132 270036 454184 270088
rect 454500 270036 454552 270088
rect 473360 270036 473412 270088
rect 525524 270036 525576 270088
rect 619640 270036 619692 270088
rect 346768 269900 346820 269952
rect 364340 269900 364392 269952
rect 364984 269900 365036 269952
rect 390560 269900 390612 269952
rect 391940 269900 391992 269952
rect 409880 269900 409932 269952
rect 412456 269900 412508 269952
rect 458180 269900 458232 269952
rect 458548 269900 458600 269952
rect 524420 269900 524472 269952
rect 531688 269900 531740 269952
rect 627920 269900 627972 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 140688 269764 140740 269816
rect 188620 269764 188672 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 119068 269628 119120 269680
rect 173348 269628 173400 269680
rect 174912 269628 174964 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 204168 269492 204220 269544
rect 136088 269356 136140 269408
rect 180892 269356 180944 269408
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 250260 269764 250312 269816
rect 266636 269764 266688 269816
rect 266820 269764 266872 269816
rect 278044 269764 278096 269816
rect 314476 269764 314528 269816
rect 318984 269764 319036 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336832 269764 336884 269816
rect 350540 269764 350592 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 374920 269764 374972 269816
rect 404360 269764 404412 269816
rect 417148 269764 417200 269816
rect 465080 269764 465132 269816
rect 466000 269764 466052 269816
rect 534356 269764 534408 269816
rect 535552 269764 535604 269816
rect 633532 269764 633584 269816
rect 236092 269628 236144 269680
rect 253756 269628 253808 269680
rect 341800 269628 341852 269680
rect 349712 269628 349764 269680
rect 393320 269628 393372 269680
rect 412640 269628 412692 269680
rect 422116 269628 422168 269680
rect 472072 269628 472124 269680
rect 474648 269628 474700 269680
rect 546500 269628 546552 269680
rect 205088 269492 205140 269544
rect 223488 269492 223540 269544
rect 388168 269492 388220 269544
rect 423036 269492 423088 269544
rect 424600 269492 424652 269544
rect 476120 269492 476172 269544
rect 476764 269492 476816 269544
rect 549904 269492 549956 269544
rect 210976 269356 211028 269408
rect 273076 269356 273128 269408
rect 277400 269356 277452 269408
rect 401692 269356 401744 269408
rect 419540 269356 419592 269408
rect 419816 269356 419868 269408
rect 462320 269356 462372 269408
rect 507952 269356 508004 269408
rect 560300 269356 560352 269408
rect 251456 269220 251508 269272
rect 258264 269220 258316 269272
rect 295340 269220 295392 269272
rect 297916 269220 297968 269272
rect 441620 269220 441672 269272
rect 460940 269220 460992 269272
rect 463516 269220 463568 269272
rect 531320 269220 531372 269272
rect 146944 269152 146996 269204
rect 153844 269152 153896 269204
rect 294144 269084 294196 269136
rect 297088 269084 297140 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 342260 269084 342312 269136
rect 345112 269084 345164 269136
rect 115848 269016 115900 269068
rect 171232 269016 171284 269068
rect 428740 269016 428792 269068
rect 475200 269016 475252 269068
rect 475384 269016 475436 269068
rect 494244 269016 494296 269068
rect 495808 269016 495860 269068
rect 576860 269016 576912 269068
rect 108948 268880 109000 268932
rect 166264 268880 166316 268932
rect 172428 268880 172480 268932
rect 204352 268880 204404 268932
rect 208216 268880 208268 268932
rect 227720 268880 227772 268932
rect 382372 268880 382424 268932
rect 411260 268880 411312 268932
rect 429568 268880 429620 268932
rect 483112 268880 483164 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 582288 268880 582340 268932
rect 600596 268880 600648 268932
rect 99288 268744 99340 268796
rect 91008 268608 91060 268660
rect 99288 268608 99340 268660
rect 110236 268744 110288 268796
rect 167920 268744 167972 268796
rect 173808 268744 173860 268796
rect 212632 268744 212684 268796
rect 215208 268744 215260 268796
rect 220820 268744 220872 268796
rect 377404 268744 377456 268796
rect 408500 268744 408552 268796
rect 416412 268744 416464 268796
rect 433340 268744 433392 268796
rect 441160 268744 441212 268796
rect 498476 268744 498528 268796
rect 500684 268744 500736 268796
rect 583852 268744 583904 268796
rect 160468 268608 160520 268660
rect 168656 268608 168708 268660
rect 208492 268608 208544 268660
rect 208676 268608 208728 268660
rect 214288 268608 214340 268660
rect 228088 268608 228140 268660
rect 250720 268608 250772 268660
rect 256700 268608 256752 268660
rect 263968 268608 264020 268660
rect 355876 268608 355928 268660
rect 367836 268608 367888 268660
rect 372344 268608 372396 268660
rect 385960 268608 386012 268660
rect 387340 268608 387392 268660
rect 418528 268608 418580 268660
rect 443920 268608 443972 268660
rect 502340 268608 502392 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 160008 268472 160060 268524
rect 200396 268472 200448 268524
rect 212448 268472 212500 268524
rect 238300 268472 238352 268524
rect 241336 268472 241388 268524
rect 256700 268472 256752 268524
rect 266452 268472 266504 268524
rect 275560 268472 275612 268524
rect 326068 268472 326120 268524
rect 331404 268472 331456 268524
rect 335176 268472 335228 268524
rect 347780 268472 347832 268524
rect 357532 268472 357584 268524
rect 379520 268472 379572 268524
rect 398748 268472 398800 268524
rect 430580 268472 430632 268524
rect 433708 268472 433760 268524
rect 488540 268472 488592 268524
rect 510712 268472 510764 268524
rect 598940 268472 598992 268524
rect 87144 268336 87196 268388
rect 152188 268336 152240 268388
rect 152740 268336 152792 268388
rect 196072 268336 196124 268388
rect 200580 268336 200632 268388
rect 231676 268336 231728 268388
rect 234804 268336 234856 268388
rect 255688 268336 255740 268388
rect 256516 268336 256568 268388
rect 270592 268336 270644 268388
rect 276204 268336 276256 268388
rect 280528 268336 280580 268388
rect 337660 268336 337712 268388
rect 351920 268336 351972 268388
rect 352564 268336 352616 268388
rect 368756 268336 368808 268388
rect 369952 268336 370004 268388
rect 397460 268336 397512 268388
rect 399760 268336 399812 268388
rect 440240 268336 440292 268388
rect 459560 268336 459612 268388
rect 517612 268336 517664 268388
rect 534724 268336 534776 268388
rect 535736 268336 535788 268388
rect 536380 268336 536432 268388
rect 634820 268336 634872 268388
rect 118608 268200 118660 268252
rect 174544 268200 174596 268252
rect 413008 268200 413060 268252
rect 459744 268200 459796 268252
rect 469496 268200 469548 268252
rect 475384 268200 475436 268252
rect 490840 268200 490892 268252
rect 569960 268200 570012 268252
rect 137008 268064 137060 268116
rect 182180 268064 182232 268116
rect 422300 268064 422352 268116
rect 443276 268064 443328 268116
rect 475200 268064 475252 268116
rect 478972 268064 479024 268116
rect 489184 268064 489236 268116
rect 567292 268064 567344 268116
rect 448612 267928 448664 267980
rect 506480 267928 506532 267980
rect 436192 267792 436244 267844
rect 491852 267792 491904 267844
rect 493324 267792 493376 267844
rect 551284 267792 551336 267844
rect 328552 267724 328604 267776
rect 337108 267724 337160 267776
rect 132408 267656 132460 267708
rect 184480 267656 184532 267708
rect 189816 267656 189868 267708
rect 197728 267656 197780 267708
rect 204168 267656 204220 267708
rect 218428 267656 218480 267708
rect 224224 267656 224276 267708
rect 229192 267656 229244 267708
rect 99288 267520 99340 267572
rect 154672 267520 154724 267572
rect 167644 267520 167696 267572
rect 186964 267520 187016 267572
rect 195244 267520 195296 267572
rect 216772 267520 216824 267572
rect 218796 267520 218848 267572
rect 226708 267520 226760 267572
rect 107660 267384 107712 267436
rect 167092 267384 167144 267436
rect 170404 267384 170456 267436
rect 95884 267248 95936 267300
rect 156420 267248 156472 267300
rect 156604 267248 156656 267300
rect 159640 267248 159692 267300
rect 160744 267248 160796 267300
rect 164608 267248 164660 267300
rect 166448 267248 166500 267300
rect 172888 267248 172940 267300
rect 186320 267384 186372 267436
rect 221740 267384 221792 267436
rect 227720 267384 227772 267436
rect 236644 267384 236696 267436
rect 340972 267384 341024 267436
rect 356060 267724 356112 267776
rect 368112 267656 368164 267708
rect 378784 267656 378836 267708
rect 380624 267656 380676 267708
rect 393320 267656 393372 267708
rect 402244 267656 402296 267708
rect 422300 267656 422352 267708
rect 430396 267656 430448 267708
rect 458824 267656 458876 267708
rect 460204 267656 460256 267708
rect 512552 267656 512604 267708
rect 514392 267656 514444 267708
rect 541624 267656 541676 267708
rect 357072 267520 357124 267572
rect 358360 267384 358412 267436
rect 360844 267384 360896 267436
rect 373264 267520 373316 267572
rect 387708 267520 387760 267572
rect 404728 267520 404780 267572
rect 429844 267520 429896 267572
rect 436744 267520 436796 267572
rect 441620 267520 441672 267572
rect 442816 267520 442868 267572
rect 485044 267520 485096 267572
rect 487160 267520 487212 267572
rect 487804 267520 487856 267572
rect 494704 267520 494756 267572
rect 501604 267520 501656 267572
rect 502432 267520 502484 267572
rect 366364 267384 366416 267436
rect 375748 267384 375800 267436
rect 389640 267384 389692 267436
rect 394792 267384 394844 267436
rect 416412 267384 416464 267436
rect 419632 267384 419684 267436
rect 446404 267384 446456 267436
rect 450268 267384 450320 267436
rect 505836 267384 505888 267436
rect 507584 267520 507636 267572
rect 576124 267520 576176 267572
rect 508412 267384 508464 267436
rect 509884 267384 509936 267436
rect 517796 267384 517848 267436
rect 86224 267112 86276 267164
rect 148048 267112 148100 267164
rect 149704 267112 149756 267164
rect 194416 267112 194468 267164
rect 199292 267112 199344 267164
rect 201868 267112 201920 267164
rect 206284 267248 206336 267300
rect 213460 267248 213512 267300
rect 217416 267248 217468 267300
rect 219900 267248 219952 267300
rect 220084 267248 220136 267300
rect 222568 267248 222620 267300
rect 223488 267248 223540 267300
rect 234160 267248 234212 267300
rect 238024 267248 238076 267300
rect 251548 267248 251600 267300
rect 261484 267248 261536 267300
rect 268936 267248 268988 267300
rect 334348 267248 334400 267300
rect 344284 267248 344336 267300
rect 360844 267248 360896 267300
rect 373080 267248 373132 267300
rect 378232 267248 378284 267300
rect 206836 267112 206888 267164
rect 207020 267112 207072 267164
rect 73804 266976 73856 267028
rect 141424 266976 141476 267028
rect 146944 266976 146996 267028
rect 189448 266976 189500 267028
rect 191104 266976 191156 267028
rect 211804 266976 211856 267028
rect 215944 267112 215996 267164
rect 220084 267112 220136 267164
rect 220820 267112 220872 267164
rect 241612 267112 241664 267164
rect 243912 267112 243964 267164
rect 254860 267112 254912 267164
rect 282828 267112 282880 267164
rect 288808 267112 288860 267164
rect 324412 267112 324464 267164
rect 330484 267112 330536 267164
rect 333520 267112 333572 267164
rect 342260 267112 342312 267164
rect 350908 267112 350960 267164
rect 359464 267112 359516 267164
rect 363328 267112 363380 267164
rect 377956 267112 378008 267164
rect 220912 266976 220964 267028
rect 222016 266976 222068 267028
rect 246580 266976 246632 267028
rect 249064 266976 249116 267028
rect 261484 266976 261536 267028
rect 276020 266976 276072 267028
rect 283840 266976 283892 267028
rect 343364 266976 343416 267028
rect 352380 266976 352432 267028
rect 353392 266976 353444 267028
rect 363604 266976 363656 267028
rect 365812 266976 365864 267028
rect 383844 267112 383896 267164
rect 389824 267248 389876 267300
rect 395344 267248 395396 267300
rect 397092 267248 397144 267300
rect 421564 267248 421616 267300
rect 426072 267248 426124 267300
rect 453304 267248 453356 267300
rect 455236 267248 455288 267300
rect 510528 267248 510580 267300
rect 512368 267248 512420 267300
rect 582288 267384 582340 267436
rect 520648 267248 520700 267300
rect 537484 267248 537536 267300
rect 539692 267248 539744 267300
rect 540888 267248 540940 267300
rect 541348 267248 541400 267300
rect 542176 267248 542228 267300
rect 542360 267248 542412 267300
rect 623044 267248 623096 267300
rect 385684 267112 385736 267164
rect 401692 267112 401744 267164
rect 414664 267112 414716 267164
rect 436744 267112 436796 267164
rect 440332 267112 440384 267164
rect 443644 267112 443696 267164
rect 445300 267112 445352 267164
rect 494704 267112 494756 267164
rect 494888 267112 494940 267164
rect 507308 267112 507360 267164
rect 508228 267112 508280 267164
rect 522396 267112 522448 267164
rect 522672 267112 522724 267164
rect 526628 267112 526680 267164
rect 532240 267112 532292 267164
rect 596824 267112 596876 267164
rect 391940 266976 391992 267028
rect 392308 266976 392360 267028
rect 418988 266976 419040 267028
rect 422944 266976 422996 267028
rect 454500 266976 454552 267028
rect 454776 266976 454828 267028
rect 459192 266976 459244 267028
rect 459376 266976 459428 267028
rect 467104 266976 467156 267028
rect 467288 266976 467340 267028
rect 469496 266976 469548 267028
rect 119804 266840 119856 266892
rect 156604 266840 156656 266892
rect 169852 266840 169904 266892
rect 132592 266704 132644 266756
rect 147220 266704 147272 266756
rect 148508 266704 148560 266756
rect 179512 266704 179564 266756
rect 198188 266840 198240 266892
rect 200212 266840 200264 266892
rect 202328 266840 202380 266892
rect 207020 266840 207072 266892
rect 219900 266840 219952 266892
rect 223396 266840 223448 266892
rect 242256 266840 242308 266892
rect 249064 266840 249116 266892
rect 251824 266840 251876 266892
rect 259000 266840 259052 266892
rect 264980 266840 265032 266892
rect 276388 266840 276440 266892
rect 285680 266840 285732 266892
rect 287980 266840 288032 266892
rect 312820 266840 312872 266892
rect 316408 266840 316460 266892
rect 321928 266840 321980 266892
rect 327080 266840 327132 266892
rect 349252 266840 349304 266892
rect 355324 266840 355376 266892
rect 393136 266840 393188 266892
rect 398748 266840 398800 266892
rect 403072 266840 403124 266892
rect 404176 266840 404228 266892
rect 405556 266840 405608 266892
rect 425704 266840 425756 266892
rect 199384 266704 199436 266756
rect 232688 266704 232740 266756
rect 239128 266704 239180 266756
rect 317788 266704 317840 266756
rect 322940 266704 322992 266756
rect 390652 266704 390704 266756
rect 395528 266704 395580 266756
rect 398104 266704 398156 266756
rect 414480 266704 414532 266756
rect 423772 266704 423824 266756
rect 424968 266704 425020 266756
rect 425428 266704 425480 266756
rect 426256 266704 426308 266756
rect 427912 266704 427964 266756
rect 428924 266704 428976 266756
rect 312360 266636 312412 266688
rect 314660 266636 314712 266688
rect 123484 266568 123536 266620
rect 150532 266568 150584 266620
rect 154028 266568 154080 266620
rect 161940 266568 161992 266620
rect 162124 266568 162176 266620
rect 162952 266568 163004 266620
rect 141608 266432 141660 266484
rect 146944 266432 146996 266484
rect 156604 266432 156656 266484
rect 162124 266432 162176 266484
rect 170404 266500 170456 266552
rect 182180 266500 182232 266552
rect 186136 266500 186188 266552
rect 161940 266296 161992 266348
rect 165068 266364 165120 266416
rect 169576 266364 169628 266416
rect 181536 266364 181588 266416
rect 182824 266364 182876 266416
rect 184204 266364 184256 266416
rect 195244 266568 195296 266620
rect 316132 266568 316184 266620
rect 320548 266568 320600 266620
rect 418804 266568 418856 266620
rect 438124 266840 438176 266892
rect 446956 266840 447008 266892
rect 456064 266840 456116 266892
rect 457720 266840 457772 266892
rect 464436 266840 464488 266892
rect 437848 266704 437900 266756
rect 452752 266704 452804 266756
rect 457444 266704 457496 266756
rect 462688 266704 462740 266756
rect 469956 266840 470008 266892
rect 470140 266840 470192 266892
rect 530676 266976 530728 267028
rect 537208 266976 537260 267028
rect 636200 266976 636252 267028
rect 473452 266840 473504 266892
rect 474372 266840 474424 266892
rect 475108 266840 475160 266892
rect 475936 266840 475988 266892
rect 465172 266704 465224 266756
rect 513748 266840 513800 266892
rect 514024 266840 514076 266892
rect 518716 266840 518768 266892
rect 518900 266840 518952 266892
rect 526444 266840 526496 266892
rect 526628 266840 526680 266892
rect 615500 266840 615552 266892
rect 483204 266704 483256 266756
rect 487160 266704 487212 266756
rect 487528 266704 487580 266756
rect 494704 266704 494756 266756
rect 467288 266568 467340 266620
rect 467564 266568 467616 266620
rect 493140 266568 493192 266620
rect 497464 266704 497516 266756
rect 499948 266704 500000 266756
rect 500868 266704 500920 266756
rect 504088 266704 504140 266756
rect 504916 266704 504968 266756
rect 506572 266704 506624 266756
rect 507768 266704 507820 266756
rect 508412 266704 508464 266756
rect 559564 266704 559616 266756
rect 258264 266500 258316 266552
rect 267280 266500 267332 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 330208 266500 330260 266552
rect 334624 266500 334676 266552
rect 395620 266500 395672 266552
rect 313648 266432 313700 266484
rect 317420 266432 317472 266484
rect 200396 266364 200448 266416
rect 202696 266364 202748 266416
rect 213184 266364 213236 266416
rect 215944 266364 215996 266416
rect 222844 266364 222896 266416
rect 224224 266364 224276 266416
rect 239496 266364 239548 266416
rect 244096 266364 244148 266416
rect 253756 266364 253808 266416
rect 256516 266364 256568 266416
rect 256700 266364 256752 266416
rect 259828 266364 259880 266416
rect 269764 266364 269816 266416
rect 272248 266364 272300 266416
rect 272892 266364 272944 266416
rect 277216 266364 277268 266416
rect 277400 266364 277452 266416
rect 282184 266364 282236 266416
rect 293960 266364 294012 266416
rect 296260 266364 296312 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 320272 266364 320324 266416
rect 324964 266364 325016 266416
rect 332692 266364 332744 266416
rect 333796 266364 333848 266416
rect 342628 266364 342680 266416
rect 343548 266364 343600 266416
rect 345112 266364 345164 266416
rect 349896 266364 349948 266416
rect 355048 266364 355100 266416
rect 356704 266364 356756 266416
rect 361672 266364 361724 266416
rect 362868 266364 362920 266416
rect 367468 266364 367520 266416
rect 368296 266364 368348 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 379888 266364 379940 266416
rect 380808 266364 380860 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387524 266364 387576 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 405004 266500 405056 266552
rect 441988 266500 442040 266552
rect 445024 266500 445076 266552
rect 421288 266432 421340 266484
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 419816 266364 419868 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 439320 266364 439372 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 446128 266364 446180 266416
rect 447784 266364 447836 266416
rect 456892 266364 456944 266416
rect 457996 266364 458048 266416
rect 466828 266364 466880 266416
rect 467748 266364 467800 266416
rect 469312 266364 469364 266416
rect 470416 266364 470468 266416
rect 469956 266228 470008 266280
rect 483204 266432 483256 266484
rect 483388 266432 483440 266484
rect 484308 266432 484360 266484
rect 485872 266432 485924 266484
rect 486976 266432 487028 266484
rect 490012 266432 490064 266484
rect 495164 266568 495216 266620
rect 494152 266432 494204 266484
rect 495348 266432 495400 266484
rect 497464 266568 497516 266620
rect 552664 266568 552716 266620
rect 514024 266432 514076 266484
rect 514852 266432 514904 266484
rect 516048 266432 516100 266484
rect 516508 266432 516560 266484
rect 517336 266432 517388 266484
rect 518992 266432 519044 266484
rect 520096 266432 520148 266484
rect 524788 266432 524840 266484
rect 525708 266432 525760 266484
rect 527272 266432 527324 266484
rect 592684 266432 592736 266484
rect 480076 266296 480128 266348
rect 554780 266296 554832 266348
rect 485044 266160 485096 266212
rect 561680 266160 561732 266212
rect 486700 266024 486752 266076
rect 564440 266024 564492 266076
rect 492496 265888 492548 265940
rect 572720 265888 572772 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 142160 265616 142212 265668
rect 142804 265616 142856 265668
rect 191840 265616 191892 265668
rect 192484 265616 192536 265668
rect 234620 265616 234672 265668
rect 235540 265616 235592 265668
rect 518164 265616 518216 265668
rect 608692 265616 608744 265668
rect 481732 265480 481784 265532
rect 557540 265480 557592 265532
rect 479248 265344 479300 265396
rect 553400 265344 553452 265396
rect 571984 261468 572036 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 563704 259428 563756 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 560944 256708 560996 256760
rect 553768 255280 553820 255332
rect 556804 255280 556856 255332
rect 35808 252832 35860 252884
rect 41328 252832 41380 252884
rect 35624 252696 35676 252748
rect 41696 252696 41748 252748
rect 35808 252560 35860 252612
rect 40684 252560 40736 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 676036 252356 676088 252408
rect 679624 252356 679676 252408
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 35808 251200 35860 251252
rect 37924 251200 37976 251252
rect 553492 251200 553544 251252
rect 555424 251200 555476 251252
rect 558184 246304 558236 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 606484 245624 606536 245676
rect 554504 244536 554556 244588
rect 559564 244536 559616 244588
rect 37924 242836 37976 242888
rect 41696 242836 41748 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 628564 241476 628616 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 671712 237804 671764 237856
rect 671896 237600 671948 237652
rect 672080 237396 672132 237448
rect 673092 237464 673144 237516
rect 671528 237260 671580 237312
rect 672724 237124 672776 237176
rect 668952 236852 669004 236904
rect 673528 236852 673580 236904
rect 673644 236444 673696 236496
rect 673752 236308 673804 236360
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 671344 236036 671396 236088
rect 668676 235900 668728 235952
rect 672080 235900 672132 235952
rect 671160 235764 671212 235816
rect 672744 235220 672796 235272
rect 674196 235424 674248 235476
rect 674426 235084 674478 235136
rect 554412 234540 554464 234592
rect 571984 234540 572036 234592
rect 668308 234540 668360 234592
rect 674288 234608 674340 234660
rect 669780 234336 669832 234388
rect 674380 234200 674432 234252
rect 675852 234472 675904 234524
rect 679808 234472 679860 234524
rect 674886 234268 674938 234320
rect 672380 233996 672432 234048
rect 674536 234064 674588 234116
rect 675852 234064 675904 234116
rect 679624 234064 679676 234116
rect 674978 233860 675030 233912
rect 675852 233792 675904 233844
rect 677876 233792 677928 233844
rect 675116 233724 675168 233776
rect 674536 233588 674588 233640
rect 672908 233452 672960 233504
rect 675208 233384 675260 233436
rect 670976 233316 671028 233368
rect 675852 233248 675904 233300
rect 683396 233248 683448 233300
rect 671712 233180 671764 233232
rect 673000 233180 673052 233232
rect 671160 232976 671212 233028
rect 674840 232976 674892 233028
rect 670240 232840 670292 232892
rect 674196 232840 674248 232892
rect 661868 232568 661920 232620
rect 675484 232568 675536 232620
rect 675852 232500 675904 232552
rect 683672 232500 683724 232552
rect 664996 232160 665048 232212
rect 673828 231956 673880 232008
rect 674840 231752 674892 231804
rect 675070 231480 675122 231532
rect 675852 231480 675904 231532
rect 677600 231480 677652 231532
rect 668124 231412 668176 231464
rect 674518 231412 674570 231464
rect 674956 231276 675008 231328
rect 674656 231140 674708 231192
rect 662328 231072 662380 231124
rect 673828 231072 673880 231124
rect 675852 231072 675904 231124
rect 678428 231072 678480 231124
rect 674732 231004 674784 231056
rect 124128 230732 124180 230784
rect 194600 230732 194652 230784
rect 97908 230596 97960 230648
rect 173992 230596 174044 230648
rect 439320 230528 439372 230580
rect 91008 230460 91060 230512
rect 168840 230460 168892 230512
rect 184112 230392 184164 230444
rect 189448 230392 189500 230444
rect 196072 230392 196124 230444
rect 198464 230392 198516 230444
rect 207664 230392 207716 230444
rect 251272 230392 251324 230444
rect 256608 230392 256660 230444
rect 297640 230392 297692 230444
rect 323584 230392 323636 230444
rect 324688 230392 324740 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443552 230392 443604 230444
rect 444472 230392 444524 230444
rect 447600 230392 447652 230444
rect 468300 230392 468352 230444
rect 469036 230392 469088 230444
rect 472164 230392 472216 230444
rect 473084 230392 473136 230444
rect 376024 230324 376076 230376
rect 380716 230324 380768 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 473452 230324 473504 230376
rect 474556 230324 474608 230376
rect 477316 230324 477368 230376
rect 480076 230324 480128 230376
rect 480536 230324 480588 230376
rect 481548 230324 481600 230376
rect 499856 230324 499908 230376
rect 501604 230324 501656 230376
rect 501788 230324 501840 230376
rect 508504 230324 508556 230376
rect 509516 230324 509568 230376
rect 518164 230324 518216 230376
rect 520464 230324 520516 230376
rect 521476 230324 521528 230376
rect 530124 230324 530176 230376
rect 531228 230324 531280 230376
rect 133788 230256 133840 230308
rect 202328 230256 202380 230308
rect 126888 230120 126940 230172
rect 197176 230120 197228 230172
rect 197452 230120 197504 230172
rect 201040 230120 201092 230172
rect 202144 230120 202196 230172
rect 240968 230256 241020 230308
rect 242532 230256 242584 230308
rect 287336 230256 287388 230308
rect 305644 230256 305696 230308
rect 334992 230256 335044 230308
rect 387340 230188 387392 230240
rect 388444 230188 388496 230240
rect 413836 230188 413888 230240
rect 420000 230188 420052 230240
rect 443828 230188 443880 230240
rect 444656 230188 444708 230240
rect 470876 230188 470928 230240
rect 471888 230188 471940 230240
rect 474096 230188 474148 230240
rect 477408 230188 477460 230240
rect 530768 230188 530820 230240
rect 543004 230392 543056 230444
rect 668860 230392 668912 230444
rect 674380 230936 674432 230988
rect 673644 230800 673696 230852
rect 533528 230256 533580 230308
rect 541256 230256 541308 230308
rect 674380 230596 674432 230648
rect 674518 230460 674570 230512
rect 674396 230256 674448 230308
rect 214380 230120 214432 230172
rect 225512 230120 225564 230172
rect 230480 230120 230532 230172
rect 277032 230120 277084 230172
rect 294604 230120 294656 230172
rect 323400 230120 323452 230172
rect 324964 230120 325016 230172
rect 350448 230120 350500 230172
rect 354864 230120 354916 230172
rect 371056 230120 371108 230172
rect 503720 230120 503772 230172
rect 512644 230120 512696 230172
rect 515312 230120 515364 230172
rect 525156 230120 525208 230172
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 486332 230052 486384 230104
rect 487068 230052 487120 230104
rect 490196 230052 490248 230104
rect 86224 229984 86276 230036
rect 155960 229984 156012 230036
rect 157064 229984 157116 230036
rect 117228 229848 117280 229900
rect 184112 229848 184164 229900
rect 184480 229848 184532 229900
rect 214380 229848 214432 229900
rect 225788 229984 225840 230036
rect 271880 229984 271932 230036
rect 300124 229984 300176 230036
rect 329840 229984 329892 230036
rect 337844 229984 337896 230036
rect 360752 229984 360804 230036
rect 465448 229984 465500 230036
rect 473728 229984 473780 230036
rect 484400 229916 484452 229968
rect 496820 229916 496872 229968
rect 220360 229848 220412 229900
rect 224040 229848 224092 229900
rect 266728 229848 266780 229900
rect 283564 229848 283616 229900
rect 318248 229848 318300 229900
rect 318432 229848 318484 229900
rect 345296 229848 345348 229900
rect 361212 229848 361264 229900
rect 378784 229848 378836 229900
rect 389916 229848 389968 229900
rect 399392 229848 399444 229900
rect 410800 229848 410852 229900
rect 417424 229848 417476 229900
rect 505652 229984 505704 230036
rect 505744 229848 505796 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 528836 229984 528888 230036
rect 533528 229984 533580 230036
rect 534632 229984 534684 230036
rect 552204 229984 552256 230036
rect 556804 229984 556856 230036
rect 571340 229984 571392 230036
rect 675852 229984 675904 230036
rect 677416 229984 677468 230036
rect 510804 229916 510856 229968
rect 511816 229916 511868 229968
rect 673920 229916 673972 229968
rect 674172 229916 674224 229968
rect 519176 229848 519228 229900
rect 529204 229848 529256 229900
rect 536564 229848 536616 229900
rect 556988 229848 557040 229900
rect 515404 229780 515456 229832
rect 675852 229848 675904 229900
rect 676772 229848 676824 229900
rect 110328 229712 110380 229764
rect 184296 229712 184348 229764
rect 185584 229712 185636 229764
rect 207480 229712 207532 229764
rect 210424 229712 210476 229764
rect 261576 229712 261628 229764
rect 270132 229712 270184 229764
rect 307944 229712 307996 229764
rect 95240 229576 95292 229628
rect 161112 229576 161164 229628
rect 161296 229576 161348 229628
rect 175096 229576 175148 229628
rect 175280 229576 175332 229628
rect 217784 229576 217836 229628
rect 251732 229576 251784 229628
rect 292488 229576 292540 229628
rect 311900 229576 311952 229628
rect 340144 229712 340196 229764
rect 345664 229712 345716 229764
rect 355600 229712 355652 229764
rect 357072 229712 357124 229764
rect 376208 229712 376260 229764
rect 380716 229712 380768 229764
rect 394240 229712 394292 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 479248 229712 479300 229764
rect 489920 229712 489972 229764
rect 494336 229712 494388 229764
rect 509884 229712 509936 229764
rect 523040 229712 523092 229764
rect 534908 229712 534960 229764
rect 538496 229712 538548 229764
rect 565636 229712 565688 229764
rect 526904 229576 526956 229628
rect 534724 229576 534776 229628
rect 448980 229508 449032 229560
rect 452200 229508 452252 229560
rect 673948 229508 674000 229560
rect 94504 229440 94556 229492
rect 145656 229440 145708 229492
rect 146208 229440 146260 229492
rect 210056 229440 210108 229492
rect 137284 229304 137336 229356
rect 143724 229304 143776 229356
rect 144184 229304 144236 229356
rect 148876 229304 148928 229356
rect 150072 229304 150124 229356
rect 215208 229440 215260 229492
rect 217324 229440 217376 229492
rect 224040 229440 224092 229492
rect 213092 229304 213144 229356
rect 256424 229440 256476 229492
rect 276664 229440 276716 229492
rect 302792 229440 302844 229492
rect 673828 229440 673880 229492
rect 450912 229372 450964 229424
rect 453028 229372 453080 229424
rect 453488 229372 453540 229424
rect 455788 229372 455840 229424
rect 261484 229304 261536 229356
rect 282184 229304 282236 229356
rect 288716 229304 288768 229356
rect 313096 229304 313148 229356
rect 517428 229304 517480 229356
rect 520280 229304 520332 229356
rect 448336 229236 448388 229288
rect 449808 229236 449860 229288
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 452844 229236 452896 229288
rect 454684 229236 454736 229288
rect 497924 229236 497976 229288
rect 500224 229236 500276 229288
rect 521108 229236 521160 229288
rect 526444 229236 526496 229288
rect 106924 229168 106976 229220
rect 166264 229168 166316 229220
rect 167644 229168 167696 229220
rect 174912 229168 174964 229220
rect 175096 229168 175148 229220
rect 185584 229168 185636 229220
rect 189724 229168 189776 229220
rect 235816 229168 235868 229220
rect 513380 229168 513432 229220
rect 519544 229168 519596 229220
rect 419632 229100 419684 229152
rect 421932 229100 421984 229152
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 446404 229100 446456 229152
rect 448520 229100 448572 229152
rect 449624 229100 449676 229152
rect 450728 229100 450780 229152
rect 451556 229100 451608 229152
rect 453304 229100 453356 229152
rect 454132 229100 454184 229152
rect 455328 229100 455380 229152
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 119988 229032 120040 229084
rect 190092 229032 190144 229084
rect 193128 229032 193180 229084
rect 246764 229032 246816 229084
rect 257712 229032 257764 229084
rect 299572 229032 299624 229084
rect 308772 229032 308824 229084
rect 336280 229032 336332 229084
rect 508228 228964 508280 229016
rect 523316 229032 523368 229084
rect 100668 228896 100720 228948
rect 174636 228896 174688 228948
rect 176384 228896 176436 228948
rect 233884 228896 233936 228948
rect 234528 228896 234580 228948
rect 278320 228896 278372 228948
rect 288072 228896 288124 228948
rect 322756 228896 322808 228948
rect 327724 228896 327776 228948
rect 337568 228896 337620 228948
rect 350172 228896 350224 228948
rect 369124 228896 369176 228948
rect 517888 228896 517940 228948
rect 540796 228896 540848 228948
rect 106188 228760 106240 228812
rect 179788 228760 179840 228812
rect 183468 228760 183520 228812
rect 239036 228760 239088 228812
rect 246304 228760 246356 228812
rect 289268 228760 289320 228812
rect 304908 228760 304960 228812
rect 333704 228760 333756 228812
rect 335268 228760 335320 228812
rect 356888 228760 356940 228812
rect 373816 228760 373868 228812
rect 387156 228760 387208 228812
rect 485044 228760 485096 228812
rect 498752 228760 498804 228812
rect 526260 228760 526312 228812
rect 550640 228760 550692 228812
rect 93768 228624 93820 228676
rect 169484 228624 169536 228676
rect 169944 228624 169996 228676
rect 228732 228624 228784 228676
rect 235816 228624 235868 228676
rect 280252 228624 280304 228676
rect 285588 228624 285640 228676
rect 318892 228624 318944 228676
rect 336556 228624 336608 228676
rect 358820 228624 358872 228676
rect 371056 228624 371108 228676
rect 385224 228624 385276 228676
rect 404176 228624 404228 228676
rect 410984 228624 411036 228676
rect 486884 228624 486936 228676
rect 500960 228624 501012 228676
rect 506296 228624 506348 228676
rect 526628 228624 526680 228676
rect 531412 228624 531464 228676
rect 558276 228624 558328 228676
rect 64144 228488 64196 228540
rect 143080 228488 143132 228540
rect 153108 228488 153160 228540
rect 215852 228488 215904 228540
rect 222016 228488 222068 228540
rect 269948 228488 270000 228540
rect 274088 228488 274140 228540
rect 309232 228488 309284 228540
rect 326896 228488 326948 228540
rect 351092 228488 351144 228540
rect 360108 228488 360160 228540
rect 376852 228488 376904 228540
rect 377772 228488 377824 228540
rect 390376 228488 390428 228540
rect 400220 228488 400272 228540
rect 407764 228488 407816 228540
rect 410984 228488 411036 228540
rect 416136 228488 416188 228540
rect 480076 228488 480128 228540
rect 489184 228488 489236 228540
rect 495348 228488 495400 228540
rect 510620 228488 510672 228540
rect 511448 228488 511500 228540
rect 531964 228488 532016 228540
rect 537852 228488 537904 228540
rect 566096 228488 566148 228540
rect 57244 228352 57296 228404
rect 141148 228352 141200 228404
rect 145932 228352 145984 228404
rect 210700 228352 210752 228404
rect 215208 228352 215260 228404
rect 266084 228352 266136 228404
rect 271788 228352 271840 228404
rect 308588 228352 308640 228404
rect 313004 228352 313056 228404
rect 340788 228352 340840 228404
rect 126704 228216 126756 228268
rect 195244 228216 195296 228268
rect 205364 228216 205416 228268
rect 257068 228216 257120 228268
rect 265624 228216 265676 228268
rect 274456 228216 274508 228268
rect 309692 228216 309744 228268
rect 327264 228216 327316 228268
rect 340144 228216 340196 228268
rect 362684 228352 362736 228404
rect 362868 228352 362920 228404
rect 379428 228352 379480 228404
rect 379244 228216 379296 228268
rect 393596 228352 393648 228404
rect 409788 228352 409840 228404
rect 415492 228352 415544 228404
rect 470232 228352 470284 228404
rect 479708 228352 479760 228404
rect 481824 228352 481876 228404
rect 494704 228352 494756 228404
rect 497280 228352 497332 228404
rect 514300 228352 514352 228404
rect 521752 228352 521804 228404
rect 545764 228352 545816 228404
rect 554044 228352 554096 228404
rect 632704 228352 632756 228404
rect 673460 229100 673512 229152
rect 673736 229100 673788 229152
rect 672816 228964 672868 229016
rect 673598 228896 673650 228948
rect 673506 228692 673558 228744
rect 672816 228488 672868 228540
rect 672816 228352 672868 228404
rect 390100 228216 390152 228268
rect 400036 228216 400088 228268
rect 133512 228080 133564 228132
rect 200396 228080 200448 228132
rect 211068 228080 211120 228132
rect 260288 228080 260340 228132
rect 398656 228080 398708 228132
rect 409052 228216 409104 228268
rect 523316 228216 523368 228268
rect 527732 228216 527784 228268
rect 669412 228216 669464 228268
rect 672356 228012 672408 228064
rect 139308 227944 139360 227996
rect 205548 227944 205600 227996
rect 252376 227944 252428 227996
rect 293132 227944 293184 227996
rect 393964 227876 394016 227928
rect 401324 227876 401376 227928
rect 402244 227876 402296 227928
rect 143448 227808 143500 227860
rect 146208 227808 146260 227860
rect 169576 227808 169628 227860
rect 169944 227808 169996 227860
rect 196716 227808 196768 227860
rect 230664 227808 230716 227860
rect 280712 227808 280764 227860
rect 284760 227808 284812 227860
rect 297364 227808 297416 227860
rect 305368 227808 305420 227860
rect 396632 227740 396684 227792
rect 397460 227740 397512 227792
rect 400772 227740 400824 227792
rect 402612 227740 402664 227792
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 672816 227808 672868 227860
rect 403256 227740 403308 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416688 227740 416740 227792
rect 420644 227740 420696 227792
rect 474740 227740 474792 227792
rect 482928 227740 482980 227792
rect 659476 227740 659528 227792
rect 665180 227740 665232 227792
rect 116952 227672 117004 227724
rect 187516 227672 187568 227724
rect 200028 227672 200080 227724
rect 251916 227672 251968 227724
rect 263416 227672 263468 227724
rect 301504 227672 301556 227724
rect 110144 227536 110196 227588
rect 182364 227536 182416 227588
rect 182824 227536 182876 227588
rect 236460 227536 236512 227588
rect 241980 227536 242032 227588
rect 285404 227536 285456 227588
rect 293776 227536 293828 227588
rect 325332 227536 325384 227588
rect 515404 227536 515456 227588
rect 524972 227536 525024 227588
rect 526444 227536 526496 227588
rect 544384 227536 544436 227588
rect 560944 227536 560996 227588
rect 568120 227536 568172 227588
rect 672816 227468 672868 227520
rect 103428 227400 103480 227452
rect 177212 227400 177264 227452
rect 81348 227264 81400 227316
rect 95240 227264 95292 227316
rect 96252 227264 96304 227316
rect 172060 227264 172112 227316
rect 173164 227264 173216 227316
rect 185584 227400 185636 227452
rect 188988 227400 189040 227452
rect 244188 227400 244240 227452
rect 251088 227400 251140 227452
rect 294420 227400 294472 227452
rect 302148 227400 302200 227452
rect 331128 227400 331180 227452
rect 333888 227400 333940 227452
rect 356244 227400 356296 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 184940 227264 184992 227316
rect 192668 227264 192720 227316
rect 198648 227264 198700 227316
rect 253204 227264 253256 227316
rect 259368 227264 259420 227316
rect 298284 227264 298336 227316
rect 308956 227264 309008 227316
rect 339500 227264 339552 227316
rect 351092 227264 351144 227316
rect 363328 227264 363380 227316
rect 363512 227264 363564 227316
rect 368480 227264 368532 227316
rect 385684 227264 385736 227316
rect 391664 227264 391716 227316
rect 477408 227264 477460 227316
rect 485044 227264 485096 227316
rect 490840 227264 490892 227316
rect 505468 227264 505520 227316
rect 506940 227264 506992 227316
rect 526352 227264 526404 227316
rect 528192 227264 528244 227316
rect 554044 227264 554096 227316
rect 68284 227128 68336 227180
rect 146392 227128 146444 227180
rect 152924 227128 152976 227180
rect 213368 227128 213420 227180
rect 224776 227128 224828 227180
rect 273812 227128 273864 227180
rect 274272 227128 274324 227180
rect 312452 227128 312504 227180
rect 319812 227128 319864 227180
rect 345848 227128 345900 227180
rect 346124 227128 346176 227180
rect 366548 227128 366600 227180
rect 369492 227128 369544 227180
rect 384580 227128 384632 227180
rect 391572 227128 391624 227180
rect 400588 227128 400640 227180
rect 401508 227128 401560 227180
rect 408408 227128 408460 227180
rect 483756 227128 483808 227180
rect 497556 227128 497608 227180
rect 498568 227128 498620 227180
rect 515772 227128 515824 227180
rect 525616 227128 525668 227180
rect 550824 227128 550876 227180
rect 671896 227196 671948 227248
rect 56508 226992 56560 227044
rect 142436 226992 142488 227044
rect 143264 226992 143316 227044
rect 208124 226992 208176 227044
rect 122748 226856 122800 226908
rect 184940 226856 184992 226908
rect 185584 226856 185636 226908
rect 226156 226992 226208 227044
rect 228732 226992 228784 227044
rect 275100 226992 275152 227044
rect 284852 226992 284904 227044
rect 320180 226992 320232 227044
rect 325516 226992 325568 227044
rect 349160 226992 349212 227044
rect 357256 226992 357308 227044
rect 374276 226992 374328 227044
rect 376668 226992 376720 227044
rect 389732 226992 389784 227044
rect 395804 226992 395856 227044
rect 406476 226992 406528 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 491484 226992 491536 227044
rect 506848 226992 506900 227044
rect 512092 226992 512144 227044
rect 533436 226992 533488 227044
rect 535276 226992 535328 227044
rect 562784 226992 562836 227044
rect 471520 226924 471572 226976
rect 479524 226924 479576 226976
rect 671344 226924 671396 226976
rect 671712 226924 671764 226976
rect 212172 226856 212224 226908
rect 262220 226856 262272 226908
rect 275652 226856 275704 226908
rect 311164 226856 311216 226908
rect 384948 226856 385000 226908
rect 395528 226856 395580 226908
rect 419448 226856 419500 226908
rect 424508 226856 424560 226908
rect 479892 226856 479944 226908
rect 491944 226856 491996 226908
rect 671712 226788 671764 226840
rect 672080 226788 672132 226840
rect 129372 226720 129424 226772
rect 197820 226720 197872 226772
rect 224592 226720 224644 226772
rect 270592 226720 270644 226772
rect 672380 226652 672432 226704
rect 150256 226584 150308 226636
rect 152924 226584 152976 226636
rect 160008 226584 160060 226636
rect 221004 226584 221056 226636
rect 671942 226584 671994 226636
rect 177212 226448 177264 226500
rect 231308 226448 231360 226500
rect 465908 226448 465960 226500
rect 469864 226448 469916 226500
rect 671820 226448 671872 226500
rect 407764 226312 407816 226364
rect 411628 226312 411680 226364
rect 135168 226244 135220 226296
rect 204260 226244 204312 226296
rect 205548 226244 205600 226296
rect 99288 226108 99340 226160
rect 175924 226108 175976 226160
rect 202696 226108 202748 226160
rect 206744 226108 206796 226160
rect 219348 226244 219400 226296
rect 267372 226244 267424 226296
rect 303252 226244 303304 226296
rect 333060 226244 333112 226296
rect 258356 226108 258408 226160
rect 286692 226108 286744 226160
rect 319536 226108 319588 226160
rect 350356 226108 350408 226160
rect 354864 226108 354916 226160
rect 501144 226108 501196 226160
rect 519268 226108 519320 226160
rect 529940 226108 529992 226160
rect 549904 226108 549956 226160
rect 672034 226108 672086 226160
rect 84108 225972 84160 226024
rect 161756 225972 161808 226024
rect 186044 225972 186096 226024
rect 241612 225972 241664 226024
rect 245292 225972 245344 226024
rect 287612 225972 287664 226024
rect 296628 225972 296680 226024
rect 329196 225972 329248 226024
rect 330392 225972 330444 226024
rect 351920 225972 351972 226024
rect 352564 225972 352616 226024
rect 358176 225972 358228 226024
rect 515956 225972 516008 226024
rect 538956 225972 539008 226024
rect 671942 225904 671994 225956
rect 70308 225836 70360 225888
rect 151452 225836 151504 225888
rect 158352 225836 158404 225888
rect 222292 225836 222344 225888
rect 239404 225836 239456 225888
rect 284116 225836 284168 225888
rect 288256 225836 288308 225888
rect 321468 225836 321520 225888
rect 324228 225836 324280 225888
rect 348516 225836 348568 225888
rect 355324 225836 355376 225888
rect 372344 225836 372396 225888
rect 495992 225836 496044 225888
rect 512460 225836 512512 225888
rect 524328 225836 524380 225888
rect 547880 225836 547932 225888
rect 555424 225836 555476 225888
rect 570788 225836 570840 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 60004 225700 60056 225752
rect 141792 225700 141844 225752
rect 141976 225700 142028 225752
rect 209412 225700 209464 225752
rect 209596 225700 209648 225752
rect 259644 225700 259696 225752
rect 264888 225700 264940 225752
rect 304724 225700 304776 225752
rect 319996 225700 320048 225752
rect 347228 225700 347280 225752
rect 349068 225700 349120 225752
rect 367192 225700 367244 225752
rect 375288 225700 375340 225752
rect 387800 225700 387852 225752
rect 388444 225700 388496 225752
rect 396448 225700 396500 225752
rect 476028 225700 476080 225752
rect 483572 225700 483624 225752
rect 489552 225700 489604 225752
rect 504180 225700 504232 225752
rect 510160 225700 510212 225752
rect 530860 225700 530912 225752
rect 533988 225700 534040 225752
rect 561496 225700 561548 225752
rect 671820 225700 671872 225752
rect 667940 225632 667992 225684
rect 62028 225564 62080 225616
rect 144368 225564 144420 225616
rect 155868 225564 155920 225616
rect 219716 225564 219768 225616
rect 220452 225564 220504 225616
rect 268016 225564 268068 225616
rect 269028 225564 269080 225616
rect 306012 225564 306064 225616
rect 306196 225564 306248 225616
rect 336924 225564 336976 225616
rect 340696 225564 340748 225616
rect 361488 225564 361540 225616
rect 365536 225564 365588 225616
rect 379796 225564 379848 225616
rect 380072 225564 380124 225616
rect 391020 225564 391072 225616
rect 391756 225564 391808 225616
rect 403532 225564 403584 225616
rect 467656 225564 467708 225616
rect 477040 225564 477092 225616
rect 481180 225564 481232 225616
rect 493692 225564 493744 225616
rect 508872 225564 508924 225616
rect 529204 225564 529256 225616
rect 529480 225564 529532 225616
rect 555884 225564 555936 225616
rect 132408 225428 132460 225480
rect 201684 225428 201736 225480
rect 206192 225428 206244 225480
rect 139124 225292 139176 225344
rect 206376 225292 206428 225344
rect 206744 225428 206796 225480
rect 254492 225428 254544 225480
rect 255228 225428 255280 225480
rect 296996 225428 297048 225480
rect 492772 225428 492824 225480
rect 508688 225428 508740 225480
rect 228088 225292 228140 225344
rect 255044 225292 255096 225344
rect 295708 225292 295760 225344
rect 671596 225292 671648 225344
rect 155684 225156 155736 225208
rect 218428 225156 218480 225208
rect 225604 225156 225656 225208
rect 246120 225156 246172 225208
rect 671482 225088 671534 225140
rect 166264 225020 166316 225072
rect 186872 225020 186924 225072
rect 195612 225020 195664 225072
rect 249340 225020 249392 225072
rect 404360 225020 404412 225072
rect 412272 225020 412324 225072
rect 463148 225020 463200 225072
rect 467472 225020 467524 225072
rect 669412 225020 669464 225072
rect 260012 224952 260064 225004
rect 264152 224952 264204 225004
rect 367652 224952 367704 225004
rect 373632 224952 373684 225004
rect 118608 224884 118660 224936
rect 185584 224884 185636 224936
rect 191472 224884 191524 224936
rect 248052 224884 248104 224936
rect 266268 224884 266320 224936
rect 303436 224884 303488 224936
rect 321468 224884 321520 224936
rect 346584 224884 346636 224936
rect 426440 224884 426492 224936
rect 426992 224884 427044 224936
rect 460572 224884 460624 224936
rect 463148 224884 463200 224936
rect 669412 224816 669464 224868
rect 112812 224748 112864 224800
rect 185860 224748 185912 224800
rect 106004 224612 106056 224664
rect 181076 224612 181128 224664
rect 181996 224612 182048 224664
rect 185216 224612 185268 224664
rect 185400 224612 185452 224664
rect 242900 224748 242952 224800
rect 271604 224748 271656 224800
rect 309876 224748 309928 224800
rect 313188 224748 313240 224800
rect 342076 224748 342128 224800
rect 186228 224612 186280 224664
rect 240324 224612 240376 224664
rect 249616 224612 249668 224664
rect 290556 224612 290608 224664
rect 294972 224612 295024 224664
rect 325976 224612 326028 224664
rect 347044 224612 347096 224664
rect 365904 224748 365956 224800
rect 670976 224680 671028 224732
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 172336 224476 172388 224528
rect 232596 224476 232648 224528
rect 233148 224476 233200 224528
rect 277676 224476 277728 224528
rect 282460 224476 282512 224528
rect 316316 224476 316368 224528
rect 317144 224476 317196 224528
rect 342996 224476 343048 224528
rect 343456 224476 343508 224528
rect 363972 224612 364024 224664
rect 499212 224612 499264 224664
rect 516784 224612 516836 224664
rect 518532 224612 518584 224664
rect 541624 224612 541676 224664
rect 363788 224476 363840 224528
rect 378140 224476 378192 224528
rect 387708 224476 387760 224528
rect 398104 224476 398156 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 505008 224476 505060 224528
rect 523040 224476 523092 224528
rect 523684 224476 523736 224528
rect 548340 224476 548392 224528
rect 666836 224408 666888 224460
rect 76564 224340 76616 224392
rect 157892 224340 157944 224392
rect 165528 224340 165580 224392
rect 227444 224340 227496 224392
rect 241152 224340 241204 224392
rect 286508 224340 286560 224392
rect 291016 224340 291068 224392
rect 324044 224340 324096 224392
rect 341984 224340 342036 224392
rect 365260 224340 365312 224392
rect 368388 224340 368440 224392
rect 382556 224340 382608 224392
rect 382924 224340 382976 224392
rect 396172 224340 396224 224392
rect 436376 224340 436428 224392
rect 436836 224340 436888 224392
rect 462504 224340 462556 224392
rect 469312 224340 469364 224392
rect 478604 224340 478656 224392
rect 490288 224340 490340 224392
rect 492128 224340 492180 224392
rect 507768 224340 507820 224392
rect 514668 224340 514720 224392
rect 535644 224340 535696 224392
rect 536012 224340 536064 224392
rect 563980 224340 564032 224392
rect 565636 224272 565688 224324
rect 568580 224272 568632 224324
rect 63408 224204 63460 224256
rect 147588 224204 147640 224256
rect 151728 224204 151780 224256
rect 217140 224204 217192 224256
rect 223488 224204 223540 224256
rect 225788 224204 225840 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 281448 224204 281500 224256
rect 317604 224204 317656 224256
rect 322296 224204 322348 224256
rect 349804 224204 349856 224256
rect 351736 224204 351788 224256
rect 369768 224204 369820 224256
rect 372436 224204 372488 224256
rect 387340 224204 387392 224256
rect 394516 224204 394568 224256
rect 404544 224204 404596 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 420828 224204 420880 224256
rect 425152 224204 425204 224256
rect 436284 224204 436336 224256
rect 437020 224204 437072 224256
rect 469588 224204 469640 224256
rect 477592 224204 477644 224256
rect 488908 224204 488960 224256
rect 502984 224204 503036 224256
rect 504364 224204 504416 224256
rect 523500 224204 523552 224256
rect 533712 224204 533764 224256
rect 561312 224204 561364 224256
rect 563704 224136 563756 224188
rect 568948 224136 569000 224188
rect 606300 224136 606352 224188
rect 115848 224068 115900 224120
rect 188804 224068 188856 224120
rect 189908 224068 189960 224120
rect 212632 224068 212684 224120
rect 216588 224068 216640 224120
rect 264428 224068 264480 224120
rect 275836 224068 275888 224120
rect 288716 224068 288768 224120
rect 415032 224000 415084 224052
rect 419632 224000 419684 224052
rect 489920 224000 489972 224052
rect 491116 224000 491168 224052
rect 535644 224000 535696 224052
rect 536656 224000 536708 224052
rect 567844 224000 567896 224052
rect 670930 224136 670982 224188
rect 122564 223932 122616 223984
rect 193956 223932 194008 223984
rect 200764 223932 200816 223984
rect 222936 223932 222988 223984
rect 226156 223932 226208 223984
rect 272524 223932 272576 223984
rect 289084 223864 289136 223916
rect 294788 223864 294840 223916
rect 512460 223864 512512 223916
rect 606300 223864 606352 223916
rect 616880 224000 616932 224052
rect 630956 223864 631008 223916
rect 139952 223796 140004 223848
rect 171416 223796 171468 223848
rect 174912 223796 174964 223848
rect 235172 223796 235224 223848
rect 496820 223728 496872 223780
rect 497372 223728 497424 223780
rect 567844 223728 567896 223780
rect 568580 223728 568632 223780
rect 627920 223728 627972 223780
rect 185584 223660 185636 223712
rect 191012 223660 191064 223712
rect 227628 223660 227680 223712
rect 273168 223660 273220 223712
rect 491116 223592 491168 223644
rect 629852 223592 629904 223644
rect 654968 223592 655020 223644
rect 655612 223592 655664 223644
rect 87972 223524 88024 223576
rect 164976 223524 165028 223576
rect 166448 223524 166500 223576
rect 192024 223524 192076 223576
rect 194508 223524 194560 223576
rect 247408 223524 247460 223576
rect 253572 223524 253624 223576
rect 293500 223524 293552 223576
rect 307024 223524 307076 223576
rect 315672 223524 315724 223576
rect 416504 223524 416556 223576
rect 422208 223524 422260 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 102048 223388 102100 223440
rect 178500 223388 178552 223440
rect 197268 223388 197320 223440
rect 249984 223388 250036 223440
rect 267556 223388 267608 223440
rect 307300 223388 307352 223440
rect 322848 223388 322900 223440
rect 332416 223388 332468 223440
rect 520280 223388 520332 223440
rect 539968 223388 540020 223440
rect 78588 223252 78640 223304
rect 157248 223252 157300 223304
rect 159364 223252 159416 223304
rect 181720 223252 181772 223304
rect 191656 223252 191708 223304
rect 244832 223252 244884 223304
rect 261852 223252 261904 223304
rect 300860 223252 300912 223304
rect 315856 223252 315908 223304
rect 341432 223252 341484 223304
rect 342168 223252 342220 223304
rect 362040 223252 362092 223304
rect 366732 223252 366784 223304
rect 382004 223252 382056 223304
rect 406752 223252 406804 223304
rect 414848 223252 414900 223304
rect 513104 223252 513156 223304
rect 534540 223252 534592 223304
rect 541256 223252 541308 223304
rect 554872 223252 554924 223304
rect 81164 223116 81216 223168
rect 159824 223116 159876 223168
rect 168288 223116 168340 223168
rect 226800 223116 226852 223168
rect 248236 223116 248288 223168
rect 291844 223116 291896 223168
rect 300768 223116 300820 223168
rect 330116 223116 330168 223168
rect 336372 223116 336424 223168
rect 359740 223116 359792 223168
rect 366916 223116 366968 223168
rect 383936 223116 383988 223168
rect 477960 223116 478012 223168
rect 489460 223116 489512 223168
rect 496636 223116 496688 223168
rect 513564 223116 513616 223168
rect 519820 223116 519872 223168
rect 542360 223116 542412 223168
rect 552204 223116 552256 223168
rect 561680 223116 561732 223168
rect 75828 222980 75880 223032
rect 154672 222980 154724 223032
rect 164056 222980 164108 223032
rect 224224 222980 224276 223032
rect 238668 222980 238720 223032
rect 282828 222980 282880 223032
rect 292488 222980 292540 223032
rect 326620 222980 326672 223032
rect 329748 222980 329800 223032
rect 353668 222980 353720 223032
rect 355968 222980 356020 223032
rect 375564 222980 375616 223032
rect 382096 222980 382148 223032
rect 392952 222980 393004 223032
rect 483112 222980 483164 223032
rect 496084 222980 496136 223032
rect 502432 222980 502484 223032
rect 521016 222980 521068 223032
rect 527548 222980 527600 223032
rect 553308 222980 553360 223032
rect 68928 222844 68980 222896
rect 149520 222844 149572 222896
rect 154212 222844 154264 222896
rect 216220 222844 216272 222896
rect 217876 222844 217928 222896
rect 268660 222844 268712 222896
rect 278412 222844 278464 222896
rect 313740 222844 313792 222896
rect 315672 222844 315724 222896
rect 344652 222844 344704 222896
rect 346308 222844 346360 222896
rect 367468 222844 367520 222896
rect 386328 222844 386380 222896
rect 398288 222844 398340 222896
rect 398472 222844 398524 222896
rect 405832 222844 405884 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467288 222844 467340 222896
rect 475384 222844 475436 222896
rect 476672 222844 476724 222896
rect 487804 222844 487856 222896
rect 488264 222844 488316 222896
rect 503168 222844 503220 222896
rect 507584 222844 507636 222896
rect 527548 222844 527600 222896
rect 532424 222844 532476 222896
rect 559012 222844 559064 222896
rect 559564 222844 559616 222896
rect 633716 222844 633768 222896
rect 131028 222708 131080 222760
rect 196072 222708 196124 222760
rect 208032 222708 208084 222760
rect 260932 222708 260984 222760
rect 290832 222708 290884 222760
rect 321836 222708 321888 222760
rect 503352 222708 503404 222760
rect 521844 222708 521896 222760
rect 558644 222708 558696 222760
rect 568764 222708 568816 222760
rect 146116 222572 146168 222624
rect 211988 222572 212040 222624
rect 213828 222572 213880 222624
rect 262864 222572 262916 222624
rect 561680 222572 561732 222624
rect 562140 222572 562192 222624
rect 563152 222572 563204 222624
rect 565452 222572 565504 222624
rect 567108 222572 567160 222624
rect 567660 222572 567712 222624
rect 571616 222572 571668 222624
rect 134984 222436 135036 222488
rect 197452 222436 197504 222488
rect 203892 222436 203944 222488
rect 254860 222436 254912 222488
rect 482928 222436 482980 222488
rect 593972 222436 594024 222488
rect 244096 222300 244148 222352
rect 286048 222300 286100 222352
rect 556068 222300 556120 222352
rect 557356 222300 557408 222352
rect 626540 222300 626592 222352
rect 550824 222164 550876 222216
rect 111156 222096 111208 222148
rect 182548 222096 182600 222148
rect 184020 222096 184072 222148
rect 239220 222096 239272 222148
rect 282644 222096 282696 222148
rect 283564 222096 283616 222148
rect 283748 222096 283800 222148
rect 314844 222096 314896 222148
rect 386880 222096 386932 222148
rect 389916 222096 389968 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468668 222096 468720 222148
rect 563152 222164 563204 222216
rect 628196 222164 628248 222216
rect 558368 222096 558420 222148
rect 560760 222096 560812 222148
rect 561312 222096 561364 222148
rect 563014 222096 563066 222148
rect 543004 222028 543056 222080
rect 104532 221960 104584 222012
rect 177396 221960 177448 222012
rect 194784 221960 194836 222012
rect 250168 221960 250220 222012
rect 258080 221960 258132 222012
rect 269212 221960 269264 222012
rect 270040 221960 270092 222012
rect 306564 221960 306616 222012
rect 330576 221960 330628 222012
rect 345664 221960 345716 222012
rect 556068 221960 556120 222012
rect 556252 221960 556304 222012
rect 559564 221960 559616 222012
rect 562324 221960 562376 222012
rect 571432 221960 571484 222012
rect 571616 221960 571668 222012
rect 577688 221960 577740 222012
rect 596272 221960 596324 222012
rect 597008 221960 597060 222012
rect 101220 221824 101272 221876
rect 175464 221824 175516 221876
rect 189172 221824 189224 221876
rect 245016 221824 245068 221876
rect 252560 221824 252612 221876
rect 258632 221824 258684 221876
rect 266820 221824 266872 221876
rect 297180 221824 297232 221876
rect 60648 221688 60700 221740
rect 94412 221688 94464 221740
rect 94596 221688 94648 221740
rect 169760 221688 169812 221740
rect 177396 221688 177448 221740
rect 234160 221688 234212 221740
rect 247132 221688 247184 221740
rect 253388 221688 253440 221740
rect 260196 221688 260248 221740
rect 298560 221824 298612 221876
rect 306564 221824 306616 221876
rect 335452 221824 335504 221876
rect 344652 221824 344704 221876
rect 364524 221824 364576 221876
rect 512644 221824 512696 221876
rect 522580 221824 522632 221876
rect 525156 221824 525208 221876
rect 537484 221824 537536 221876
rect 547144 221824 547196 221876
rect 559840 221824 559892 221876
rect 562784 221824 562836 221876
rect 610532 221824 610584 221876
rect 298284 221688 298336 221740
rect 328552 221688 328604 221740
rect 331404 221688 331456 221740
rect 353852 221688 353904 221740
rect 362040 221688 362092 221740
rect 376024 221688 376076 221740
rect 73896 221552 73948 221604
rect 86224 221552 86276 221604
rect 91284 221552 91336 221604
rect 167092 221552 167144 221604
rect 178224 221552 178276 221604
rect 237380 221552 237432 221604
rect 238852 221552 238904 221604
rect 248604 221552 248656 221604
rect 250260 221552 250312 221604
rect 291384 221552 291436 221604
rect 84660 221416 84712 221468
rect 161480 221416 161532 221468
rect 161664 221416 161716 221468
rect 224408 221416 224460 221468
rect 234344 221416 234396 221468
rect 121092 221280 121144 221332
rect 190644 221280 190696 221332
rect 201408 221280 201460 221332
rect 255412 221280 255464 221332
rect 277584 221416 277636 221468
rect 283748 221416 283800 221468
rect 284024 221416 284076 221468
rect 289912 221416 289964 221468
rect 296444 221416 296496 221468
rect 327540 221552 327592 221604
rect 328092 221552 328144 221604
rect 351276 221552 351328 221604
rect 353300 221552 353352 221604
rect 369952 221552 370004 221604
rect 370504 221552 370556 221604
rect 382740 221688 382792 221740
rect 475752 221688 475804 221740
rect 486148 221688 486200 221740
rect 487068 221688 487120 221740
rect 500040 221688 500092 221740
rect 501604 221688 501656 221740
rect 517704 221688 517756 221740
rect 522856 221688 522908 221740
rect 546592 221688 546644 221740
rect 548340 221688 548392 221740
rect 553032 221688 553084 221740
rect 553308 221688 553360 221740
rect 608600 221688 608652 221740
rect 382740 221552 382792 221604
rect 394884 221552 394936 221604
rect 396816 221552 396868 221604
rect 407304 221552 407356 221604
rect 469036 221552 469088 221604
rect 474556 221552 474608 221604
rect 485504 221552 485556 221604
rect 499396 221552 499448 221604
rect 500224 221552 500276 221604
rect 517520 221552 517572 221604
rect 518164 221552 518216 221604
rect 530032 221552 530084 221604
rect 531228 221552 531280 221604
rect 556528 221552 556580 221604
rect 556988 221552 557040 221604
rect 564900 221552 564952 221604
rect 567660 221552 567712 221604
rect 567844 221552 567896 221604
rect 596272 221552 596324 221604
rect 596456 221552 596508 221604
rect 607312 221552 607364 221604
rect 297180 221416 297232 221468
rect 281724 221280 281776 221332
rect 292304 221280 292356 221332
rect 299940 221280 299992 221332
rect 302424 221416 302476 221468
rect 334072 221416 334124 221468
rect 334992 221416 335044 221468
rect 357532 221416 357584 221468
rect 357900 221416 357952 221468
rect 374552 221416 374604 221468
rect 375472 221416 375524 221468
rect 386512 221416 386564 221468
rect 390284 221416 390336 221468
rect 401692 221416 401744 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 473084 221416 473136 221468
rect 481180 221416 481232 221468
rect 483756 221416 483808 221468
rect 538772 221416 538824 221468
rect 540888 221416 540940 221468
rect 605472 221416 605524 221468
rect 606484 221416 606536 221468
rect 633440 221416 633492 221468
rect 303804 221280 303856 221332
rect 534908 221280 534960 221332
rect 546776 221280 546828 221332
rect 148416 221144 148468 221196
rect 214104 221144 214156 221196
rect 214288 221144 214340 221196
rect 263140 221144 263192 221196
rect 374000 221144 374052 221196
rect 381084 221144 381136 221196
rect 542360 221144 542412 221196
rect 543280 221144 543332 221196
rect 552848 221212 552900 221264
rect 558184 221212 558236 221264
rect 558368 221212 558420 221264
rect 596456 221212 596508 221264
rect 596640 221212 596692 221264
rect 607496 221212 607548 221264
rect 140964 221008 141016 221060
rect 205824 221008 205876 221060
rect 222568 221008 222620 221060
rect 270868 221008 270920 221060
rect 545764 221008 545816 221060
rect 552848 220940 552900 220992
rect 553032 220940 553084 220992
rect 596640 220940 596692 220992
rect 597008 221076 597060 221128
rect 606944 221076 606996 221128
rect 606208 220940 606260 220992
rect 172612 220872 172664 220924
rect 199476 220872 199528 220924
rect 227904 220872 227956 220924
rect 276112 220872 276164 220924
rect 420644 220804 420696 220856
rect 423864 220804 423916 220856
rect 456708 220804 456760 220856
rect 462136 220804 462188 220856
rect 558184 220804 558236 220856
rect 567844 220804 567896 220856
rect 577688 220804 577740 220856
rect 628380 220804 628432 220856
rect 107844 220736 107896 220788
rect 179972 220736 180024 220788
rect 187332 220736 187384 220788
rect 241796 220736 241848 220788
rect 261024 220736 261076 220788
rect 301688 220736 301740 220788
rect 313832 220736 313884 220788
rect 320364 220736 320416 220788
rect 339224 220736 339276 220788
rect 342444 220736 342496 220788
rect 414204 220736 414256 220788
rect 418344 220736 418396 220788
rect 465724 220736 465776 220788
rect 469588 220736 469640 220788
rect 471888 220736 471940 220788
rect 477868 220736 477920 220788
rect 552480 220736 552532 220788
rect 455328 220668 455380 220720
rect 458824 220668 458876 220720
rect 568028 220736 568080 220788
rect 577320 220736 577372 220788
rect 563060 220668 563112 220720
rect 66444 220600 66496 220652
rect 144092 220600 144144 220652
rect 144276 220600 144328 220652
rect 208584 220600 208636 220652
rect 216312 220600 216364 220652
rect 217324 220600 217376 220652
rect 217508 220600 217560 220652
rect 265072 220600 265124 220652
rect 280068 220600 280120 220652
rect 314016 220600 314068 220652
rect 318156 220600 318208 220652
rect 343824 220600 343876 220652
rect 508504 220600 508556 220652
rect 520188 220600 520240 220652
rect 521476 220600 521528 220652
rect 544108 220600 544160 220652
rect 553676 220532 553728 220584
rect 86316 220464 86368 220516
rect 164332 220464 164384 220516
rect 180708 220464 180760 220516
rect 76380 220328 76432 220380
rect 156144 220328 156196 220380
rect 170772 220328 170824 220380
rect 229100 220328 229152 220380
rect 232688 220464 232740 220516
rect 238024 220464 238076 220516
rect 240324 220464 240376 220516
rect 283104 220464 283156 220516
rect 283380 220464 283432 220516
rect 316592 220464 316644 220516
rect 328920 220464 328972 220516
rect 354680 220464 354732 220516
rect 79692 220192 79744 220244
rect 158904 220192 158956 220244
rect 161940 220192 161992 220244
rect 73068 220056 73120 220108
rect 153752 220056 153804 220108
rect 157524 220056 157576 220108
rect 218704 220056 218756 220108
rect 220820 220192 220872 220244
rect 233424 220192 233476 220244
rect 235632 220328 235684 220380
rect 243084 220328 243136 220380
rect 246948 220328 247000 220380
rect 288532 220328 288584 220380
rect 309876 220328 309928 220380
rect 338120 220328 338172 220380
rect 343640 220328 343692 220380
rect 347872 220328 347924 220380
rect 352932 220328 352984 220380
rect 371424 220328 371476 220380
rect 372252 220328 372304 220380
rect 385408 220464 385460 220516
rect 488080 220464 488132 220516
rect 501880 220464 501932 220516
rect 519544 220464 519596 220516
rect 534356 220464 534408 220516
rect 534724 220464 534776 220516
rect 552480 220464 552532 220516
rect 572076 220600 572128 220652
rect 605288 220600 605340 220652
rect 608968 220600 609020 220652
rect 563428 220464 563480 220516
rect 565452 220464 565504 220516
rect 565636 220464 565688 220516
rect 566372 220464 566424 220516
rect 566832 220464 566884 220516
rect 606484 220464 606536 220516
rect 493968 220328 494020 220380
rect 236644 220192 236696 220244
rect 237012 220192 237064 220244
rect 280436 220192 280488 220244
rect 299112 220192 299164 220244
rect 331220 220192 331272 220244
rect 338028 220192 338080 220244
rect 359004 220192 359056 220244
rect 361120 220192 361172 220244
rect 377036 220192 377088 220244
rect 378048 220192 378100 220244
rect 388628 220192 388680 220244
rect 432236 220192 432288 220244
rect 434812 220192 434864 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 468852 220192 468904 220244
rect 476212 220192 476264 220244
rect 481548 220192 481600 220244
rect 492772 220192 492824 220244
rect 495164 220192 495216 220244
rect 500408 220328 500460 220380
rect 515128 220328 515180 220380
rect 517152 220328 517204 220380
rect 539232 220328 539284 220380
rect 553124 220328 553176 220380
rect 554228 220328 554280 220380
rect 555424 220328 555476 220380
rect 566556 220328 566608 220380
rect 427912 220124 427964 220176
rect 428740 220124 428792 220176
rect 221280 220056 221332 220108
rect 230204 220056 230256 220108
rect 275284 220056 275336 220108
rect 276848 220056 276900 220108
rect 311348 220056 311400 220108
rect 311532 220056 311584 220108
rect 338396 220056 338448 220108
rect 342720 220056 342772 220108
rect 352380 220056 352432 220108
rect 354404 220056 354456 220108
rect 372804 220056 372856 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 473268 220056 473320 220108
rect 482008 220056 482060 220108
rect 482744 220056 482796 220108
rect 495256 220056 495308 220108
rect 509332 220192 509384 220244
rect 536932 220192 536984 220244
rect 558828 220192 558880 220244
rect 559380 220192 559432 220244
rect 606300 220328 606352 220380
rect 510988 220056 511040 220108
rect 511816 220056 511868 220108
rect 531688 220056 531740 220108
rect 534356 220056 534408 220108
rect 535000 220056 535052 220108
rect 114468 219920 114520 219972
rect 185032 219920 185084 219972
rect 200580 219920 200632 219972
rect 252744 219920 252796 219972
rect 256884 219920 256936 219972
rect 295984 219920 296036 219972
rect 529020 219852 529072 219904
rect 542544 219852 542596 219904
rect 556252 219920 556304 219972
rect 577320 220056 577372 220108
rect 611360 220056 611412 220108
rect 621112 220056 621164 220108
rect 636476 220056 636528 220108
rect 653404 220056 653456 220108
rect 676496 220056 676548 220108
rect 677048 220056 677100 220108
rect 568304 219988 568356 220040
rect 574468 219988 574520 220040
rect 559564 219920 559616 219972
rect 622492 219852 622544 219904
rect 127716 219784 127768 219836
rect 195428 219784 195480 219836
rect 207204 219784 207256 219836
rect 257252 219784 257304 219836
rect 288440 219784 288492 219836
rect 310704 219784 310756 219836
rect 555792 219784 555844 219836
rect 558460 219784 558512 219836
rect 558828 219784 558880 219836
rect 546776 219716 546828 219768
rect 547420 219716 547472 219768
rect 555424 219716 555476 219768
rect 563428 219716 563480 219768
rect 564348 219716 564400 219768
rect 568580 219716 568632 219768
rect 568764 219716 568816 219768
rect 605656 219716 605708 219768
rect 606484 219716 606536 219768
rect 624332 219716 624384 219768
rect 137652 219648 137704 219700
rect 203156 219648 203208 219700
rect 236184 219648 236236 219700
rect 261484 219648 261536 219700
rect 558828 219648 558880 219700
rect 559380 219648 559432 219700
rect 563796 219648 563848 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 539968 219580 540020 219632
rect 558368 219580 558420 219632
rect 179420 219512 179472 219564
rect 231952 219512 232004 219564
rect 270776 219512 270828 219564
rect 279240 219512 279292 219564
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 70584 219376 70636 219428
rect 149060 219376 149112 219428
rect 149244 219376 149296 219428
rect 150256 219376 150308 219428
rect 152556 219376 152608 219428
rect 153108 219376 153160 219428
rect 155040 219376 155092 219428
rect 155960 219376 156012 219428
rect 156144 219376 156196 219428
rect 162860 219376 162912 219428
rect 165804 219376 165856 219428
rect 173164 219376 173216 219428
rect 179052 219376 179104 219428
rect 182824 219376 182876 219428
rect 183192 219376 183244 219428
rect 199292 219376 199344 219428
rect 199752 219376 199804 219428
rect 203064 219376 203116 219428
rect 204720 219376 204772 219428
rect 205640 219376 205692 219428
rect 209688 219376 209740 219428
rect 210332 219376 210384 219428
rect 212816 219376 212868 219428
rect 252560 219376 252612 219428
rect 254400 219376 254452 219428
rect 255320 219376 255372 219428
rect 272432 219376 272484 219428
rect 297364 219376 297416 219428
rect 312360 219376 312412 219428
rect 313280 219376 313332 219428
rect 323124 219376 323176 219428
rect 324228 219376 324280 219428
rect 324780 219376 324832 219428
rect 325516 219376 325568 219428
rect 326436 219376 326488 219428
rect 326896 219376 326948 219428
rect 63960 219240 64012 219292
rect 65524 219240 65576 219292
rect 113640 219240 113692 219292
rect 166264 219240 166316 219292
rect 192944 219240 192996 219292
rect 233884 219240 233936 219292
rect 237840 219240 237892 219292
rect 239404 219240 239456 219292
rect 252744 219240 252796 219292
rect 87144 219104 87196 219156
rect 106924 219104 106976 219156
rect 107108 219104 107160 219156
rect 159364 219104 159416 219156
rect 163320 219104 163372 219156
rect 59820 218968 59872 219020
rect 137284 218968 137336 219020
rect 143724 218968 143776 219020
rect 160744 218968 160796 219020
rect 162492 218968 162544 219020
rect 168932 218968 168984 219020
rect 169944 219104 169996 219156
rect 196624 219104 196676 219156
rect 203064 219104 203116 219156
rect 247132 219104 247184 219156
rect 259184 219240 259236 219292
rect 292304 219240 292356 219292
rect 307392 219240 307444 219292
rect 184204 218968 184256 219020
rect 186504 218968 186556 219020
rect 235632 218968 235684 219020
rect 246120 218968 246172 219020
rect 284024 218968 284076 219020
rect 300584 219104 300636 219156
rect 322848 219104 322900 219156
rect 323952 219240 324004 219292
rect 324964 219240 325016 219292
rect 327724 219376 327776 219428
rect 341340 219376 341392 219428
rect 342260 219376 342312 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 354588 219376 354640 219428
rect 355324 219376 355376 219428
rect 373632 219376 373684 219428
rect 378048 219376 378100 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 403440 219376 403492 219428
rect 404360 219376 404412 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 432052 219512 432104 219564
rect 558644 219512 558696 219564
rect 563520 219580 563572 219632
rect 676220 219648 676272 219700
rect 678428 219648 678480 219700
rect 605288 219580 605340 219632
rect 606300 219580 606352 219632
rect 622676 219580 622728 219632
rect 428280 219376 428332 219428
rect 438216 219376 438268 219428
rect 438860 219376 438912 219428
rect 439872 219376 439924 219428
rect 440332 219376 440384 219428
rect 527732 219376 527784 219428
rect 528284 219376 528336 219428
rect 548156 219376 548208 219428
rect 552664 219376 552716 219428
rect 563014 219444 563066 219496
rect 327264 219240 327316 219292
rect 342720 219240 342772 219292
rect 358728 219240 358780 219292
rect 363788 219240 363840 219292
rect 479708 219240 479760 219292
rect 480352 219240 480404 219292
rect 533712 219240 533764 219292
rect 534448 219240 534500 219292
rect 547880 219240 547932 219292
rect 549076 219240 549128 219292
rect 549904 219240 549956 219292
rect 553860 219308 553912 219360
rect 325608 219104 325660 219156
rect 330392 219104 330444 219156
rect 363696 219104 363748 219156
rect 374000 219104 374052 219156
rect 419172 219104 419224 219156
rect 422668 219104 422720 219156
rect 466092 219104 466144 219156
rect 472900 219104 472952 219156
rect 531964 219104 532016 219156
rect 532516 219104 532568 219156
rect 534264 219104 534316 219156
rect 537484 219104 537536 219156
rect 539692 219104 539744 219156
rect 544384 219104 544436 219156
rect 545028 219104 545080 219156
rect 548156 219104 548208 219156
rect 563704 219444 563756 219496
rect 564164 219444 564216 219496
rect 625160 219444 625212 219496
rect 605656 219308 605708 219360
rect 608784 219308 608836 219360
rect 289084 218968 289136 219020
rect 294144 218968 294196 219020
rect 309692 218968 309744 219020
rect 314016 218968 314068 219020
rect 339224 218968 339276 219020
rect 340512 218968 340564 219020
rect 351092 218968 351144 219020
rect 370320 218968 370372 219020
rect 375472 218968 375524 219020
rect 383568 218968 383620 219020
rect 388444 218968 388496 219020
rect 505100 218968 505152 219020
rect 83832 218832 83884 218884
rect 156144 218832 156196 218884
rect 92940 218696 92992 218748
rect 93768 218696 93820 218748
rect 100392 218696 100444 218748
rect 146944 218696 146996 218748
rect 149060 218696 149112 218748
rect 153200 218696 153252 218748
rect 153384 218696 153436 218748
rect 167644 218832 167696 218884
rect 173256 218832 173308 218884
rect 210884 218832 210936 218884
rect 232872 218832 232924 218884
rect 270776 218832 270828 218884
rect 285864 218832 285916 218884
rect 313832 218832 313884 218884
rect 166632 218696 166684 218748
rect 169760 218696 169812 218748
rect 171416 218696 171468 218748
rect 175924 218696 175976 218748
rect 176292 218696 176344 218748
rect 189724 218696 189776 218748
rect 63132 218628 63184 218680
rect 68284 218628 68336 218680
rect 93768 218560 93820 218612
rect 139952 218560 140004 218612
rect 140136 218560 140188 218612
rect 143724 218560 143776 218612
rect 146760 218560 146812 218612
rect 189908 218560 189960 218612
rect 68744 218288 68796 218340
rect 72424 218288 72476 218340
rect 120264 218288 120316 218340
rect 166448 218424 166500 218476
rect 168104 218424 168156 218476
rect 171048 218424 171100 218476
rect 172152 218424 172204 218476
rect 177212 218424 177264 218476
rect 179880 218424 179932 218476
rect 232688 218696 232740 218748
rect 233884 218696 233936 218748
rect 238852 218696 238904 218748
rect 239496 218696 239548 218748
rect 280712 218696 280764 218748
rect 291660 218696 291712 218748
rect 323584 218696 323636 218748
rect 198924 218560 198976 218612
rect 200028 218560 200080 218612
rect 201868 218560 201920 218612
rect 206192 218560 206244 218612
rect 206376 218560 206428 218612
rect 212816 218560 212868 218612
rect 213000 218560 213052 218612
rect 260012 218560 260064 218612
rect 262680 218560 262732 218612
rect 276572 218560 276624 218612
rect 279240 218560 279292 218612
rect 307024 218560 307076 218612
rect 320640 218560 320692 218612
rect 343640 218832 343692 218884
rect 347136 218832 347188 218884
rect 363512 218832 363564 218884
rect 392676 218832 392728 218884
rect 400772 218832 400824 218884
rect 401784 218832 401836 218884
rect 407764 218832 407816 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 499580 218832 499632 218884
rect 505284 218832 505336 218884
rect 534080 218968 534132 219020
rect 548708 218968 548760 219020
rect 563428 219240 563480 219292
rect 572444 219240 572496 219292
rect 572628 219240 572680 219292
rect 575664 219240 575716 219292
rect 591396 219172 591448 219224
rect 594156 219172 594208 219224
rect 554872 219104 554924 219156
rect 556896 219104 556948 219156
rect 587348 219104 587400 219156
rect 566740 218968 566792 219020
rect 518900 218900 518952 218952
rect 519452 218900 519504 218952
rect 524788 218900 524840 218952
rect 528468 218900 528520 218952
rect 534448 218832 534500 218884
rect 553676 218832 553728 218884
rect 553860 218832 553912 218884
rect 558184 218832 558236 218884
rect 559840 218832 559892 218884
rect 563014 218832 563066 218884
rect 563152 218832 563204 218884
rect 572260 218968 572312 219020
rect 572444 218968 572496 219020
rect 575848 218968 575900 219020
rect 567108 218832 567160 218884
rect 597744 218968 597796 219020
rect 587164 218832 587216 218884
rect 596824 218832 596876 218884
rect 519084 218764 519136 218816
rect 524420 218764 524472 218816
rect 533896 218764 533948 218816
rect 333704 218696 333756 218748
rect 352564 218696 352616 218748
rect 353760 218696 353812 218748
rect 367652 218696 367704 218748
rect 376944 218696 376996 218748
rect 385684 218696 385736 218748
rect 386052 218696 386104 218748
rect 396632 218696 396684 218748
rect 402612 218696 402664 218748
rect 409052 218696 409104 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 482928 218696 482980 218748
rect 485320 218696 485372 218748
rect 502800 218696 502852 218748
rect 503168 218696 503220 218748
rect 388536 218560 388588 218612
rect 393964 218560 394016 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 474740 218560 474792 218612
rect 482836 218560 482888 218612
rect 505284 218696 505336 218748
rect 505744 218696 505796 218748
rect 534080 218696 534132 218748
rect 548708 218696 548760 218748
rect 556896 218696 556948 218748
rect 550640 218560 550692 218612
rect 551560 218560 551612 218612
rect 552664 218560 552716 218612
rect 618168 218696 618220 218748
rect 558184 218560 558236 218612
rect 587164 218560 587216 218612
rect 587348 218560 587400 218612
rect 611544 218560 611596 218612
rect 196440 218424 196492 218476
rect 207664 218424 207716 218476
rect 210884 218424 210936 218476
rect 220820 218424 220872 218476
rect 225972 218424 226024 218476
rect 265624 218424 265676 218476
rect 265992 218424 266044 218476
rect 272432 218424 272484 218476
rect 272616 218424 272668 218476
rect 288440 218424 288492 218476
rect 500040 218424 500092 218476
rect 500224 218424 500276 218476
rect 604368 218424 604420 218476
rect 458180 218356 458232 218408
rect 136824 218288 136876 218340
rect 139492 218288 139544 218340
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 64144 218152 64196 218204
rect 67272 218152 67324 218204
rect 71044 218152 71096 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 130200 218152 130252 218204
rect 172612 218288 172664 218340
rect 174084 218288 174136 218340
rect 179420 218288 179472 218340
rect 190644 218288 190696 218340
rect 191656 218288 191708 218340
rect 192300 218288 192352 218340
rect 193128 218288 193180 218340
rect 193956 218288 194008 218340
rect 194508 218288 194560 218340
rect 198096 218288 198148 218340
rect 198648 218288 198700 218340
rect 199292 218288 199344 218340
rect 202052 218288 202104 218340
rect 203064 218288 203116 218340
rect 213184 218288 213236 218340
rect 219624 218288 219676 218340
rect 258080 218288 258132 218340
rect 365352 218288 365404 218340
rect 370504 218288 370556 218340
rect 426624 218288 426676 218340
rect 429568 218288 429620 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 510160 218288 510212 218340
rect 616144 218288 616196 218340
rect 142620 218152 142672 218204
rect 143264 218152 143316 218204
rect 145104 218152 145156 218204
rect 146116 218152 146168 218204
rect 159180 218152 159232 218204
rect 160008 218152 160060 218204
rect 160836 218152 160888 218204
rect 161940 218152 161992 218204
rect 164976 218152 165028 218204
rect 165528 218152 165580 218204
rect 167460 218152 167512 218204
rect 168288 218152 168340 218204
rect 169116 218152 169168 218204
rect 169576 218152 169628 218204
rect 169760 218152 169812 218204
rect 201868 218152 201920 218204
rect 202236 218152 202288 218204
rect 202696 218152 202748 218204
rect 208860 218152 208912 218204
rect 209504 218152 209556 218204
rect 210516 218152 210568 218204
rect 211068 218152 211120 218204
rect 211344 218152 211396 218204
rect 214288 218152 214340 218204
rect 214656 218152 214708 218204
rect 215208 218152 215260 218204
rect 215484 218152 215536 218204
rect 216588 218152 216640 218204
rect 218796 218152 218848 218204
rect 219348 218152 219400 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 60004 218016 60056 218068
rect 61476 218016 61528 218068
rect 62028 218016 62080 218068
rect 62304 218016 62356 218068
rect 63408 218016 63460 218068
rect 65616 218016 65668 218068
rect 66904 218016 66956 218068
rect 68100 218016 68152 218068
rect 68928 218016 68980 218068
rect 69756 218016 69808 218068
rect 70308 218016 70360 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 80520 218016 80572 218068
rect 81440 218016 81492 218068
rect 82176 218016 82228 218068
rect 82728 218016 82780 218068
rect 83004 218016 83056 218068
rect 84108 218016 84160 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 90456 218016 90508 218068
rect 91008 218016 91060 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 111984 218016 112036 218068
rect 112812 218016 112864 218068
rect 115296 218016 115348 218068
rect 115848 218016 115900 218068
rect 116124 218016 116176 218068
rect 116952 218016 117004 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 123576 218016 123628 218068
rect 124128 218016 124180 218068
rect 126060 218016 126112 218068
rect 126704 218016 126756 218068
rect 131856 218016 131908 218068
rect 132408 218016 132460 218068
rect 132684 218016 132736 218068
rect 133512 218016 133564 218068
rect 134340 218016 134392 218068
rect 134984 218016 135036 218068
rect 135996 218016 136048 218068
rect 136548 218016 136600 218068
rect 138480 218016 138532 218068
rect 139124 218016 139176 218068
rect 139492 218016 139544 218068
rect 171416 218016 171468 218068
rect 171600 218016 171652 218068
rect 172336 218016 172388 218068
rect 175740 218016 175792 218068
rect 176476 218016 176528 218068
rect 181536 218016 181588 218068
rect 181996 218016 182048 218068
rect 182364 218016 182416 218068
rect 183468 218016 183520 218068
rect 184848 218016 184900 218068
rect 185492 218016 185544 218068
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 188160 218016 188212 218068
rect 189172 218016 189224 218068
rect 189816 218016 189868 218068
rect 225604 218152 225656 218204
rect 249432 218152 249484 218204
rect 251732 218152 251784 218204
rect 289176 218152 289228 218204
rect 294604 218152 294656 218204
rect 297456 218152 297508 218204
rect 300124 218152 300176 218204
rect 304080 218152 304132 218204
rect 305644 218152 305696 218204
rect 332232 218152 332284 218204
rect 334992 218152 335044 218204
rect 338856 218152 338908 218204
rect 340144 218152 340196 218204
rect 348792 218152 348844 218204
rect 353300 218152 353352 218204
rect 368664 218152 368716 218204
rect 372252 218152 372304 218204
rect 375104 218152 375156 218204
rect 380072 218152 380124 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 394332 218152 394384 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 428464 218152 428516 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 435732 218152 435784 218204
rect 436836 218152 436888 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 498660 218152 498712 218204
rect 503628 218152 503680 218204
rect 505284 218152 505336 218204
rect 605748 218152 605800 218204
rect 648252 218152 648304 218204
rect 654784 218152 654836 218204
rect 221280 218016 221332 218068
rect 222568 218016 222620 218068
rect 222936 218016 222988 218068
rect 223488 218016 223540 218068
rect 223764 218016 223816 218068
rect 224592 218016 224644 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 227076 218016 227128 218068
rect 227628 218016 227680 218068
rect 229560 218016 229612 218068
rect 230480 218016 230532 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 233700 218016 233752 218068
rect 234620 218016 234672 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 244464 218016 244516 218068
rect 246304 218016 246356 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249616 218016 249668 218068
rect 251916 218016 251968 218068
rect 252376 218016 252428 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 258540 218016 258592 218068
rect 259368 218016 259420 218068
rect 264336 218016 264388 218068
rect 264888 218016 264940 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 268476 218016 268528 218068
rect 269028 218016 269080 218068
rect 269304 218016 269356 218068
rect 270224 218016 270276 218068
rect 270960 218016 271012 218068
rect 271604 218016 271656 218068
rect 273444 218016 273496 218068
rect 274088 218016 274140 218068
rect 275100 218016 275152 218068
rect 275652 218016 275704 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282460 218016 282512 218068
rect 284208 218016 284260 218068
rect 284852 218016 284904 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288072 218016 288124 218068
rect 290004 218016 290056 218068
rect 290832 218016 290884 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 295800 218016 295852 218068
rect 296720 218016 296772 218068
rect 299940 218016 299992 218068
rect 300768 218016 300820 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 308220 218016 308272 218068
rect 308772 218016 308824 218068
rect 310704 218016 310756 218068
rect 311808 218016 311860 218068
rect 314844 218016 314896 218068
rect 315856 218016 315908 218068
rect 316500 218016 316552 218068
rect 317144 218016 317196 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 319996 218016 320048 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335268 218016 335320 218068
rect 335544 218016 335596 218068
rect 336372 218016 336424 218068
rect 337200 218016 337252 218068
rect 337844 218016 337896 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 342996 218016 343048 218068
rect 343456 218016 343508 218068
rect 345480 218016 345532 218068
rect 346400 218016 346452 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 351276 218016 351328 218068
rect 351736 218016 351788 218068
rect 352104 218016 352156 218068
rect 354404 218016 354456 218068
rect 355416 218016 355468 218068
rect 355968 218016 356020 218068
rect 356244 218016 356296 218068
rect 357256 218016 357308 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361304 218016 361356 218068
rect 364524 218016 364576 218068
rect 365536 218016 365588 218068
rect 366180 218016 366232 218068
rect 366732 218016 366784 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372436 218016 372488 218068
rect 372804 218016 372856 218068
rect 373816 218016 373868 218068
rect 374460 218016 374512 218068
rect 375288 218016 375340 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 380256 218016 380308 218068
rect 380716 218016 380768 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 384396 218016 384448 218068
rect 384948 218016 385000 218068
rect 385224 218016 385276 218068
rect 386328 218016 386380 218068
rect 389364 218016 389416 218068
rect 390100 218016 390152 218068
rect 391020 218016 391072 218068
rect 391572 218016 391624 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 398472 218016 398524 218068
rect 400956 218016 401008 218068
rect 401508 218016 401560 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 418344 218016 418396 218068
rect 419448 218016 419500 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 434904 218016 434956 218068
rect 436284 218016 436336 218068
rect 436468 218016 436520 218068
rect 437756 218016 437808 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 483572 218016 483624 218068
rect 486976 218016 487028 218068
rect 519452 218016 519504 218068
rect 520188 218016 520240 218068
rect 524788 218016 524840 218068
rect 539692 218016 539744 218068
rect 563014 218016 563066 218068
rect 573180 218016 573232 218068
rect 582288 218016 582340 218068
rect 655428 218016 655480 218068
rect 656164 218016 656216 218068
rect 518900 217880 518952 217932
rect 524604 217880 524656 217932
rect 514944 217744 514996 217796
rect 518716 217744 518768 217796
rect 518900 217744 518952 217796
rect 534080 217948 534132 218000
rect 538404 217948 538456 218000
rect 538956 217948 539008 218000
rect 539508 217948 539560 218000
rect 563152 217948 563204 218000
rect 568304 217948 568356 218000
rect 568672 217948 568724 218000
rect 572168 217948 572220 218000
rect 572306 217948 572358 218000
rect 525984 217812 526036 217864
rect 526720 217812 526772 217864
rect 534172 217812 534224 217864
rect 563244 217812 563296 217864
rect 563428 217812 563480 217864
rect 567568 217812 567620 217864
rect 572720 217812 572772 217864
rect 610072 217812 610124 217864
rect 528284 217676 528336 217728
rect 539048 217676 539100 217728
rect 539508 217676 539560 217728
rect 568120 217676 568172 217728
rect 572076 217676 572128 217728
rect 572260 217676 572312 217728
rect 572720 217676 572772 217728
rect 573088 217676 573140 217728
rect 577320 217676 577372 217728
rect 582104 217676 582156 217728
rect 586888 217676 586940 217728
rect 592040 217676 592092 217728
rect 594984 217676 595036 217728
rect 605748 217676 605800 217728
rect 615040 217676 615092 217728
rect 517704 217608 517756 217660
rect 518348 217472 518400 217524
rect 519084 217472 519136 217524
rect 526720 217540 526772 217592
rect 128544 217404 128596 217456
rect 199108 217404 199160 217456
rect 534172 217404 534224 217456
rect 535920 217336 535972 217388
rect 538680 217336 538732 217388
rect 103658 217200 103710 217252
rect 178408 217268 178460 217320
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 477592 217200 477644 217252
rect 478742 217200 478794 217252
rect 510620 217200 510672 217252
rect 511862 217200 511914 217252
rect 523040 217200 523092 217252
rect 524282 217200 524334 217252
rect 533344 217200 533396 217252
rect 596640 217404 596692 217456
rect 602068 217540 602120 217592
rect 613384 217540 613436 217592
rect 602344 217404 602396 217456
rect 604368 217404 604420 217456
rect 614120 217404 614172 217456
rect 539048 217268 539100 217320
rect 603080 217268 603132 217320
rect 612740 217268 612792 217320
rect 629392 217268 629444 217320
rect 539048 217132 539100 217184
rect 604552 217132 604604 217184
rect 523454 217064 523506 217116
rect 575480 216996 575532 217048
rect 577320 216996 577372 217048
rect 605104 216996 605156 217048
rect 582380 216860 582432 216912
rect 592040 216860 592092 216912
rect 596640 216860 596692 216912
rect 604000 216860 604052 216912
rect 618168 216656 618220 216708
rect 623872 216656 623924 216708
rect 597744 216044 597796 216096
rect 626080 216044 626132 216096
rect 596824 215908 596876 215960
rect 625252 215908 625304 215960
rect 577044 215840 577096 215892
rect 582564 215840 582616 215892
rect 594616 215568 594668 215620
rect 598480 215568 598532 215620
rect 596180 215296 596232 215348
rect 596824 215296 596876 215348
rect 611544 215296 611596 215348
rect 614488 215296 614540 215348
rect 676036 215092 676088 215144
rect 677600 215092 677652 215144
rect 575848 214956 575900 215008
rect 612280 214956 612332 215008
rect 574468 214820 574520 214872
rect 612832 214820 612884 214872
rect 675852 214820 675904 214872
rect 677324 214820 677376 214872
rect 575664 214684 575716 214736
rect 622308 214684 622360 214736
rect 628564 214684 628616 214736
rect 632888 214684 632940 214736
rect 652852 214684 652904 214736
rect 661684 214684 661736 214736
rect 574100 214548 574152 214600
rect 607312 214548 607364 214600
rect 607864 214548 607916 214600
rect 608784 214548 608836 214600
rect 609520 214548 609572 214600
rect 621112 214548 621164 214600
rect 621664 214548 621716 214600
rect 622492 214548 622544 214600
rect 623320 214548 623372 214600
rect 627920 214548 627972 214600
rect 628840 214548 628892 214600
rect 636292 214548 636344 214600
rect 639604 214548 639656 214600
rect 648436 214548 648488 214600
rect 658924 214548 658976 214600
rect 627184 214412 627236 214464
rect 35808 213936 35860 213988
rect 41696 213936 41748 213988
rect 627736 213936 627788 213988
rect 631600 213936 631652 213988
rect 637580 213868 637632 213920
rect 638224 213868 638276 213920
rect 645492 213868 645544 213920
rect 646136 213868 646188 213920
rect 648620 213868 648672 213920
rect 649264 213868 649316 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 638040 213732 638092 213784
rect 641168 213732 641220 213784
rect 660948 213732 661000 213784
rect 663064 213732 663116 213784
rect 641628 213596 641680 213648
rect 650644 213596 650696 213648
rect 651840 213596 651892 213648
rect 657544 213596 657596 213648
rect 676036 213596 676088 213648
rect 676956 213596 677008 213648
rect 635556 213460 635608 213512
rect 652392 213460 652444 213512
rect 663156 213460 663208 213512
rect 665824 213460 665876 213512
rect 575480 213324 575532 213376
rect 601792 213324 601844 213376
rect 640248 213324 640300 213376
rect 660764 213324 660816 213376
rect 574284 213188 574336 213240
rect 615592 213188 615644 213240
rect 642180 213188 642232 213240
rect 664168 213120 664220 213172
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 632704 212712 632756 212764
rect 634360 212712 634412 212764
rect 658740 212712 658792 212764
rect 659476 212712 659528 212764
rect 600320 212372 600372 212424
rect 601240 212372 601292 212424
rect 35624 211284 35676 211336
rect 41696 211284 41748 211336
rect 578240 211284 578292 211336
rect 580448 211284 580500 211336
rect 35808 211148 35860 211200
rect 41696 211148 41748 211200
rect 600504 211012 600556 211064
rect 600872 211012 600924 211064
rect 619640 211012 619692 211064
rect 620008 211012 620060 211064
rect 35808 209788 35860 209840
rect 41328 209788 41380 209840
rect 579252 209788 579304 209840
rect 581736 209788 581788 209840
rect 581552 208564 581604 208616
rect 632152 209516 632204 209568
rect 652024 209516 652076 209568
rect 652208 209516 652260 209568
rect 666836 209516 666888 209568
rect 666652 209040 666704 209092
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 580448 207612 580500 207664
rect 589464 207612 589516 207664
rect 581736 206252 581788 206304
rect 589648 206252 589700 206304
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 667940 199180 667992 199232
rect 670792 199180 670844 199232
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 667940 194284 667992 194336
rect 670792 194284 670844 194336
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 667940 189388 667992 189440
rect 670792 189388 670844 189440
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 669228 184492 669280 184544
rect 669780 184492 669832 184544
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 667940 174700 667992 174752
rect 670240 174700 670292 174752
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 667940 169668 667992 169720
rect 670056 169668 670108 169720
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 675852 162528 675904 162580
rect 681004 162528 681056 162580
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580448 151784 580500 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 668308 150220 668360 150272
rect 670792 150220 670844 150272
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 579252 145256 579304 145308
rect 585140 145256 585192 145308
rect 585968 144916 586020 144968
rect 589464 144916 589516 144968
rect 579528 144644 579580 144696
rect 584404 144644 584456 144696
rect 584588 143556 584640 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 583024 140768 583076 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580448 140700 580500 140752
rect 580264 139408 580316 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579068 136824 579120 136876
rect 585968 136824 586020 136876
rect 585784 136620 585836 136672
rect 589464 136620 589516 136672
rect 584404 135260 584456 135312
rect 589464 135260 589516 135312
rect 579528 135124 579580 135176
rect 588544 135124 588596 135176
rect 580632 131724 580684 131776
rect 590292 131724 590344 131776
rect 578884 131248 578936 131300
rect 589464 131248 589516 131300
rect 579068 131112 579120 131164
rect 584588 131112 584640 131164
rect 579160 128256 579212 128308
rect 587164 128256 587216 128308
rect 587624 127168 587676 127220
rect 589464 127168 589516 127220
rect 579068 126216 579120 126268
rect 587624 126216 587676 126268
rect 579528 125332 579580 125384
rect 583024 125332 583076 125384
rect 583208 124856 583260 124908
rect 589648 124856 589700 124908
rect 578332 124108 578384 124160
rect 580264 124108 580316 124160
rect 580448 122816 580500 122868
rect 589464 122816 589516 122868
rect 581828 122068 581880 122120
rect 590108 122068 590160 122120
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 579528 121388 579580 121440
rect 585784 121388 585836 121440
rect 667940 120096 667992 120148
rect 670148 120096 670200 120148
rect 584588 118668 584640 118720
rect 589464 118668 589516 118720
rect 578700 118532 578752 118584
rect 584404 118532 584456 118584
rect 668032 118532 668084 118584
rect 670332 118532 670384 118584
rect 585968 117308 586020 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 678244 117240 678296 117292
rect 578700 117172 578752 117224
rect 580632 117172 580684 117224
rect 585784 115948 585836 116000
rect 589464 115948 589516 116000
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 584404 113160 584456 113212
rect 589464 113160 589516 113212
rect 579160 113024 579212 113076
rect 588728 113024 588780 113076
rect 588544 111800 588596 111852
rect 590384 111800 590436 111852
rect 581644 111052 581696 111104
rect 589924 111052 589976 111104
rect 583024 109692 583076 109744
rect 589372 109692 589424 109744
rect 578884 108944 578936 108996
rect 581828 108944 581880 108996
rect 581276 107652 581328 107704
rect 589464 107652 589516 107704
rect 666560 106088 666612 106140
rect 666836 106088 666888 106140
rect 670700 106088 670752 106140
rect 579344 105136 579396 105188
rect 581276 105136 581328 105188
rect 581828 104864 581880 104916
rect 589464 104864 589516 104916
rect 580264 104116 580316 104168
rect 589648 104116 589700 104168
rect 578332 103300 578384 103352
rect 583208 103300 583260 103352
rect 578516 102076 578568 102128
rect 580448 102076 580500 102128
rect 587164 100716 587216 100768
rect 590292 100716 590344 100768
rect 624792 100104 624844 100156
rect 668400 100104 668452 100156
rect 580448 99968 580500 100020
rect 590108 99968 590160 100020
rect 594064 99968 594116 100020
rect 667940 99968 667992 100020
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 579160 99220 579212 99272
rect 581644 99220 581696 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 627552 98880 627604 98932
rect 640708 98880 640760 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98744 647200 98796
rect 661960 98744 662012 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 631416 98200 631468 98252
rect 642180 98132 642232 98184
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 629760 97928 629812 97980
rect 645124 97996 645176 98048
rect 653956 97928 654008 97980
rect 655060 97928 655112 97980
rect 628288 97792 628340 97844
rect 631416 97792 631468 97844
rect 631600 97792 631652 97844
rect 637764 97792 637816 97844
rect 644296 97792 644348 97844
rect 658832 97792 658884 97844
rect 591304 97656 591356 97708
rect 598204 97656 598256 97708
rect 620192 97656 620244 97708
rect 625988 97656 626040 97708
rect 626816 97656 626868 97708
rect 639236 97656 639288 97708
rect 643008 97656 643060 97708
rect 658004 97656 658056 97708
rect 658188 97656 658240 97708
rect 663064 97656 663116 97708
rect 626172 97520 626224 97572
rect 631600 97520 631652 97572
rect 631968 97520 632020 97572
rect 648620 97520 648672 97572
rect 650368 97520 650420 97572
rect 658280 97520 658332 97572
rect 659200 97520 659252 97572
rect 663892 97520 663944 97572
rect 612648 97384 612700 97436
rect 620284 97384 620336 97436
rect 623136 97384 623188 97436
rect 632060 97384 632112 97436
rect 632704 97384 632756 97436
rect 650276 97384 650328 97436
rect 651840 97384 651892 97436
rect 659568 97384 659620 97436
rect 659936 97384 659988 97436
rect 665364 97384 665416 97436
rect 605472 97248 605524 97300
rect 613384 97248 613436 97300
rect 621664 97248 621716 97300
rect 629300 97248 629352 97300
rect 633256 97248 633308 97300
rect 650552 97248 650604 97300
rect 656808 97180 656860 97232
rect 661408 97180 661460 97232
rect 634728 97112 634780 97164
rect 649080 97112 649132 97164
rect 658004 97044 658056 97096
rect 660120 97044 660172 97096
rect 624608 96976 624660 97028
rect 635004 96976 635056 97028
rect 638592 96976 638644 97028
rect 647792 96976 647844 97028
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 610624 96908 610676 96960
rect 611084 96908 611136 96960
rect 614028 96908 614080 96960
rect 614764 96908 614816 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 660672 96908 660724 96960
rect 663248 96908 663300 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 634176 96840 634228 96892
rect 647976 96840 648028 96892
rect 613568 96772 613620 96824
rect 614028 96772 614080 96824
rect 655244 96772 655296 96824
rect 662512 96772 662564 96824
rect 639052 96568 639104 96620
rect 640340 96568 640392 96620
rect 640524 96568 640576 96620
rect 648436 96568 648488 96620
rect 653312 96568 653364 96620
rect 665180 96568 665232 96620
rect 640064 96432 640116 96484
rect 652024 96432 652076 96484
rect 652576 96432 652628 96484
rect 664168 96432 664220 96484
rect 631232 96296 631284 96348
rect 647148 96296 647200 96348
rect 648896 96296 648948 96348
rect 664352 96296 664404 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 641536 96024 641588 96076
rect 663708 96024 663760 96076
rect 577504 95888 577556 95940
rect 600412 95888 600464 95940
rect 609152 95888 609204 95940
rect 621664 95888 621716 95940
rect 644848 95888 644900 95940
rect 648068 95888 648120 95940
rect 648436 95888 648488 95940
rect 664536 95888 664588 95940
rect 645768 95752 645820 95804
rect 652208 95752 652260 95804
rect 646412 95616 646464 95668
rect 653404 95616 653456 95668
rect 640340 95412 640392 95464
rect 643468 95412 643520 95464
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 579528 95004 579580 95056
rect 584588 95004 584640 95056
rect 648160 95344 648212 95396
rect 656164 95752 656216 95804
rect 647884 95140 647936 95192
rect 648068 95140 648120 95192
rect 650000 95140 650052 95192
rect 648804 95004 648856 95056
rect 607680 94596 607732 94648
rect 620928 94596 620980 94648
rect 606944 94460 606996 94512
rect 623044 94460 623096 94512
rect 648436 93848 648488 93900
rect 654784 93848 654836 93900
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 651288 93508 651340 93560
rect 655428 93508 655480 93560
rect 579160 93372 579212 93424
rect 585968 93372 586020 93424
rect 611084 93100 611136 93152
rect 618536 93100 618588 93152
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 616604 91740 616656 91792
rect 626264 91740 626316 91792
rect 578516 91672 578568 91724
rect 585784 91672 585836 91724
rect 647700 91672 647752 91724
rect 654692 91672 654744 91724
rect 618168 91128 618220 91180
rect 611268 90992 611320 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 648804 90652 648856 90704
rect 655428 90652 655480 90704
rect 620928 89632 620980 89684
rect 626448 89632 626500 89684
rect 581644 88952 581696 89004
rect 601700 88952 601752 89004
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 578516 88272 578568 88324
rect 588544 88272 588596 88324
rect 618168 88272 618220 88324
rect 625620 88272 625672 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 623044 88136 623096 88188
rect 626448 88136 626500 88188
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 659568 86912 659620 86964
rect 663248 86912 663300 86964
rect 652208 86844 652260 86896
rect 657728 86844 657780 86896
rect 647884 86708 647936 86760
rect 661408 86708 661460 86760
rect 652024 86572 652076 86624
rect 660120 86572 660172 86624
rect 656164 86436 656216 86488
rect 660672 86436 660724 86488
rect 618536 86300 618588 86352
rect 626448 86300 626500 86352
rect 654876 86300 654928 86352
rect 662512 86300 662564 86352
rect 653404 86164 653456 86216
rect 657176 86164 657228 86216
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 579068 85416 579120 85468
rect 581828 85416 581880 85468
rect 621664 85348 621716 85400
rect 625252 85348 625304 85400
rect 608508 84124 608560 84176
rect 626448 84124 626500 84176
rect 579528 83988 579580 84040
rect 583024 83988 583076 84040
rect 578516 82560 578568 82612
rect 584404 82560 584456 82612
rect 628748 80928 628800 80980
rect 642456 80928 642508 80980
rect 615408 80792 615460 80844
rect 646136 80792 646188 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 612648 79432 612700 79484
rect 645952 79432 646004 79484
rect 584404 79296 584456 79348
rect 589924 79296 589976 79348
rect 614764 79296 614816 79348
rect 648712 79296 648764 79348
rect 578516 78412 578568 78464
rect 580264 78412 580316 78464
rect 633440 78208 633492 78260
rect 645308 78208 645360 78260
rect 631048 78072 631100 78124
rect 643100 78072 643152 78124
rect 614028 77936 614080 77988
rect 647240 77936 647292 77988
rect 628472 77392 628524 77444
rect 632796 77392 632848 77444
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 616788 76644 616840 76696
rect 646504 76644 646556 76696
rect 579344 76508 579396 76560
rect 666560 76508 666612 76560
rect 621664 75896 621716 75948
rect 628472 75896 628524 75948
rect 620284 75420 620336 75472
rect 648896 75420 648948 75472
rect 607128 75284 607180 75336
rect 646320 75284 646372 75336
rect 613384 75148 613436 75200
rect 662604 75148 662656 75200
rect 579528 73108 579580 73160
rect 587164 73108 587216 73160
rect 578516 71544 578568 71596
rect 584404 71544 584456 71596
rect 584404 68280 584456 68332
rect 604460 68280 604512 68332
rect 579528 66240 579580 66292
rect 623044 66240 623096 66292
rect 579528 64812 579580 64864
rect 594064 64812 594116 64864
rect 579528 62024 579580 62076
rect 612004 62024 612056 62076
rect 579528 60664 579580 60716
rect 624424 60664 624476 60716
rect 579068 58760 579120 58812
rect 597560 58760 597612 58812
rect 577688 58624 577740 58676
rect 603080 58624 603132 58676
rect 574928 57332 574980 57384
rect 600504 57332 600556 57384
rect 575480 57196 575532 57248
rect 601884 57196 601936 57248
rect 578516 56516 578568 56568
rect 621664 56516 621716 56568
rect 574744 55972 574796 56024
rect 598940 55972 598992 56024
rect 574560 55836 574612 55888
rect 599124 55836 599176 55888
rect 577504 55156 577556 55208
rect 462136 53592 462188 53644
rect 591304 55020 591356 55072
rect 596456 54884 596508 54936
rect 596272 54748 596324 54800
rect 463332 53592 463384 53644
rect 464068 53592 464120 53644
rect 464988 53592 465040 53644
rect 465908 53592 465960 53644
rect 625988 54612 626040 54664
rect 625804 54476 625856 54528
rect 580448 54340 580500 54392
rect 579068 54204 579120 54256
rect 574560 54068 574612 54120
rect 467932 53592 467984 53644
rect 468576 53592 468628 53644
rect 468760 53592 468812 53644
rect 461308 53456 461360 53508
rect 574928 53932 574980 53984
rect 49148 53320 49200 53372
rect 129188 53320 129240 53372
rect 463148 53320 463200 53372
rect 50344 53184 50396 53236
rect 130384 53184 130436 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 465448 53116 465500 53168
rect 468576 53116 468628 53168
rect 46204 53048 46256 53100
rect 129004 53048 129056 53100
rect 460066 52776 460118 52828
rect 467932 52912 467984 52964
rect 464206 52776 464258 52828
rect 468760 52776 468812 52828
rect 48964 51960 49016 52012
rect 129556 51960 129608 52012
rect 47584 51824 47636 51876
rect 129372 51824 129424 51876
rect 46388 51688 46440 51740
rect 130568 51688 130620 51740
rect 145380 51688 145432 51740
rect 306012 51688 306064 51740
rect 50528 50464 50580 50516
rect 128728 50464 128780 50516
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 128544 50328 128596 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 51724 49104 51776 49156
rect 128912 49104 128964 49156
rect 47768 48968 47820 49020
rect 131028 48968 131080 49020
rect 128912 47812 128964 47864
rect 131580 47812 131632 47864
rect 128728 47676 128780 47728
rect 132040 47676 132092 47728
rect 623044 46452 623096 46504
rect 661592 46452 661644 46504
rect 129556 45024 129608 45076
rect 129372 44752 129424 44804
rect 131580 44752 131632 44804
rect 129188 44616 129240 44668
rect 129004 44480 129056 44532
rect 132040 44480 132092 44532
rect 132408 44412 132460 44464
rect 130568 44276 130620 44328
rect 128544 44140 128596 44192
rect 132224 44140 132276 44192
rect 130384 44004 130436 44056
rect 131028 43868 131080 43920
rect 43444 42780 43496 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 439596 43596 439648 43648
rect 441620 43596 441672 43648
rect 310428 42712 310480 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 463056 42712 463108 42764
rect 404452 42304 404504 42356
rect 405556 42304 405608 42356
rect 420736 42304 420788 42356
rect 427084 42304 427136 42356
rect 662420 42173 662472 42225
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 427084 41420 427136 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 428002 1006904 428058 1006913
rect 428002 1006839 428004 1006848
rect 428056 1006839 428058 1006848
rect 504546 1006904 504602 1006913
rect 559654 1006904 559710 1006913
rect 504546 1006839 504548 1006848
rect 428004 1006810 428056 1006816
rect 504600 1006839 504602 1006848
rect 516968 1006868 517020 1006874
rect 504548 1006810 504600 1006816
rect 516968 1006810 517020 1006816
rect 556988 1006868 557040 1006874
rect 559654 1006839 559656 1006848
rect 556988 1006810 557040 1006816
rect 559708 1006839 559710 1006848
rect 559656 1006810 559708 1006816
rect 428370 1006768 428426 1006777
rect 505374 1006768 505430 1006777
rect 428370 1006703 428372 1006712
rect 428424 1006703 428426 1006712
rect 434444 1006732 434496 1006738
rect 428372 1006674 428424 1006680
rect 505374 1006703 505376 1006712
rect 434444 1006674 434496 1006680
rect 505428 1006703 505430 1006712
rect 515404 1006732 515456 1006738
rect 505376 1006674 505428 1006680
rect 515404 1006674 515456 1006680
rect 357716 1006664 357768 1006670
rect 152922 1006632 152978 1006641
rect 145564 1006596 145616 1006602
rect 308126 1006632 308182 1006641
rect 152922 1006567 152924 1006576
rect 145564 1006538 145616 1006544
rect 152976 1006567 152978 1006576
rect 300124 1006596 300176 1006602
rect 152924 1006538 152976 1006544
rect 308126 1006567 308128 1006576
rect 300124 1006538 300176 1006544
rect 308180 1006567 308182 1006576
rect 357714 1006632 357716 1006641
rect 371884 1006664 371936 1006670
rect 357768 1006632 357770 1006641
rect 371884 1006606 371936 1006612
rect 357714 1006567 357770 1006576
rect 308128 1006538 308180 1006544
rect 103978 1006496 104034 1006505
rect 94504 1006460 94556 1006466
rect 103978 1006431 103980 1006440
rect 94504 1006402 94556 1006408
rect 104032 1006431 104034 1006440
rect 103980 1006402 104032 1006408
rect 93308 1006188 93360 1006194
rect 93308 1006130 93360 1006136
rect 93124 1006052 93176 1006058
rect 93124 1005994 93176 1006000
rect 92664 1003944 92716 1003950
rect 92664 1003886 92716 1003892
rect 92480 998708 92532 998714
rect 92480 998650 92532 998656
rect 92296 998436 92348 998442
rect 92296 998378 92348 998384
rect 92308 997914 92336 998378
rect 92308 997886 92428 997914
rect 74446 996976 74502 996985
rect 74446 996911 74502 996920
rect 74630 996976 74686 996985
rect 74630 996911 74686 996920
rect 74460 994566 74488 996911
rect 74644 994702 74672 996911
rect 80426 995752 80482 995761
rect 80178 995710 80426 995738
rect 84658 995752 84714 995761
rect 84502 995710 84658 995738
rect 80426 995687 80482 995696
rect 87878 995752 87934 995761
rect 87538 995710 87878 995738
rect 84658 995687 84714 995696
rect 88982 995752 89038 995761
rect 88734 995710 88982 995738
rect 87878 995687 87934 995696
rect 89626 995752 89682 995761
rect 89378 995710 89626 995738
rect 88982 995687 89038 995696
rect 89626 995687 89682 995696
rect 92400 995602 92428 997886
rect 92032 995574 92428 995602
rect 77942 995480 77998 995489
rect 77036 995217 77064 995452
rect 77694 995438 77942 995466
rect 90270 995480 90326 995489
rect 77942 995415 77998 995424
rect 77022 995208 77078 995217
rect 77022 995143 77078 995152
rect 78324 994838 78352 995452
rect 78312 994832 78364 994838
rect 78312 994774 78364 994780
rect 74632 994696 74684 994702
rect 74632 994638 74684 994644
rect 74448 994560 74500 994566
rect 74448 994502 74500 994508
rect 73160 994288 73212 994294
rect 73160 994230 73212 994236
rect 51724 993200 51776 993206
rect 51724 993142 51776 993148
rect 50344 993064 50396 993070
rect 50344 993006 50396 993012
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 44824 990140 44876 990146
rect 44824 990082 44876 990088
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 968833 42196 969272
rect 42154 968824 42210 968833
rect 42154 968759 42210 968768
rect 42182 968034 42564 968062
rect 41984 967201 42012 967405
rect 41970 967192 42026 967201
rect 41970 967127 42026 967136
rect 42338 966784 42394 966793
rect 42182 966742 42338 966770
rect 42338 966719 42394 966728
rect 42536 966014 42564 968034
rect 43456 966793 43484 975666
rect 43810 968824 43866 968833
rect 43810 968759 43866 968768
rect 43442 966784 43498 966793
rect 43442 966719 43498 966728
rect 42536 965986 42656 966014
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42444 963937 42472 964362
rect 42430 963928 42486 963937
rect 42430 963863 42486 963872
rect 42182 963711 42472 963739
rect 42444 963393 42472 963711
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42338 963112 42394 963121
rect 42182 963070 42338 963098
rect 42338 963047 42394 963056
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 41786 959103 41842 959112
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 42076 957953 42104 958188
rect 42062 957944 42118 957953
rect 42062 957879 42118 957888
rect 42182 956338 42380 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 42260 953594 42288 955182
rect 41708 953566 42288 953594
rect 28538 952912 28594 952921
rect 28538 952847 28594 952856
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28552 942721 28580 952847
rect 41708 952474 41736 953566
rect 36544 952468 36596 952474
rect 36544 952410 36596 952416
rect 41696 952468 41748 952474
rect 41696 952410 41748 952416
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35820 942750 35848 943055
rect 35808 942744 35860 942750
rect 28538 942712 28594 942721
rect 35808 942686 35860 942692
rect 28538 942647 28594 942656
rect 35806 941896 35862 941905
rect 35806 941831 35862 941840
rect 35820 941390 35848 941831
rect 35808 941384 35860 941390
rect 35808 941326 35860 941332
rect 35806 940264 35862 940273
rect 35806 940199 35862 940208
rect 35820 939894 35848 940199
rect 35808 939888 35860 939894
rect 35808 939830 35860 939836
rect 36556 938471 36584 952410
rect 42352 952354 42380 956338
rect 42628 956354 42656 965986
rect 43166 963384 43222 963393
rect 43166 963319 43222 963328
rect 42798 963112 42854 963121
rect 42798 963047 42854 963056
rect 42628 956326 42748 956354
rect 42720 953594 42748 956326
rect 41708 952326 42380 952354
rect 42536 953566 42748 953594
rect 42812 953594 42840 963047
rect 42812 953566 42932 953594
rect 41708 952270 41736 952326
rect 37924 952264 37976 952270
rect 41696 952264 41748 952270
rect 37924 952206 37976 952212
rect 39302 952232 39358 952241
rect 37936 939049 37964 952206
rect 41696 952206 41748 952212
rect 39302 952167 39358 952176
rect 38476 941384 38528 941390
rect 38476 941326 38528 941332
rect 37922 939040 37978 939049
rect 37922 938975 37978 938984
rect 36542 938462 36598 938471
rect 36542 938397 36598 938406
rect 38488 937582 38516 941326
rect 38476 937576 38528 937582
rect 38476 937518 38528 937524
rect 39316 937417 39344 952167
rect 41602 951960 41658 951969
rect 41602 951895 41658 951904
rect 40038 951824 40094 951833
rect 40038 951759 40094 951768
rect 39488 939888 39540 939894
rect 39488 939830 39540 939836
rect 39500 938194 39528 939830
rect 39488 938188 39540 938194
rect 39488 938130 39540 938136
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 40052 934391 40080 951759
rect 41418 951688 41474 951697
rect 41418 951623 41474 951632
rect 40406 943800 40462 943809
rect 40406 943735 40462 943744
rect 40420 942750 40448 943735
rect 40408 942744 40460 942750
rect 40408 942686 40460 942692
rect 41432 938641 41460 951623
rect 41616 944353 41644 951895
rect 42536 949454 42564 953566
rect 41708 949426 42564 949454
rect 41708 946694 41736 949426
rect 41708 946666 41920 946694
rect 41892 945314 41920 946666
rect 41800 945286 41920 945314
rect 41602 944344 41658 944353
rect 41602 944279 41658 944288
rect 41800 940250 41828 945286
rect 42246 943800 42302 943809
rect 42246 943735 42302 943744
rect 41616 940222 41828 940250
rect 41418 938632 41474 938641
rect 41418 938567 41474 938576
rect 41616 938346 41644 940222
rect 41524 938318 41644 938346
rect 41524 937122 41552 938318
rect 41696 938188 41748 938194
rect 41696 938130 41748 938136
rect 41708 938074 41736 938130
rect 41708 938046 42196 938074
rect 41696 937576 41748 937582
rect 41748 937536 42012 937564
rect 41696 937518 41748 937524
rect 41524 937094 41920 937122
rect 40038 934382 40094 934391
rect 40038 934317 40094 934326
rect 41328 934380 41380 934386
rect 41328 934322 41380 934328
rect 41696 934380 41748 934386
rect 41892 934368 41920 937094
rect 41748 934340 41920 934368
rect 41696 934322 41748 934328
rect 41340 932929 41368 934322
rect 41326 932920 41382 932929
rect 41326 932855 41382 932864
rect 41984 930134 42012 937536
rect 42168 937122 42196 938046
rect 41800 930106 42012 930134
rect 42076 937094 42196 937122
rect 42076 930134 42104 937094
rect 42260 935785 42288 943735
rect 42246 935776 42302 935785
rect 42246 935711 42302 935720
rect 42904 934153 42932 953566
rect 43180 934969 43208 963319
rect 43444 961920 43496 961926
rect 43444 961862 43496 961868
rect 43456 952921 43484 961862
rect 43626 958760 43682 958769
rect 43626 958695 43682 958704
rect 43442 952912 43498 952921
rect 43442 952847 43498 952856
rect 43640 936193 43668 958695
rect 43824 937009 43852 968759
rect 44638 964744 44694 964753
rect 44638 964679 44694 964688
rect 44270 963928 44326 963937
rect 44270 963863 44326 963872
rect 43810 937000 43866 937009
rect 43810 936935 43866 936944
rect 43626 936184 43682 936193
rect 43626 936119 43682 936128
rect 43166 934960 43222 934969
rect 43166 934895 43222 934904
rect 42890 934144 42946 934153
rect 42890 934079 42946 934088
rect 44284 933745 44312 963863
rect 44454 941080 44510 941089
rect 44454 941015 44510 941024
rect 44270 933736 44326 933745
rect 44270 933671 44326 933680
rect 43626 933328 43682 933337
rect 43626 933263 43682 933272
rect 42076 930106 42288 930134
rect 41800 911849 41828 930106
rect 42260 911985 42288 930106
rect 42246 911976 42302 911985
rect 42246 911911 42302 911920
rect 41786 911840 41842 911849
rect 41786 911775 41842 911784
rect 42936 892256 42992 892265
rect 42936 892191 42992 892200
rect 43074 891984 43130 891993
rect 43074 891919 43076 891928
rect 43128 891919 43130 891928
rect 43076 891890 43128 891896
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817086 35848 817255
rect 35808 817080 35860 817086
rect 35808 817022 35860 817028
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 815658 35848 816439
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814298 35848 814807
rect 41432 814298 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815674 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815658 41644 815674
rect 41524 815652 41656 815658
rect 41524 815646 41604 815652
rect 41604 815594 41656 815600
rect 43074 815280 43130 815289
rect 43074 815215 43130 815224
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41420 814292 41472 814298
rect 41420 814234 41472 814240
rect 41142 813240 41198 813249
rect 41142 813175 41198 813184
rect 40958 812424 41014 812433
rect 40958 812359 41014 812368
rect 39302 811608 39358 811617
rect 39302 811543 39358 811552
rect 33046 811200 33102 811209
rect 33046 811135 33102 811144
rect 33060 802466 33088 811135
rect 33048 802460 33100 802466
rect 33048 802402 33100 802408
rect 39316 801718 39344 811543
rect 40972 805361 41000 812359
rect 41156 805633 41184 813175
rect 41326 812832 41382 812841
rect 41326 812767 41382 812776
rect 41340 810762 41368 812767
rect 41328 810756 41380 810762
rect 41328 810698 41380 810704
rect 41696 810756 41748 810762
rect 41696 810698 41748 810704
rect 41708 810642 41736 810698
rect 41708 810614 42104 810642
rect 42076 808694 42104 810614
rect 42522 809024 42578 809033
rect 42522 808959 42578 808968
rect 42076 808666 42472 808694
rect 41786 808344 41842 808353
rect 41786 808279 41842 808288
rect 41142 805624 41198 805633
rect 41142 805559 41198 805568
rect 40958 805352 41014 805361
rect 40958 805287 41014 805296
rect 41800 805089 41828 808279
rect 42246 806712 42302 806721
rect 42246 806647 42302 806656
rect 41786 805080 41842 805089
rect 41786 805015 41842 805024
rect 41696 802460 41748 802466
rect 41696 802402 41748 802408
rect 41708 802346 41736 802402
rect 41708 802318 41828 802346
rect 39304 801712 39356 801718
rect 41604 801712 41656 801718
rect 39304 801654 39356 801660
rect 41602 801680 41604 801689
rect 41656 801680 41658 801689
rect 41602 801615 41658 801624
rect 41800 800329 41828 802318
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 806647
rect 42444 804554 42472 808666
rect 42182 798238 42288 798266
rect 42352 804526 42472 804554
rect 42352 797619 42380 804526
rect 42536 804409 42564 808959
rect 42522 804400 42578 804409
rect 42522 804335 42578 804344
rect 42706 801680 42762 801689
rect 42706 801615 42762 801624
rect 42522 799640 42578 799649
rect 42522 799575 42578 799584
rect 42182 797591 42380 797619
rect 42536 796974 42564 799575
rect 42720 799490 42748 801615
rect 42628 799462 42748 799490
rect 42628 797619 42656 799462
rect 42628 797591 42748 797619
rect 42182 796946 42564 796974
rect 42522 796784 42578 796793
rect 42522 796719 42578 796728
rect 41970 796104 42026 796113
rect 41970 796039 42026 796048
rect 42246 796104 42302 796113
rect 42246 796039 42302 796048
rect 41984 795765 42012 796039
rect 42260 794894 42288 796039
rect 42536 794894 42564 796719
rect 42720 794894 42748 797591
rect 42168 794866 42288 794894
rect 42352 794866 42564 794894
rect 42628 794866 42748 794894
rect 42168 794580 42196 794866
rect 42352 794458 42380 794866
rect 42260 794430 42380 794458
rect 42260 794186 42288 794430
rect 42430 794336 42486 794345
rect 42430 794271 42486 794280
rect 42168 794158 42288 794186
rect 42168 793900 42196 794158
rect 42444 793302 42472 794271
rect 42182 793274 42472 793302
rect 42628 792758 42656 794866
rect 42182 792730 42656 792758
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42614 792296 42670 792305
rect 42614 792231 42670 792240
rect 42430 791752 42486 791761
rect 42430 791687 42486 791696
rect 42168 790622 42288 790650
rect 42168 790228 42196 790622
rect 42154 790120 42210 790129
rect 42154 790055 42210 790064
rect 42168 789616 42196 790055
rect 42168 788990 42288 789018
rect 42168 788936 42196 788990
rect 42260 788950 42288 788990
rect 42444 788950 42472 791687
rect 42628 790129 42656 792231
rect 42614 790120 42670 790129
rect 42614 790055 42670 790064
rect 42260 788922 42472 788950
rect 41786 788624 41842 788633
rect 41786 788559 41842 788568
rect 42706 788624 42762 788633
rect 42706 788559 42762 788568
rect 41800 788392 41828 788559
rect 42246 787944 42302 787953
rect 42246 787879 42302 787888
rect 42260 786570 42288 787879
rect 42182 786542 42288 786570
rect 42062 786448 42118 786457
rect 42062 786383 42118 786392
rect 42076 785944 42104 786383
rect 41786 785632 41842 785641
rect 41786 785567 41842 785576
rect 41800 785264 41828 785567
rect 42720 779714 42748 788559
rect 41708 779686 42748 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 772886 35848 773463
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 43088 772449 43116 815215
rect 43258 810384 43314 810393
rect 43258 810319 43314 810328
rect 43272 791761 43300 810319
rect 43442 807664 43498 807673
rect 43442 807599 43498 807608
rect 43456 804554 43484 807599
rect 43456 804526 43576 804554
rect 43258 791752 43314 791761
rect 43258 791687 43314 791696
rect 43074 772440 43130 772449
rect 43074 772375 43130 772384
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768874 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35532 768984
rect 35584 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 39304 769004 39356 769010
rect 35532 768946 35584 768952
rect 35348 768868 35400 768874
rect 35348 768810 35400 768816
rect 35820 768738 35848 768975
rect 39304 768946 39356 768952
rect 35808 768732 35860 768738
rect 35808 768674 35860 768680
rect 35622 768224 35678 768233
rect 35622 768159 35678 768168
rect 31022 767816 31078 767825
rect 31022 767751 31078 767760
rect 31036 759694 31064 767751
rect 35636 767378 35664 768159
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35624 767372 35676 767378
rect 35624 767314 35676 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 31024 759688 31076 759694
rect 31024 759630 31076 759636
rect 35176 758334 35204 766935
rect 35806 763328 35862 763337
rect 35806 763263 35808 763272
rect 35860 763263 35862 763272
rect 35808 763234 35860 763240
rect 36556 759121 36584 767450
rect 37924 763292 37976 763298
rect 37924 763234 37976 763240
rect 36542 759112 36598 759121
rect 36542 759047 36598 759056
rect 35164 758328 35216 758334
rect 35164 758270 35216 758276
rect 37936 757790 37964 763234
rect 37924 757784 37976 757790
rect 39316 757761 39344 768946
rect 40408 768868 40460 768874
rect 40408 768810 40460 768816
rect 40420 763745 40448 768810
rect 40592 768732 40644 768738
rect 40592 768674 40644 768680
rect 40604 764153 40632 768674
rect 41328 767372 41380 767378
rect 41328 767314 41380 767320
rect 41340 765377 41368 767314
rect 42798 766728 42854 766737
rect 42798 766663 42854 766672
rect 41326 765368 41382 765377
rect 41326 765303 41382 765312
rect 42614 765368 42670 765377
rect 42614 765303 42670 765312
rect 42628 765218 42656 765303
rect 42628 765190 42748 765218
rect 40590 764144 40646 764153
rect 40590 764079 40646 764088
rect 42522 764144 42578 764153
rect 42522 764079 42578 764088
rect 40406 763736 40462 763745
rect 40406 763671 40462 763680
rect 42338 763736 42394 763745
rect 42338 763671 42394 763680
rect 41512 759688 41564 759694
rect 41512 759630 41564 759636
rect 40590 758432 40646 758441
rect 40590 758367 40592 758376
rect 40644 758367 40646 758376
rect 40592 758338 40644 758344
rect 41524 758146 41552 759630
rect 42352 758849 42380 763671
rect 42536 763154 42564 764079
rect 42536 763126 42656 763154
rect 42338 758840 42394 758849
rect 42338 758775 42394 758784
rect 42338 758432 42394 758441
rect 42394 758390 42564 758418
rect 42338 758367 42394 758376
rect 41524 758118 42288 758146
rect 41604 757784 41656 757790
rect 37924 757726 37976 757732
rect 39302 757752 39358 757761
rect 41656 757732 41828 757738
rect 41604 757726 41828 757732
rect 41616 757710 41828 757726
rect 39302 757687 39358 757696
rect 41800 757081 41828 757710
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42260 756254 42288 758118
rect 42168 756226 42288 756254
rect 41878 755440 41934 755449
rect 41878 755375 41934 755384
rect 41892 755072 41920 755375
rect 42154 754624 42210 754633
rect 42154 754559 42210 754568
rect 42168 754392 42196 754559
rect 42062 754216 42118 754225
rect 42062 754151 42118 754160
rect 42076 753780 42104 754151
rect 42338 753944 42394 753953
rect 42338 753879 42394 753888
rect 42352 753522 42380 753879
rect 42352 753494 42472 753522
rect 42168 753466 42472 753494
rect 42168 753409 42196 753466
rect 42154 753400 42210 753409
rect 42154 753335 42210 753344
rect 41970 752992 42026 753001
rect 41970 752927 42026 752936
rect 41984 752556 42012 752927
rect 42536 752570 42564 758390
rect 42260 752542 42564 752570
rect 42260 752434 42288 752542
rect 42076 752406 42288 752434
rect 42430 752448 42486 752457
rect 42076 752162 42104 752406
rect 42628 752434 42656 763126
rect 42486 752406 42656 752434
rect 42430 752383 42486 752392
rect 42076 752134 42288 752162
rect 42260 751890 42288 752134
rect 42720 752026 42748 765190
rect 42812 753494 42840 766663
rect 43350 764688 43406 764697
rect 43350 764623 43406 764632
rect 43166 763056 43222 763065
rect 43166 762991 43222 763000
rect 42812 753466 42932 753494
rect 42904 752185 42932 753466
rect 42890 752176 42946 752185
rect 42890 752111 42946 752120
rect 42720 751998 43116 752026
rect 42260 751862 42380 751890
rect 42154 751768 42210 751777
rect 42154 751703 42210 751712
rect 42168 751369 42196 751703
rect 41786 751088 41842 751097
rect 41786 751023 41842 751032
rect 41800 750720 41828 751023
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42154 749728 42210 749737
rect 42154 749663 42210 749672
rect 42168 749529 42196 749663
rect 42062 749184 42118 749193
rect 42118 749142 42288 749170
rect 42062 749119 42118 749128
rect 42260 747062 42288 749142
rect 42182 747034 42288 747062
rect 42154 746872 42210 746881
rect 42154 746807 42210 746816
rect 42168 746401 42196 746807
rect 42352 745770 42380 751862
rect 42890 749728 42946 749737
rect 43088 749714 43116 751998
rect 42946 749686 43116 749714
rect 42890 749663 42946 749672
rect 42182 745742 42380 745770
rect 42154 745512 42210 745521
rect 42154 745447 42210 745456
rect 42168 745212 42196 745447
rect 42706 745240 42762 745249
rect 42536 745198 42706 745226
rect 42338 744968 42394 744977
rect 42338 744903 42394 744912
rect 42352 743730 42380 744903
rect 42168 743702 42380 743730
rect 42168 743376 42196 743702
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42536 742710 42564 745198
rect 42706 745175 42762 745184
rect 42798 744424 42854 744433
rect 42260 742682 42564 742710
rect 42628 744382 42798 744410
rect 42628 742098 42656 744382
rect 42798 744359 42854 744368
rect 42890 742792 42946 742801
rect 42890 742727 42946 742736
rect 42182 742070 42656 742098
rect 42904 734174 42932 742727
rect 43180 736934 43208 762991
rect 43364 753953 43392 764623
rect 43350 753944 43406 753953
rect 43350 753879 43406 753888
rect 42720 734146 42932 734174
rect 43088 736906 43208 736934
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42720 731414 42748 734146
rect 41708 731386 42748 731414
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35820 730114 35848 730895
rect 41708 730114 41736 731386
rect 35808 730108 35860 730114
rect 35808 730050 35860 730056
rect 41696 730108 41748 730114
rect 41696 730050 41748 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41142 726064 41198 726073
rect 41142 725999 41198 726008
rect 33782 725248 33838 725257
rect 33782 725183 33838 725192
rect 31666 724432 31722 724441
rect 31666 724367 31722 724376
rect 31680 715465 31708 724367
rect 33796 715562 33824 725183
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 34518 724024 34574 724033
rect 34518 723959 34574 723968
rect 34532 715698 34560 723959
rect 36556 717398 36584 724775
rect 40682 723208 40738 723217
rect 40682 723143 40738 723152
rect 38750 720352 38806 720361
rect 38750 720287 38806 720296
rect 36544 717392 36596 717398
rect 36544 717334 36596 717340
rect 34520 715692 34572 715698
rect 34520 715634 34572 715640
rect 33784 715556 33836 715562
rect 33784 715498 33836 715504
rect 31666 715456 31722 715465
rect 31666 715391 31722 715400
rect 38764 714241 38792 720287
rect 40314 715728 40370 715737
rect 40314 715663 40370 715672
rect 40328 715562 40356 715663
rect 40316 715556 40368 715562
rect 40316 715498 40368 715504
rect 40696 714241 40724 723143
rect 41156 721777 41184 725999
rect 41340 725966 41368 726407
rect 41328 725960 41380 725966
rect 41328 725902 41380 725908
rect 41696 725960 41748 725966
rect 41748 725908 42012 725914
rect 41696 725902 42012 725908
rect 41708 725886 42012 725902
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724538 41368 725591
rect 41328 724532 41380 724538
rect 41328 724474 41380 724480
rect 41696 724532 41748 724538
rect 41696 724474 41748 724480
rect 41142 721768 41198 721777
rect 41708 721754 41736 724474
rect 41984 721754 42012 725886
rect 41708 721726 41920 721754
rect 41984 721726 42656 721754
rect 41142 721703 41198 721712
rect 41420 717392 41472 717398
rect 41420 717334 41472 717340
rect 41432 714241 41460 717334
rect 41696 715692 41748 715698
rect 41696 715634 41748 715640
rect 41708 715193 41736 715634
rect 41694 715184 41750 715193
rect 41694 715119 41750 715128
rect 41892 714649 41920 721726
rect 42062 715728 42118 715737
rect 42062 715663 42118 715672
rect 41878 714640 41934 714649
rect 41878 714575 41934 714584
rect 42076 714377 42104 715663
rect 42628 715306 42656 721726
rect 42628 715278 42932 715306
rect 42706 715184 42762 715193
rect 42706 715119 42762 715128
rect 42430 714640 42486 714649
rect 42430 714575 42486 714584
rect 42062 714368 42118 714377
rect 42062 714303 42118 714312
rect 38750 714232 38806 714241
rect 38750 714167 38806 714176
rect 40682 714232 40738 714241
rect 40682 714167 40738 714176
rect 41418 714232 41474 714241
rect 41418 714167 41474 714176
rect 41786 713552 41842 713561
rect 41786 713487 41842 713496
rect 41800 713048 41828 713487
rect 42246 713280 42302 713289
rect 42246 713215 42302 713224
rect 41786 712192 41842 712201
rect 41786 712127 41842 712136
rect 41800 711824 41828 712127
rect 42260 711226 42288 713215
rect 42182 711198 42288 711226
rect 42246 711104 42302 711113
rect 42246 711039 42302 711048
rect 42260 710682 42288 711039
rect 42168 710654 42288 710682
rect 42168 710561 42196 710654
rect 42444 710575 42472 714575
rect 42720 714105 42748 715119
rect 42706 714096 42762 714105
rect 42706 714031 42762 714040
rect 42614 713280 42670 713289
rect 42904 713266 42932 715278
rect 42670 713238 42932 713266
rect 42614 713215 42670 713224
rect 42444 710547 42564 710575
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 42062 709064 42118 709073
rect 42118 709022 42288 709050
rect 42062 708999 42118 709008
rect 41786 708520 41842 708529
rect 41786 708455 41842 708464
rect 41800 708152 41828 708455
rect 42062 707840 42118 707849
rect 42062 707775 42118 707784
rect 42076 707540 42104 707775
rect 42260 707418 42288 709022
rect 42168 707390 42288 707418
rect 42168 706860 42196 707390
rect 42246 706752 42302 706761
rect 42246 706687 42302 706696
rect 42260 706602 42288 706687
rect 42260 706574 42380 706602
rect 41970 706480 42026 706489
rect 41970 706415 42026 706424
rect 41984 706316 42012 706415
rect 42352 706194 42380 706574
rect 42352 706166 42472 706194
rect 42246 705256 42302 705265
rect 42246 705191 42302 705200
rect 42260 704585 42288 705191
rect 42246 704576 42302 704585
rect 42246 704511 42302 704520
rect 42444 704018 42472 706166
rect 42076 703990 42472 704018
rect 42076 703868 42104 703990
rect 42154 703488 42210 703497
rect 42154 703423 42210 703432
rect 42168 703188 42196 703423
rect 42536 703066 42564 710547
rect 42706 710016 42762 710025
rect 42706 709951 42762 709960
rect 42444 703038 42564 703066
rect 42062 702808 42118 702817
rect 42062 702743 42118 702752
rect 42076 702576 42104 702743
rect 42168 701978 42196 702032
rect 42444 701978 42472 703038
rect 42720 702817 42748 709951
rect 42706 702808 42762 702817
rect 42706 702743 42762 702752
rect 42614 702400 42670 702409
rect 42614 702335 42670 702344
rect 42168 701950 42472 701978
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 41786 699816 41842 699825
rect 41786 699751 41842 699760
rect 41800 699516 41828 699751
rect 42628 698918 42656 702335
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 41418 689344 41474 689353
rect 41418 689279 41474 689288
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35622 687304 35678 687313
rect 35820 687274 35848 687647
rect 41432 687274 41460 689279
rect 35622 687239 35678 687248
rect 35808 687268 35860 687274
rect 35808 687210 35860 687216
rect 41420 687268 41472 687274
rect 41420 687210 41472 687216
rect 35806 683632 35862 683641
rect 35806 683567 35862 683576
rect 35820 683398 35848 683567
rect 35808 683392 35860 683398
rect 35808 683334 35860 683340
rect 41512 683324 41564 683330
rect 41512 683266 41564 683272
rect 35806 683224 35862 683233
rect 35806 683159 35808 683168
rect 35860 683159 35862 683168
rect 35808 683130 35860 683136
rect 35438 682816 35494 682825
rect 35438 682751 35494 682760
rect 35452 681766 35480 682751
rect 35622 682408 35678 682417
rect 35622 682343 35678 682352
rect 35636 681902 35664 682343
rect 35808 682032 35860 682038
rect 35806 682000 35808 682009
rect 36544 682032 36596 682038
rect 35860 682000 35862 682009
rect 36544 681974 36596 681980
rect 35806 681935 35862 681944
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35440 681760 35492 681766
rect 35440 681702 35492 681708
rect 32402 681592 32458 681601
rect 32402 681527 32458 681536
rect 31022 681184 31078 681193
rect 31022 681119 31078 681128
rect 31036 671401 31064 681119
rect 32416 672790 32444 681527
rect 35622 680776 35678 680785
rect 35622 680711 35678 680720
rect 35636 674150 35664 680711
rect 35624 674144 35676 674150
rect 35624 674086 35676 674092
rect 36556 673198 36584 681974
rect 40960 681760 41012 681766
rect 40960 681702 41012 681708
rect 37186 677104 37242 677113
rect 37186 677039 37242 677048
rect 36544 673192 36596 673198
rect 36544 673134 36596 673140
rect 32404 672784 32456 672790
rect 32404 672726 32456 672732
rect 31022 671392 31078 671401
rect 31022 671327 31078 671336
rect 37200 671022 37228 677039
rect 40972 676025 41000 681702
rect 41524 677634 41552 683266
rect 41696 683188 41748 683194
rect 41696 683130 41748 683136
rect 41708 681986 41736 683130
rect 41708 681958 42012 681986
rect 41696 681896 41748 681902
rect 41694 681864 41696 681873
rect 41748 681864 41750 681873
rect 41694 681799 41750 681808
rect 41984 681714 42012 681958
rect 42614 681864 42670 681873
rect 42614 681799 42670 681808
rect 41984 681686 42564 681714
rect 41786 677648 41842 677657
rect 41524 677606 41786 677634
rect 41786 677583 41842 677592
rect 40958 676016 41014 676025
rect 40958 675951 41014 675960
rect 39672 674144 39724 674150
rect 39672 674086 39724 674092
rect 39684 671945 39712 674086
rect 42536 673577 42564 681686
rect 42628 678974 42656 681799
rect 42890 679960 42946 679969
rect 42890 679895 42946 679904
rect 42904 678974 42932 679895
rect 42628 678946 42748 678974
rect 42904 678946 43024 678974
rect 42522 673568 42578 673577
rect 42522 673503 42578 673512
rect 40592 673192 40644 673198
rect 40590 673160 40592 673169
rect 40644 673160 40646 673169
rect 40590 673095 40646 673104
rect 42338 673160 42394 673169
rect 42394 673118 42656 673146
rect 42338 673095 42394 673104
rect 41696 672784 41748 672790
rect 41748 672732 41920 672738
rect 41696 672726 41920 672732
rect 41708 672710 41920 672726
rect 39670 671936 39726 671945
rect 39670 671871 39726 671880
rect 37188 671016 37240 671022
rect 40132 671016 40184 671022
rect 37188 670958 37240 670964
rect 40130 670984 40132 670993
rect 40184 670984 40186 670993
rect 40130 670919 40186 670928
rect 41892 670834 41920 672710
rect 42338 671936 42394 671945
rect 42394 671894 42564 671922
rect 42338 671871 42394 671880
rect 42154 670984 42210 670993
rect 42210 670942 42380 670970
rect 42154 670919 42210 670928
rect 41892 670806 42288 670834
rect 42168 669746 42196 669868
rect 42260 669746 42288 670806
rect 42168 669718 42288 669746
rect 42352 668658 42380 670942
rect 42182 668630 42380 668658
rect 42062 668264 42118 668273
rect 42062 668199 42118 668208
rect 42076 668032 42104 668199
rect 42246 667856 42302 667865
rect 42246 667791 42302 667800
rect 42260 667366 42288 667791
rect 42182 667338 42288 667366
rect 42246 667040 42302 667049
rect 42246 666975 42302 666984
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 41786 665408 41842 665417
rect 41786 665343 41842 665352
rect 41800 664972 41828 665343
rect 42260 664339 42288 666975
rect 42536 666554 42564 671894
rect 42182 664311 42288 664339
rect 42352 666526 42564 666554
rect 41786 664184 41842 664193
rect 41786 664119 41842 664128
rect 41800 663680 41828 664119
rect 42352 663377 42380 666526
rect 42338 663368 42394 663377
rect 42338 663303 42394 663312
rect 42628 663150 42656 673118
rect 42720 668046 42748 678946
rect 42996 669314 43024 678946
rect 42904 669286 43024 669314
rect 42720 668018 42840 668046
rect 42812 667842 42840 668018
rect 42182 663122 42656 663150
rect 42720 667814 42840 667842
rect 42430 662960 42486 662969
rect 42430 662895 42486 662904
rect 42062 662824 42118 662833
rect 42118 662782 42288 662810
rect 42062 662759 42118 662768
rect 42260 661042 42288 662782
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42444 660022 42472 662895
rect 42182 659994 42472 660022
rect 42154 659832 42210 659841
rect 42154 659767 42210 659776
rect 42168 659357 42196 659767
rect 42720 659025 42748 667814
rect 42904 666641 42932 669286
rect 42890 666632 42946 666641
rect 42890 666567 42946 666576
rect 42154 659016 42210 659025
rect 42154 658951 42210 658960
rect 42706 659016 42762 659025
rect 42706 658951 42762 658960
rect 42168 658784 42196 658951
rect 42614 658608 42670 658617
rect 42614 658543 42670 658552
rect 42430 658336 42486 658345
rect 42430 658271 42486 658280
rect 41970 657384 42026 657393
rect 41970 657319 42026 657328
rect 41984 656948 42012 657319
rect 42444 656350 42472 658271
rect 42182 656322 42472 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42628 655670 42656 658543
rect 42260 655642 42656 655670
rect 42614 655480 42670 655489
rect 42614 655415 42670 655424
rect 42628 654134 42656 655415
rect 41708 654106 42656 654134
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35820 644502 35848 644671
rect 41708 644502 41736 654106
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 41696 644496 41748 644502
rect 41696 644438 41748 644444
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35346 639840 35402 639849
rect 35346 639775 35402 639784
rect 35360 639130 35388 639775
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35348 639124 35400 639130
rect 35348 639066 35400 639072
rect 35544 638994 35572 639367
rect 35820 639266 35848 639367
rect 35808 639260 35860 639266
rect 35808 639202 35860 639208
rect 40040 639260 40092 639266
rect 40040 639202 40092 639208
rect 35532 638988 35584 638994
rect 35532 638930 35584 638936
rect 36544 638988 36596 638994
rect 36544 638930 36596 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 33782 638208 33838 638217
rect 33782 638143 33838 638152
rect 33796 629950 33824 638143
rect 35820 637634 35848 638551
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 36556 630737 36584 638930
rect 40052 638625 40080 639202
rect 41696 639124 41748 639130
rect 41696 639066 41748 639072
rect 41708 639010 41736 639066
rect 41708 638982 42012 639010
rect 40038 638616 40094 638625
rect 40038 638551 40094 638560
rect 41786 638208 41842 638217
rect 41786 638143 41842 638152
rect 41328 637628 41380 637634
rect 41800 637605 41828 638143
rect 41328 637570 41380 637576
rect 41786 637596 41842 637605
rect 41340 634814 41368 637570
rect 41786 637531 41842 637540
rect 41340 634786 41460 634814
rect 36542 630728 36598 630737
rect 36542 630663 36598 630672
rect 41432 630057 41460 634786
rect 41418 630048 41474 630057
rect 41984 630034 42012 638982
rect 42890 636304 42946 636313
rect 42890 636239 42946 636248
rect 42522 633856 42578 633865
rect 42522 633791 42578 633800
rect 41984 630006 42472 630034
rect 41418 629983 41474 629992
rect 33784 629944 33836 629950
rect 33784 629886 33836 629892
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42444 625954 42472 630006
rect 42260 625926 42472 625954
rect 42062 625832 42118 625841
rect 42062 625767 42118 625776
rect 42076 625464 42104 625767
rect 42260 625546 42288 625926
rect 42536 625841 42564 633791
rect 42706 630048 42762 630057
rect 42706 629983 42762 629992
rect 42522 625832 42578 625841
rect 42522 625767 42578 625776
rect 42260 625518 42472 625546
rect 42168 624838 42288 624866
rect 42168 624784 42196 624838
rect 42260 624798 42288 624838
rect 42444 624798 42472 625518
rect 42260 624770 42472 624798
rect 42430 624200 42486 624209
rect 42182 624158 42430 624186
rect 42430 624135 42486 624144
rect 42720 623914 42748 629983
rect 42904 625154 42932 636239
rect 42628 623886 42748 623914
rect 42812 625126 42932 625154
rect 42246 623792 42302 623801
rect 42246 623727 42302 623736
rect 42430 623792 42486 623801
rect 42430 623727 42486 623736
rect 42260 623642 42288 623727
rect 42260 623614 42380 623642
rect 42062 623384 42118 623393
rect 42062 623319 42118 623328
rect 42076 622948 42104 623319
rect 42352 621806 42380 623614
rect 42168 621738 42196 621792
rect 42260 621778 42380 621806
rect 42260 621738 42288 621778
rect 42168 621710 42288 621738
rect 42444 621330 42472 623727
rect 42260 621302 42472 621330
rect 42260 621126 42288 621302
rect 42182 621098 42288 621126
rect 42062 620936 42118 620945
rect 42062 620871 42118 620880
rect 42076 620500 42104 620871
rect 42628 620242 42656 623886
rect 42812 623801 42840 625126
rect 42798 623792 42854 623801
rect 42798 623727 42854 623736
rect 42076 620214 42656 620242
rect 42076 619956 42104 620214
rect 42246 620120 42302 620129
rect 42246 620055 42302 620064
rect 42260 617454 42288 620055
rect 42706 619848 42762 619857
rect 42706 619783 42762 619792
rect 42522 619576 42578 619585
rect 42522 619511 42578 619520
rect 42536 618882 42564 619511
rect 42352 618854 42564 618882
rect 42352 618254 42380 618854
rect 42522 618760 42578 618769
rect 42522 618695 42578 618704
rect 42352 618226 42472 618254
rect 42182 617426 42288 617454
rect 42444 616842 42472 618226
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42536 616434 42564 618695
rect 42352 616406 42564 616434
rect 42352 616162 42380 616406
rect 42182 616134 42380 616162
rect 42430 616040 42486 616049
rect 42430 615975 42486 615984
rect 41786 615768 41842 615777
rect 41786 615703 41842 615712
rect 41800 615604 41828 615703
rect 42444 614122 42472 615975
rect 42168 614094 42472 614122
rect 42168 613768 42196 614094
rect 42154 613592 42210 613601
rect 42154 613527 42210 613536
rect 42168 613121 42196 613527
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 42720 610722 42748 619783
rect 43088 612377 43116 736906
rect 43350 633448 43406 633457
rect 43350 633383 43406 633392
rect 43074 612368 43130 612377
rect 43074 612303 43130 612312
rect 43364 611017 43392 633383
rect 43548 621014 43576 804526
rect 43456 620986 43576 621014
rect 43456 612626 43484 620986
rect 43640 612746 43668 933263
rect 43810 932104 43866 932113
rect 43810 932039 43866 932048
rect 43628 612740 43680 612746
rect 43628 612682 43680 612688
rect 43824 612678 43852 932039
rect 44086 892800 44142 892809
rect 44086 892735 44088 892744
rect 44140 892735 44142 892744
rect 44088 892706 44140 892712
rect 44086 892528 44142 892537
rect 44086 892463 44142 892472
rect 44100 891886 44128 892463
rect 44088 891880 44140 891886
rect 44088 891822 44140 891828
rect 44468 815697 44496 941015
rect 44652 935377 44680 964679
rect 44836 941497 44864 990082
rect 46296 946008 46348 946014
rect 46296 945950 46348 945956
rect 46308 943537 46336 945950
rect 46294 943528 46350 943537
rect 46294 943463 46350 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44638 935368 44694 935377
rect 44638 935303 44694 935312
rect 47596 891993 47624 991714
rect 48964 991636 49016 991642
rect 48964 991578 49016 991584
rect 48976 942313 49004 991578
rect 48962 942304 49018 942313
rect 48962 942239 49018 942248
rect 50356 940681 50384 993006
rect 50342 940672 50398 940681
rect 50342 940607 50398 940616
rect 51736 939865 51764 993142
rect 55864 992928 55916 992934
rect 55864 992870 55916 992876
rect 54484 991500 54536 991506
rect 54484 991442 54536 991448
rect 53288 988780 53340 988786
rect 53288 988722 53340 988728
rect 51722 939856 51778 939865
rect 51722 939791 51778 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44914 816096 44970 816105
rect 44914 816031 44970 816040
rect 44454 815688 44510 815697
rect 44454 815623 44510 815632
rect 44638 814464 44694 814473
rect 44638 814399 44694 814408
rect 44178 807936 44234 807945
rect 44178 807871 44234 807880
rect 43994 806304 44050 806313
rect 43994 806239 44050 806248
rect 43812 612672 43864 612678
rect 43456 612598 43622 612626
rect 43812 612614 43864 612620
rect 43594 612338 43622 612598
rect 44008 612542 44036 806239
rect 44192 796385 44220 807871
rect 44178 796376 44234 796385
rect 44178 796311 44234 796320
rect 44178 772848 44234 772857
rect 44178 772783 44234 772792
rect 44192 730153 44220 772783
rect 44454 772032 44510 772041
rect 44454 771967 44510 771976
rect 44178 730144 44234 730153
rect 44178 730079 44234 730088
rect 44270 729736 44326 729745
rect 44270 729671 44326 729680
rect 44284 728634 44312 729671
rect 44468 729337 44496 771967
rect 44652 771633 44680 814399
rect 44928 810642 44956 816031
rect 45466 813648 45522 813657
rect 45466 813583 45522 813592
rect 45098 810792 45154 810801
rect 45098 810727 45154 810736
rect 44928 810614 45048 810642
rect 44822 809568 44878 809577
rect 44822 809503 44878 809512
rect 44836 797745 44864 809503
rect 44822 797736 44878 797745
rect 44822 797671 44878 797680
rect 44824 793620 44876 793626
rect 44824 793562 44876 793568
rect 44638 771624 44694 771633
rect 44638 771559 44694 771568
rect 44638 771216 44694 771225
rect 44638 771151 44694 771160
rect 44454 729328 44510 729337
rect 44454 729263 44510 729272
rect 44284 728606 44404 728634
rect 44178 722800 44234 722809
rect 44178 722735 44234 722744
rect 44192 707849 44220 722735
rect 44178 707840 44234 707849
rect 44178 707775 44234 707784
rect 44376 686905 44404 728606
rect 44652 728521 44680 771151
rect 44836 731377 44864 793562
rect 45020 773265 45048 810614
rect 45112 808694 45140 810727
rect 45282 809976 45338 809985
rect 45282 809911 45338 809920
rect 45296 808694 45324 809911
rect 45112 808666 45232 808694
rect 45296 808666 45416 808694
rect 45204 794894 45232 808666
rect 45388 794894 45416 808666
rect 45112 794866 45232 794894
rect 45296 794866 45416 794894
rect 45112 792134 45140 794866
rect 45296 792305 45324 794866
rect 45282 792296 45338 792305
rect 45282 792231 45338 792240
rect 45112 792106 45232 792134
rect 45204 786457 45232 792106
rect 45190 786448 45246 786457
rect 45190 786383 45246 786392
rect 45006 773256 45062 773265
rect 45006 773191 45062 773200
rect 45480 770817 45508 813583
rect 45466 770808 45522 770817
rect 45466 770743 45522 770752
rect 45006 770400 45062 770409
rect 45006 770335 45062 770344
rect 44822 731368 44878 731377
rect 44822 731303 44878 731312
rect 44638 728512 44694 728521
rect 44638 728447 44694 728456
rect 44822 728104 44878 728113
rect 44822 728039 44878 728048
rect 44638 727288 44694 727297
rect 44638 727223 44694 727232
rect 44362 686896 44418 686905
rect 44362 686831 44418 686840
rect 44362 686488 44418 686497
rect 44362 686423 44418 686432
rect 44178 684856 44234 684865
rect 44178 684791 44234 684800
rect 44192 642297 44220 684791
rect 44376 643657 44404 686423
rect 44652 684457 44680 727223
rect 44836 685273 44864 728039
rect 45020 727705 45048 770335
rect 45190 766320 45246 766329
rect 45190 766255 45246 766264
rect 45204 754905 45232 766255
rect 45190 754896 45246 754905
rect 45190 754831 45246 754840
rect 46216 754225 46244 870810
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 46938 764416 46994 764425
rect 46938 764351 46994 764360
rect 46202 754216 46258 754225
rect 46202 754151 46258 754160
rect 45190 728920 45246 728929
rect 45190 728855 45246 728864
rect 45006 727696 45062 727705
rect 45006 727631 45062 727640
rect 45006 723616 45062 723625
rect 45006 723551 45062 723560
rect 45020 705265 45048 723551
rect 45006 705256 45062 705265
rect 45006 705191 45062 705200
rect 45204 686089 45232 728855
rect 45558 721168 45614 721177
rect 45558 721103 45614 721112
rect 45190 686080 45246 686089
rect 45190 686015 45246 686024
rect 45190 685672 45246 685681
rect 45190 685607 45246 685616
rect 44822 685264 44878 685273
rect 44822 685199 44878 685208
rect 44638 684448 44694 684457
rect 44638 684383 44694 684392
rect 45006 684040 45062 684049
rect 45006 683975 45062 683984
rect 44546 680368 44602 680377
rect 44546 680303 44602 680312
rect 44560 662969 44588 680303
rect 44730 679552 44786 679561
rect 44730 679487 44786 679496
rect 44744 667049 44772 679487
rect 44730 667040 44786 667049
rect 44730 666975 44786 666984
rect 44546 662960 44602 662969
rect 44546 662895 44602 662904
rect 44362 643648 44418 643657
rect 44362 643583 44418 643592
rect 44822 643376 44878 643385
rect 44822 643311 44878 643320
rect 44638 642560 44694 642569
rect 44638 642495 44694 642504
rect 44178 642288 44234 642297
rect 44178 642223 44234 642232
rect 44270 636576 44326 636585
rect 44270 636511 44326 636520
rect 44284 623393 44312 636511
rect 44454 635760 44510 635769
rect 44454 635695 44510 635704
rect 44270 623384 44326 623393
rect 44270 623319 44326 623328
rect 44468 620129 44496 635695
rect 44454 620120 44510 620129
rect 44454 620055 44510 620064
rect 43996 612536 44048 612542
rect 43996 612478 44048 612484
rect 43718 612368 43774 612377
rect 43582 612332 43634 612338
rect 43718 612303 43720 612312
rect 43582 612274 43634 612280
rect 43772 612303 43774 612312
rect 43720 612274 43772 612280
rect 43350 611008 43406 611017
rect 43350 610943 43406 610952
rect 44086 611008 44142 611017
rect 44086 610943 44142 610952
rect 44270 611008 44326 611017
rect 44270 610943 44272 610952
rect 44100 610858 44128 610943
rect 44324 610943 44326 610952
rect 44272 610914 44324 610920
rect 44100 610842 44419 610858
rect 44100 610836 44431 610842
rect 44100 610830 44379 610836
rect 44379 610778 44431 610784
rect 44502 610768 44554 610774
rect 42720 610716 44502 610722
rect 42720 610710 44554 610716
rect 42720 610694 44542 610710
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 44652 599729 44680 642495
rect 44836 600545 44864 643311
rect 45020 641481 45048 683975
rect 45204 643113 45232 685607
rect 45190 643104 45246 643113
rect 45190 643039 45246 643048
rect 45006 641472 45062 641481
rect 45006 641407 45062 641416
rect 45374 641200 45430 641209
rect 45374 641135 45430 641144
rect 45190 640928 45246 640937
rect 45190 640863 45246 640872
rect 45006 635352 45062 635361
rect 45006 635287 45062 635296
rect 45020 620945 45048 635287
rect 45006 620936 45062 620945
rect 45006 620871 45062 620880
rect 44822 600536 44878 600545
rect 44822 600471 44878 600480
rect 44822 600128 44878 600137
rect 44822 600063 44878 600072
rect 44638 599720 44694 599729
rect 44638 599655 44694 599664
rect 44638 598496 44694 598505
rect 44638 598431 44694 598440
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 41326 596864 41382 596873
rect 41326 596799 41382 596808
rect 41340 596086 41368 596799
rect 41328 596080 41380 596086
rect 41142 596048 41198 596057
rect 41328 596022 41380 596028
rect 41604 596080 41656 596086
rect 41604 596022 41656 596028
rect 41142 595983 41198 595992
rect 33046 595640 33102 595649
rect 33046 595575 33102 595584
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595575
rect 35162 595232 35218 595241
rect 35162 595167 35218 595176
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 35176 585954 35204 595167
rect 40682 594824 40738 594833
rect 41156 594794 41184 595983
rect 41616 595898 41644 596022
rect 41616 595870 42104 595898
rect 40682 594759 40738 594768
rect 41144 594788 41196 594794
rect 40500 592340 40552 592346
rect 40500 592282 40552 592288
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 585993 39988 590679
rect 40512 589665 40540 592282
rect 40498 589656 40554 589665
rect 40498 589591 40554 589600
rect 40132 587172 40184 587178
rect 40132 587114 40184 587120
rect 39946 585984 40002 585993
rect 35164 585948 35216 585954
rect 39946 585919 40002 585928
rect 35164 585890 35216 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 39396 585812 39448 585818
rect 39396 585754 39448 585760
rect 39408 584633 39436 585754
rect 40144 584905 40172 587114
rect 40130 584896 40186 584905
rect 40130 584831 40186 584840
rect 40696 584633 40724 594759
rect 41144 594730 41196 594736
rect 41696 594788 41748 594794
rect 41696 594730 41748 594736
rect 41708 594561 41736 594730
rect 41694 594552 41750 594561
rect 41694 594487 41750 594496
rect 41786 593600 41842 593609
rect 41616 593558 41786 593586
rect 41616 593298 41644 593558
rect 41786 593535 41842 593544
rect 40868 593292 40920 593298
rect 40868 593234 40920 593240
rect 41604 593292 41656 593298
rect 41604 593234 41656 593240
rect 39394 584624 39450 584633
rect 39394 584559 39450 584568
rect 40682 584624 40738 584633
rect 40880 584594 40908 593234
rect 41786 593192 41842 593201
rect 41432 593150 41786 593178
rect 41432 589529 41460 593150
rect 41786 593127 41842 593136
rect 41786 592784 41842 592793
rect 41616 592742 41786 592770
rect 41616 592346 41644 592742
rect 41786 592719 41842 592728
rect 41878 592376 41934 592385
rect 41604 592340 41656 592346
rect 41878 592311 41934 592320
rect 41604 592282 41656 592288
rect 41418 589520 41474 589529
rect 41418 589455 41474 589464
rect 41892 589393 41920 592311
rect 42076 592034 42104 595870
rect 42522 594552 42578 594561
rect 42522 594487 42578 594496
rect 42536 592034 42564 594487
rect 42798 594008 42854 594017
rect 42798 593943 42854 593952
rect 42812 593858 42840 593943
rect 42812 593830 42932 593858
rect 42076 592006 42196 592034
rect 41878 589384 41934 589393
rect 41878 589319 41934 589328
rect 42168 589274 42196 592006
rect 42444 592006 42564 592034
rect 42444 589274 42472 592006
rect 42168 589246 42380 589274
rect 42444 589246 42840 589274
rect 42352 586378 42380 589246
rect 42352 586350 42564 586378
rect 42338 585984 42394 585993
rect 41696 585948 41748 585954
rect 42338 585919 42394 585928
rect 41696 585890 41748 585896
rect 41708 585834 41736 585890
rect 41708 585806 42288 585834
rect 40682 584559 40738 584568
rect 40868 584588 40920 584594
rect 40868 584530 40920 584536
rect 41604 584588 41656 584594
rect 41604 584530 41656 584536
rect 41616 584474 41644 584530
rect 41616 584446 41828 584474
rect 41800 584361 41828 584446
rect 41786 584352 41842 584361
rect 41786 584287 41842 584296
rect 42260 583454 42288 585806
rect 42182 583426 42288 583454
rect 42352 583250 42380 585919
rect 42260 583222 42380 583250
rect 42260 582263 42288 583222
rect 42182 582235 42288 582263
rect 42536 582162 42564 586350
rect 42168 582134 42564 582162
rect 42168 581604 42196 582134
rect 42430 582040 42486 582049
rect 42430 581975 42486 581984
rect 41984 580825 42012 580961
rect 41970 580816 42026 580825
rect 41970 580751 42026 580760
rect 42246 580816 42302 580825
rect 42246 580751 42302 580760
rect 41970 580272 42026 580281
rect 41970 580207 42026 580216
rect 41984 579768 42012 580207
rect 42260 578626 42288 580751
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 41786 578232 41842 578241
rect 41786 578167 41842 578176
rect 41800 577932 41828 578167
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42444 577130 42472 581975
rect 42812 581618 42840 589246
rect 42628 581590 42840 581618
rect 42628 581482 42656 581590
rect 42260 577102 42472 577130
rect 42536 581454 42656 581482
rect 42260 576994 42288 577102
rect 42168 576966 42288 576994
rect 42168 576708 42196 576966
rect 42338 576736 42394 576745
rect 42338 576671 42394 576680
rect 42062 576600 42118 576609
rect 42118 576558 42288 576586
rect 42062 576535 42118 576544
rect 42260 574274 42288 576558
rect 42182 574246 42288 574274
rect 42154 573880 42210 573889
rect 42154 573815 42210 573824
rect 42168 573580 42196 573815
rect 42352 572982 42380 576671
rect 42536 576042 42564 581454
rect 42706 581360 42762 581369
rect 42706 581295 42762 581304
rect 42720 576745 42748 581295
rect 42706 576736 42762 576745
rect 42706 576671 42762 576680
rect 42182 572954 42380 572982
rect 42444 576014 42564 576042
rect 42444 572438 42472 576014
rect 42904 575634 42932 593830
rect 42720 575606 42932 575634
rect 42720 573889 42748 575606
rect 42706 573880 42762 573889
rect 42706 573815 42762 573824
rect 42614 573336 42670 573345
rect 42614 573271 42670 573280
rect 42168 572370 42196 572424
rect 42260 572410 42472 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42628 572234 42656 573271
rect 42352 572206 42656 572234
rect 42352 571010 42380 572206
rect 42522 572112 42578 572121
rect 42522 572047 42578 572056
rect 42076 570982 42380 571010
rect 42076 570588 42104 570982
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42536 569514 42564 572047
rect 42076 569486 42564 569514
rect 42076 569296 42104 569486
rect 42338 569256 42394 569265
rect 42338 569191 42394 569200
rect 42352 567194 42380 569191
rect 41524 567166 42380 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41326 558104 41382 558113
rect 41326 558039 41382 558048
rect 41340 557598 41368 558039
rect 41524 557598 41552 567166
rect 41328 557592 41380 557598
rect 41328 557534 41380 557540
rect 41512 557592 41564 557598
rect 41512 557534 41564 557540
rect 41326 554840 41382 554849
rect 41326 554775 41328 554784
rect 41380 554775 41382 554784
rect 41696 554804 41748 554810
rect 41328 554746 41380 554752
rect 42996 554792 43024 596935
rect 44178 591968 44234 591977
rect 44178 591903 44234 591912
rect 43442 590336 43498 590345
rect 43442 590271 43498 590280
rect 41748 554764 43024 554792
rect 41696 554746 41748 554752
rect 41234 553408 41290 553417
rect 40972 553366 41234 553394
rect 32402 551984 32458 551993
rect 32402 551919 32458 551928
rect 31758 548142 31814 548151
rect 31758 548077 31814 548086
rect 31772 547874 31800 548077
rect 31760 547868 31812 547874
rect 31760 547810 31812 547816
rect 32416 543046 32444 551919
rect 40972 550610 41000 553366
rect 41234 553343 41290 553352
rect 41142 552800 41198 552809
rect 41142 552735 41198 552744
rect 41156 552158 41184 552735
rect 42890 552392 42946 552401
rect 42890 552327 42946 552336
rect 41144 552152 41196 552158
rect 41144 552094 41196 552100
rect 41604 552152 41656 552158
rect 41604 552094 41656 552100
rect 41616 551970 41644 552094
rect 41786 551984 41842 551993
rect 41616 551942 41786 551970
rect 41786 551919 41842 551928
rect 41786 551168 41842 551177
rect 41786 551103 41842 551112
rect 41800 550634 41828 551103
rect 40972 550582 41460 550610
rect 40774 550352 40830 550361
rect 40774 550287 40830 550296
rect 40592 549432 40644 549438
rect 40592 549374 40644 549380
rect 38292 547868 38344 547874
rect 38292 547810 38344 547816
rect 32404 543040 32456 543046
rect 32404 542982 32456 542988
rect 38304 542366 38332 547810
rect 40604 545465 40632 549374
rect 40788 545737 40816 550287
rect 41234 549536 41290 549545
rect 41234 549471 41290 549480
rect 41248 549302 41276 549471
rect 41236 549296 41288 549302
rect 41236 549238 41288 549244
rect 41234 548142 41290 548151
rect 41234 548077 41290 548086
rect 40774 545728 40830 545737
rect 40774 545663 40830 545672
rect 40590 545456 40646 545465
rect 40590 545391 40646 545400
rect 41432 543734 41460 550582
rect 41708 550606 41828 550634
rect 41708 550202 41736 550606
rect 41878 550216 41934 550225
rect 41708 550174 41878 550202
rect 41878 550151 41934 550160
rect 41786 549944 41842 549953
rect 41616 549902 41786 549930
rect 41616 549438 41644 549902
rect 41786 549879 41842 549888
rect 41604 549432 41656 549438
rect 41604 549374 41656 549380
rect 41696 549296 41748 549302
rect 41748 549256 42840 549284
rect 41696 549238 41748 549244
rect 41694 548176 41750 548185
rect 41694 548111 41696 548120
rect 41748 548111 41750 548120
rect 41696 548082 41748 548088
rect 41432 543706 42472 543734
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 38292 542360 38344 542366
rect 38292 542302 38344 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538438 42472 543706
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42168 538370 42196 538424
rect 42260 538410 42472 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42168 537798 42288 537826
rect 42168 537744 42196 537798
rect 42260 537758 42288 537798
rect 42628 537758 42656 540223
rect 42260 537730 42656 537758
rect 42522 537432 42578 537441
rect 42522 537367 42578 537376
rect 41786 537024 41842 537033
rect 41786 536959 41842 536968
rect 42062 537024 42118 537033
rect 42062 536959 42118 536968
rect 41800 536588 41828 536959
rect 42076 536874 42104 536959
rect 42076 536846 42288 536874
rect 42260 535378 42288 536846
rect 42182 535350 42288 535378
rect 41786 535256 41842 535265
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42536 534290 42564 537367
rect 42812 535650 42840 549256
rect 42352 534262 42564 534290
rect 42628 535622 42840 535650
rect 42352 534086 42380 534262
rect 42182 534058 42380 534086
rect 42154 533896 42210 533905
rect 42154 533831 42210 533840
rect 42168 533528 42196 533831
rect 42628 532794 42656 535622
rect 42904 534177 42932 552327
rect 43074 550216 43130 550225
rect 43074 550151 43130 550160
rect 42890 534168 42946 534177
rect 42890 534103 42946 534112
rect 43088 534074 43116 550151
rect 42352 532766 42656 532794
rect 42996 534046 43116 534074
rect 42352 531314 42380 532766
rect 42522 532672 42578 532681
rect 42522 532607 42578 532616
rect 42168 531286 42380 531314
rect 42168 531045 42196 531286
rect 42536 531026 42564 532607
rect 42996 531434 43024 534046
rect 42352 530998 42564 531026
rect 42720 531406 43024 531434
rect 42352 530890 42380 530998
rect 42260 530862 42380 530890
rect 42260 530414 42288 530862
rect 42182 530386 42288 530414
rect 42720 529938 42748 531406
rect 42260 529910 42748 529938
rect 42260 529771 42288 529910
rect 42182 529743 42288 529771
rect 42430 529816 42486 529825
rect 42430 529751 42486 529760
rect 42246 529544 42302 529553
rect 42246 529479 42302 529488
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42260 527762 42288 529479
rect 42168 527734 42288 527762
rect 42168 527340 42196 527734
rect 42444 526742 42472 529751
rect 42706 529136 42762 529145
rect 42182 526714 42472 526742
rect 42536 529094 42706 529122
rect 42536 526091 42564 529094
rect 42706 529071 42762 529080
rect 42182 526063 42564 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40958 425640 41014 425649
rect 40958 425575 41014 425584
rect 33690 424416 33746 424425
rect 33690 424351 33746 424360
rect 33704 416226 33732 424351
rect 40972 421274 41000 425575
rect 41340 425066 41368 425983
rect 41328 425060 41380 425066
rect 41328 425002 41380 425008
rect 41696 425060 41748 425066
rect 41696 425002 41748 425008
rect 41708 424946 41736 425002
rect 41708 424918 42012 424946
rect 41326 424008 41382 424017
rect 41326 423943 41382 423952
rect 41340 423842 41368 423943
rect 41786 423872 41842 423881
rect 41328 423836 41380 423842
rect 41328 423778 41380 423784
rect 41604 423836 41656 423842
rect 41656 423816 41786 423824
rect 41656 423807 41842 423816
rect 41656 423796 41828 423807
rect 41604 423778 41656 423784
rect 41326 422376 41382 422385
rect 41786 422376 41842 422385
rect 41326 422311 41328 422320
rect 41380 422311 41382 422320
rect 41604 422340 41656 422346
rect 41328 422282 41380 422288
rect 41656 422320 41786 422328
rect 41656 422311 41842 422320
rect 41656 422300 41828 422311
rect 41604 422282 41656 422288
rect 41786 421288 41842 421297
rect 40972 421246 41786 421274
rect 41786 421223 41842 421232
rect 41326 421152 41382 421161
rect 41326 421087 41382 421096
rect 41340 420986 41368 421087
rect 41786 421016 41842 421025
rect 41328 420980 41380 420986
rect 41328 420922 41380 420928
rect 41604 420980 41656 420986
rect 41656 420960 41786 420968
rect 41656 420951 41842 420960
rect 41656 420940 41828 420951
rect 41604 420922 41656 420928
rect 41984 418154 42012 424918
rect 42798 423872 42854 423881
rect 42798 423807 42854 423816
rect 42154 422784 42210 422793
rect 42154 422719 42210 422728
rect 42168 418849 42196 422719
rect 42338 421968 42394 421977
rect 42338 421903 42394 421912
rect 42154 418840 42210 418849
rect 42154 418775 42210 418784
rect 42352 418577 42380 421903
rect 42522 419928 42578 419937
rect 42522 419863 42578 419872
rect 42338 418568 42394 418577
rect 42338 418503 42394 418512
rect 41984 418126 42472 418154
rect 33692 416220 33744 416226
rect 33692 416162 33744 416168
rect 41696 416220 41748 416226
rect 41696 416162 41748 416168
rect 41708 416106 41736 416162
rect 41708 416078 42288 416106
rect 42260 413114 42288 416078
rect 42444 415394 42472 418126
rect 42168 413086 42288 413114
rect 42352 415366 42472 415394
rect 42536 415394 42564 419863
rect 42536 415366 42656 415394
rect 42168 412624 42196 413086
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42352 411074 42380 415366
rect 42628 411913 42656 415366
rect 42614 411904 42670 411913
rect 42614 411839 42670 411848
rect 42168 411046 42380 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42430 407144 42486 407153
rect 42182 407102 42430 407130
rect 42430 407079 42486 407088
rect 42430 406872 42486 406881
rect 42430 406807 42486 406816
rect 42444 406518 42472 406807
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42182 402138 42472 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42444 400217 42472 402138
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423807
rect 43166 422376 43222 422385
rect 43166 422311 43222 422320
rect 42982 421016 43038 421025
rect 42982 420951 43038 420960
rect 42996 407833 43024 420951
rect 42982 407824 43038 407833
rect 42982 407759 43038 407768
rect 43180 407153 43208 422311
rect 43166 407144 43222 407153
rect 43166 407079 43222 407088
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41340 387654 41552 387682
rect 41142 387152 41198 387161
rect 41142 387087 41144 387096
rect 41196 387087 41198 387096
rect 41144 387058 41196 387064
rect 41340 386753 41368 387654
rect 41524 386753 41552 387654
rect 41708 387122 41920 387138
rect 41696 387116 41920 387122
rect 41748 387110 41920 387116
rect 41696 387058 41748 387064
rect 41892 387025 41920 387110
rect 41878 387016 41934 387025
rect 41878 386951 41934 386960
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 41326 383072 41382 383081
rect 41326 383007 41382 383016
rect 41142 382664 41198 382673
rect 41142 382599 41198 382608
rect 41156 382294 41184 382599
rect 41340 382430 41368 383007
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41696 382424 41748 382430
rect 41748 382384 42840 382412
rect 41696 382366 41748 382372
rect 41144 382288 41196 382294
rect 40222 382256 40278 382265
rect 41144 382230 41196 382236
rect 41696 382288 41748 382294
rect 41748 382248 41920 382276
rect 41696 382230 41748 382236
rect 40222 382191 40278 382200
rect 40038 381848 40094 381857
rect 40038 381783 40094 381792
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 35820 379409 35848 379510
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 40052 376553 40080 381783
rect 40236 376961 40264 382191
rect 41326 381032 41382 381041
rect 41326 380967 41382 380976
rect 41340 378593 41368 380967
rect 41696 379568 41748 379574
rect 41696 379510 41748 379516
rect 41892 379514 41920 382248
rect 41708 379409 41736 379510
rect 41892 379486 42564 379514
rect 41694 379400 41750 379409
rect 41694 379335 41750 379344
rect 41326 378584 41382 378593
rect 41326 378519 41382 378528
rect 42338 378584 42394 378593
rect 42338 378519 42394 378528
rect 40222 376952 40278 376961
rect 40222 376887 40278 376896
rect 42352 376754 42380 378519
rect 42352 376726 42472 376754
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 40038 376544 40094 376553
rect 40038 376479 40094 376488
rect 28906 376136 28962 376145
rect 28906 376071 28962 376080
rect 28920 371890 28948 376071
rect 35820 376038 35848 376479
rect 35808 376032 35860 376038
rect 35808 375974 35860 375980
rect 39580 376032 39632 376038
rect 39580 375974 39632 375980
rect 39592 375737 39620 375974
rect 39578 375728 39634 375737
rect 39578 375663 39634 375672
rect 41694 371920 41750 371929
rect 28908 371884 28960 371890
rect 41694 371855 41696 371864
rect 28908 371826 28960 371832
rect 41748 371855 41750 371864
rect 41696 371826 41748 371832
rect 42444 369458 42472 376726
rect 42182 369430 42472 369458
rect 41786 368656 41842 368665
rect 41786 368591 41842 368600
rect 41800 368249 41828 368591
rect 42536 367622 42564 379486
rect 42182 367594 42564 367622
rect 42430 367024 42486 367033
rect 42182 366968 42430 366975
rect 42182 366959 42486 366968
rect 42182 366947 42472 366959
rect 42430 365800 42486 365809
rect 42182 365758 42430 365786
rect 42430 365735 42486 365744
rect 41800 364313 41828 364548
rect 41786 364304 41842 364313
rect 41786 364239 41842 364248
rect 42182 363922 42472 363950
rect 41786 363624 41842 363633
rect 41786 363559 41842 363568
rect 41800 363256 41828 363559
rect 41878 362944 41934 362953
rect 41878 362879 41934 362888
rect 41892 362712 41920 362879
rect 42444 361593 42472 363922
rect 42430 361584 42486 361593
rect 42430 361519 42486 361528
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 42182 358958 42472 358986
rect 42062 358728 42118 358737
rect 42062 358663 42118 358672
rect 42076 358428 42104 358663
rect 42444 357377 42472 358958
rect 42430 357368 42486 357377
rect 42430 357303 42486 357312
rect 42812 356674 42840 382384
rect 43456 379514 43484 590271
rect 44192 581097 44220 591903
rect 44178 581088 44234 581097
rect 44178 581023 44234 581032
rect 44652 555665 44680 598431
rect 44836 557297 44864 600063
rect 45006 599312 45062 599321
rect 45006 599247 45062 599256
rect 44822 557288 44878 557297
rect 44822 557223 44878 557232
rect 45020 556481 45048 599247
rect 45204 598097 45232 640863
rect 45388 598913 45416 641135
rect 45572 611522 45600 721103
rect 46110 719944 46166 719953
rect 46110 719879 46166 719888
rect 45742 676696 45798 676705
rect 45742 676631 45798 676640
rect 45560 611516 45612 611522
rect 45560 611458 45612 611464
rect 45756 611318 45784 676631
rect 45926 637800 45982 637809
rect 45926 637735 45982 637744
rect 45940 613601 45968 637735
rect 45926 613592 45982 613601
rect 45926 613527 45982 613536
rect 46124 611726 46152 719879
rect 46294 636984 46350 636993
rect 46294 636919 46350 636928
rect 46308 619585 46336 636919
rect 46478 626648 46534 626657
rect 46478 626583 46534 626592
rect 46492 624209 46520 626583
rect 46478 624200 46534 624209
rect 46478 624135 46534 624144
rect 46294 619576 46350 619585
rect 46294 619511 46350 619520
rect 46952 611930 46980 764351
rect 47596 712201 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47582 712192 47638 712201
rect 47582 712127 47638 712136
rect 47214 677920 47270 677929
rect 47214 677855 47270 677864
rect 46940 611924 46992 611930
rect 46940 611866 46992 611872
rect 46112 611720 46164 611726
rect 46112 611662 46164 611668
rect 45744 611312 45796 611318
rect 45744 611254 45796 611260
rect 47228 611017 47256 677855
rect 48976 669361 49004 767314
rect 50356 730561 50384 805938
rect 53116 799649 53144 923238
rect 53300 892537 53328 988722
rect 53286 892528 53342 892537
rect 53286 892463 53342 892472
rect 54496 892265 54524 991442
rect 55876 892809 55904 992870
rect 73172 983634 73200 994230
rect 80716 994158 80744 995452
rect 81360 994430 81388 995452
rect 82004 994702 82032 995452
rect 85040 994945 85068 995452
rect 85698 995438 86080 995466
rect 85026 994936 85082 994945
rect 85026 994871 85082 994880
rect 81992 994696 82044 994702
rect 81992 994638 82044 994644
rect 85488 994696 85540 994702
rect 85488 994638 85540 994644
rect 85500 994430 85528 994638
rect 81348 994424 81400 994430
rect 81348 994366 81400 994372
rect 85488 994424 85540 994430
rect 85488 994366 85540 994372
rect 85672 994424 85724 994430
rect 86052 994401 86080 995438
rect 86328 995217 86356 995452
rect 90022 995438 90270 995466
rect 91218 995438 91692 995466
rect 90270 995415 90326 995424
rect 91664 995330 91692 995438
rect 92032 995330 92060 995574
rect 92492 995489 92520 998650
rect 92676 995761 92704 1003886
rect 92848 999796 92900 999802
rect 92848 999738 92900 999744
rect 92662 995752 92718 995761
rect 92662 995687 92718 995696
rect 92664 995580 92716 995586
rect 92664 995522 92716 995528
rect 92478 995480 92534 995489
rect 92478 995415 92534 995424
rect 91664 995302 92060 995330
rect 86314 995208 86370 995217
rect 86314 995143 86370 995152
rect 92676 994945 92704 995522
rect 92662 994936 92718 994945
rect 92662 994871 92718 994880
rect 92860 994401 92888 999738
rect 93136 995217 93164 1005994
rect 93320 998714 93348 1006130
rect 93492 1001224 93544 1001230
rect 93492 1001166 93544 1001172
rect 93308 998708 93360 998714
rect 93308 998650 93360 998656
rect 93308 997756 93360 997762
rect 93308 997698 93360 997704
rect 93320 996441 93348 997698
rect 93504 997257 93532 1001166
rect 93490 997248 93546 997257
rect 93490 997183 93546 997192
rect 94516 996985 94544 1006402
rect 101126 1006360 101182 1006369
rect 94688 1006324 94740 1006330
rect 101126 1006295 101128 1006304
rect 94688 1006266 94740 1006272
rect 101180 1006295 101182 1006304
rect 144276 1006324 144328 1006330
rect 101128 1006266 101180 1006272
rect 144276 1006266 144328 1006272
rect 94502 996976 94558 996985
rect 94502 996911 94558 996920
rect 94700 996713 94728 1006266
rect 98274 1006224 98330 1006233
rect 98274 1006159 98276 1006168
rect 98328 1006159 98330 1006168
rect 107658 1006224 107714 1006233
rect 107658 1006159 107660 1006168
rect 98276 1006130 98328 1006136
rect 107712 1006159 107714 1006168
rect 124864 1006188 124916 1006194
rect 107660 1006130 107712 1006136
rect 124864 1006130 124916 1006136
rect 144092 1006188 144144 1006194
rect 144092 1006130 144144 1006136
rect 99470 1006088 99526 1006097
rect 104806 1006088 104862 1006097
rect 99470 1006023 99472 1006032
rect 99524 1006023 99526 1006032
rect 102784 1006052 102836 1006058
rect 99472 1005994 99524 1006000
rect 104806 1006023 104808 1006032
rect 102784 1005994 102836 1006000
rect 104860 1006023 104862 1006032
rect 108486 1006088 108542 1006097
rect 108486 1006023 108488 1006032
rect 104808 1005994 104860 1006000
rect 108540 1006023 108542 1006032
rect 108488 1005994 108540 1006000
rect 101494 1002552 101550 1002561
rect 98644 1002516 98696 1002522
rect 101494 1002487 101496 1002496
rect 98644 1002458 98696 1002464
rect 101548 1002487 101550 1002496
rect 101496 1002458 101548 1002464
rect 97264 1002380 97316 1002386
rect 97264 1002322 97316 1002328
rect 95884 1002244 95936 1002250
rect 95884 1002186 95936 1002192
rect 94686 996704 94742 996713
rect 94686 996639 94742 996648
rect 93306 996432 93362 996441
rect 93306 996367 93362 996376
rect 93308 996260 93360 996266
rect 93308 996202 93360 996208
rect 93320 996033 93348 996202
rect 93306 996024 93362 996033
rect 93306 995959 93362 995968
rect 93122 995208 93178 995217
rect 93122 995143 93178 995152
rect 85672 994366 85724 994372
rect 86038 994392 86094 994401
rect 85684 994158 85712 994366
rect 86038 994327 86094 994336
rect 92846 994392 92902 994401
rect 92846 994327 92902 994336
rect 80704 994152 80756 994158
rect 80704 994094 80756 994100
rect 85672 994152 85724 994158
rect 85672 994094 85724 994100
rect 89720 990276 89772 990282
rect 89720 990218 89772 990224
rect 89732 985402 89760 990218
rect 95896 988786 95924 1002186
rect 96068 1001972 96120 1001978
rect 96068 1001914 96120 1001920
rect 96080 991778 96108 1001914
rect 97276 994566 97304 1002322
rect 97448 1002108 97500 1002114
rect 97448 1002050 97500 1002056
rect 97460 995586 97488 1002050
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 98000 1000544 98052 1000550
rect 98000 1000486 98052 1000492
rect 98012 998442 98040 1000486
rect 98000 998436 98052 998442
rect 98000 998378 98052 998384
rect 97448 995580 97500 995586
rect 97448 995522 97500 995528
rect 98656 994702 98684 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100484 1002380 100536 1002386
rect 100300 1002322 100352 1002328
rect 100484 1002322 100536 1002328
rect 99102 1002280 99158 1002289
rect 99102 1002215 99104 1002224
rect 99156 1002215 99158 1002224
rect 100024 1002244 100076 1002250
rect 99104 1002186 99156 1002192
rect 100024 1002186 100076 1002192
rect 98828 1001972 98880 1001978
rect 98828 1001914 98880 1001920
rect 98840 999802 98868 1001914
rect 98828 999796 98880 999802
rect 98828 999738 98880 999744
rect 98644 994696 98696 994702
rect 98644 994638 98696 994644
rect 97264 994560 97316 994566
rect 97264 994502 97316 994508
rect 100036 994430 100064 1002186
rect 100298 1002144 100354 1002153
rect 100298 1002079 100300 1002088
rect 100352 1002079 100354 1002088
rect 100300 1002050 100352 1002056
rect 100496 1000550 100524 1002322
rect 101954 1002280 102010 1002289
rect 101954 1002215 101956 1002224
rect 102008 1002215 102010 1002224
rect 101956 1002186 102008 1002192
rect 101588 1002108 101640 1002114
rect 101588 1002050 101640 1002056
rect 101126 1002008 101182 1002017
rect 101126 1001943 101128 1001952
rect 101180 1001943 101182 1001952
rect 101404 1001972 101456 1001978
rect 101128 1001914 101180 1001920
rect 101404 1001914 101456 1001920
rect 100484 1000544 100536 1000550
rect 100484 1000486 100536 1000492
rect 101416 995217 101444 1001914
rect 101600 1001230 101628 1002050
rect 102322 1002008 102378 1002017
rect 102322 1001943 102324 1001952
rect 102376 1001943 102378 1001952
rect 102324 1001914 102376 1001920
rect 101588 1001224 101640 1001230
rect 101588 1001166 101640 1001172
rect 101402 995208 101458 995217
rect 101402 995143 101458 995152
rect 102796 994838 102824 1005994
rect 104808 1003944 104860 1003950
rect 104806 1003912 104808 1003921
rect 104860 1003912 104862 1003921
rect 104806 1003847 104862 1003856
rect 106830 1002688 106886 1002697
rect 106830 1002623 106832 1002632
rect 106884 1002623 106886 1002632
rect 109500 1002652 109552 1002658
rect 106832 1002594 106884 1002600
rect 109500 1002594 109552 1002600
rect 108026 1002552 108082 1002561
rect 108026 1002487 108028 1002496
rect 108080 1002487 108082 1002496
rect 108028 1002458 108080 1002464
rect 103150 1002416 103206 1002425
rect 103150 1002351 103152 1002360
rect 103204 1002351 103206 1002360
rect 106830 1002416 106886 1002425
rect 106830 1002351 106832 1002360
rect 103152 1002322 103204 1002328
rect 106884 1002351 106886 1002360
rect 109040 1002380 109092 1002386
rect 106832 1002322 106884 1002328
rect 109040 1002322 109092 1002328
rect 106002 1002280 106058 1002289
rect 108854 1002280 108910 1002289
rect 106002 1002215 106004 1002224
rect 106056 1002215 106058 1002224
rect 108304 1002244 108356 1002250
rect 106004 1002186 106056 1002192
rect 108854 1002215 108856 1002224
rect 108304 1002186 108356 1002192
rect 108908 1002215 108910 1002224
rect 108856 1002186 108908 1002192
rect 103150 1002144 103206 1002153
rect 103150 1002079 103152 1002088
rect 103204 1002079 103206 1002088
rect 105634 1002144 105690 1002153
rect 105634 1002079 105636 1002088
rect 103152 1002050 103204 1002056
rect 105688 1002079 105690 1002088
rect 107752 1002108 107804 1002114
rect 105636 1002050 105688 1002056
rect 107752 1002050 107804 1002056
rect 103978 1002008 104034 1002017
rect 103532 1001966 103978 1001994
rect 103532 997762 103560 1001966
rect 103978 1001943 104034 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 103520 997756 103572 997762
rect 103520 997698 103572 997704
rect 106924 996804 106976 996810
rect 106924 996746 106976 996752
rect 103888 996396 103940 996402
rect 103888 996338 103940 996344
rect 102784 994832 102836 994838
rect 102784 994774 102836 994780
rect 103900 994430 103928 996338
rect 100024 994424 100076 994430
rect 100024 994366 100076 994372
rect 103888 994424 103940 994430
rect 103888 994366 103940 994372
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 988780 95936 988786
rect 95884 988722 95936 988728
rect 106936 986610 106964 996746
rect 107764 993206 107792 1002050
rect 108120 1001972 108172 1001978
rect 108120 1001914 108172 1001920
rect 107752 993200 107804 993206
rect 107752 993142 107804 993148
rect 108132 993070 108160 1001914
rect 108316 997626 108344 1002186
rect 108854 1002008 108910 1002017
rect 108854 1001943 108856 1001952
rect 108908 1001943 108910 1001952
rect 108856 1001914 108908 1001920
rect 108304 997620 108356 997626
rect 108304 997562 108356 997568
rect 108120 993064 108172 993070
rect 108120 993006 108172 993012
rect 109052 990146 109080 1002322
rect 109512 997762 109540 1002594
rect 110696 1002516 110748 1002522
rect 110696 1002458 110748 1002464
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 110512 1001972 110564 1001978
rect 110512 1001914 110564 1001920
rect 109500 997756 109552 997762
rect 109500 997698 109552 997704
rect 110524 996810 110552 1001914
rect 110512 996804 110564 996810
rect 110512 996746 110564 996752
rect 110708 991642 110736 1002458
rect 111892 1002244 111944 1002250
rect 111892 1002186 111944 1002192
rect 111904 994294 111932 1002186
rect 112076 1002108 112128 1002114
rect 112076 1002050 112128 1002056
rect 111892 994288 111944 994294
rect 111892 994230 111944 994236
rect 110696 991636 110748 991642
rect 110696 991578 110748 991584
rect 112088 990282 112116 1002050
rect 116308 997756 116360 997762
rect 116308 997698 116360 997704
rect 116320 996985 116348 997698
rect 117228 997620 117280 997626
rect 117228 997562 117280 997568
rect 117240 997257 117268 997562
rect 117226 997248 117282 997257
rect 117226 997183 117282 997192
rect 116306 996976 116362 996985
rect 116306 996911 116362 996920
rect 124876 995081 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 126256 996305 126284 1005994
rect 144104 1001894 144132 1006130
rect 143828 1001866 144132 1001894
rect 144288 1001894 144316 1006266
rect 144288 1001866 144408 1001894
rect 126242 996296 126298 996305
rect 126242 996231 126298 996240
rect 136468 995858 136496 995860
rect 143828 995858 143856 1001866
rect 144184 998436 144236 998442
rect 144184 998378 144236 998384
rect 144000 997756 144052 997762
rect 144000 997698 144052 997704
rect 144012 996985 144040 997698
rect 143998 996976 144054 996985
rect 143998 996911 144054 996920
rect 144000 996396 144052 996402
rect 144000 996338 144052 996344
rect 136456 995852 136508 995858
rect 136456 995794 136508 995800
rect 143816 995852 143868 995858
rect 143816 995794 143868 995800
rect 131854 995752 131910 995761
rect 131606 995710 131854 995738
rect 131854 995687 131910 995696
rect 132958 995752 133014 995761
rect 140410 995752 140466 995761
rect 133014 995710 133446 995738
rect 140162 995710 140410 995738
rect 132958 995687 133014 995696
rect 141054 995752 141110 995761
rect 140806 995710 141054 995738
rect 140410 995687 140466 995696
rect 144012 995738 144040 996338
rect 144196 995897 144224 998378
rect 144182 995888 144238 995897
rect 144182 995823 144238 995832
rect 141054 995687 141110 995696
rect 143460 995710 144040 995738
rect 141790 995616 141846 995625
rect 141450 995574 141790 995602
rect 141790 995551 141846 995560
rect 137374 995480 137430 995489
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994702 128492 995452
rect 128452 994696 128504 994702
rect 128452 994638 128504 994644
rect 129108 994430 129136 995452
rect 129752 994838 129780 995452
rect 129740 994832 129792 994838
rect 132144 994809 132172 995452
rect 132802 995438 133184 995466
rect 132406 995344 132462 995353
rect 132406 995279 132462 995288
rect 129740 994774 129792 994780
rect 132130 994800 132186 994809
rect 132130 994735 132186 994744
rect 132420 994566 132448 995279
rect 132408 994560 132460 994566
rect 132408 994502 132460 994508
rect 121736 994424 121788 994430
rect 121736 994366 121788 994372
rect 129096 994424 129148 994430
rect 129096 994366 129148 994372
rect 112076 990276 112128 990282
rect 112076 990218 112128 990224
rect 109040 990140 109092 990146
rect 109040 990082 109092 990088
rect 105820 986604 105872 986610
rect 105820 986546 105872 986552
rect 106924 986604 106976 986610
rect 106924 986546 106976 986552
rect 89640 985374 89760 985402
rect 73172 983606 73462 983634
rect 89640 983620 89668 985374
rect 105832 983620 105860 986546
rect 121748 983634 121776 994366
rect 133156 993721 133184 995438
rect 135916 994401 135944 995452
rect 137126 995438 137374 995466
rect 137374 995415 137430 995424
rect 135902 994392 135958 994401
rect 135902 994327 135958 994336
rect 137558 994120 137614 994129
rect 137558 994055 137560 994064
rect 137612 994055 137614 994064
rect 137560 994026 137612 994032
rect 137756 993993 137784 995452
rect 138966 995438 139348 995466
rect 142646 995438 143028 995466
rect 139320 995058 139348 995438
rect 143000 995330 143028 995438
rect 143460 995330 143488 995710
rect 143000 995302 143488 995330
rect 139320 995030 139440 995058
rect 139216 994220 139268 994226
rect 139216 994162 139268 994168
rect 137742 993984 137798 993993
rect 137742 993919 137798 993928
rect 139228 993721 139256 994162
rect 139412 993721 139440 995030
rect 144380 994809 144408 1001866
rect 144828 997620 144880 997626
rect 144828 997562 144880 997568
rect 144840 997257 144868 997562
rect 144826 997248 144882 997257
rect 144826 997183 144882 997192
rect 144826 996568 144882 996577
rect 144826 996503 144828 996512
rect 144880 996503 144882 996512
rect 144828 996474 144880 996480
rect 144366 994800 144422 994809
rect 144366 994735 144422 994744
rect 144550 994800 144606 994809
rect 144550 994735 144606 994744
rect 142158 994528 142214 994537
rect 141804 994486 142158 994514
rect 141804 994090 141832 994486
rect 142158 994463 142214 994472
rect 141974 994392 142030 994401
rect 141974 994327 142030 994336
rect 141792 994084 141844 994090
rect 141792 994026 141844 994032
rect 133142 993712 133198 993721
rect 133142 993647 133198 993656
rect 139214 993712 139270 993721
rect 139214 993647 139270 993656
rect 139398 993712 139454 993721
rect 141988 993698 142016 994327
rect 144564 994226 144592 994735
rect 144552 994220 144604 994226
rect 144552 994162 144604 994168
rect 145576 993993 145604 1006538
rect 152094 1006496 152150 1006505
rect 145748 1006460 145800 1006466
rect 152094 1006431 152096 1006440
rect 145748 1006402 145800 1006408
rect 152148 1006431 152150 1006440
rect 157430 1006496 157486 1006505
rect 157430 1006431 157432 1006440
rect 152096 1006402 152148 1006408
rect 157484 1006431 157486 1006440
rect 166264 1006460 166316 1006466
rect 157432 1006402 157484 1006408
rect 166264 1006402 166316 1006408
rect 171784 1006460 171836 1006466
rect 171784 1006402 171836 1006408
rect 145760 996169 145788 1006402
rect 158258 1006360 158314 1006369
rect 158258 1006295 158260 1006304
rect 158312 1006295 158314 1006304
rect 158260 1006266 158312 1006272
rect 151266 1006224 151322 1006233
rect 151266 1006159 151268 1006168
rect 151320 1006159 151322 1006168
rect 153750 1006224 153806 1006233
rect 153750 1006159 153752 1006168
rect 151268 1006130 151320 1006136
rect 153804 1006159 153806 1006168
rect 160282 1006224 160338 1006233
rect 166276 1006194 166304 1006402
rect 160282 1006159 160284 1006168
rect 153752 1006130 153804 1006136
rect 160336 1006159 160338 1006168
rect 164884 1006188 164936 1006194
rect 160284 1006130 160336 1006136
rect 164884 1006130 164936 1006136
rect 166264 1006188 166316 1006194
rect 166264 1006130 166316 1006136
rect 147126 1006088 147182 1006097
rect 147126 1006023 147182 1006032
rect 148874 1006088 148930 1006097
rect 148874 1006023 148876 1006032
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145746 996160 145802 996169
rect 145746 996095 145802 996104
rect 142342 993984 142398 993993
rect 142342 993919 142398 993928
rect 145562 993984 145618 993993
rect 145562 993919 145618 993928
rect 142158 993712 142214 993721
rect 141988 993670 142158 993698
rect 139398 993647 139454 993656
rect 142158 993647 142214 993656
rect 142356 993449 142384 993919
rect 142342 993440 142398 993449
rect 142342 993375 142398 993384
rect 146956 992934 146984 1001914
rect 147140 995625 147168 1006023
rect 148928 1006023 148930 1006032
rect 150070 1006088 150126 1006097
rect 150070 1006023 150072 1006032
rect 148876 1005994 148928 1006000
rect 150124 1006023 150126 1006032
rect 159454 1006088 159510 1006097
rect 159454 1006023 159456 1006032
rect 150072 1005994 150124 1006000
rect 159508 1006023 159510 1006032
rect 159456 1005994 159508 1006000
rect 152922 1005136 152978 1005145
rect 149888 1005100 149940 1005106
rect 152922 1005071 152924 1005080
rect 149888 1005042 149940 1005048
rect 152976 1005071 152978 1005080
rect 158626 1005136 158682 1005145
rect 158626 1005071 158628 1005080
rect 152924 1005042 152976 1005048
rect 158680 1005071 158682 1005080
rect 162124 1005100 162176 1005106
rect 158628 1005042 158680 1005048
rect 162124 1005042 162176 1005048
rect 149704 1004828 149756 1004834
rect 149704 1004770 149756 1004776
rect 148508 1002380 148560 1002386
rect 148508 1002322 148560 1002328
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 147126 995616 147182 995625
rect 147126 995551 147182 995560
rect 146944 992928 146996 992934
rect 146944 992870 146996 992876
rect 138296 991636 138348 991642
rect 138296 991578 138348 991584
rect 121748 983606 122130 983634
rect 138308 983620 138336 991578
rect 148336 991506 148364 1002050
rect 148520 994265 148548 1002322
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149716 994566 149744 1004770
rect 149900 994809 149928 1005042
rect 153750 1005000 153806 1005009
rect 151084 1004964 151136 1004970
rect 153750 1004935 153752 1004944
rect 151084 1004906 151136 1004912
rect 153804 1004935 153806 1004944
rect 153752 1004906 153804 1004912
rect 150898 1002416 150954 1002425
rect 150898 1002351 150900 1002360
rect 150952 1002351 150954 1002360
rect 150900 1002322 150952 1002328
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 150440 996532 150492 996538
rect 150440 996474 150492 996480
rect 149886 994800 149942 994809
rect 149886 994735 149942 994744
rect 149704 994560 149756 994566
rect 149704 994502 149756 994508
rect 150452 994294 150480 996474
rect 151096 994430 151124 1004906
rect 151726 1004864 151782 1004873
rect 151726 1004799 151728 1004808
rect 151780 1004799 151782 1004808
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 151728 1004770 151780 1004776
rect 160704 1004799 160706 1004808
rect 160652 1004770 160704 1004776
rect 154118 1004728 154174 1004737
rect 151268 1004692 151320 1004698
rect 154118 1004663 154120 1004672
rect 151268 1004634 151320 1004640
rect 154172 1004663 154174 1004672
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 154120 1004634 154172 1004640
rect 161164 1004663 161166 1004672
rect 161112 1004634 161164 1004640
rect 151280 996402 151308 1004634
rect 155774 1002280 155830 1002289
rect 153844 1002244 153896 1002250
rect 155774 1002215 155776 1002224
rect 153844 1002186 153896 1002192
rect 155828 1002215 155830 1002224
rect 156602 1002280 156658 1002289
rect 156602 1002215 156604 1002224
rect 155776 1002186 155828 1002192
rect 156656 1002215 156658 1002224
rect 158720 1002244 158772 1002250
rect 156604 1002186 156656 1002192
rect 158720 1002186 158772 1002192
rect 152464 1001972 152516 1001978
rect 152464 1001914 152516 1001920
rect 151268 996396 151320 996402
rect 151268 996338 151320 996344
rect 151084 994424 151136 994430
rect 151084 994366 151136 994372
rect 150440 994288 150492 994294
rect 148506 994256 148562 994265
rect 150440 994230 150492 994236
rect 148506 994191 148562 994200
rect 152476 993993 152504 1001914
rect 153856 994702 153884 1002186
rect 154578 1002008 154634 1002017
rect 154578 1001943 154580 1001952
rect 154632 1001943 154634 1001952
rect 154946 1002008 155002 1002017
rect 155774 1002008 155830 1002017
rect 154946 1001943 154948 1001952
rect 154580 1001914 154632 1001920
rect 155000 1001943 155002 1001952
rect 155236 1001966 155774 1001994
rect 154948 1001914 155000 1001920
rect 155236 998442 155264 1001966
rect 156602 1002008 156658 1002017
rect 155774 1001943 155830 1001952
rect 155972 1001966 156602 1001994
rect 155224 998436 155276 998442
rect 155224 998378 155276 998384
rect 155130 995616 155186 995625
rect 155130 995551 155186 995560
rect 155144 995081 155172 995551
rect 155130 995072 155186 995081
rect 155130 995007 155186 995016
rect 155972 994838 156000 1001966
rect 157798 1002008 157854 1002017
rect 156602 1001943 156658 1001952
rect 157340 1001972 157392 1001978
rect 157798 1001943 157800 1001952
rect 157340 1001914 157392 1001920
rect 157852 1001943 157854 1001952
rect 157800 1001914 157852 1001920
rect 155960 994832 156012 994838
rect 155960 994774 156012 994780
rect 153844 994696 153896 994702
rect 153844 994638 153896 994644
rect 157352 994537 157380 1001914
rect 158732 997626 158760 1002186
rect 160100 1001972 160152 1001978
rect 160100 1001914 160152 1001920
rect 160112 997762 160140 1001914
rect 162136 997762 162164 1005042
rect 163136 1004828 163188 1004834
rect 163136 1004770 163188 1004776
rect 162952 1004692 163004 1004698
rect 162952 1004634 163004 1004640
rect 160100 997756 160152 997762
rect 160100 997698 160152 997704
rect 162124 997756 162176 997762
rect 162124 997698 162176 997704
rect 158720 997620 158772 997626
rect 158720 997562 158772 997568
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 157338 994528 157394 994537
rect 157338 994463 157394 994472
rect 152462 993984 152518 993993
rect 152462 993919 152518 993928
rect 148324 991500 148376 991506
rect 148324 991442 148376 991448
rect 160756 985726 160784 997154
rect 163148 991642 163176 1004770
rect 163136 991636 163188 991642
rect 163136 991578 163188 991584
rect 164896 990894 164924 1006130
rect 170312 997756 170364 997762
rect 170312 997698 170364 997704
rect 170324 997257 170352 997698
rect 170310 997248 170366 997257
rect 170310 997183 170366 997192
rect 171796 996130 171824 1006402
rect 210054 1006360 210110 1006369
rect 204904 1006324 204956 1006330
rect 254122 1006360 254178 1006369
rect 210054 1006295 210056 1006304
rect 204904 1006266 204956 1006272
rect 210108 1006295 210110 1006304
rect 249248 1006324 249300 1006330
rect 210056 1006266 210108 1006272
rect 254122 1006295 254124 1006304
rect 249248 1006266 249300 1006272
rect 254176 1006295 254178 1006304
rect 298928 1006324 298980 1006330
rect 254124 1006266 254176 1006272
rect 298928 1006266 298980 1006272
rect 175924 1006188 175976 1006194
rect 175924 1006130 175976 1006136
rect 172334 996296 172390 996305
rect 172334 996231 172390 996240
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 169392 995988 169444 995994
rect 169392 995930 169444 995936
rect 171508 995988 171560 995994
rect 171508 995930 171560 995936
rect 169404 994770 169432 995930
rect 170680 995852 170732 995858
rect 170680 995794 170732 995800
rect 169392 994764 169444 994770
rect 169392 994706 169444 994712
rect 170692 994498 170720 995794
rect 171048 995580 171100 995586
rect 171048 995522 171100 995528
rect 170864 994881 170916 994887
rect 170864 994823 170916 994829
rect 170680 994492 170732 994498
rect 170680 994434 170732 994440
rect 170876 993682 170904 994823
rect 171060 994634 171088 995522
rect 171520 995223 171548 995930
rect 171692 995852 171744 995858
rect 171692 995794 171744 995800
rect 171704 995335 171732 995794
rect 171692 995329 171744 995335
rect 171692 995271 171744 995277
rect 171508 995217 171560 995223
rect 171508 995159 171560 995165
rect 172348 995110 172376 996231
rect 172336 995104 172388 995110
rect 175936 995081 175964 1006130
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 198372 1006052 198424 1006058
rect 201038 1006023 201040 1006032
rect 198372 1005994 198424 1006000
rect 201092 1006023 201094 1006032
rect 201040 1005994 201092 1006000
rect 177316 995994 177344 1005994
rect 195152 1002108 195204 1002114
rect 195152 1002050 195204 1002056
rect 195164 1001894 195192 1002050
rect 195072 1001866 195192 1001894
rect 195072 996985 195100 1001866
rect 195888 1001836 195940 1001842
rect 195888 1001778 195940 1001784
rect 195520 998436 195572 998442
rect 195520 998378 195572 998384
rect 195336 997960 195388 997966
rect 195256 997908 195336 997914
rect 195256 997902 195388 997908
rect 195256 997886 195376 997902
rect 195058 996976 195114 996985
rect 195058 996911 195114 996920
rect 177304 995988 177356 995994
rect 177304 995930 177356 995936
rect 183834 995752 183890 995761
rect 183540 995710 183834 995738
rect 183834 995687 183890 995696
rect 188802 995616 188858 995625
rect 188508 995574 188802 995602
rect 190458 995616 190514 995625
rect 190348 995574 190458 995602
rect 188802 995551 188858 995560
rect 190458 995551 190514 995560
rect 194876 995512 194928 995518
rect 179860 995438 180196 995466
rect 180504 995438 180656 995466
rect 181148 995438 181484 995466
rect 182988 995438 183324 995466
rect 184184 995438 184704 995466
rect 172336 995046 172388 995052
rect 175922 995072 175978 995081
rect 175922 995007 175978 995016
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 171048 994628 171100 994634
rect 171048 994570 171100 994576
rect 171244 993818 171272 994823
rect 180168 994809 180196 995438
rect 180628 995110 180656 995438
rect 180616 995104 180668 995110
rect 180616 995046 180668 995052
rect 181456 994974 181484 995438
rect 181444 994968 181496 994974
rect 181444 994910 181496 994916
rect 180154 994800 180210 994809
rect 180154 994735 180210 994744
rect 183296 994265 183324 995438
rect 184676 995058 184704 995438
rect 184814 995246 184842 995452
rect 187312 995438 187648 995466
rect 187864 995438 188200 995466
rect 189152 995438 189488 995466
rect 191544 995438 191788 995466
rect 192188 995438 192524 995466
rect 192832 995438 193168 995466
rect 194028 995438 194364 995466
rect 195256 995466 195284 997886
rect 194876 995454 194928 995460
rect 184802 995240 184854 995246
rect 184802 995182 184854 995188
rect 184676 995030 184980 995058
rect 183282 994256 183338 994265
rect 183282 994191 183338 994200
rect 184952 994158 184980 995030
rect 187620 994537 187648 995438
rect 188172 995353 188200 995438
rect 189460 995382 189488 995438
rect 189448 995376 189500 995382
rect 188158 995344 188214 995353
rect 189448 995318 189500 995324
rect 188158 995279 188214 995288
rect 187606 994528 187662 994537
rect 187606 994463 187662 994472
rect 191760 994362 191788 995438
rect 192496 995353 192524 995438
rect 193140 995382 193168 995438
rect 192944 995376 192996 995382
rect 192482 995344 192538 995353
rect 192482 995279 192538 995288
rect 192942 995344 192944 995353
rect 193128 995376 193180 995382
rect 192996 995344 192998 995353
rect 193128 995318 193180 995324
rect 192942 995279 192998 995288
rect 194336 995246 194364 995438
rect 194888 995330 194916 995454
rect 194520 995302 194916 995330
rect 195164 995438 195284 995466
rect 194140 995240 194192 995246
rect 194140 995182 194192 995188
rect 194324 995240 194376 995246
rect 194324 995182 194376 995188
rect 194152 995058 194180 995182
rect 194520 995058 194548 995302
rect 194152 995030 194548 995058
rect 191748 994356 191800 994362
rect 191748 994298 191800 994304
rect 186504 994288 186556 994294
rect 186504 994230 186556 994236
rect 184940 994152 184992 994158
rect 184940 994094 184992 994100
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 170864 993676 170916 993682
rect 170864 993618 170916 993624
rect 164884 990888 164936 990894
rect 164884 990830 164936 990836
rect 170772 990888 170824 990894
rect 170772 990830 170824 990836
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 154500 983620 154528 985662
rect 170784 983620 170812 990830
rect 186516 983634 186544 994230
rect 195164 993818 195192 995438
rect 195532 995246 195560 998378
rect 195704 997688 195756 997694
rect 195704 997630 195756 997636
rect 195716 996441 195744 997630
rect 195702 996432 195758 996441
rect 195702 996367 195758 996376
rect 195704 996260 195756 996266
rect 195704 996202 195756 996208
rect 195520 995240 195572 995246
rect 195520 995182 195572 995188
rect 195152 993812 195204 993818
rect 195152 993754 195204 993760
rect 195716 993682 195744 996202
rect 195900 995353 195928 1001778
rect 196624 998708 196676 998714
rect 196624 998650 196676 998656
rect 196072 997824 196124 997830
rect 196072 997766 196124 997772
rect 196084 995382 196112 997766
rect 196072 995376 196124 995382
rect 195886 995344 195942 995353
rect 196072 995318 196124 995324
rect 195886 995279 195942 995288
rect 196636 994158 196664 998650
rect 196808 998300 196860 998306
rect 196808 998242 196860 998248
rect 196624 994152 196676 994158
rect 196624 994094 196676 994100
rect 196820 993993 196848 998242
rect 198384 997830 198412 1005994
rect 203340 1002244 203392 1002250
rect 203340 1002186 203392 1002192
rect 202694 1002008 202750 1002017
rect 202694 1001943 202696 1001952
rect 202748 1001943 202750 1001952
rect 202696 1001914 202748 1001920
rect 200856 998572 200908 998578
rect 200856 998514 200908 998520
rect 199384 998096 199436 998102
rect 199384 998038 199436 998044
rect 198372 997824 198424 997830
rect 198372 997766 198424 997772
rect 197360 996940 197412 996946
rect 197360 996882 197412 996888
rect 197372 995518 197400 996882
rect 199396 996402 199424 998038
rect 200672 997960 200724 997966
rect 200670 997928 200672 997937
rect 200724 997928 200726 997937
rect 200670 997863 200726 997872
rect 200868 997754 200896 998514
rect 202694 998336 202750 998345
rect 202694 998271 202696 998280
rect 202748 998271 202750 998280
rect 202696 998242 202748 998248
rect 202144 998164 202196 998170
rect 202144 998106 202196 998112
rect 201868 998096 201920 998102
rect 201866 998064 201868 998073
rect 201920 998064 201922 998073
rect 201866 997999 201922 998008
rect 201040 997892 201092 997898
rect 201040 997834 201092 997840
rect 201052 997754 201080 997834
rect 200776 997726 200896 997754
rect 200960 997726 201080 997754
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 199384 996396 199436 996402
rect 199384 996338 199436 996344
rect 200776 995625 200804 997726
rect 200960 996946 200988 997726
rect 200948 996940 201000 996946
rect 200948 996882 201000 996888
rect 200948 996328 201000 996334
rect 200948 996270 201000 996276
rect 200762 995616 200818 995625
rect 200762 995551 200818 995560
rect 197360 995512 197412 995518
rect 197360 995454 197412 995460
rect 200960 994974 200988 996270
rect 202156 995110 202184 998106
rect 202328 998028 202380 998034
rect 202328 997970 202380 997976
rect 202340 995897 202368 997970
rect 202326 995888 202382 995897
rect 202326 995823 202382 995832
rect 202144 995104 202196 995110
rect 202144 995046 202196 995052
rect 200948 994968 201000 994974
rect 200948 994910 201000 994916
rect 203352 994537 203380 1002186
rect 203522 1002144 203578 1002153
rect 203522 1002079 203524 1002088
rect 203576 1002079 203578 1002088
rect 203524 1002050 203576 1002056
rect 204168 1001972 204220 1001978
rect 204168 1001914 204220 1001920
rect 203890 998608 203946 998617
rect 203890 998543 203892 998552
rect 203944 998543 203946 998552
rect 203892 998514 203944 998520
rect 204180 998442 204208 1001914
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 204168 998436 204220 998442
rect 204168 998378 204220 998384
rect 204718 998064 204774 998073
rect 204718 997999 204720 998008
rect 204772 997999 204774 998008
rect 204720 997970 204772 997976
rect 203522 997928 203578 997937
rect 203522 997863 203524 997872
rect 203576 997863 203578 997872
rect 203524 997834 203576 997840
rect 204916 997286 204944 1006266
rect 210422 1006224 210478 1006233
rect 210422 1006159 210424 1006168
rect 210476 1006159 210478 1006168
rect 228364 1006188 228416 1006194
rect 210424 1006130 210476 1006136
rect 228364 1006130 228416 1006136
rect 247040 1006188 247092 1006194
rect 247040 1006130 247092 1006136
rect 208398 1006088 208454 1006097
rect 208398 1006023 208400 1006032
rect 208452 1006023 208454 1006032
rect 208400 1005994 208452 1006000
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 207570 1004864 207626 1004873
rect 211250 1004864 211306 1004873
rect 207570 1004799 207572 1004808
rect 207624 1004799 207626 1004808
rect 209780 1004828 209832 1004834
rect 207572 1004770 207624 1004776
rect 211250 1004799 211252 1004808
rect 209780 1004770 209832 1004776
rect 211304 1004799 211306 1004808
rect 211252 1004770 211304 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 209228 1004634 209280 1004640
rect 206374 1002280 206430 1002289
rect 206374 1002215 206376 1002224
rect 206428 1002215 206430 1002224
rect 206376 1002186 206428 1002192
rect 206742 1002144 206798 1002153
rect 206742 1002079 206744 1002088
rect 206796 1002079 206798 1002088
rect 208400 1002108 208452 1002114
rect 206744 1002050 206796 1002056
rect 208400 1002050 208452 1002056
rect 205546 1002008 205602 1002017
rect 207202 1002008 207258 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 206284 1001972 206336 1001978
rect 205548 1001914 205600 1001920
rect 206284 1001914 206336 1001920
rect 207032 1001966 207202 1001994
rect 205546 998200 205602 998209
rect 205546 998135 205548 998144
rect 205600 998135 205602 998144
rect 205548 998106 205600 998112
rect 204904 997280 204956 997286
rect 204904 997222 204956 997228
rect 206296 996334 206324 1001914
rect 206284 996328 206336 996334
rect 206284 996270 206336 996276
rect 207032 994809 207060 1001966
rect 207202 1001943 207258 1001952
rect 207570 1002008 207626 1002017
rect 207570 1001943 207572 1001952
rect 207624 1001943 207626 1001952
rect 207572 1001914 207624 1001920
rect 207018 994800 207074 994809
rect 207018 994735 207074 994744
rect 203338 994528 203394 994537
rect 203338 994463 203394 994472
rect 197360 994356 197412 994362
rect 197360 994298 197412 994304
rect 196806 993984 196862 993993
rect 196806 993919 196862 993928
rect 195704 993676 195756 993682
rect 195704 993618 195756 993624
rect 197372 992934 197400 994298
rect 208412 994265 208440 1002050
rect 209792 997762 209820 1004770
rect 211160 1004692 211212 1004698
rect 211160 1004634 211212 1004640
rect 210882 1002416 210938 1002425
rect 210882 1002351 210884 1002360
rect 210936 1002351 210938 1002360
rect 210884 1002322 210936 1002328
rect 210882 1002144 210938 1002153
rect 210882 1002079 210884 1002088
rect 210936 1002079 210938 1002088
rect 210884 1002050 210936 1002056
rect 209780 997756 209832 997762
rect 209780 997698 209832 997704
rect 211172 996130 211200 1004634
rect 211816 996130 211844 1004906
rect 215944 1004828 215996 1004834
rect 215944 1004770 215996 1004776
rect 212538 1004728 212594 1004737
rect 212538 1004663 212540 1004672
rect 212592 1004663 212594 1004672
rect 212540 1004634 212592 1004640
rect 213184 1002380 213236 1002386
rect 213184 1002322 213236 1002328
rect 212540 1002108 212592 1002114
rect 212540 1002050 212592 1002056
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212080 1001914 212132 1001920
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211804 996124 211856 996130
rect 211804 996066 211856 996072
rect 212552 995994 212580 1002050
rect 212540 995988 212592 995994
rect 212540 995930 212592 995936
rect 213196 995858 213224 1002322
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213184 995852 213236 995858
rect 213184 995794 213236 995800
rect 208398 994256 208454 994265
rect 208398 994191 208454 994200
rect 213932 993070 213960 1001914
rect 202880 993064 202932 993070
rect 202880 993006 202932 993012
rect 213920 993064 213972 993070
rect 213920 993006 213972 993012
rect 197360 992928 197412 992934
rect 197360 992870 197412 992876
rect 202892 983634 202920 993006
rect 215956 985998 215984 1004770
rect 217324 1004692 217376 1004698
rect 217324 1004634 217376 1004640
rect 217336 986678 217364 1004634
rect 228376 995382 228404 1006130
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 229006 997792 229062 997801
rect 229006 997727 229062 997736
rect 229374 997792 229430 997801
rect 229374 997727 229430 997736
rect 228822 997248 228878 997257
rect 228822 997183 228878 997192
rect 228364 995376 228416 995382
rect 228364 995318 228416 995324
rect 228836 993954 228864 997183
rect 229020 994974 229048 997727
rect 229190 997248 229246 997257
rect 229190 997183 229246 997192
rect 229008 994968 229060 994974
rect 229008 994910 229060 994916
rect 229204 994362 229232 997183
rect 229192 994356 229244 994362
rect 229192 994298 229244 994304
rect 228824 993948 228876 993954
rect 228824 993890 228876 993896
rect 229388 993682 229416 997727
rect 229756 995994 229784 1005994
rect 246580 997756 246632 997762
rect 246580 997698 246632 997704
rect 229744 995988 229796 995994
rect 229744 995930 229796 995936
rect 239586 995752 239642 995761
rect 239292 995710 239586 995738
rect 242070 995752 242126 995761
rect 241776 995710 242070 995738
rect 239586 995687 239642 995696
rect 242070 995687 242126 995696
rect 246212 995580 246264 995586
rect 246212 995522 246264 995528
rect 240046 995480 240102 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 994226 231624 995438
rect 231584 994220 231636 994226
rect 231584 994162 231636 994168
rect 232240 993818 232268 995438
rect 232884 995110 232912 995438
rect 234080 995438 234416 995466
rect 234968 995438 235304 995466
rect 235612 995438 235948 995466
rect 236256 995438 236592 995466
rect 232872 995104 232924 995110
rect 232872 995046 232924 995052
rect 234080 994362 234108 995438
rect 235276 994537 235304 995438
rect 235262 994528 235318 994537
rect 235262 994463 235318 994472
rect 234068 994356 234120 994362
rect 234068 994298 234120 994304
rect 235920 994090 235948 995438
rect 236564 994809 236592 995438
rect 238404 995438 238740 995466
rect 239936 995438 240046 995466
rect 236550 994800 236606 994809
rect 236550 994735 236606 994744
rect 237472 994220 237524 994226
rect 237472 994162 237524 994168
rect 235908 994084 235960 994090
rect 235908 994026 235960 994032
rect 237484 993818 237512 994162
rect 232228 993812 232280 993818
rect 232228 993754 232280 993760
rect 237472 993812 237524 993818
rect 237472 993754 237524 993760
rect 238404 993682 238432 995438
rect 243266 995480 243322 995489
rect 240580 995438 240916 995466
rect 242972 995438 243266 995466
rect 240046 995415 240102 995424
rect 240888 994265 240916 995438
rect 243616 995438 243952 995466
rect 243266 995415 243322 995424
rect 243924 995217 243952 995438
rect 244246 995246 244274 995452
rect 245456 995438 245608 995466
rect 245580 995382 245608 995438
rect 245292 995376 245344 995382
rect 245292 995318 245344 995324
rect 245568 995376 245620 995382
rect 245568 995318 245620 995324
rect 244234 995240 244286 995246
rect 243910 995208 243966 995217
rect 244234 995182 244286 995188
rect 243910 995143 243966 995152
rect 245304 994838 245332 995318
rect 246224 994974 246252 995522
rect 246592 995382 246620 997698
rect 247052 995761 247080 1006130
rect 247408 998436 247460 998442
rect 247408 998378 247460 998384
rect 247224 998300 247276 998306
rect 247224 998242 247276 998248
rect 247038 995752 247094 995761
rect 247038 995687 247094 995696
rect 246764 995444 246816 995450
rect 246764 995386 246816 995392
rect 246580 995376 246632 995382
rect 246580 995318 246632 995324
rect 246212 994968 246264 994974
rect 246212 994910 246264 994916
rect 245292 994832 245344 994838
rect 245292 994774 245344 994780
rect 243176 994764 243228 994770
rect 243176 994706 243228 994712
rect 240874 994256 240930 994265
rect 240874 994191 240930 994200
rect 243188 993818 243216 994706
rect 246776 994537 246804 995386
rect 247236 995246 247264 998242
rect 247224 995240 247276 995246
rect 247420 995217 247448 998378
rect 249064 998164 249116 998170
rect 249064 998106 249116 998112
rect 247776 997892 247828 997898
rect 247776 997834 247828 997840
rect 247592 996260 247644 996266
rect 247592 996202 247644 996208
rect 247224 995182 247276 995188
rect 247406 995208 247462 995217
rect 247406 995143 247462 995152
rect 247604 994838 247632 996202
rect 247592 994832 247644 994838
rect 247592 994774 247644 994780
rect 246762 994528 246818 994537
rect 246762 994463 246818 994472
rect 247788 993818 247816 997834
rect 249076 994265 249104 998106
rect 249260 996033 249288 1006266
rect 255318 1006224 255374 1006233
rect 255318 1006159 255320 1006168
rect 255372 1006159 255374 1006168
rect 261850 1006224 261906 1006233
rect 261850 1006159 261852 1006168
rect 255320 1006130 255372 1006136
rect 261904 1006159 261906 1006168
rect 279424 1006188 279476 1006194
rect 261852 1006130 261904 1006136
rect 279424 1006130 279476 1006136
rect 252466 1006088 252522 1006097
rect 251088 1006052 251140 1006058
rect 252466 1006023 252468 1006032
rect 251088 1005994 251140 1006000
rect 252520 1006023 252522 1006032
rect 260194 1006088 260250 1006097
rect 260194 1006023 260196 1006032
rect 252468 1005994 252520 1006000
rect 260248 1006023 260250 1006032
rect 260196 1005994 260248 1006000
rect 251100 998306 251128 1005994
rect 263046 1005136 263102 1005145
rect 263046 1005071 263048 1005080
rect 263100 1005071 263102 1005080
rect 268384 1005100 268436 1005106
rect 263048 1005042 263100 1005048
rect 268384 1005042 268436 1005048
rect 256146 1002688 256202 1002697
rect 253480 1002652 253532 1002658
rect 256146 1002623 256148 1002632
rect 253480 1002594 253532 1002600
rect 256200 1002623 256202 1002632
rect 261022 1002688 261078 1002697
rect 261022 1002623 261024 1002632
rect 256148 1002594 256200 1002600
rect 261076 1002623 261078 1002632
rect 264244 1002652 264296 1002658
rect 261024 1002594 261076 1002600
rect 264244 1002594 264296 1002600
rect 251916 1002516 251968 1002522
rect 251916 1002458 251968 1002464
rect 251456 1002244 251508 1002250
rect 251456 1002186 251508 1002192
rect 251088 998300 251140 998306
rect 251088 998242 251140 998248
rect 250444 998028 250496 998034
rect 250444 997970 250496 997976
rect 250456 997257 250484 997970
rect 250442 997248 250498 997257
rect 250442 997183 250498 997192
rect 249246 996024 249302 996033
rect 249246 995959 249302 995968
rect 251468 994809 251496 1002186
rect 251928 996418 251956 1002458
rect 253020 1002380 253072 1002386
rect 253020 1002322 253072 1002328
rect 252466 997928 252522 997937
rect 252466 997863 252468 997872
rect 252520 997863 252522 997872
rect 252468 997834 252520 997840
rect 251652 996390 251956 996418
rect 251652 996305 251680 996390
rect 251638 996296 251694 996305
rect 251638 996231 251694 996240
rect 251454 994800 251510 994809
rect 251454 994735 251510 994744
rect 249062 994256 249118 994265
rect 249062 994191 249118 994200
rect 253032 994090 253060 1002322
rect 253294 998064 253350 998073
rect 253294 997999 253296 998008
rect 253348 997999 253350 998008
rect 253296 997970 253348 997976
rect 253492 995450 253520 1002594
rect 255318 1002552 255374 1002561
rect 255318 1002487 255320 1002496
rect 255372 1002487 255374 1002496
rect 255320 1002458 255372 1002464
rect 261024 1002448 261076 1002454
rect 256146 1002416 256202 1002425
rect 256146 1002351 256148 1002360
rect 256200 1002351 256202 1002360
rect 261022 1002416 261024 1002425
rect 263692 1002448 263744 1002454
rect 261076 1002416 261078 1002425
rect 263692 1002390 263744 1002396
rect 261022 1002351 261078 1002360
rect 256148 1002322 256200 1002328
rect 262680 1002312 262732 1002318
rect 254490 1002280 254546 1002289
rect 254490 1002215 254492 1002224
rect 254544 1002215 254546 1002224
rect 262678 1002280 262680 1002289
rect 262732 1002280 262734 1002289
rect 262678 1002215 262734 1002224
rect 254492 1002186 254544 1002192
rect 263508 1002040 263560 1002046
rect 263506 1002008 263508 1002017
rect 263560 1002008 263562 1002017
rect 263506 1001943 263562 1001952
rect 256700 999184 256752 999190
rect 258172 999184 258224 999190
rect 256700 999126 256752 999132
rect 258170 999152 258172 999161
rect 258224 999152 258226 999161
rect 253662 998200 253718 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 256332 998164 256384 998170
rect 253664 998106 253716 998112
rect 256332 998106 256384 998112
rect 254584 997960 254636 997966
rect 254584 997902 254636 997908
rect 253480 995444 253532 995450
rect 253480 995386 253532 995392
rect 253204 994764 253256 994770
rect 253204 994706 253256 994712
rect 253020 994084 253072 994090
rect 253020 994026 253072 994032
rect 253216 993954 253244 994706
rect 254596 994226 254624 997902
rect 254952 997824 255004 997830
rect 254780 997772 254952 997778
rect 254780 997766 255004 997772
rect 254780 997762 254992 997766
rect 254768 997756 254992 997762
rect 254820 997750 254992 997756
rect 254768 997698 254820 997704
rect 256344 995586 256372 998106
rect 256516 997960 256568 997966
rect 256514 997928 256516 997937
rect 256568 997928 256570 997937
rect 256514 997863 256570 997872
rect 256332 995580 256384 995586
rect 256332 995522 256384 995528
rect 256712 994362 256740 999126
rect 258170 999087 258226 999096
rect 258998 998472 259054 998481
rect 258998 998407 259000 998416
rect 259052 998407 259054 998416
rect 259000 998378 259052 998384
rect 257342 998200 257398 998209
rect 257342 998135 257344 998144
rect 257396 998135 257398 998144
rect 257344 998106 257396 998112
rect 257344 997960 257396 997966
rect 259000 997960 259052 997966
rect 257344 997902 257396 997908
rect 258998 997928 259000 997937
rect 259828 997960 259880 997966
rect 259052 997928 259054 997937
rect 256976 997824 257028 997830
rect 256974 997792 256976 997801
rect 257028 997792 257030 997801
rect 256974 997727 257030 997736
rect 257356 995110 257384 997902
rect 258998 997863 259054 997872
rect 259826 997928 259828 997937
rect 262312 997960 262364 997966
rect 259880 997928 259882 997937
rect 262312 997902 262364 997908
rect 259826 997863 259882 997872
rect 258172 997824 258224 997830
rect 258170 997792 258172 997801
rect 259460 997824 259512 997830
rect 258224 997792 258226 997801
rect 260196 997824 260248 997830
rect 259460 997766 259512 997772
rect 260194 997792 260196 997801
rect 260248 997792 260250 997801
rect 258170 997727 258226 997736
rect 257344 995104 257396 995110
rect 257344 995046 257396 995052
rect 259472 994770 259500 997766
rect 261850 997792 261906 997801
rect 260194 997727 260250 997736
rect 261312 997736 261850 997754
rect 261312 997727 261906 997736
rect 261312 997726 261892 997727
rect 261312 995858 261340 997726
rect 262324 995994 262352 997902
rect 262496 997824 262548 997830
rect 262496 997766 262548 997772
rect 262508 996130 262536 997766
rect 263704 996266 263732 1002390
rect 263876 1002176 263928 1002182
rect 263874 1002144 263876 1002153
rect 263928 1002144 263930 1002153
rect 263874 1002079 263930 1002088
rect 263692 996260 263744 996266
rect 263692 996202 263744 996208
rect 262496 996124 262548 996130
rect 262496 996066 262548 996072
rect 264256 995994 264284 1002594
rect 265808 1002312 265860 1002318
rect 265808 1002254 265860 1002260
rect 265624 1002040 265676 1002046
rect 265624 1001982 265676 1001988
rect 262312 995988 262364 995994
rect 262312 995930 262364 995936
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 261300 995852 261352 995858
rect 261300 995794 261352 995800
rect 259460 994764 259512 994770
rect 259460 994706 259512 994712
rect 256700 994356 256752 994362
rect 256700 994298 256752 994304
rect 254584 994220 254636 994226
rect 254584 994162 254636 994168
rect 253204 993948 253256 993954
rect 253204 993890 253256 993896
rect 243176 993812 243228 993818
rect 243176 993754 243228 993760
rect 247776 993812 247828 993818
rect 247776 993754 247828 993760
rect 229376 993676 229428 993682
rect 229376 993618 229428 993624
rect 238392 993676 238444 993682
rect 238392 993618 238444 993624
rect 251456 992928 251508 992934
rect 251456 992870 251508 992876
rect 217324 986672 217376 986678
rect 217324 986614 217376 986620
rect 219440 986672 219492 986678
rect 219440 986614 219492 986620
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 186516 983606 186990 983634
rect 202892 983606 203182 983634
rect 219452 983620 219480 986614
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 992870
rect 265636 990894 265664 1001982
rect 265820 996130 265848 1002254
rect 267004 1002176 267056 1002182
rect 267004 1002118 267056 1002124
rect 265808 996124 265860 996130
rect 265808 996066 265860 996072
rect 267016 991506 267044 1002118
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1005042
rect 279436 995081 279464 1006130
rect 280804 1006052 280856 1006058
rect 280804 1005994 280856 1006000
rect 298744 1006052 298796 1006058
rect 298744 1005994 298796 1006000
rect 280816 995353 280844 1005994
rect 298756 1001894 298784 1005994
rect 298756 1001866 298876 1001894
rect 298466 999152 298522 999161
rect 298466 999087 298522 999096
rect 298282 998472 298338 998481
rect 298282 998407 298338 998416
rect 298098 998064 298154 998073
rect 298098 997999 298154 998008
rect 282734 995752 282790 995761
rect 290646 995752 290702 995761
rect 282790 995710 282854 995738
rect 290306 995710 290646 995738
rect 282734 995687 282790 995696
rect 294786 995752 294842 995761
rect 294538 995710 294786 995738
rect 290646 995687 290702 995696
rect 294786 995687 294842 995696
rect 295062 995752 295118 995761
rect 298112 995738 298140 997999
rect 298296 997914 298324 998407
rect 295118 995710 295182 995738
rect 297836 995710 298140 995738
rect 298204 997886 298324 997914
rect 295062 995687 295118 995696
rect 290462 995616 290518 995625
rect 290518 995574 290858 995602
rect 290462 995551 290518 995560
rect 280802 995344 280858 995353
rect 280802 995279 280858 995288
rect 283484 995246 283512 995452
rect 283472 995240 283524 995246
rect 283472 995182 283524 995188
rect 279422 995072 279478 995081
rect 279422 995007 279478 995016
rect 284128 994974 284156 995452
rect 285968 995110 285996 995452
rect 285956 995104 286008 995110
rect 285956 995046 286008 995052
rect 284116 994968 284168 994974
rect 284116 994910 284168 994916
rect 286520 994226 286548 995452
rect 287164 994838 287192 995452
rect 287822 995438 288112 995466
rect 291502 995438 291884 995466
rect 292146 995438 292528 995466
rect 287152 994832 287204 994838
rect 287152 994774 287204 994780
rect 287704 994628 287756 994634
rect 287704 994570 287756 994576
rect 287716 994362 287744 994570
rect 288084 994537 288112 995438
rect 291856 994809 291884 995438
rect 292304 995376 292356 995382
rect 292302 995344 292304 995353
rect 292500 995353 292528 995438
rect 292356 995344 292358 995353
rect 292302 995279 292358 995288
rect 292486 995344 292542 995353
rect 292486 995279 292542 995288
rect 291842 994800 291898 994809
rect 291842 994735 291898 994744
rect 289544 994696 289596 994702
rect 289544 994638 289596 994644
rect 288070 994528 288126 994537
rect 288070 994463 288126 994472
rect 287704 994356 287756 994362
rect 287704 994298 287756 994304
rect 289556 994226 289584 994638
rect 293328 994537 293356 995452
rect 295826 995438 296208 995466
rect 297022 995438 297404 995466
rect 296180 995382 296208 995438
rect 295984 995376 296036 995382
rect 295706 995344 295762 995353
rect 295984 995318 296036 995324
rect 296168 995376 296220 995382
rect 296718 995344 296774 995353
rect 296168 995318 296220 995324
rect 295706 995279 295762 995288
rect 295720 995058 295748 995279
rect 295996 995194 296024 995318
rect 296364 995302 296718 995330
rect 296364 995194 296392 995302
rect 297376 995330 297404 995438
rect 297836 995330 297864 995710
rect 298204 995602 298232 997886
rect 297376 995302 297864 995330
rect 297928 995574 298232 995602
rect 296718 995279 296774 995288
rect 297928 995194 297956 995574
rect 298480 995382 298508 999087
rect 298650 996704 298706 996713
rect 298650 996639 298706 996648
rect 298468 995376 298520 995382
rect 298468 995318 298520 995324
rect 295996 995166 296392 995194
rect 296640 995166 297956 995194
rect 296640 995058 296668 995166
rect 295720 995030 296668 995058
rect 296720 994832 296772 994838
rect 296772 994780 296852 994786
rect 296720 994774 296852 994780
rect 296732 994758 296852 994774
rect 293314 994528 293370 994537
rect 293314 994463 293370 994472
rect 296824 994430 296852 994758
rect 298664 994537 298692 996639
rect 298650 994528 298706 994537
rect 298650 994463 298706 994472
rect 296812 994424 296864 994430
rect 296812 994366 296864 994372
rect 298848 994294 298876 1001866
rect 298940 996010 298968 1006266
rect 299480 1006188 299532 1006194
rect 299480 1006130 299532 1006136
rect 299492 1001994 299520 1006130
rect 299662 1002688 299718 1002697
rect 299662 1002623 299718 1002632
rect 299308 1001966 299520 1001994
rect 299308 997801 299336 1001966
rect 299294 997792 299350 997801
rect 299112 997756 299164 997762
rect 299294 997727 299350 997736
rect 299112 997698 299164 997704
rect 299124 997257 299152 997698
rect 299110 997248 299166 997257
rect 299110 997183 299166 997192
rect 299676 996985 299704 1002623
rect 299662 996976 299718 996985
rect 299662 996911 299718 996920
rect 299386 996432 299442 996441
rect 299386 996367 299388 996376
rect 299440 996367 299442 996376
rect 299388 996338 299440 996344
rect 298940 995994 299336 996010
rect 298940 995988 299348 995994
rect 298940 995982 299296 995988
rect 299296 995930 299348 995936
rect 300136 995246 300164 1006538
rect 359740 1006528 359792 1006534
rect 359738 1006496 359740 1006505
rect 370504 1006528 370556 1006534
rect 359792 1006496 359794 1006505
rect 370504 1006470 370556 1006476
rect 359738 1006431 359794 1006440
rect 358542 1006360 358598 1006369
rect 311808 1006324 311860 1006330
rect 358542 1006295 358544 1006304
rect 311808 1006266 311860 1006272
rect 358596 1006295 358598 1006304
rect 358544 1006266 358596 1006272
rect 306102 1006224 306158 1006233
rect 306102 1006159 306104 1006168
rect 306156 1006159 306158 1006168
rect 306104 1006130 306156 1006136
rect 311820 1006097 311848 1006266
rect 361394 1006224 361450 1006233
rect 361394 1006159 361396 1006168
rect 361448 1006159 361450 1006168
rect 367008 1006188 367060 1006194
rect 361396 1006130 361448 1006136
rect 367008 1006130 367060 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301504 1002108 301556 1002114
rect 301504 1002050 301556 1002056
rect 301516 1001894 301544 1002050
rect 301332 1001866 301544 1001894
rect 300124 995240 300176 995246
rect 300124 995182 300176 995188
rect 301332 994566 301360 1001866
rect 301700 999161 301728 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 354862 1006088 354918 1006097
rect 314658 1006023 314660 1006032
rect 304080 1005994 304132 1006000
rect 314712 1006023 314714 1006032
rect 319444 1006052 319496 1006058
rect 314660 1005994 314712 1006000
rect 354862 1006023 354918 1006032
rect 319444 1005994 319496 1006000
rect 304080 1005848 304132 1005854
rect 304078 1005816 304080 1005825
rect 304132 1005816 304134 1005825
rect 304078 1005751 304134 1005760
rect 313830 1005000 313886 1005009
rect 313830 1004935 313832 1004944
rect 313884 1004935 313886 1004944
rect 316040 1004964 316092 1004970
rect 313832 1004906 313884 1004912
rect 316040 1004906 316092 1004912
rect 314658 1004864 314714 1004873
rect 314658 1004799 314660 1004808
rect 314712 1004799 314714 1004808
rect 314660 1004770 314712 1004776
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 303250 1002688 303306 1002697
rect 303250 1002623 303252 1002632
rect 303304 1002623 303306 1002632
rect 306930 1002688 306986 1002697
rect 306930 1002623 306932 1002632
rect 303252 1002594 303304 1002600
rect 306984 1002623 306986 1002632
rect 306932 1002594 306984 1002600
rect 304906 1002144 304962 1002153
rect 304906 1002079 304908 1002088
rect 304960 1002079 304962 1002088
rect 304908 1002050 304960 1002056
rect 310150 1002008 310206 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 311900 1001972 311952 1001978
rect 310152 1001914 310204 1001920
rect 311900 1001914 311952 1001920
rect 301686 999152 301742 999161
rect 301686 999087 301742 999096
rect 303068 998640 303120 998646
rect 308956 998640 309008 998646
rect 303068 998582 303120 998588
rect 308954 998608 308956 998617
rect 309008 998608 309010 998617
rect 303080 998073 303108 998582
rect 308954 998543 309010 998552
rect 303252 998504 303304 998510
rect 303250 998472 303252 998481
rect 305276 998504 305328 998510
rect 303304 998472 303306 998481
rect 303250 998407 303306 998416
rect 305274 998472 305276 998481
rect 305328 998472 305330 998481
rect 305274 998407 305330 998416
rect 307298 998336 307354 998345
rect 304264 998300 304316 998306
rect 307298 998271 307300 998280
rect 304264 998242 304316 998248
rect 307352 998271 307354 998280
rect 307300 998242 307352 998248
rect 303066 998064 303122 998073
rect 302884 998028 302936 998034
rect 303066 997999 303122 998008
rect 302884 997970 302936 997976
rect 301502 996160 301558 996169
rect 301502 996095 301558 996104
rect 301516 995625 301544 996095
rect 301502 995616 301558 995625
rect 301502 995551 301558 995560
rect 302896 994809 302924 997970
rect 303252 996736 303304 996742
rect 303250 996704 303252 996713
rect 303304 996704 303306 996713
rect 303250 996639 303306 996648
rect 302882 994800 302938 994809
rect 302882 994735 302938 994744
rect 301320 994560 301372 994566
rect 301320 994502 301372 994508
rect 304276 994430 304304 998242
rect 306930 998200 306986 998209
rect 304448 998164 304500 998170
rect 306930 998135 306932 998144
rect 304448 998106 304500 998112
rect 306984 998135 306986 998144
rect 306932 998106 306984 998112
rect 304460 996742 304488 998106
rect 306102 998064 306158 998073
rect 308954 998064 309010 998073
rect 306102 997999 306104 998008
rect 306156 997999 306158 998008
rect 307024 998028 307076 998034
rect 306104 997970 306156 997976
rect 308954 997999 308956 998008
rect 307024 997970 307076 997976
rect 309008 997999 309010 998008
rect 308956 997970 309008 997976
rect 305644 997892 305696 997898
rect 305644 997834 305696 997840
rect 304448 996736 304500 996742
rect 304448 996678 304500 996684
rect 305656 994702 305684 997834
rect 307036 995625 307064 997970
rect 307758 997928 307814 997937
rect 310610 997928 310666 997937
rect 307758 997863 307760 997872
rect 307812 997863 307814 997872
rect 308404 997892 308456 997898
rect 307760 997834 307812 997840
rect 310610 997863 310612 997872
rect 308404 997834 308456 997840
rect 310664 997863 310666 997872
rect 310612 997834 310664 997840
rect 307022 995616 307078 995625
rect 307022 995551 307078 995560
rect 308416 994974 308444 997834
rect 309782 997792 309838 997801
rect 309152 997736 309782 997754
rect 311912 997762 311940 1001914
rect 309152 997727 309838 997736
rect 311900 997756 311952 997762
rect 309152 997726 309824 997727
rect 309152 995110 309180 997726
rect 311900 997698 311952 997704
rect 316052 996130 316080 1004906
rect 316684 1004828 316736 1004834
rect 316684 1004770 316736 1004776
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 309140 995104 309192 995110
rect 309140 995046 309192 995052
rect 308404 994968 308456 994974
rect 308404 994910 308456 994916
rect 305644 994696 305696 994702
rect 305644 994638 305696 994644
rect 304264 994424 304316 994430
rect 304264 994366 304316 994372
rect 298836 994288 298888 994294
rect 298836 994230 298888 994236
rect 316406 994256 316462 994265
rect 286508 994220 286560 994226
rect 286508 994162 286560 994168
rect 289544 994220 289596 994226
rect 316406 994191 316462 994200
rect 289544 994162 289596 994168
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994191
rect 316696 992934 316724 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316684 992928 316736 992934
rect 316684 992870 316736 992876
rect 318076 991506 318104 1004634
rect 318064 991500 318116 991506
rect 318064 991442 318116 991448
rect 319456 990146 319484 1005994
rect 354876 1005310 354904 1006023
rect 363420 1005984 363472 1005990
rect 363418 1005952 363420 1005961
rect 363472 1005952 363474 1005961
rect 363418 1005887 363474 1005896
rect 367020 1005718 367048 1006130
rect 367008 1005712 367060 1005718
rect 367008 1005654 367060 1005660
rect 360568 1005576 360620 1005582
rect 360566 1005544 360568 1005553
rect 360620 1005544 360622 1005553
rect 360566 1005479 360622 1005488
rect 358544 1005440 358596 1005446
rect 358542 1005408 358544 1005417
rect 358596 1005408 358598 1005417
rect 358542 1005343 358598 1005352
rect 354864 1005304 354916 1005310
rect 354864 1005246 354916 1005252
rect 356518 1005136 356574 1005145
rect 354404 1005100 354456 1005106
rect 356518 1005071 356520 1005080
rect 354404 1005042 354456 1005048
rect 356572 1005071 356574 1005080
rect 361394 1005136 361450 1005145
rect 361394 1005071 361396 1005080
rect 356520 1005042 356572 1005048
rect 361448 1005071 361450 1005080
rect 364892 1005100 364944 1005106
rect 361396 1005042 361448 1005048
rect 364892 1005042 364944 1005048
rect 353208 1004964 353260 1004970
rect 353208 1004906 353260 1004912
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998578 351868 1001914
rect 353220 1001230 353248 1004906
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998572 351880 998578
rect 351828 998514 351880 998520
rect 354416 998442 354444 1005042
rect 355690 1005000 355746 1005009
rect 355690 1004935 355692 1004944
rect 355744 1004935 355746 1004944
rect 355692 1004906 355744 1004912
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 356888 1003944 356940 1003950
rect 356886 1003912 356888 1003921
rect 356940 1003912 356942 1003921
rect 356886 1003847 356942 1003856
rect 359370 1002552 359426 1002561
rect 358728 1002516 358780 1002522
rect 359370 1002487 359372 1002496
rect 358728 1002458 358780 1002464
rect 359424 1002487 359426 1002496
rect 359372 1002458 359424 1002464
rect 357346 1002416 357402 1002425
rect 357346 1002351 357348 1002360
rect 357400 1002351 357402 1002360
rect 357348 1002322 357400 1002328
rect 357714 1002280 357770 1002289
rect 357714 1002215 357716 1002224
rect 357768 1002215 357770 1002224
rect 357716 1002186 357768 1002192
rect 355690 1002008 355746 1002017
rect 355690 1001943 355692 1001952
rect 355744 1001943 355746 1001952
rect 356704 1001972 356756 1001978
rect 355692 1001914 355744 1001920
rect 356704 1001914 356756 1001920
rect 354404 998436 354456 998442
rect 354404 998378 354456 998384
rect 356716 994498 356744 1001914
rect 358740 995042 358768 1002458
rect 359464 1002380 359516 1002386
rect 359464 1002322 359516 1002328
rect 359476 1001366 359504 1002322
rect 360844 1002244 360896 1002250
rect 360844 1002186 360896 1002192
rect 360566 1002144 360622 1002153
rect 360566 1002079 360568 1002088
rect 360620 1002079 360622 1002088
rect 360568 1002050 360620 1002056
rect 360198 1002008 360254 1002017
rect 360198 1001943 360200 1001952
rect 360252 1001943 360254 1001952
rect 360200 1001914 360252 1001920
rect 359464 1001360 359516 1001366
rect 359464 1001302 359516 1001308
rect 360856 997626 360884 1002186
rect 363604 1002108 363656 1002114
rect 363604 1002050 363656 1002056
rect 362224 1001972 362276 1001978
rect 362224 1001914 362276 1001920
rect 360844 997620 360896 997626
rect 360844 997562 360896 997568
rect 360200 996396 360252 996402
rect 360200 996338 360252 996344
rect 358728 995036 358780 995042
rect 358728 994978 358780 994984
rect 356704 994492 356756 994498
rect 356704 994434 356756 994440
rect 360212 994294 360240 996338
rect 362236 995314 362264 1001914
rect 362224 995308 362276 995314
rect 362224 995250 362276 995256
rect 363616 994906 363644 1002050
rect 364904 995858 364932 1005042
rect 365260 1004828 365312 1004834
rect 365260 1004770 365312 1004776
rect 365076 1002312 365128 1002318
rect 365074 1002280 365076 1002289
rect 365128 1002280 365130 1002289
rect 365074 1002215 365130 1002224
rect 365076 1002040 365128 1002046
rect 365074 1002008 365076 1002017
rect 365128 1002008 365130 1002017
rect 365074 1001943 365130 1001952
rect 365272 997762 365300 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365904 1002176 365956 1002182
rect 365902 1002144 365904 1002153
rect 365956 1002144 365958 1002153
rect 365902 1002079 365958 1002088
rect 365260 997756 365312 997762
rect 365260 997698 365312 997704
rect 366376 995994 366404 1004634
rect 367928 1002312 367980 1002318
rect 367928 1002254 367980 1002260
rect 367744 1002040 367796 1002046
rect 367744 1001982 367796 1001988
rect 366364 995988 366416 995994
rect 366364 995930 366416 995936
rect 364892 995852 364944 995858
rect 364892 995794 364944 995800
rect 363604 994900 363656 994906
rect 363604 994842 363656 994848
rect 360200 994288 360252 994294
rect 360200 994230 360252 994236
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 349160 991500 349212 991506
rect 349160 991442 349212 991448
rect 319444 990140 319496 990146
rect 319444 990082 319496 990088
rect 332968 990140 333020 990146
rect 332968 990082 333020 990088
rect 316420 983606 316802 983634
rect 332980 983620 333008 990082
rect 349172 983620 349200 991442
rect 364996 983634 365024 992870
rect 367756 991506 367784 1001982
rect 367940 992934 367968 1002254
rect 369124 1002176 369176 1002182
rect 369124 1002118 369176 1002124
rect 367928 992928 367980 992934
rect 367928 992870 367980 992876
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 369136 990146 369164 1002118
rect 370516 998850 370544 1006470
rect 370504 998844 370556 998850
rect 370504 998786 370556 998792
rect 371896 998306 371924 1006606
rect 422668 1006528 422720 1006534
rect 422668 1006470 422720 1006476
rect 426532 1006528 426584 1006534
rect 426532 1006470 426584 1006476
rect 431682 1006496 431738 1006505
rect 377404 1006324 377456 1006330
rect 377404 1006266 377456 1006272
rect 373264 1005440 373316 1005446
rect 373264 1005382 373316 1005388
rect 372712 1001360 372764 1001366
rect 372712 1001302 372764 1001308
rect 371884 998300 371936 998306
rect 371884 998242 371936 998248
rect 372528 997756 372580 997762
rect 372528 997698 372580 997704
rect 372344 997620 372396 997626
rect 372344 997562 372396 997568
rect 372356 996441 372384 997562
rect 372540 996985 372568 997698
rect 372526 996976 372582 996985
rect 372526 996911 372582 996920
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 372724 994634 372752 1001302
rect 372988 998300 373040 998306
rect 372988 998242 373040 998248
rect 373000 995081 373028 998242
rect 373276 996169 373304 1005382
rect 374644 1005304 374696 1005310
rect 374644 1005246 374696 1005252
rect 374656 998306 374684 1005246
rect 375380 1003944 375432 1003950
rect 375380 1003886 375432 1003892
rect 374644 998300 374696 998306
rect 374644 998242 374696 998248
rect 373262 996160 373318 996169
rect 373262 996095 373318 996104
rect 375392 995353 375420 1003886
rect 377416 997966 377444 1006266
rect 402244 1006188 402296 1006194
rect 402244 1006130 402296 1006136
rect 382924 1006052 382976 1006058
rect 382924 1005994 382976 1006000
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 380164 1005712 380216 1005718
rect 380164 1005654 380216 1005660
rect 378784 1005576 378836 1005582
rect 378784 1005518 378836 1005524
rect 378048 998844 378100 998850
rect 378048 998786 378100 998792
rect 377404 997960 377456 997966
rect 377404 997902 377456 997908
rect 375378 995344 375434 995353
rect 375378 995279 375434 995288
rect 372986 995072 373042 995081
rect 372986 995007 373042 995016
rect 372712 994628 372764 994634
rect 372712 994570 372764 994576
rect 378060 994537 378088 998786
rect 378796 997830 378824 1005518
rect 379152 998300 379204 998306
rect 379152 998242 379204 998248
rect 378784 997824 378836 997830
rect 378784 997766 378836 997772
rect 379164 994770 379192 998242
rect 380176 996713 380204 1005654
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 380162 996704 380218 996713
rect 380162 996639 380218 996648
rect 380912 995178 380940 1001166
rect 382280 998572 382332 998578
rect 382280 998514 382332 998520
rect 382292 996033 382320 998514
rect 382936 996130 382964 1005994
rect 399944 1001972 399996 1001978
rect 399944 1001914 399996 1001920
rect 383568 998436 383620 998442
rect 383568 998378 383620 998384
rect 383200 997960 383252 997966
rect 383200 997902 383252 997908
rect 382924 996124 382976 996130
rect 382924 996066 382976 996072
rect 382278 996024 382334 996033
rect 382278 995959 382334 995968
rect 383212 995586 383240 997902
rect 383384 997824 383436 997830
rect 383384 997766 383436 997772
rect 383396 997098 383424 997766
rect 383580 997257 383608 998378
rect 399956 997914 399984 1001914
rect 399956 997886 400168 997914
rect 399944 997756 399996 997762
rect 399944 997698 399996 997704
rect 383566 997248 383622 997257
rect 383566 997183 383622 997192
rect 383396 997070 383700 997098
rect 383474 996704 383530 996713
rect 383474 996639 383530 996648
rect 383200 995580 383252 995586
rect 383200 995522 383252 995528
rect 383488 995450 383516 996639
rect 383476 995444 383528 995450
rect 383476 995386 383528 995392
rect 383672 995330 383700 997070
rect 399956 996985 399984 997698
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 388166 995752 388222 995761
rect 388222 995710 388378 995738
rect 388166 995687 388222 995696
rect 385052 995586 385342 995602
rect 385040 995580 385342 995586
rect 385092 995574 385342 995580
rect 385040 995522 385092 995528
rect 392398 995480 392454 995489
rect 384316 995438 384698 995466
rect 385696 995450 385986 995466
rect 385684 995444 385986 995450
rect 384316 995330 384344 995438
rect 385736 995438 385986 995444
rect 385684 995386 385736 995392
rect 383672 995302 384344 995330
rect 387812 995314 387840 995452
rect 387800 995308 387852 995314
rect 387800 995250 387852 995256
rect 380900 995172 380952 995178
rect 380900 995114 380952 995120
rect 389008 995081 389036 995452
rect 389376 995438 389666 995466
rect 389376 995353 389404 995438
rect 389362 995344 389418 995353
rect 389362 995279 389418 995288
rect 388994 995072 389050 995081
rect 388994 995007 389050 995016
rect 379152 994764 379204 994770
rect 379152 994706 379204 994712
rect 392136 994537 392164 995452
rect 394974 995480 395030 995489
rect 392454 995438 392702 995466
rect 392398 995415 392454 995424
rect 393332 994634 393360 995452
rect 393320 994628 393372 994634
rect 393320 994570 393372 994576
rect 378046 994528 378102 994537
rect 378046 994463 378102 994472
rect 392122 994528 392178 994537
rect 393976 994498 394004 995452
rect 395030 995438 395186 995466
rect 396382 995438 396672 995466
rect 394974 995415 395030 995424
rect 396644 995382 396672 995438
rect 396632 995376 396684 995382
rect 396632 995318 396684 995324
rect 397012 994906 397040 995452
rect 397000 994900 397052 994906
rect 397000 994842 397052 994848
rect 397656 994770 397684 995452
rect 398852 995042 398880 995452
rect 400140 995382 400168 997886
rect 400876 995994 400904 1005994
rect 400864 995988 400916 995994
rect 400864 995930 400916 995936
rect 402256 995858 402284 1006130
rect 422680 1006097 422708 1006470
rect 425336 1006392 425388 1006398
rect 425336 1006334 425388 1006340
rect 422666 1006088 422722 1006097
rect 425348 1006058 425376 1006334
rect 425518 1006088 425574 1006097
rect 422666 1006023 422722 1006032
rect 425336 1006052 425388 1006058
rect 425518 1006023 425520 1006032
rect 425336 1005994 425388 1006000
rect 425572 1006023 425574 1006032
rect 425520 1005994 425572 1006000
rect 426346 1005816 426402 1005825
rect 426346 1005751 426348 1005760
rect 426400 1005751 426402 1005760
rect 426348 1005722 426400 1005728
rect 426348 1005576 426400 1005582
rect 426346 1005544 426348 1005553
rect 426400 1005544 426402 1005553
rect 426346 1005479 426402 1005488
rect 423496 1005304 423548 1005310
rect 423494 1005272 423496 1005281
rect 423548 1005272 423550 1005281
rect 423494 1005207 423550 1005216
rect 423494 1005000 423550 1005009
rect 422208 1004964 422260 1004970
rect 423494 1004935 423496 1004944
rect 422208 1004906 422260 1004912
rect 423548 1004935 423550 1004944
rect 423496 1004906 423548 1004912
rect 420828 1004828 420880 1004834
rect 420828 1004770 420880 1004776
rect 419448 1002108 419500 1002114
rect 419448 1002050 419500 1002056
rect 402244 995852 402296 995858
rect 402244 995794 402296 995800
rect 415950 995752 416006 995761
rect 415950 995687 416006 995696
rect 415964 995586 415992 995687
rect 415952 995580 416004 995586
rect 415952 995522 416004 995528
rect 400128 995376 400180 995382
rect 400128 995318 400180 995324
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 419460 994974 419488 1002050
rect 419448 994968 419500 994974
rect 419448 994910 419500 994916
rect 397644 994764 397696 994770
rect 397644 994706 397696 994712
rect 420840 994702 420868 1004770
rect 422220 1002590 422248 1004906
rect 422666 1004864 422722 1004873
rect 422666 1004799 422668 1004808
rect 422720 1004799 422722 1004808
rect 422668 1004770 422720 1004776
rect 424324 1002856 424376 1002862
rect 424322 1002824 424324 1002833
rect 424376 1002824 424378 1002833
rect 424322 1002759 424378 1002768
rect 426544 1002726 426572 1006470
rect 431682 1006431 431684 1006440
rect 431736 1006431 431738 1006440
rect 431684 1006402 431736 1006408
rect 431684 1006256 431736 1006262
rect 429198 1006224 429254 1006233
rect 429198 1006159 429200 1006168
rect 429252 1006159 429254 1006168
rect 431682 1006224 431684 1006233
rect 431736 1006224 431738 1006233
rect 431682 1006159 431738 1006168
rect 429200 1006130 429252 1006136
rect 429200 1006052 429252 1006058
rect 429200 1005994 429252 1006000
rect 429212 1004086 429240 1005994
rect 430856 1005984 430908 1005990
rect 430854 1005952 430856 1005961
rect 430908 1005952 430910 1005961
rect 430854 1005887 430910 1005896
rect 434456 1005446 434484 1006674
rect 506202 1006496 506258 1006505
rect 506202 1006431 506204 1006440
rect 506256 1006431 506258 1006440
rect 506204 1006402 506256 1006408
rect 464988 1006324 465040 1006330
rect 464988 1006266 465040 1006272
rect 440884 1005780 440936 1005786
rect 440884 1005722 440936 1005728
rect 430028 1005440 430080 1005446
rect 430026 1005408 430028 1005417
rect 431960 1005440 432012 1005446
rect 430080 1005408 430082 1005417
rect 431960 1005382 432012 1005388
rect 434444 1005440 434496 1005446
rect 434444 1005382 434496 1005388
rect 430026 1005343 430082 1005352
rect 430026 1005136 430082 1005145
rect 430026 1005071 430028 1005080
rect 430080 1005071 430082 1005080
rect 430028 1005042 430080 1005048
rect 431222 1005000 431278 1005009
rect 431222 1004935 431224 1004944
rect 431276 1004935 431278 1004944
rect 431224 1004906 431276 1004912
rect 429200 1004080 429252 1004086
rect 429200 1004022 429252 1004028
rect 427176 1003944 427228 1003950
rect 427174 1003912 427176 1003921
rect 427228 1003912 427230 1003921
rect 427174 1003847 427230 1003856
rect 426532 1002720 426584 1002726
rect 426532 1002662 426584 1002668
rect 422208 1002584 422260 1002590
rect 422208 1002526 422260 1002532
rect 427728 1002584 427780 1002590
rect 427728 1002526 427780 1002532
rect 421470 1002144 421526 1002153
rect 421470 1002079 421472 1002088
rect 421524 1002079 421526 1002088
rect 427542 1002144 427598 1002153
rect 427542 1002079 427544 1002088
rect 421472 1002050 421524 1002056
rect 427596 1002079 427598 1002088
rect 427544 1002050 427596 1002056
rect 424322 1002008 424378 1002017
rect 422300 1001972 422352 1001978
rect 422300 1001914 422352 1001920
rect 423404 1001972 423456 1001978
rect 424322 1001943 424324 1001952
rect 423404 1001914 423456 1001920
rect 424376 1001943 424378 1001952
rect 425150 1002008 425206 1002017
rect 425150 1001943 425206 1001952
rect 425518 1002008 425574 1002017
rect 425518 1001943 425520 1001952
rect 424324 1001914 424376 1001920
rect 422312 997626 422340 1001914
rect 423416 1001230 423444 1001914
rect 423404 1001224 423456 1001230
rect 423404 1001166 423456 1001172
rect 422300 997620 422352 997626
rect 422300 997562 422352 997568
rect 425164 995110 425192 1001943
rect 425572 1001943 425574 1001952
rect 425520 1001914 425572 1001920
rect 427740 998578 427768 1002526
rect 431972 1002402 432000 1005382
rect 432604 1005100 432656 1005106
rect 432604 1005042 432656 1005048
rect 431926 1002374 432000 1002402
rect 428370 1002280 428426 1002289
rect 428370 1002215 428372 1002224
rect 428424 1002215 428426 1002224
rect 431408 1002244 431460 1002250
rect 428372 1002186 428424 1002192
rect 431408 1002186 431460 1002192
rect 429936 1002108 429988 1002114
rect 429936 1002050 429988 1002056
rect 429198 1002008 429254 1002017
rect 428464 1001972 428516 1001978
rect 429198 1001943 429200 1001952
rect 428464 1001914 428516 1001920
rect 429252 1001943 429254 1001952
rect 429200 1001914 429252 1001920
rect 428476 1001502 428504 1001914
rect 428464 1001496 428516 1001502
rect 428464 1001438 428516 1001444
rect 427728 998572 427780 998578
rect 427728 998514 427780 998520
rect 429948 998442 429976 1002050
rect 431224 1001972 431276 1001978
rect 431224 1001914 431276 1001920
rect 429936 998436 429988 998442
rect 429936 998378 429988 998384
rect 431236 997626 431264 1001914
rect 431420 1001366 431448 1002186
rect 431926 1002130 431954 1002374
rect 432050 1002280 432106 1002289
rect 432050 1002215 432052 1002224
rect 432104 1002215 432106 1002224
rect 432052 1002186 432104 1002192
rect 431926 1002102 432000 1002130
rect 431408 1001360 431460 1001366
rect 431408 1001302 431460 1001308
rect 431972 997762 432000 1002102
rect 432616 997762 432644 1005042
rect 433524 1004964 433576 1004970
rect 433524 1004906 433576 1004912
rect 433338 1002144 433394 1002153
rect 433338 1002079 433340 1002088
rect 433392 1002079 433394 1002088
rect 433340 1002050 433392 1002056
rect 432878 1002008 432934 1002017
rect 432878 1001943 432880 1001952
rect 432932 1001943 432934 1001952
rect 432880 1001914 432932 1001920
rect 431960 997756 432012 997762
rect 431960 997698 432012 997704
rect 432604 997756 432656 997762
rect 432604 997698 432656 997704
rect 426256 997620 426308 997626
rect 426256 997562 426308 997568
rect 431224 997620 431276 997626
rect 431224 997562 431276 997568
rect 425152 995104 425204 995110
rect 425152 995046 425204 995052
rect 420828 994696 420880 994702
rect 420828 994638 420880 994644
rect 392122 994463 392178 994472
rect 393964 994492 394016 994498
rect 393964 994434 394016 994440
rect 426268 994294 426296 997562
rect 433536 996130 433564 1004906
rect 435548 1002244 435600 1002250
rect 435548 1002186 435600 1002192
rect 435364 1002108 435416 1002114
rect 435364 1002050 435416 1002056
rect 433524 996124 433576 996130
rect 433524 996066 433576 996072
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 426256 994288 426308 994294
rect 426256 994230 426308 994236
rect 369124 990140 369176 990146
rect 369124 990082 369176 990088
rect 381188 983634 381216 994230
rect 429936 992928 429988 992934
rect 429936 992870 429988 992876
rect 397828 991500 397880 991506
rect 397828 991442 397880 991448
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 991442
rect 414112 990140 414164 990146
rect 414112 990082 414164 990088
rect 414124 983620 414152 990082
rect 429948 983634 429976 992870
rect 435376 991506 435404 1002050
rect 435560 992934 435588 1002186
rect 436744 1001972 436796 1001978
rect 436744 1001914 436796 1001920
rect 435548 992928 435600 992934
rect 435548 992870 435600 992876
rect 435364 991500 435416 991506
rect 435364 991442 435416 991448
rect 436756 985998 436784 1001914
rect 440896 999122 440924 1005722
rect 443644 1005576 443696 1005582
rect 443644 1005518 443696 1005524
rect 440884 999116 440936 999122
rect 440884 999058 440936 999064
rect 443656 998714 443684 1005518
rect 458824 1005440 458876 1005446
rect 458824 1005382 458876 1005388
rect 456064 1005304 456116 1005310
rect 456064 1005246 456116 1005252
rect 446404 1004080 446456 1004086
rect 446404 1004022 446456 1004028
rect 446416 1001638 446444 1004022
rect 449164 1002720 449216 1002726
rect 449164 1002662 449216 1002668
rect 446404 1001632 446456 1001638
rect 446404 1001574 446456 1001580
rect 446404 1001496 446456 1001502
rect 446404 1001438 446456 1001444
rect 444288 999116 444340 999122
rect 444288 999058 444340 999064
rect 443644 998708 443696 998714
rect 443644 998650 443696 998656
rect 439872 997756 439924 997762
rect 439872 997698 439924 997704
rect 439688 997620 439740 997626
rect 439688 997562 439740 997568
rect 439700 996985 439728 997562
rect 439884 997257 439912 997698
rect 439870 997248 439926 997257
rect 439870 997183 439926 997192
rect 444300 997082 444328 999058
rect 444288 997076 444340 997082
rect 444288 997018 444340 997024
rect 439686 996976 439742 996985
rect 439686 996911 439742 996920
rect 446416 994809 446444 1001438
rect 449176 995625 449204 1002662
rect 456076 1001894 456104 1005246
rect 456076 1001866 456288 1001894
rect 453212 1001632 453264 1001638
rect 453212 1001574 453264 1001580
rect 453224 996305 453252 1001574
rect 456064 998572 456116 998578
rect 456064 998514 456116 998520
rect 456076 998306 456104 998514
rect 456064 998300 456116 998306
rect 456064 998242 456116 998248
rect 453210 996296 453266 996305
rect 453210 996231 453266 996240
rect 449162 995616 449218 995625
rect 449162 995551 449218 995560
rect 456260 994838 456288 1001866
rect 458836 998209 458864 1005382
rect 464804 1003944 464856 1003950
rect 464804 1003886 464856 1003892
rect 461860 1001360 461912 1001366
rect 461860 1001302 461912 1001308
rect 461124 998300 461176 998306
rect 461124 998242 461176 998248
rect 458822 998200 458878 998209
rect 458822 998135 458878 998144
rect 456248 994832 456300 994838
rect 446402 994800 446458 994809
rect 456248 994774 456300 994780
rect 446402 994735 446458 994744
rect 461136 994537 461164 998242
rect 461872 997898 461900 1001302
rect 464816 998578 464844 1003886
rect 465000 1003338 465028 1006266
rect 508226 1006224 508282 1006233
rect 471244 1006188 471296 1006194
rect 508226 1006159 508228 1006168
rect 471244 1006130 471296 1006136
rect 508280 1006159 508282 1006168
rect 508228 1006130 508280 1006136
rect 469864 1006052 469916 1006058
rect 469864 1005994 469916 1006000
rect 464988 1003332 465040 1003338
rect 464988 1003274 465040 1003280
rect 464988 1002584 465040 1002590
rect 464988 1002526 465040 1002532
rect 464804 998572 464856 998578
rect 464804 998514 464856 998520
rect 461860 997892 461912 997898
rect 461860 997834 461912 997840
rect 463884 997892 463936 997898
rect 463884 997834 463936 997840
rect 461122 994528 461178 994537
rect 461122 994463 461178 994472
rect 463896 994430 463924 997834
rect 465000 997762 465028 1002526
rect 466460 1001224 466512 1001230
rect 466460 1001166 466512 1001172
rect 464988 997756 465040 997762
rect 466472 997754 466500 1001166
rect 466472 997726 466592 997754
rect 464988 997698 465040 997704
rect 466564 994430 466592 997726
rect 469876 995625 469904 1005994
rect 471060 997756 471112 997762
rect 471060 997698 471112 997704
rect 470508 997076 470560 997082
rect 470508 997018 470560 997024
rect 469862 995616 469918 995625
rect 469862 995551 469918 995560
rect 470520 994566 470548 997018
rect 470508 994560 470560 994566
rect 470508 994502 470560 994508
rect 463884 994424 463936 994430
rect 463884 994366 463936 994372
rect 466552 994424 466604 994430
rect 466552 994366 466604 994372
rect 446128 994288 446180 994294
rect 446128 994230 446180 994236
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 994230
rect 471072 994158 471100 997698
rect 471256 995081 471284 1006130
rect 498842 1006088 498898 1006097
rect 498108 1006052 498160 1006058
rect 498842 1006023 498844 1006032
rect 498108 1005994 498160 1006000
rect 498896 1006023 498898 1006032
rect 509054 1006088 509110 1006097
rect 509054 1006023 509056 1006032
rect 498844 1005994 498896 1006000
rect 509108 1006023 509110 1006032
rect 509056 1005994 509108 1006000
rect 472440 1003332 472492 1003338
rect 472440 1003274 472492 1003280
rect 472256 998572 472308 998578
rect 472256 998514 472308 998520
rect 472072 998436 472124 998442
rect 472072 998378 472124 998384
rect 471242 995072 471298 995081
rect 471242 995007 471298 995016
rect 471244 994832 471296 994838
rect 471244 994774 471296 994780
rect 471060 994152 471112 994158
rect 471060 994094 471112 994100
rect 471256 994022 471284 994774
rect 472084 994265 472112 998378
rect 472268 996033 472296 998514
rect 472452 998458 472480 1003274
rect 496728 1001972 496780 1001978
rect 496728 1001914 496780 1001920
rect 496740 1001230 496768 1001914
rect 496728 1001224 496780 1001230
rect 496728 1001166 496780 1001172
rect 472624 998708 472676 998714
rect 472624 998650 472676 998656
rect 472636 998594 472664 998650
rect 472636 998566 472756 998594
rect 472452 998430 472664 998458
rect 472438 998200 472494 998209
rect 472438 998135 472494 998144
rect 472452 996577 472480 998135
rect 472438 996568 472494 996577
rect 472438 996503 472494 996512
rect 472254 996024 472310 996033
rect 472254 995959 472310 995968
rect 472438 995616 472494 995625
rect 472636 995586 472664 998430
rect 472728 995738 472756 998566
rect 488908 997756 488960 997762
rect 488908 997698 488960 997704
rect 488920 997257 488948 997698
rect 489092 997620 489144 997626
rect 489092 997562 489144 997568
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 489104 996985 489132 997562
rect 489090 996976 489146 996985
rect 489090 996911 489146 996920
rect 489550 996704 489606 996713
rect 489550 996639 489606 996648
rect 490102 996704 490158 996713
rect 490102 996639 490158 996648
rect 472898 995752 472954 995761
rect 472728 995710 472898 995738
rect 472898 995687 472954 995696
rect 474002 995752 474058 995761
rect 476946 995752 477002 995761
rect 474058 995710 474306 995738
rect 474002 995687 474058 995696
rect 480810 995752 480866 995761
rect 477002 995710 477342 995738
rect 476946 995687 477002 995696
rect 485594 995752 485650 995761
rect 480866 995710 481114 995738
rect 485346 995710 485594 995738
rect 480810 995687 480866 995696
rect 485594 995687 485650 995696
rect 474738 995616 474794 995625
rect 473372 995586 473662 995602
rect 472438 995551 472494 995560
rect 472624 995580 472676 995586
rect 472452 994838 472480 995551
rect 472624 995522 472676 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 478326 995616 478382 995625
rect 474794 995574 474950 995602
rect 477986 995574 478326 995602
rect 474738 995551 474794 995560
rect 478326 995551 478382 995560
rect 480258 995616 480314 995625
rect 480258 995551 480314 995560
rect 473360 995522 473412 995528
rect 476072 995072 476128 995081
rect 475948 995030 476072 995058
rect 475948 994838 475976 995030
rect 476072 995007 476128 995016
rect 472440 994832 472492 994838
rect 472440 994774 472492 994780
rect 475936 994832 475988 994838
rect 475936 994774 475988 994780
rect 476120 994832 476172 994838
rect 476120 994774 476172 994780
rect 476132 994650 476160 994774
rect 475672 994622 476160 994650
rect 475672 994566 475700 994622
rect 475660 994560 475712 994566
rect 475660 994502 475712 994508
rect 475936 994560 475988 994566
rect 475936 994502 475988 994508
rect 475752 994424 475804 994430
rect 475948 994412 475976 994502
rect 475804 994384 475976 994412
rect 476074 994424 476126 994430
rect 475752 994366 475804 994372
rect 476040 994372 476074 994378
rect 476040 994366 476126 994372
rect 476040 994350 476114 994366
rect 472070 994256 472126 994265
rect 472070 994191 472126 994200
rect 476040 994158 476068 994350
rect 476776 994265 476804 995452
rect 478248 995438 478630 995466
rect 478248 995353 478276 995438
rect 478234 995344 478290 995353
rect 478234 995279 478290 995288
rect 480272 994809 480300 995551
rect 480258 994800 480314 994809
rect 480258 994735 480314 994744
rect 476762 994256 476818 994265
rect 476762 994191 476818 994200
rect 481652 994158 481680 995452
rect 482296 994158 482324 995452
rect 482664 995438 482954 995466
rect 482664 994537 482692 995438
rect 484136 995110 484164 995452
rect 484124 995104 484176 995110
rect 484124 995046 484176 995052
rect 485228 994832 485280 994838
rect 485228 994774 485280 994780
rect 482650 994528 482706 994537
rect 482650 994463 482706 994472
rect 485240 994430 485268 994774
rect 485228 994424 485280 994430
rect 485228 994366 485280 994372
rect 476028 994152 476080 994158
rect 476028 994094 476080 994100
rect 481640 994152 481692 994158
rect 481640 994094 481692 994100
rect 482284 994152 482336 994158
rect 482284 994094 482336 994100
rect 485976 994022 486004 995452
rect 486620 994838 486648 995452
rect 486608 994832 486660 994838
rect 486608 994774 486660 994780
rect 487816 994430 487844 995452
rect 487804 994424 487856 994430
rect 487804 994366 487856 994372
rect 489564 994158 489592 996639
rect 489736 995172 489788 995178
rect 489736 995114 489788 995120
rect 489920 995172 489972 995178
rect 489920 995114 489972 995120
rect 489748 994838 489776 995114
rect 489736 994832 489788 994838
rect 489736 994774 489788 994780
rect 489932 994294 489960 995114
rect 490116 994566 490144 996639
rect 494702 996432 494758 996441
rect 494702 996367 494758 996376
rect 494716 995586 494744 996367
rect 494704 995580 494756 995586
rect 494704 995522 494756 995528
rect 490104 994560 490156 994566
rect 490104 994502 490156 994508
rect 498120 994430 498148 1005994
rect 514024 1005984 514076 1005990
rect 514024 1005926 514076 1005932
rect 502156 1005440 502208 1005446
rect 502154 1005408 502156 1005417
rect 502208 1005408 502210 1005417
rect 502154 1005343 502210 1005352
rect 499672 1005304 499724 1005310
rect 499670 1005272 499672 1005281
rect 499724 1005272 499726 1005281
rect 499670 1005207 499726 1005216
rect 507030 1005000 507086 1005009
rect 507030 1004935 507032 1004944
rect 507084 1004935 507086 1004944
rect 509700 1004964 509752 1004970
rect 507032 1004906 507084 1004912
rect 509700 1004906 509752 1004912
rect 507858 1004864 507914 1004873
rect 507858 1004799 507860 1004808
rect 507912 1004799 507914 1004808
rect 507860 1004770 507912 1004776
rect 501326 1004728 501382 1004737
rect 499304 1004692 499356 1004698
rect 501326 1004663 501328 1004672
rect 499304 1004634 499356 1004640
rect 501380 1004663 501382 1004672
rect 501328 1004634 501380 1004640
rect 498474 1002008 498530 1002017
rect 498474 1001943 498476 1001952
rect 498528 1001943 498530 1001952
rect 498476 1001914 498528 1001920
rect 499316 998850 499344 1004634
rect 505376 1004624 505428 1004630
rect 505374 1004592 505376 1004601
rect 505428 1004592 505430 1004601
rect 505374 1004527 505430 1004536
rect 505008 1003944 505060 1003950
rect 505006 1003912 505008 1003921
rect 505060 1003912 505062 1003921
rect 505006 1003847 505062 1003856
rect 504180 1002720 504232 1002726
rect 504178 1002688 504180 1002697
rect 504232 1002688 504234 1002697
rect 504178 1002623 504234 1002632
rect 501696 1002584 501748 1002590
rect 501694 1002552 501696 1002561
rect 501748 1002552 501750 1002561
rect 501694 1002487 501750 1002496
rect 503350 1002416 503406 1002425
rect 500316 1002380 500368 1002386
rect 503350 1002351 503352 1002360
rect 500316 1002322 500368 1002328
rect 503404 1002351 503406 1002360
rect 503352 1002322 503404 1002328
rect 499580 1001972 499632 1001978
rect 499580 1001914 499632 1001920
rect 499304 998844 499356 998850
rect 499304 998786 499356 998792
rect 499592 998714 499620 1001914
rect 499580 998708 499632 998714
rect 499580 998650 499632 998656
rect 500328 998578 500356 1002322
rect 500498 1002280 500554 1002289
rect 500498 1002215 500500 1002224
rect 500552 1002215 500554 1002224
rect 502984 1002244 503036 1002250
rect 500500 1002186 500552 1002192
rect 502984 1002186 503036 1002192
rect 500498 1002008 500554 1002017
rect 502154 1002008 502210 1002017
rect 500498 1001943 500500 1001952
rect 500552 1001943 500554 1001952
rect 500960 1001972 501012 1001978
rect 500500 1001914 500552 1001920
rect 502154 1001943 502156 1001952
rect 500960 1001914 501012 1001920
rect 502208 1001943 502210 1001952
rect 502522 1002008 502578 1002017
rect 502522 1001943 502524 1001952
rect 502156 1001914 502208 1001920
rect 502576 1001943 502578 1001952
rect 502524 1001914 502576 1001920
rect 500316 998572 500368 998578
rect 500316 998514 500368 998520
rect 500972 998442 501000 1001914
rect 500960 998436 501012 998442
rect 500960 998378 501012 998384
rect 502996 994838 503024 1002186
rect 503350 1002144 503406 1002153
rect 503350 1002079 503352 1002088
rect 503404 1002079 503406 1002088
rect 505744 1002108 505796 1002114
rect 503352 1002050 503404 1002056
rect 505744 1002050 505796 1002056
rect 504364 1001972 504416 1001978
rect 504364 1001914 504416 1001920
rect 504376 999802 504404 1001914
rect 504364 999796 504416 999802
rect 504364 999738 504416 999744
rect 505756 997082 505784 1002050
rect 506202 1002008 506258 1002017
rect 507398 1002008 507454 1002017
rect 506258 1001966 506520 1001994
rect 506202 1001943 506258 1001952
rect 506492 997626 506520 1001966
rect 507454 1001966 507900 1001994
rect 507398 1001943 507454 1001952
rect 507872 997762 507900 1001966
rect 509712 997762 509740 1004906
rect 510068 1004828 510120 1004834
rect 510068 1004770 510120 1004776
rect 509882 1002280 509938 1002289
rect 509882 1002215 509884 1002224
rect 509936 1002215 509938 1002224
rect 509884 1002186 509936 1002192
rect 510080 1001894 510108 1004770
rect 510252 1004624 510304 1004630
rect 509988 1001866 510108 1001894
rect 510172 1004572 510252 1004578
rect 510172 1004566 510304 1004572
rect 510172 1004550 510292 1004566
rect 507860 997756 507912 997762
rect 507860 997698 507912 997704
rect 509700 997756 509752 997762
rect 509700 997698 509752 997704
rect 509988 997626 510016 1001866
rect 510172 1001774 510200 1004550
rect 512828 1002244 512880 1002250
rect 512828 1002186 512880 1002192
rect 510342 1002144 510398 1002153
rect 510342 1002079 510344 1002088
rect 510396 1002079 510398 1002088
rect 512644 1002108 512696 1002114
rect 510344 1002050 510396 1002056
rect 512644 1002050 512696 1002056
rect 510160 1001768 510212 1001774
rect 510160 1001710 510212 1001716
rect 506480 997620 506532 997626
rect 506480 997562 506532 997568
rect 509976 997620 510028 997626
rect 509976 997562 510028 997568
rect 505744 997076 505796 997082
rect 505744 997018 505796 997024
rect 503810 995616 503866 995625
rect 503810 995551 503866 995560
rect 511080 995580 511132 995586
rect 503824 995081 503852 995551
rect 511080 995522 511132 995528
rect 503810 995072 503866 995081
rect 503810 995007 503866 995016
rect 502984 994832 503036 994838
rect 502984 994774 503036 994780
rect 498108 994424 498160 994430
rect 498108 994366 498160 994372
rect 489920 994288 489972 994294
rect 489920 994230 489972 994236
rect 489552 994152 489604 994158
rect 489552 994094 489604 994100
rect 471244 994016 471296 994022
rect 471244 993958 471296 993964
rect 485964 994016 486016 994022
rect 485964 993958 486016 993964
rect 494704 992928 494756 992934
rect 494704 992870 494756 992876
rect 478972 991500 479024 991506
rect 478972 991442 479024 991448
rect 462780 985992 462832 985998
rect 462780 985934 462832 985940
rect 429948 983606 430330 983634
rect 446140 983606 446522 983634
rect 462792 983620 462820 985934
rect 478984 983620 479012 991442
rect 494716 983634 494744 992870
rect 511092 983634 511120 995522
rect 512656 991506 512684 1002050
rect 512840 992934 512868 1002186
rect 512828 992928 512880 992934
rect 512828 992870 512880 992876
rect 512644 991500 512696 991506
rect 512644 991442 512696 991448
rect 514036 985998 514064 1005926
rect 515416 995110 515444 1006674
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 516796 1001894 516824 1005246
rect 516520 1001866 516824 1001894
rect 515404 995104 515456 995110
rect 515404 995046 515456 995052
rect 516520 993682 516548 1001866
rect 516692 1001768 516744 1001774
rect 516692 1001710 516744 1001716
rect 516704 998617 516732 1001710
rect 516980 999122 517008 1006810
rect 554318 1006768 554374 1006777
rect 554318 1006703 554320 1006712
rect 554372 1006703 554374 1006712
rect 554320 1006674 554372 1006680
rect 555974 1006496 556030 1006505
rect 555974 1006431 555976 1006440
rect 556028 1006431 556030 1006440
rect 555976 1006402 556028 1006408
rect 520924 1006324 520976 1006330
rect 520924 1006266 520976 1006272
rect 518164 1005440 518216 1005446
rect 518164 1005382 518216 1005388
rect 517520 1003944 517572 1003950
rect 517520 1003886 517572 1003892
rect 516968 999116 517020 999122
rect 516968 999058 517020 999064
rect 517532 998850 517560 1003886
rect 516876 998844 516928 998850
rect 516876 998786 516928 998792
rect 517520 998844 517572 998850
rect 517520 998786 517572 998792
rect 516690 998608 516746 998617
rect 516690 998543 516746 998552
rect 516692 997756 516744 997762
rect 516692 997698 516744 997704
rect 516704 997257 516732 997698
rect 516690 997248 516746 997257
rect 516690 997183 516746 997192
rect 516888 995625 516916 998786
rect 517520 998708 517572 998714
rect 517520 998650 517572 998656
rect 517060 997620 517112 997626
rect 517060 997562 517112 997568
rect 517072 996985 517100 997562
rect 517058 996976 517114 996985
rect 517058 996911 517114 996920
rect 516874 995616 516930 995625
rect 516874 995551 516930 995560
rect 517532 994537 517560 998650
rect 518176 995858 518204 1005382
rect 518900 1002720 518952 1002726
rect 518900 1002662 518952 1002668
rect 518912 999258 518940 1002662
rect 519820 999796 519872 999802
rect 519820 999738 519872 999744
rect 518900 999252 518952 999258
rect 518900 999194 518952 999200
rect 519832 996305 519860 999738
rect 520188 999116 520240 999122
rect 520188 999058 520240 999064
rect 520004 997076 520056 997082
rect 520004 997018 520056 997024
rect 519818 996296 519874 996305
rect 519818 996231 519874 996240
rect 518164 995852 518216 995858
rect 518164 995794 518216 995800
rect 520016 994566 520044 997018
rect 520200 995081 520228 999058
rect 520936 995897 520964 1006266
rect 550270 1006088 550326 1006097
rect 522304 1006052 522356 1006058
rect 522304 1005994 522356 1006000
rect 549168 1006052 549220 1006058
rect 550270 1006023 550272 1006032
rect 549168 1005994 549220 1006000
rect 550324 1006023 550326 1006032
rect 553950 1006088 554006 1006097
rect 553950 1006023 553952 1006032
rect 550272 1005994 550324 1006000
rect 554004 1006023 554006 1006032
rect 556160 1006052 556212 1006058
rect 553952 1005994 554004 1006000
rect 556160 1005994 556212 1006000
rect 522316 996305 522344 1005994
rect 523316 1002584 523368 1002590
rect 523316 1002526 523368 1002532
rect 523328 1001894 523356 1002526
rect 523236 1001866 523356 1001894
rect 522764 1001224 522816 1001230
rect 522764 1001166 522816 1001172
rect 522302 996296 522358 996305
rect 522302 996231 522358 996240
rect 520922 995888 520978 995897
rect 520922 995823 520978 995832
rect 520186 995072 520242 995081
rect 520186 995007 520242 995016
rect 520004 994560 520056 994566
rect 517518 994528 517574 994537
rect 520004 994502 520056 994508
rect 517518 994463 517574 994472
rect 522776 993818 522804 1001166
rect 522948 998572 523000 998578
rect 522948 998514 523000 998520
rect 522960 995353 522988 998514
rect 522946 995344 523002 995353
rect 522946 995279 523002 995288
rect 523236 994265 523264 1001866
rect 524052 999252 524104 999258
rect 524052 999194 524104 999200
rect 523684 998844 523736 998850
rect 523684 998786 523736 998792
rect 523406 998608 523462 998617
rect 523406 998543 523462 998552
rect 523420 995081 523448 998543
rect 523696 995586 523724 998786
rect 523868 998436 523920 998442
rect 523868 998378 523920 998384
rect 523880 996033 523908 998378
rect 524064 997801 524092 999194
rect 524050 997792 524106 997801
rect 524050 997727 524106 997736
rect 540520 997688 540572 997694
rect 540520 997630 540572 997636
rect 540336 997416 540388 997422
rect 540336 997358 540388 997364
rect 540348 997257 540376 997358
rect 540334 997248 540390 997257
rect 540334 997183 540390 997192
rect 540532 996985 540560 997630
rect 540518 996976 540574 996985
rect 540518 996911 540574 996920
rect 523866 996024 523922 996033
rect 523866 995959 523922 995968
rect 524052 995852 524104 995858
rect 524052 995794 524104 995800
rect 523684 995580 523736 995586
rect 523684 995522 523736 995528
rect 523406 995072 523462 995081
rect 523406 995007 523462 995016
rect 524064 994294 524092 995794
rect 532238 995752 532294 995761
rect 532294 995710 532542 995738
rect 532238 995687 532294 995696
rect 529846 995616 529902 995625
rect 524800 995586 525090 995602
rect 524788 995580 525090 995586
rect 524840 995574 525090 995580
rect 528572 995574 528770 995602
rect 524788 995522 524840 995528
rect 525352 995438 525734 995466
rect 526088 995438 526378 995466
rect 527928 995438 528218 995466
rect 525352 995353 525380 995438
rect 525338 995344 525394 995353
rect 525338 995279 525394 995288
rect 526088 995081 526116 995438
rect 527928 995081 527956 995438
rect 528572 995353 528600 995574
rect 536930 995616 536986 995625
rect 529902 995574 530058 995602
rect 536774 995574 536930 995602
rect 529846 995551 529902 995560
rect 536930 995551 536986 995560
rect 528940 995438 529414 995466
rect 528940 995353 528968 995438
rect 528558 995344 528614 995353
rect 528558 995279 528614 995288
rect 528926 995344 528982 995353
rect 528926 995279 528982 995288
rect 526074 995072 526130 995081
rect 526074 995007 526130 995016
rect 527914 995072 527970 995081
rect 527914 995007 527970 995016
rect 526534 994800 526590 994809
rect 526534 994735 526590 994744
rect 524052 994288 524104 994294
rect 523222 994256 523278 994265
rect 526548 994265 526576 994735
rect 533080 994537 533108 995452
rect 533724 994809 533752 995452
rect 534368 994838 534396 995452
rect 534356 994832 534408 994838
rect 533710 994800 533766 994809
rect 534356 994774 534408 994780
rect 533710 994735 533766 994744
rect 533066 994528 533122 994537
rect 533066 994463 533122 994472
rect 535564 994294 535592 995452
rect 537404 995110 537432 995452
rect 537392 995104 537444 995110
rect 537392 995046 537444 995052
rect 538048 994430 538076 995452
rect 539244 994566 539272 995452
rect 539232 994560 539284 994566
rect 539232 994502 539284 994508
rect 538036 994424 538088 994430
rect 538036 994366 538088 994372
rect 535552 994288 535604 994294
rect 524052 994230 524104 994236
rect 526534 994256 526590 994265
rect 523222 994191 523278 994200
rect 535552 994230 535604 994236
rect 526534 994191 526590 994200
rect 522764 993812 522816 993818
rect 522764 993754 522816 993760
rect 516508 993676 516560 993682
rect 516508 993618 516560 993624
rect 549180 993546 549208 1005994
rect 556172 1005582 556200 1005994
rect 556160 1005576 556212 1005582
rect 556160 1005518 556212 1005524
rect 551468 1005440 551520 1005446
rect 551466 1005408 551468 1005417
rect 551520 1005408 551522 1005417
rect 551466 1005343 551522 1005352
rect 551468 1005168 551520 1005174
rect 551466 1005136 551468 1005145
rect 551520 1005136 551522 1005145
rect 551466 1005071 551522 1005080
rect 556802 1005000 556858 1005009
rect 556802 1004935 556804 1004944
rect 556856 1004935 556858 1004944
rect 556804 1004906 556856 1004912
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 552296 1003944 552348 1003950
rect 552294 1003912 552296 1003921
rect 552348 1003912 552350 1003921
rect 552294 1003847 552350 1003856
rect 554778 1002280 554834 1002289
rect 554608 1002238 554778 1002266
rect 552294 1002144 552350 1002153
rect 552294 1002079 552296 1002088
rect 552348 1002079 552350 1002088
rect 552296 1002050 552348 1002056
rect 554318 1002008 554374 1002017
rect 553308 1001972 553360 1001978
rect 554374 1001966 554544 1001994
rect 554318 1001943 554374 1001952
rect 553308 1001914 553360 1001920
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 553122 998064 553178 998073
rect 550548 998028 550600 998034
rect 553122 997999 553124 998008
rect 550548 997970 550600 997976
rect 553176 997999 553178 998008
rect 553124 997970 553176 997976
rect 550560 997082 550588 997970
rect 551744 997824 551796 997830
rect 553124 997824 553176 997830
rect 551744 997766 551796 997772
rect 553122 997792 553124 997801
rect 553176 997792 553178 997801
rect 550548 997076 550600 997082
rect 550548 997018 550600 997024
rect 549168 993540 549220 993546
rect 549168 993482 549220 993488
rect 551756 993410 551784 997766
rect 553122 997727 553178 997736
rect 553320 996334 553348 1001914
rect 554516 997558 554544 1001966
rect 554608 1001894 554636 1002238
rect 554778 1002215 554834 1002224
rect 555424 1002108 555476 1002114
rect 555424 1002050 555476 1002056
rect 555146 1002008 555202 1002017
rect 555146 1001943 555148 1001952
rect 555200 1001943 555202 1001952
rect 555148 1001914 555200 1001920
rect 554608 1001866 554728 1001894
rect 554504 997552 554556 997558
rect 554504 997494 554556 997500
rect 554700 997218 554728 1001866
rect 555436 998102 555464 1002050
rect 555424 998096 555476 998102
rect 555424 998038 555476 998044
rect 557000 997694 557028 1006810
rect 562324 1006732 562376 1006738
rect 562324 1006674 562376 1006680
rect 557170 1006224 557226 1006233
rect 557170 1006159 557172 1006168
rect 557224 1006159 557226 1006168
rect 557172 1006130 557224 1006136
rect 562336 1006058 562364 1006674
rect 566464 1006460 566516 1006466
rect 566464 1006402 566516 1006408
rect 562324 1006052 562376 1006058
rect 562324 1005994 562376 1006000
rect 558920 1004964 558972 1004970
rect 558920 1004906 558972 1004912
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002144 558054 1002153
rect 557998 1002079 558000 1002088
rect 558052 1002079 558054 1002088
rect 558000 1002050 558052 1002056
rect 558196 999802 558224 1004770
rect 558932 1004086 558960 1004906
rect 559564 1004692 559616 1004698
rect 559564 1004634 559616 1004640
rect 558920 1004080 558972 1004086
rect 558920 1004022 558972 1004028
rect 558826 1002552 558882 1002561
rect 558826 1002487 558828 1002496
rect 558880 1002487 558882 1002496
rect 558828 1002458 558880 1002464
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 558184 999796 558236 999802
rect 558184 999738 558236 999744
rect 557172 998096 557224 998102
rect 557170 998064 557172 998073
rect 557224 998064 557226 998073
rect 557170 997999 557226 998008
rect 556988 997688 557040 997694
rect 556988 997630 557040 997636
rect 554688 997212 554740 997218
rect 554688 997154 554740 997160
rect 553308 996328 553360 996334
rect 553308 996270 553360 996276
rect 552662 995616 552718 995625
rect 552662 995551 552718 995560
rect 552676 995081 552704 995551
rect 552662 995072 552718 995081
rect 552662 995007 552718 995016
rect 551744 993404 551796 993410
rect 551744 993346 551796 993352
rect 527272 992928 527324 992934
rect 527272 992870 527324 992876
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 527284 983634 527312 992870
rect 559576 991506 559604 1004634
rect 562508 1002516 562560 1002522
rect 562508 1002458 562560 1002464
rect 560850 1002416 560906 1002425
rect 560850 1002351 560852 1002360
rect 560904 1002351 560906 1002360
rect 560852 1002322 560904 1002328
rect 560022 1002280 560078 1002289
rect 560022 1002215 560024 1002224
rect 560076 1002215 560078 1002224
rect 562324 1002244 562376 1002250
rect 560024 1002186 560076 1002192
rect 562324 1002186 562376 1002192
rect 560850 1002144 560906 1002153
rect 560668 1002108 560720 1002114
rect 560850 1002079 560852 1002088
rect 560668 1002050 560720 1002056
rect 560904 1002079 560906 1002088
rect 560852 1002050 560904 1002056
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 560312 997422 560340 1001914
rect 560680 1001894 560708 1002050
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 560680 1001866 560984 1001894
rect 560300 997416 560352 997422
rect 560300 997358 560352 997364
rect 543832 991500 543884 991506
rect 543832 991442 543884 991448
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 494716 983606 495190 983634
rect 511092 983606 511474 983634
rect 527284 983606 527666 983634
rect 543844 983620 543872 991442
rect 560956 990282 560984 1001866
rect 560944 990276 560996 990282
rect 560944 990218 560996 990224
rect 562336 990146 562364 1002186
rect 562520 992934 562548 1002458
rect 565268 1002380 565320 1002386
rect 565268 1002322 565320 1002328
rect 565084 1002108 565136 1002114
rect 565084 1002050 565136 1002056
rect 563704 1001972 563756 1001978
rect 563704 1001914 563756 1001920
rect 563716 993070 563744 1001914
rect 563704 993064 563756 993070
rect 563704 993006 563756 993012
rect 562508 992928 562560 992934
rect 562508 992870 562560 992876
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 565096 986134 565124 1002050
rect 565084 986128 565136 986134
rect 565084 986070 565136 986076
rect 565280 985998 565308 1002322
rect 566476 997694 566504 1006402
rect 567844 1006188 567896 1006194
rect 567844 1006130 567896 1006136
rect 566464 997688 566516 997694
rect 566464 997630 566516 997636
rect 567856 994566 567884 1006130
rect 573364 1006052 573416 1006058
rect 573364 1005994 573416 1006000
rect 570604 1005576 570656 1005582
rect 570604 1005518 570656 1005524
rect 569224 1005440 569276 1005446
rect 569224 1005382 569276 1005388
rect 568120 999796 568172 999802
rect 568120 999738 568172 999744
rect 568132 995110 568160 999738
rect 568948 997212 569000 997218
rect 568948 997154 569000 997160
rect 568120 995104 568172 995110
rect 568120 995046 568172 995052
rect 568960 994974 568988 997154
rect 568212 994968 568264 994974
rect 568212 994910 568264 994916
rect 568948 994968 569000 994974
rect 568948 994910 569000 994916
rect 567844 994560 567896 994566
rect 567844 994502 567896 994508
rect 568224 993721 568252 994910
rect 569236 994838 569264 1005382
rect 570616 996946 570644 1005518
rect 571984 1004080 572036 1004086
rect 571984 1004022 572036 1004028
rect 570604 996940 570656 996946
rect 570604 996882 570656 996888
rect 569224 994832 569276 994838
rect 569224 994774 569276 994780
rect 571996 994430 572024 1004022
rect 572628 1003944 572680 1003950
rect 572628 1003886 572680 1003892
rect 572640 997218 572668 1003886
rect 573376 997422 573404 1005994
rect 574744 1005304 574796 1005310
rect 574744 1005246 574796 1005252
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 573364 997416 573416 997422
rect 573364 997358 573416 997364
rect 572628 997212 572680 997218
rect 572628 997154 572680 997160
rect 571984 994424 572036 994430
rect 571984 994366 572036 994372
rect 574112 994090 574140 1001166
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 574756 993954 574784 1005246
rect 591488 998096 591540 998102
rect 591488 998038 591540 998044
rect 625712 998096 625764 998102
rect 625712 998038 625764 998044
rect 591120 997960 591172 997966
rect 591120 997902 591172 997908
rect 591132 997558 591160 997902
rect 591304 997824 591356 997830
rect 591304 997766 591356 997772
rect 591120 997552 591172 997558
rect 591120 997494 591172 997500
rect 591316 997422 591344 997766
rect 591500 997694 591528 998038
rect 625528 997960 625580 997966
rect 625528 997902 625580 997908
rect 625344 997824 625396 997830
rect 625344 997766 625396 997772
rect 591488 997688 591540 997694
rect 591488 997630 591540 997636
rect 591304 997416 591356 997422
rect 591304 997358 591356 997364
rect 623688 997212 623740 997218
rect 623688 997154 623740 997160
rect 620100 997076 620152 997082
rect 620100 997018 620152 997024
rect 599950 996976 600006 996985
rect 590568 996940 590620 996946
rect 599950 996911 600006 996920
rect 590568 996882 590620 996888
rect 590580 996713 590608 996882
rect 590566 996704 590622 996713
rect 590566 996639 590622 996648
rect 599964 996441 599992 996911
rect 591302 996432 591358 996441
rect 591302 996367 591358 996376
rect 599950 996432 600006 996441
rect 599950 996367 600006 996376
rect 618166 996432 618222 996441
rect 618166 996367 618222 996376
rect 590566 995072 590622 995081
rect 590566 995007 590622 995016
rect 590580 994702 590608 995007
rect 590568 994696 590620 994702
rect 590568 994638 590620 994644
rect 591316 994566 591344 996367
rect 618180 996266 618208 996367
rect 618168 996260 618220 996266
rect 618168 996202 618220 996208
rect 620112 996033 620140 997018
rect 623700 996033 623728 997154
rect 620098 996024 620154 996033
rect 620098 995959 620154 995968
rect 623686 996024 623742 996033
rect 623686 995959 623742 995968
rect 625356 994702 625384 997766
rect 625540 995489 625568 997902
rect 625724 995586 625752 998038
rect 635186 995752 635242 995761
rect 635242 995710 635536 995738
rect 635186 995687 635242 995696
rect 626552 995586 626888 995602
rect 625712 995580 625764 995586
rect 625712 995522 625764 995528
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 626540 995522 626592 995528
rect 625526 995480 625582 995489
rect 625526 995415 625582 995424
rect 627182 995480 627238 995489
rect 627918 995480 627974 995489
rect 627238 995438 627532 995466
rect 627182 995415 627238 995424
rect 631506 995480 631562 995489
rect 627974 995438 628176 995466
rect 629680 995438 630016 995466
rect 630232 995438 630568 995466
rect 631212 995438 631364 995466
rect 627918 995415 627974 995424
rect 629680 995110 629708 995438
rect 629668 995104 629720 995110
rect 629668 995046 629720 995052
rect 630232 994702 630260 995438
rect 631336 995330 631364 995438
rect 633990 995480 634046 995489
rect 631562 995438 631856 995466
rect 631506 995415 631562 995424
rect 634726 995480 634782 995489
rect 634046 995438 634340 995466
rect 633990 995415 634046 995424
rect 634782 995438 634892 995466
rect 635844 995438 636180 995466
rect 637040 995438 637376 995466
rect 638572 995438 638908 995466
rect 634726 995415 634782 995424
rect 631690 995344 631746 995353
rect 631336 995302 631690 995330
rect 631690 995279 631746 995288
rect 635844 994838 635872 995438
rect 635832 994832 635884 994838
rect 635832 994774 635884 994780
rect 625344 994696 625396 994702
rect 625344 994638 625396 994644
rect 630220 994696 630272 994702
rect 630220 994638 630272 994644
rect 591304 994560 591356 994566
rect 591304 994502 591356 994508
rect 574744 993948 574796 993954
rect 574744 993890 574796 993896
rect 568210 993712 568266 993721
rect 568210 993647 568266 993656
rect 637040 993410 637068 995438
rect 638880 995042 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640996 995438 641056 995466
rect 638868 995036 638920 995042
rect 638868 994978 638920 994984
rect 639064 994430 639092 995438
rect 639052 994424 639104 994430
rect 639052 994366 639104 994372
rect 639524 993546 639552 995438
rect 640800 995036 640852 995042
rect 640800 994978 640852 994984
rect 639512 993540 639564 993546
rect 639512 993482 639564 993488
rect 637028 993404 637080 993410
rect 637028 993346 637080 993352
rect 608600 993064 608652 993070
rect 608600 993006 608652 993012
rect 576306 990992 576362 991001
rect 576306 990927 576362 990936
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565268 985992 565320 985998
rect 565268 985934 565320 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 990927
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608612 983634 608640 993006
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 608612 983606 608810 983634
rect 624988 983620 625016 985934
rect 640812 983634 640840 994978
rect 640996 994906 641024 995438
rect 660578 995072 660634 995081
rect 641720 995036 641772 995042
rect 660578 995007 660580 995016
rect 641720 994978 641772 994984
rect 660632 995007 660634 995016
rect 640984 994900 641036 994906
rect 640984 994842 641036 994848
rect 641732 993721 641760 994978
rect 660580 994977 660632 994983
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993818 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660764 993812 660816 993818
rect 660764 993754 660816 993760
rect 641718 993712 641774 993721
rect 660960 993682 660988 994502
rect 641718 993647 641774 993656
rect 660948 993676 661000 993682
rect 660948 993618 661000 993624
rect 660304 992928 660356 992934
rect 660304 992870 660356 992876
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 660316 937281 660344 992870
rect 668584 990276 668636 990282
rect 668584 990218 668636 990224
rect 667204 975724 667256 975730
rect 667204 975666 667256 975672
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660302 937272 660358 937281
rect 660302 937207 660358 937216
rect 661696 937038 661724 957743
rect 663064 948116 663116 948122
rect 663064 948058 663116 948064
rect 663076 941769 663104 948058
rect 663062 941760 663118 941769
rect 663062 941695 663118 941704
rect 665836 939865 665864 961862
rect 667216 947345 667244 975666
rect 667202 947336 667258 947345
rect 667202 947271 667258 947280
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 668596 937825 668624 990218
rect 669964 990140 670016 990146
rect 669964 990082 670016 990088
rect 669976 938777 670004 990082
rect 675680 966521 675708 966723
rect 675666 966512 675722 966521
rect 675666 966447 675722 966456
rect 674300 966062 675418 966090
rect 673366 962840 673422 962849
rect 673366 962775 673422 962784
rect 673182 958216 673238 958225
rect 673182 958151 673238 958160
rect 672998 952232 673054 952241
rect 672998 952167 673054 952176
rect 669962 938768 670018 938777
rect 669962 938703 670018 938712
rect 671802 938360 671858 938369
rect 671802 938295 671858 938304
rect 668582 937816 668638 937825
rect 668582 937751 668638 937760
rect 671434 937544 671490 937553
rect 671434 937479 671490 937488
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 663064 921868 663116 921874
rect 663064 921810 663116 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 55862 892800 55918 892809
rect 55862 892735 55918 892744
rect 54482 892256 54538 892265
rect 54482 892191 54538 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62762 858664 62818 858673
rect 62762 858599 62818 858608
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799640 53158 799649
rect 53102 799575 53158 799584
rect 54496 774353 54524 844562
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 55876 772857 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62120 793600
rect 62172 793591 62174 793600
rect 62120 793562 62172 793568
rect 62776 788633 62804 858599
rect 651470 856352 651526 856361
rect 651470 856287 651526 856296
rect 651484 852174 651512 856287
rect 651472 852168 651524 852174
rect 651472 852110 651524 852116
rect 651838 843024 651894 843033
rect 651838 842959 651894 842968
rect 651852 841838 651880 842959
rect 651840 841832 651892 841838
rect 651840 841774 651892 841780
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 55862 772848 55918 772857
rect 55862 772783 55918 772792
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 669352 49018 669361
rect 48962 669287 49018 669296
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47398 638208 47454 638217
rect 47398 638143 47454 638152
rect 47412 618769 47440 638143
rect 47398 618760 47454 618769
rect 47398 618695 47454 618704
rect 47214 611008 47270 611017
rect 47214 610943 47270 610952
rect 45374 598904 45430 598913
rect 45374 598839 45430 598848
rect 45190 598088 45246 598097
rect 45190 598023 45246 598032
rect 47596 580553 47624 662390
rect 50356 626657 50384 714818
rect 51736 691393 51764 753510
rect 62776 743073 62804 780399
rect 652390 776656 652446 776665
rect 652390 776591 652446 776600
rect 652404 775606 652432 776591
rect 652392 775600 652444 775606
rect 652392 775542 652444 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 652022 736808 652078 736817
rect 652022 736743 652078 736752
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 54484 647896 54536 647902
rect 54484 647838 54536 647844
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 50342 626648 50398 626657
rect 50342 626583 50398 626592
rect 48964 623824 49016 623830
rect 48964 623766 49016 623772
rect 48976 601361 49004 623766
rect 51736 601769 51764 636210
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 48962 601352 49018 601361
rect 48962 601287 49018 601296
rect 54496 600953 54524 647838
rect 55876 643249 55904 701014
rect 62776 689489 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 651470 710288 651526 710297
rect 651470 710223 651526 710232
rect 651484 709374 651512 710223
rect 651472 709368 651524 709374
rect 651472 709310 651524 709316
rect 651472 696992 651524 696998
rect 651470 696960 651472 696969
rect 651524 696960 651526 696969
rect 651470 696895 651526 696904
rect 62762 689480 62818 689489
rect 62762 689415 62818 689424
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 651654 683632 651710 683641
rect 651654 683567 651710 683576
rect 651668 683194 651696 683567
rect 651656 683188 651708 683194
rect 651656 683130 651708 683136
rect 62762 676152 62818 676161
rect 62762 676087 62818 676096
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 62776 656169 62804 676087
rect 651470 670440 651526 670449
rect 651470 670375 651526 670384
rect 651484 669390 651512 670375
rect 651472 669384 651524 669390
rect 651472 669326 651524 669332
rect 651470 657112 651526 657121
rect 651470 657047 651526 657056
rect 651484 656946 651512 657047
rect 651472 656940 651524 656946
rect 651472 656882 651524 656888
rect 62762 656160 62818 656169
rect 62762 656095 62818 656104
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 651562 630592 651618 630601
rect 651562 630527 651618 630536
rect 651576 628590 651604 630527
rect 651564 628584 651616 628590
rect 652036 628561 652064 736743
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 661684 815652 661736 815658
rect 661684 815594 661736 815600
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 658924 683188 658976 683194
rect 658924 683130 658976 683136
rect 651564 628526 651616 628532
rect 652022 628552 652078 628561
rect 652022 628487 652078 628496
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 54482 600944 54538 600953
rect 54482 600879 54538 600888
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 580544 47638 580553
rect 47582 580479 47638 580488
rect 48976 557705 49004 597518
rect 50344 583772 50396 583778
rect 50344 583714 50396 583720
rect 50356 558521 50384 583714
rect 50342 558512 50398 558521
rect 50342 558447 50398 558456
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 48962 557696 49018 557705
rect 48962 557631 49018 557640
rect 45558 556880 45614 556889
rect 45558 556815 45614 556824
rect 45006 556472 45062 556481
rect 45006 556407 45062 556416
rect 44914 556064 44970 556073
rect 44914 555999 44970 556008
rect 44638 555656 44694 555665
rect 44638 555591 44694 555600
rect 44730 555248 44786 555257
rect 44730 555183 44786 555192
rect 44362 554432 44418 554441
rect 44362 554367 44418 554376
rect 44178 549128 44234 549137
rect 44178 549063 44234 549072
rect 43626 548176 43682 548185
rect 43626 548111 43682 548120
rect 43640 379514 43668 548111
rect 43810 547088 43866 547097
rect 43810 547023 43866 547032
rect 43456 379486 43576 379514
rect 43640 379486 43760 379514
rect 42982 379400 43038 379409
rect 42982 379335 43038 379344
rect 42996 365809 43024 379335
rect 43350 371920 43406 371929
rect 43350 371855 43406 371864
rect 42982 365800 43038 365809
rect 42982 365735 43038 365744
rect 42536 356646 42840 356674
rect 42536 356606 42564 356646
rect 42168 356538 42196 356592
rect 42260 356578 42564 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 42430 356144 42486 356153
rect 42430 356079 42486 356088
rect 42444 355926 42472 356079
rect 42182 355898 42472 355926
rect 43364 355881 43392 371855
rect 43350 355872 43406 355881
rect 43350 355807 43406 355816
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 43548 355314 43576 379486
rect 43732 355586 43760 379486
rect 43824 355722 43852 547023
rect 44192 537441 44220 549063
rect 44178 537432 44234 537441
rect 44178 537367 44234 537376
rect 44376 431954 44404 554367
rect 44546 550760 44602 550769
rect 44546 550695 44602 550704
rect 44560 532817 44588 550695
rect 44546 532808 44602 532817
rect 44546 532743 44602 532752
rect 44192 431926 44404 431954
rect 44192 427281 44220 431926
rect 44546 429312 44602 429321
rect 44546 429247 44602 429256
rect 44362 427680 44418 427689
rect 44362 427615 44418 427624
rect 44178 427272 44234 427281
rect 44178 427207 44234 427216
rect 44178 421560 44234 421569
rect 44178 421495 44234 421504
rect 43994 419520 44050 419529
rect 43994 419455 44050 419464
rect 44008 355858 44036 419455
rect 44192 406881 44220 421495
rect 44178 406872 44234 406881
rect 44178 406807 44234 406816
rect 44376 384849 44404 427615
rect 44560 386753 44588 429247
rect 44744 428097 44772 555183
rect 44928 428913 44956 555999
rect 45098 551576 45154 551585
rect 45098 551511 45154 551520
rect 45112 529825 45140 551511
rect 45282 548720 45338 548729
rect 45282 548655 45338 548664
rect 45296 537033 45324 548655
rect 45282 537024 45338 537033
rect 45282 536959 45338 536968
rect 45098 529816 45154 529825
rect 45098 529751 45154 529760
rect 45572 429729 45600 556815
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 45558 429720 45614 429729
rect 45558 429655 45614 429664
rect 44914 428904 44970 428913
rect 44914 428839 44970 428848
rect 45006 428496 45062 428505
rect 45006 428431 45062 428440
rect 44730 428088 44786 428097
rect 44730 428023 44786 428032
rect 44822 420744 44878 420753
rect 44822 420679 44878 420688
rect 44546 386744 44602 386753
rect 44546 386679 44602 386688
rect 44638 386064 44694 386073
rect 44638 385999 44694 386008
rect 44652 385490 44680 385999
rect 44640 385484 44692 385490
rect 44640 385426 44692 385432
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44362 384840 44418 384849
rect 44362 384775 44418 384784
rect 44454 379944 44510 379953
rect 44454 379879 44510 379888
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 44284 356697 44312 377431
rect 44468 359961 44496 379879
rect 44652 379514 44680 385183
rect 44836 379514 44864 420679
rect 45020 402974 45048 428431
rect 45190 426864 45246 426873
rect 45190 426799 45246 426808
rect 45020 402946 45140 402974
rect 45112 385665 45140 402946
rect 45204 393314 45232 426799
rect 45374 423192 45430 423201
rect 45374 423127 45430 423136
rect 45388 402937 45416 423127
rect 45374 402928 45430 402937
rect 45374 402863 45430 402872
rect 45204 393286 45416 393314
rect 45098 385656 45154 385665
rect 45098 385591 45154 385600
rect 45008 385484 45060 385490
rect 45008 385426 45060 385432
rect 44652 379486 44772 379514
rect 44836 379486 44956 379514
rect 44744 360194 44772 379486
rect 44744 360166 44864 360194
rect 44454 359952 44510 359961
rect 44454 359887 44510 359896
rect 44270 356688 44326 356697
rect 44270 356623 44326 356632
rect 44008 355830 44312 355858
rect 44284 355722 44312 355830
rect 43824 355694 44220 355722
rect 44284 355706 44680 355722
rect 44284 355700 44692 355706
rect 44284 355694 44640 355700
rect 44192 355586 44220 355694
rect 44640 355642 44692 355648
rect 43732 355558 43944 355586
rect 44192 355558 44772 355586
rect 43916 355450 43944 355558
rect 43916 355422 44128 355450
rect 43548 355286 44036 355314
rect 44008 354634 44036 355286
rect 44100 354906 44128 355422
rect 44100 354890 44615 354906
rect 44100 354884 44627 354890
rect 44100 354878 44575 354884
rect 44575 354826 44627 354832
rect 44575 354680 44627 354686
rect 44008 354628 44575 354634
rect 44008 354622 44627 354628
rect 44008 354606 44615 354622
rect 44744 354498 44772 355558
rect 44836 354634 44864 360166
rect 44928 357434 44956 379486
rect 45020 360194 45048 385426
rect 45190 384432 45246 384441
rect 45190 384367 45246 384376
rect 45204 383874 45232 384367
rect 45388 384033 45416 393286
rect 45374 384024 45430 384033
rect 45374 383959 45430 383968
rect 45204 383846 45416 383874
rect 45190 383616 45246 383625
rect 45190 383551 45246 383560
rect 45204 379514 45232 383551
rect 45204 379486 45324 379514
rect 45020 360166 45232 360194
rect 44928 357406 45048 357434
rect 45020 355842 45048 357406
rect 45008 355836 45060 355842
rect 45008 355778 45060 355784
rect 44836 354606 44956 354634
rect 44744 354482 44839 354498
rect 44744 354476 44851 354482
rect 44744 354470 44799 354476
rect 44799 354418 44851 354424
rect 44686 354340 44738 354346
rect 44686 354282 44738 354288
rect 43902 354240 43958 354249
rect 44698 354226 44726 354282
rect 43958 354198 44726 354226
rect 43902 354175 43958 354184
rect 44730 353832 44786 353841
rect 44928 353818 44956 354606
rect 45204 354090 45232 360166
rect 44786 353790 44956 353818
rect 45020 354062 45232 354090
rect 44730 353767 44786 353776
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 40222 345536 40278 345545
rect 40222 345471 40278 345480
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 35806 343904 35862 343913
rect 35806 343839 35862 343848
rect 35820 343670 35848 343839
rect 40236 343670 40264 345471
rect 35808 343664 35860 343670
rect 35808 343606 35860 343612
rect 40224 343664 40276 343670
rect 40224 343606 40276 343612
rect 45020 343369 45048 354062
rect 45296 345014 45324 379486
rect 45204 344986 45324 345014
rect 45006 343360 45062 343369
rect 45006 343295 45062 343304
rect 45204 340921 45232 344986
rect 45388 341737 45416 383846
rect 45558 380352 45614 380361
rect 45558 380287 45614 380296
rect 45572 357377 45600 380287
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 426456 46994 426465
rect 46938 426391 46994 426400
rect 46952 399809 46980 426391
rect 47122 423600 47178 423609
rect 47122 423535 47178 423544
rect 47136 400217 47164 423535
rect 47122 400208 47178 400217
rect 47122 400143 47178 400152
rect 46938 399800 46994 399809
rect 46938 399735 46994 399744
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 46938 380760 46994 380769
rect 46938 380695 46994 380704
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 46388 362976 46440 362982
rect 46388 362918 46440 362924
rect 45558 357368 45614 357377
rect 45558 357303 45614 357312
rect 45650 356688 45706 356697
rect 45480 356646 45650 356674
rect 45480 353274 45508 356646
rect 45650 356623 45706 356632
rect 45926 355872 45982 355881
rect 45652 355836 45704 355842
rect 45926 355807 45982 355816
rect 45652 355778 45704 355784
rect 45664 354074 45692 355778
rect 45652 354068 45704 354074
rect 45652 354010 45704 354016
rect 45940 353802 45968 355807
rect 45928 353796 45980 353802
rect 45928 353738 45980 353744
rect 45480 353258 45600 353274
rect 45480 353252 45612 353258
rect 45480 353246 45560 353252
rect 45560 353194 45612 353200
rect 45374 341728 45430 341737
rect 45374 341663 45430 341672
rect 45466 341320 45522 341329
rect 45466 341255 45522 341264
rect 45190 340912 45246 340921
rect 45190 340847 45246 340856
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 36636 339516 36688 339522
rect 36636 339458 36688 339464
rect 36648 336569 36676 339458
rect 36634 336560 36690 336569
rect 36634 336495 36690 336504
rect 42798 334656 42854 334665
rect 42798 334591 42854 334600
rect 43074 334656 43130 334665
rect 43074 334591 43130 334600
rect 41602 334520 41658 334529
rect 41602 334455 41658 334464
rect 41616 333713 41644 334455
rect 41602 333704 41658 333713
rect 41602 333639 41658 333648
rect 41786 326768 41842 326777
rect 41786 326703 41842 326712
rect 41800 326264 41828 326703
rect 42812 325694 42840 334591
rect 42812 325666 42932 325694
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41878 324864 41934 324873
rect 41878 324799 41934 324808
rect 41892 324428 41920 324799
rect 42182 323734 42564 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42536 321473 42564 323734
rect 42522 321464 42578 321473
rect 42522 321399 42578 321408
rect 42182 321354 42288 321382
rect 42260 321201 42288 321354
rect 42246 321192 42302 321201
rect 42246 321127 42302 321136
rect 42430 320920 42486 320929
rect 42430 320855 42486 320864
rect 42444 320739 42472 320855
rect 42182 320711 42472 320739
rect 42904 320090 42932 325666
rect 43088 322833 43116 334591
rect 44178 334384 44234 334393
rect 44178 334319 44234 334328
rect 43258 333704 43314 333713
rect 43258 333639 43314 333648
rect 43074 322824 43130 322833
rect 43074 322759 43130 322768
rect 43272 321201 43300 333639
rect 43258 321192 43314 321201
rect 43258 321127 43314 321136
rect 44192 320929 44220 334319
rect 44178 320920 44234 320929
rect 44178 320855 44234 320864
rect 42182 320062 42932 320090
rect 41786 319968 41842 319977
rect 41786 319903 41842 319912
rect 41800 319532 41828 319903
rect 42246 317520 42302 317529
rect 42246 317455 42302 317464
rect 42260 317059 42288 317455
rect 42182 317031 42288 317059
rect 41786 316704 41842 316713
rect 41786 316639 41842 316648
rect 41800 316404 41828 316639
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 42154 315480 42210 315489
rect 42154 315415 42210 315424
rect 42168 315180 42196 315415
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42154 312352 42210 312361
rect 42154 312287 42210 312296
rect 42168 312052 42196 312287
rect 44546 311536 44602 311545
rect 44546 311471 44602 311480
rect 44362 311264 44418 311273
rect 44362 311199 44418 311208
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 44376 299305 44404 311199
rect 44560 300121 44588 311471
rect 44546 300112 44602 300121
rect 44546 300047 44602 300056
rect 44638 299704 44694 299713
rect 44638 299639 44694 299648
rect 44362 299296 44418 299305
rect 44362 299231 44418 299240
rect 42890 298072 42946 298081
rect 42890 298007 42946 298016
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 37922 294808 37978 294817
rect 37922 294743 37978 294752
rect 37936 284782 37964 294743
rect 41800 292777 41828 296783
rect 42062 296032 42118 296041
rect 42062 295967 42118 295976
rect 41786 292768 41842 292777
rect 41786 292703 41842 292712
rect 42076 292369 42104 295967
rect 42062 292360 42118 292369
rect 42062 292295 42118 292304
rect 42246 291136 42302 291145
rect 42246 291071 42302 291080
rect 42062 290456 42118 290465
rect 42062 290391 42118 290400
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 284986 41368 290255
rect 42076 289921 42104 290391
rect 42260 289921 42288 291071
rect 42062 289912 42118 289921
rect 42062 289847 42118 289856
rect 42246 289912 42302 289921
rect 42246 289847 42302 289856
rect 41708 284986 42472 285002
rect 41328 284980 41380 284986
rect 41328 284922 41380 284928
rect 41696 284980 42472 284986
rect 41748 284974 42472 284980
rect 41696 284922 41748 284928
rect 37924 284776 37976 284782
rect 37924 284718 37976 284724
rect 41696 284776 41748 284782
rect 41748 284724 42288 284730
rect 41696 284718 42288 284724
rect 41708 284702 42288 284718
rect 42260 283506 42288 284702
rect 42168 283478 42288 283506
rect 42168 283045 42196 283478
rect 42444 281874 42472 284974
rect 42182 281846 42472 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42430 278695 42486 278704
rect 42430 278216 42486 278225
rect 42168 278066 42196 278188
rect 42260 278174 42430 278202
rect 42260 278066 42288 278174
rect 42430 278151 42486 278160
rect 42168 278038 42288 278066
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 41800 277508 41828 277879
rect 42338 277672 42394 277681
rect 42338 277607 42394 277616
rect 42154 277400 42210 277409
rect 42154 277335 42210 277344
rect 42168 276896 42196 277335
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42062 273456 42118 273465
rect 42062 273391 42118 273400
rect 42076 273224 42104 273391
rect 42062 272912 42118 272921
rect 42062 272847 42118 272856
rect 42076 272544 42104 272847
rect 42352 272014 42380 277607
rect 42182 271986 42380 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 42430 270464 42486 270473
rect 42430 270399 42486 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 270399
rect 42182 269507 42472 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 35806 259992 35862 260001
rect 35806 259927 35862 259936
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35820 258369 35848 259927
rect 35806 258360 35862 258369
rect 35806 258295 35862 258304
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42904 255241 42932 298007
rect 43258 297256 43314 297265
rect 43258 297191 43314 297200
rect 43074 293584 43130 293593
rect 43074 293519 43130 293528
rect 43088 273465 43116 293519
rect 43074 273456 43130 273465
rect 43074 273391 43130 273400
rect 42890 255232 42946 255241
rect 42890 255167 42946 255176
rect 42890 254824 42946 254833
rect 42890 254759 42946 254768
rect 35806 253464 35862 253473
rect 35806 253399 35862 253408
rect 35622 253056 35678 253065
rect 35622 252991 35678 253000
rect 35636 252754 35664 252991
rect 35820 252890 35848 253399
rect 35808 252884 35860 252890
rect 35808 252826 35860 252832
rect 41328 252884 41380 252890
rect 41328 252826 41380 252832
rect 35624 252748 35676 252754
rect 35624 252690 35676 252696
rect 35806 252648 35862 252657
rect 35806 252583 35808 252592
rect 35860 252583 35862 252592
rect 40684 252612 40736 252618
rect 35808 252554 35860 252560
rect 40684 252554 40736 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 37924 251252 37976 251258
rect 37924 251194 37976 251200
rect 37936 242894 37964 251194
rect 37924 242888 37976 242894
rect 37924 242830 37976 242836
rect 40696 242593 40724 252554
rect 41340 252249 41368 252826
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 41326 252240 41382 252249
rect 41326 252175 41382 252184
rect 41708 248414 41736 252690
rect 42522 252240 42578 252249
rect 42522 252175 42578 252184
rect 41708 248386 42288 248414
rect 41696 242888 41748 242894
rect 41694 242856 41696 242865
rect 41748 242856 41750 242865
rect 41694 242791 41750 242800
rect 40682 242584 40738 242593
rect 40682 242519 40738 242528
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42076 238513 42104 238649
rect 42062 238504 42118 238513
rect 42062 238439 42118 238448
rect 42260 238014 42288 248386
rect 42536 238762 42564 252175
rect 42706 242856 42762 242865
rect 42706 242791 42762 242800
rect 42536 238734 42656 238762
rect 42182 237986 42288 238014
rect 42628 237538 42656 238734
rect 42536 237510 42656 237538
rect 42536 237425 42564 237510
rect 42522 237416 42578 237425
rect 42522 237351 42578 237360
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42182 234314 42472 234342
rect 42246 234152 42302 234161
rect 42246 234087 42302 234096
rect 42260 233695 42288 234087
rect 42182 233667 42288 233695
rect 42154 233336 42210 233345
rect 42154 233271 42210 233280
rect 42168 233104 42196 233271
rect 42444 232529 42472 234314
rect 42430 232520 42486 232529
rect 42430 232455 42486 232464
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 42154 230480 42210 230489
rect 42154 230415 42210 230424
rect 42168 229976 42196 230415
rect 42430 229392 42486 229401
rect 42182 229350 42430 229378
rect 42430 229327 42486 229336
rect 42720 229094 42748 242791
rect 42904 229094 42932 254759
rect 43272 254425 43300 297191
rect 43442 294400 43498 294409
rect 43442 294335 43498 294344
rect 43456 270473 43484 294335
rect 44362 293992 44418 294001
rect 44362 293927 44418 293936
rect 43626 293176 43682 293185
rect 43626 293111 43682 293120
rect 43640 279857 43668 293111
rect 43810 291952 43866 291961
rect 43810 291887 43866 291896
rect 43626 279848 43682 279857
rect 43626 279783 43682 279792
rect 43824 277409 43852 291887
rect 44178 291544 44234 291553
rect 44178 291479 44234 291488
rect 44192 278225 44220 291479
rect 44178 278216 44234 278225
rect 44178 278151 44234 278160
rect 43810 277400 43866 277409
rect 43810 277335 43866 277344
rect 44376 272921 44404 293927
rect 44362 272912 44418 272921
rect 44362 272847 44418 272856
rect 43442 270464 43498 270473
rect 43442 270399 43498 270408
rect 44652 256873 44680 299639
rect 45190 298888 45246 298897
rect 45190 298823 45246 298832
rect 45006 295216 45062 295225
rect 45006 295151 45062 295160
rect 44822 291952 44878 291961
rect 44822 291887 44878 291896
rect 44638 256864 44694 256873
rect 44638 256799 44694 256808
rect 43626 256456 43682 256465
rect 43626 256391 43682 256400
rect 43442 255640 43498 255649
rect 43442 255575 43498 255584
rect 43258 254416 43314 254425
rect 43258 254351 43314 254360
rect 43074 250336 43130 250345
rect 43074 250271 43130 250280
rect 43088 230489 43116 250271
rect 43258 242584 43314 242593
rect 43258 242519 43314 242528
rect 43074 230480 43130 230489
rect 43074 230415 43130 230424
rect 42536 229066 42748 229094
rect 42812 229066 42932 229094
rect 42536 228834 42564 229066
rect 42182 228806 42564 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 41694 224496 41750 224505
rect 41694 224431 41750 224440
rect 28538 222864 28594 222873
rect 28538 222799 28594 222808
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 28552 214305 28580 222799
rect 28538 214296 28594 214305
rect 28538 214231 28594 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 41708 213994 41736 224431
rect 42812 219434 42840 229066
rect 43272 225729 43300 242519
rect 43258 225720 43314 225729
rect 43258 225655 43314 225664
rect 42812 219406 42932 219434
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 35622 212256 35678 212265
rect 35622 212191 35678 212200
rect 35636 211342 35664 212191
rect 42904 212129 42932 219406
rect 43456 212945 43484 255575
rect 43640 213761 43668 256391
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43810 249112 43866 249121
rect 43810 249047 43866 249056
rect 43824 231849 43852 249047
rect 43810 231840 43866 231849
rect 43810 231775 43866 231784
rect 43626 213752 43682 213761
rect 43626 213687 43682 213696
rect 43442 212936 43498 212945
rect 43442 212871 43498 212880
rect 42890 212120 42946 212129
rect 42890 212055 42946 212064
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35624 211336 35676 211342
rect 35624 211278 35676 211284
rect 35820 211206 35848 211375
rect 41696 211336 41748 211342
rect 44192 211313 44220 253943
rect 44362 251968 44418 251977
rect 44362 251903 44418 251912
rect 44376 233345 44404 251903
rect 44546 248704 44602 248713
rect 44546 248639 44602 248648
rect 44560 234161 44588 248639
rect 44546 234152 44602 234161
rect 44546 234087 44602 234096
rect 44362 233336 44418 233345
rect 44362 233271 44418 233280
rect 44836 214985 44864 291887
rect 45020 276593 45048 295151
rect 45006 276584 45062 276593
rect 45006 276519 45062 276528
rect 45204 273254 45232 298823
rect 45480 298489 45508 341255
rect 45834 340096 45890 340105
rect 45834 340031 45890 340040
rect 45650 339280 45706 339289
rect 45650 339215 45706 339224
rect 45664 312361 45692 339215
rect 45848 313721 45876 340031
rect 46018 338872 46074 338881
rect 46018 338807 46074 338816
rect 46032 315489 46060 338807
rect 46204 336796 46256 336802
rect 46204 336738 46256 336744
rect 46018 315480 46074 315489
rect 46018 315415 46074 315424
rect 45834 313712 45890 313721
rect 45834 313647 45890 313656
rect 45650 312352 45706 312361
rect 45650 312287 45706 312296
rect 45466 298480 45522 298489
rect 45466 298415 45522 298424
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 45480 291961 45508 298114
rect 45466 291952 45522 291961
rect 45466 291887 45522 291896
rect 45112 273226 45232 273254
rect 45112 256057 45140 273226
rect 46216 260001 46244 336738
rect 46400 303113 46428 362918
rect 46952 356153 46980 380695
rect 47122 379128 47178 379137
rect 47122 379063 47178 379072
rect 47136 361593 47164 379063
rect 47122 361584 47178 361593
rect 47122 361519 47178 361528
rect 46938 356144 46994 356153
rect 46938 356079 46994 356088
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46386 303104 46442 303113
rect 46386 303039 46442 303048
rect 46202 259992 46258 260001
rect 46202 259927 46258 259936
rect 45098 256048 45154 256057
rect 45098 255983 45154 255992
rect 45558 251152 45614 251161
rect 45558 251087 45614 251096
rect 45006 248296 45062 248305
rect 45006 248231 45062 248240
rect 45020 235929 45048 248231
rect 45006 235920 45062 235929
rect 45006 235855 45062 235864
rect 45572 226681 45600 251087
rect 45834 250744 45890 250753
rect 45834 250679 45890 250688
rect 45848 229401 45876 250679
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 232529 46060 249455
rect 46202 247888 46258 247897
rect 46202 247823 46258 247832
rect 46018 232520 46074 232529
rect 46018 232455 46074 232464
rect 45834 229392 45890 229401
rect 45834 229327 45890 229336
rect 45558 226672 45614 226681
rect 45558 226607 45614 226616
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 44178 211304 44234 211313
rect 41748 211284 41920 211290
rect 41696 211278 41920 211284
rect 41708 211262 41920 211278
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 41696 211200 41748 211206
rect 41696 211142 41748 211148
rect 35808 209840 35860 209846
rect 35806 209808 35808 209817
rect 41328 209840 41380 209846
rect 35860 209808 35862 209817
rect 41328 209782 41380 209788
rect 35806 209743 35862 209752
rect 41340 205737 41368 209782
rect 41708 209001 41736 211142
rect 41694 208992 41750 209001
rect 41694 208927 41750 208936
rect 41326 205728 41382 205737
rect 41326 205663 41382 205672
rect 41142 204096 41198 204105
rect 41142 204031 41198 204040
rect 41156 200705 41184 204031
rect 41326 203688 41382 203697
rect 41326 203623 41382 203632
rect 41340 202201 41368 203623
rect 41326 202192 41382 202201
rect 41326 202127 41382 202136
rect 41892 201521 41920 211262
rect 44178 211239 44234 211248
rect 44178 210488 44234 210497
rect 44178 210423 44234 210432
rect 42798 209672 42854 209681
rect 42798 209607 42854 209616
rect 41878 201512 41934 201521
rect 41878 201447 41934 201456
rect 41142 200696 41198 200705
rect 41142 200631 41198 200640
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 41786 195800 41842 195809
rect 41786 195735 41842 195744
rect 41800 195432 41828 195735
rect 42246 195392 42302 195401
rect 42246 195327 42302 195336
rect 41970 195120 42026 195129
rect 41970 195055 42026 195064
rect 41984 194820 42012 195055
rect 42260 193225 42288 195327
rect 42246 193216 42302 193225
rect 42246 193151 42302 193160
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41786 187232 41842 187241
rect 41786 187167 41842 187176
rect 41800 186796 41828 187167
rect 42062 186416 42118 186425
rect 42062 186351 42118 186360
rect 42076 186184 42104 186351
rect 42154 185872 42210 185881
rect 42154 185807 42210 185816
rect 42168 185605 42196 185807
rect 42430 184920 42486 184929
rect 42430 184855 42486 184864
rect 42444 183779 42472 184855
rect 42182 183751 42472 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42812 182491 42840 209607
rect 43258 208040 43314 208049
rect 43258 207975 43314 207984
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 183161 43300 207975
rect 43626 206816 43682 206825
rect 43626 206751 43682 206760
rect 43442 200696 43498 200705
rect 43442 200631 43498 200640
rect 43258 183152 43314 183161
rect 43258 183087 43314 183096
rect 42182 182463 42840 182491
rect 43456 42838 43484 200631
rect 43640 193225 43668 206751
rect 43810 205320 43866 205329
rect 43810 205255 43866 205264
rect 43626 193216 43682 193225
rect 43626 193151 43682 193160
rect 43824 190505 43852 205255
rect 43994 204912 44050 204921
rect 43994 204847 44050 204856
rect 44008 191729 44036 204847
rect 43994 191720 44050 191729
rect 43994 191655 44050 191664
rect 43810 190496 43866 190505
rect 43810 190431 43866 190440
rect 44192 184929 44220 210423
rect 44546 208584 44602 208593
rect 44546 208519 44602 208528
rect 44362 206000 44418 206009
rect 44362 205935 44418 205944
rect 44376 187649 44404 205935
rect 44560 189961 44588 208519
rect 44822 204504 44878 204513
rect 44822 204439 44878 204448
rect 44546 189952 44602 189961
rect 44546 189887 44602 189896
rect 44362 187640 44418 187649
rect 44362 187575 44418 187584
rect 44178 184920 44234 184929
rect 44178 184855 44234 184864
rect 44836 74534 44864 204439
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 247823
rect 46938 247072 46994 247081
rect 46938 247007 46994 247016
rect 46952 238513 46980 247007
rect 46938 238504 46994 238513
rect 46938 238439 46994 238448
rect 46386 203552 46442 203561
rect 46386 203487 46442 203496
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 46400 51746 46428 203487
rect 47596 51882 47624 333095
rect 47780 300529 47808 389234
rect 48976 386889 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 48962 386880 49018 386889
rect 48962 386815 49018 386824
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51724 375420 51776 375426
rect 51724 375362 51776 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47584 51876 47636 51882
rect 47584 51818 47636 51824
rect 46388 51740 46440 51746
rect 46388 51682 46440 51688
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 47780 49026 47808 247415
rect 47950 213344 48006 213353
rect 47950 213279 48006 213288
rect 47964 190505 47992 213279
rect 48134 210896 48190 210905
rect 48134 210831 48190 210840
rect 48148 194449 48176 210831
rect 48134 194440 48190 194449
rect 48134 194375 48190 194384
rect 47950 190496 48006 190505
rect 47950 190431 48006 190440
rect 48976 52018 49004 334047
rect 51736 301345 51764 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 652390 590744 652446 590753
rect 652390 590679 652392 590688
rect 652444 590679 652446 590688
rect 652392 590650 652444 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 658936 579737 658964 683130
rect 660316 625297 660344 763166
rect 661696 673169 661724 815594
rect 663076 760481 663104 921810
rect 665824 909492 665876 909498
rect 665824 909434 665876 909440
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868737 664484 881826
rect 664442 868728 664498 868737
rect 664442 868663 664498 868672
rect 664444 852168 664496 852174
rect 664444 852110 664496 852116
rect 663062 760472 663118 760481
rect 663062 760407 663118 760416
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 663076 689353 663104 723114
rect 664456 716553 664484 852110
rect 665836 761569 665864 909434
rect 670976 895688 671028 895694
rect 670976 895630 671028 895636
rect 670606 876888 670662 876897
rect 670606 876823 670662 876832
rect 669226 876344 669282 876353
rect 669226 876279 669282 876288
rect 668858 872264 668914 872273
rect 668858 872199 668914 872208
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666282 778424 666338 778433
rect 666282 778359 666338 778368
rect 665822 761560 665878 761569
rect 665822 761495 665878 761504
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 661682 673160 661738 673169
rect 661682 673095 661738 673104
rect 661684 669384 661736 669390
rect 661684 669326 661736 669332
rect 661696 643793 661724 669326
rect 663064 656940 663116 656946
rect 663064 656882 663116 656888
rect 661682 643784 661738 643793
rect 661682 643719 661738 643728
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 660316 599593 660344 616830
rect 661684 603152 661736 603158
rect 661684 603094 661736 603100
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 658922 579728 658978 579737
rect 658922 579663 658978 579672
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 658936 554033 658964 563042
rect 658922 554024 658978 554033
rect 658922 553959 658978 553968
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 652574 497720 652630 497729
rect 652574 497655 652630 497664
rect 652588 494766 652616 497655
rect 652576 494760 652628 494766
rect 652576 494702 652628 494708
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62946 415440 63002 415449
rect 62946 415375 63002 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 53288 322992 53340 322998
rect 53288 322934 53340 322940
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 49146 290456 49202 290465
rect 49146 290391 49202 290400
rect 49160 53378 49188 290391
rect 50342 290184 50398 290193
rect 50342 290119 50398 290128
rect 49606 208992 49662 209001
rect 49606 208927 49662 208936
rect 49422 201512 49478 201521
rect 49422 201447 49478 201456
rect 49436 192409 49464 201447
rect 49620 196489 49648 208927
rect 49606 196480 49662 196489
rect 49606 196415 49662 196424
rect 49422 192400 49478 192409
rect 49422 192335 49478 192344
rect 49148 53372 49200 53378
rect 49148 53314 49200 53320
rect 50356 53242 50384 290119
rect 51722 289912 51778 289921
rect 51722 289847 51778 289856
rect 50526 246528 50582 246537
rect 50526 246463 50582 246472
rect 50344 53236 50396 53242
rect 50344 53178 50396 53184
rect 48964 52012 49016 52018
rect 48964 51954 49016 51960
rect 50540 50522 50568 246463
rect 50528 50516 50580 50522
rect 50528 50458 50580 50464
rect 51736 49162 51764 289847
rect 53300 257553 53328 322934
rect 54484 310548 54536 310554
rect 54484 310490 54536 310496
rect 53286 257544 53342 257553
rect 53286 257479 53342 257488
rect 54496 222873 54524 310490
rect 55876 278769 55904 401610
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 62776 267073 62804 350231
rect 62960 345681 62988 415375
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 651838 364848 651894 364857
rect 651838 364783 651894 364792
rect 651852 364410 651880 364783
rect 651840 364404 651892 364410
rect 651840 364346 651892 364352
rect 652390 351656 652446 351665
rect 652390 351591 652446 351600
rect 652404 350606 652432 351591
rect 652392 350600 652444 350606
rect 652392 350542 652444 350548
rect 62946 345672 63002 345681
rect 62946 345607 63002 345616
rect 652022 338328 652078 338337
rect 652022 338263 652078 338272
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 651484 310554 651512 311743
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62946 285152 63002 285161
rect 62946 285087 63002 285096
rect 62762 267064 62818 267073
rect 62762 266999 62818 267008
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 54482 222864 54538 222873
rect 54482 222799 54538 222808
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 60004 225752 60056 225758
rect 60004 225694 60056 225700
rect 58990 224224 59046 224233
rect 58990 224159 59046 224168
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217274 59032 224159
rect 59820 219020 59872 219026
rect 59820 218962 59872 218968
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218962
rect 60016 218074 60044 225694
rect 62028 225616 62080 225622
rect 62028 225558 62080 225564
rect 60648 221740 60700 221746
rect 60648 221682 60700 221688
rect 60004 218068 60056 218074
rect 60004 218010 60056 218016
rect 60660 217274 60688 221682
rect 62040 218074 62068 225558
rect 62960 224505 62988 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 272542 65932 277780
rect 67022 277766 67588 277794
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 67560 270094 67588 277766
rect 68204 271318 68232 277780
rect 68192 271312 68244 271318
rect 68192 271254 68244 271260
rect 67548 270088 67600 270094
rect 67548 270030 67600 270036
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274718 71820 277780
rect 71780 274712 71832 274718
rect 71780 274654 71832 274660
rect 72988 271182 73016 277780
rect 74092 274718 74120 277780
rect 73804 274712 73856 274718
rect 73804 274654 73856 274660
rect 74080 274712 74132 274718
rect 74080 274654 74132 274660
rect 72976 271176 73028 271182
rect 72976 271118 73028 271124
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 73816 267034 73844 274654
rect 75288 274106 75316 277780
rect 76484 275466 76512 277780
rect 76472 275460 76524 275466
rect 76472 275402 76524 275408
rect 77208 274712 77260 274718
rect 77208 274654 77260 274660
rect 75276 274100 75328 274106
rect 75276 274042 75328 274048
rect 75920 270088 75972 270094
rect 75920 270030 75972 270036
rect 75932 267073 75960 270030
rect 77220 269958 77248 274654
rect 77680 273970 77708 277780
rect 77668 273964 77720 273970
rect 77668 273906 77720 273912
rect 78876 270366 78904 277780
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 270094 80100 277780
rect 81268 274990 81296 277780
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 82372 272678 82400 277780
rect 82360 272672 82412 272678
rect 82360 272614 82412 272620
rect 83568 271046 83596 277780
rect 84778 277766 85528 277794
rect 83556 271040 83608 271046
rect 83556 270982 83608 270988
rect 85500 270230 85528 277766
rect 85960 275602 85988 277780
rect 85948 275596 86000 275602
rect 85948 275538 86000 275544
rect 86224 274984 86276 274990
rect 86224 274926 86276 274932
rect 85488 270224 85540 270230
rect 85488 270166 85540 270172
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 77208 269952 77260 269958
rect 77208 269894 77260 269900
rect 86236 267170 86264 274926
rect 87156 268394 87184 277780
rect 88352 275874 88380 277780
rect 88340 275868 88392 275874
rect 88340 275810 88392 275816
rect 89548 271454 89576 277780
rect 90666 277766 91048 277794
rect 91862 277766 92428 277794
rect 89536 271448 89588 271454
rect 89536 271390 89588 271396
rect 91020 268666 91048 277766
rect 91008 268660 91060 268666
rect 91008 268602 91060 268608
rect 92400 268530 92428 277766
rect 93044 274378 93072 277780
rect 93032 274372 93084 274378
rect 93032 274314 93084 274320
rect 94240 272814 94268 277780
rect 95436 274242 95464 277780
rect 96632 275738 96660 277780
rect 96620 275732 96672 275738
rect 96620 275674 96672 275680
rect 97736 274378 97764 277780
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 101338 277766 102088 277794
rect 95884 274372 95936 274378
rect 95884 274314 95936 274320
rect 97724 274372 97776 274378
rect 97724 274314 97776 274320
rect 95424 274236 95476 274242
rect 95424 274178 95476 274184
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 87144 268388 87196 268394
rect 87144 268330 87196 268336
rect 95896 267306 95924 274314
rect 99300 268802 99328 277766
rect 100680 270502 100708 277766
rect 100668 270496 100720 270502
rect 100668 270438 100720 270444
rect 102060 269793 102088 277766
rect 102520 272950 102548 277780
rect 103716 276010 103744 277780
rect 103704 276004 103756 276010
rect 103704 275946 103756 275952
rect 102508 272944 102560 272950
rect 102508 272886 102560 272892
rect 104912 271726 104940 277780
rect 104900 271720 104952 271726
rect 104900 271662 104952 271668
rect 106016 271590 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 271584 106056 271590
rect 106004 271526 106056 271532
rect 102046 269784 102102 269793
rect 102046 269719 102102 269728
rect 99288 268796 99340 268802
rect 99288 268738 99340 268744
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 99300 267578 99328 268602
rect 107580 267734 107608 277766
rect 108960 268938 108988 277766
rect 108948 268932 109000 268938
rect 108948 268874 109000 268880
rect 110248 268802 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 111996 273086 112024 277780
rect 111984 273080 112036 273086
rect 111984 273022 112036 273028
rect 113192 270774 113220 277780
rect 114296 274514 114324 277780
rect 115506 277766 115888 277794
rect 114284 274508 114336 274514
rect 114284 274450 114336 274456
rect 113180 270768 113232 270774
rect 113180 270710 113232 270716
rect 115860 269074 115888 277766
rect 116688 272270 116716 277780
rect 117898 277766 118648 277794
rect 116676 272264 116728 272270
rect 116676 272206 116728 272212
rect 115848 269068 115900 269074
rect 115848 269010 115900 269016
rect 110236 268796 110288 268802
rect 110236 268738 110288 268744
rect 118620 268258 118648 277766
rect 119080 269686 119108 277780
rect 120276 274650 120304 277780
rect 120264 274644 120316 274650
rect 120264 274586 120316 274592
rect 121380 271862 121408 277780
rect 122590 277766 122788 277794
rect 121368 271856 121420 271862
rect 121368 271798 121420 271804
rect 122760 270502 122788 277766
rect 123772 271046 123800 277780
rect 124968 273698 124996 277780
rect 126178 277766 126928 277794
rect 124956 273692 125008 273698
rect 124956 273634 125008 273640
rect 123484 271040 123536 271046
rect 123484 270982 123536 270988
rect 123760 271040 123812 271046
rect 123760 270982 123812 270988
rect 119804 270496 119856 270502
rect 119804 270438 119856 270444
rect 122748 270496 122800 270502
rect 122748 270438 122800 270444
rect 119068 269680 119120 269686
rect 119068 269622 119120 269628
rect 118608 268252 118660 268258
rect 118608 268194 118660 268200
rect 107580 267706 107700 267734
rect 99288 267572 99340 267578
rect 99288 267514 99340 267520
rect 107672 267442 107700 267706
rect 107660 267436 107712 267442
rect 107660 267378 107712 267384
rect 95884 267300 95936 267306
rect 95884 267242 95936 267248
rect 86224 267164 86276 267170
rect 86224 267106 86276 267112
rect 75918 267064 75974 267073
rect 73804 267028 73856 267034
rect 75918 266999 75974 267008
rect 73804 266970 73856 266976
rect 119816 266898 119844 270438
rect 119804 266892 119856 266898
rect 119804 266834 119856 266840
rect 123496 266626 123524 270982
rect 126900 269550 126928 277766
rect 127360 272406 127388 277780
rect 128556 273222 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 130856 273834 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 273828 130896 273834
rect 130844 273770 130896 273776
rect 128544 273216 128596 273222
rect 128544 273158 128596 273164
rect 127348 272400 127400 272406
rect 127348 272342 127400 272348
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 132420 267714 132448 277766
rect 133800 270366 133828 277766
rect 134444 270910 134472 277780
rect 135640 275058 135668 277780
rect 136850 277766 137048 277794
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136088 274916 136140 274922
rect 136088 274858 136140 274864
rect 134432 270904 134484 270910
rect 134432 270846 134484 270852
rect 132592 270360 132644 270366
rect 132592 270302 132644 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 132408 267708 132460 267714
rect 132408 267650 132460 267656
rect 132604 266762 132632 270302
rect 136100 269414 136128 274858
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 136088 269408 136140 269414
rect 136088 269350 136140 269356
rect 132592 266756 132644 266762
rect 132592 266698 132644 266704
rect 123484 266620 123536 266626
rect 123484 266562 123536 266568
rect 136836 264330 136864 272478
rect 137020 268122 137048 277766
rect 137940 272542 137968 277780
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 139136 271318 139164 277780
rect 140346 277766 140728 277794
rect 141542 277766 141832 277794
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 138480 271312 138532 271318
rect 138480 271254 138532 271260
rect 139124 271312 139176 271318
rect 139124 271254 139176 271260
rect 137008 268116 137060 268122
rect 137008 268058 137060 268064
rect 138110 267064 138166 267073
rect 138110 266999 138166 267008
rect 136836 264302 137310 264330
rect 138124 264316 138152 266999
rect 138492 264330 138520 271254
rect 139768 269816 139820 269822
rect 139768 269758 139820 269764
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 140148 264330 140176 275266
rect 140700 269822 140728 277766
rect 141804 271318 141832 277766
rect 142724 274922 142752 277780
rect 143934 277766 144132 277794
rect 145038 277766 145328 277794
rect 143264 275460 143316 275466
rect 143264 275402 143316 275408
rect 142712 274916 142764 274922
rect 142712 274858 142764 274864
rect 142160 274100 142212 274106
rect 142160 274042 142212 274048
rect 141608 271312 141660 271318
rect 141608 271254 141660 271260
rect 141792 271312 141844 271318
rect 141792 271254 141844 271260
rect 140688 269816 140740 269822
rect 140688 269758 140740 269764
rect 141424 267028 141476 267034
rect 141424 266970 141476 266976
rect 140148 264302 140622 264330
rect 141436 264316 141464 266970
rect 141620 266490 141648 271254
rect 141608 266484 141660 266490
rect 141608 266426 141660 266432
rect 142172 265674 142200 274042
rect 143276 271182 143304 275402
rect 142344 271176 142396 271182
rect 142344 271118 142396 271124
rect 143264 271176 143316 271182
rect 143264 271118 143316 271124
rect 142160 265668 142212 265674
rect 142160 265610 142212 265616
rect 142356 265554 142384 271118
rect 144104 269958 144132 277766
rect 145300 273970 145328 277766
rect 146220 274786 146248 277780
rect 146944 275868 146996 275874
rect 146944 275810 146996 275816
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145104 273964 145156 273970
rect 145104 273906 145156 273912
rect 145288 273964 145340 273970
rect 145288 273906 145340 273912
rect 144368 271176 144420 271182
rect 144368 271118 144420 271124
rect 143908 269952 143960 269958
rect 143908 269894 143960 269900
rect 144092 269952 144144 269958
rect 144092 269894 144144 269900
rect 142804 265668 142856 265674
rect 142804 265610 142856 265616
rect 142264 265526 142384 265554
rect 142264 264316 142292 265526
rect 142816 264330 142844 265610
rect 142816 264302 143106 264330
rect 143920 264316 143948 269894
rect 144380 264330 144408 271118
rect 145116 264330 145144 273906
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 144380 264302 144762 264330
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 146956 269210 146984 275810
rect 147416 274106 147444 277780
rect 148612 275466 148640 277780
rect 149808 275874 149836 277780
rect 149796 275868 149848 275874
rect 149796 275810 149848 275816
rect 150808 275596 150860 275602
rect 150808 275538 150860 275544
rect 148600 275460 148652 275466
rect 148600 275402 148652 275408
rect 149704 274780 149756 274786
rect 149704 274722 149756 274728
rect 147404 274100 147456 274106
rect 147404 274042 147456 274048
rect 148416 273692 148468 273698
rect 148416 273634 148468 273640
rect 148232 272672 148284 272678
rect 148232 272614 148284 272620
rect 146944 269204 146996 269210
rect 146944 269146 146996 269152
rect 148244 267734 148272 272614
rect 148428 267734 148456 273634
rect 149428 270224 149480 270230
rect 149428 270166 149480 270172
rect 148244 267706 148364 267734
rect 148428 267706 148548 267734
rect 148048 267164 148100 267170
rect 148048 267106 148100 267112
rect 146944 267028 146996 267034
rect 146944 266970 146996 266976
rect 146956 266490 146984 266970
rect 147220 266756 147272 266762
rect 147220 266698 147272 266704
rect 146944 266484 146996 266490
rect 146944 266426 146996 266432
rect 147232 264316 147260 266698
rect 148060 264316 148088 267106
rect 148336 264466 148364 267706
rect 148520 266762 148548 267706
rect 148508 266756 148560 266762
rect 148508 266698 148560 266704
rect 148336 264438 148456 264466
rect 148428 264330 148456 264438
rect 149440 264330 149468 270166
rect 149716 267170 149744 274722
rect 150820 267734 150848 275538
rect 151004 274786 151032 277780
rect 150992 274780 151044 274786
rect 150992 274722 151044 274728
rect 152200 272134 152228 277780
rect 152740 274780 152792 274786
rect 152740 274722 152792 274728
rect 152188 272128 152240 272134
rect 152188 272070 152240 272076
rect 152372 271448 152424 271454
rect 152372 271390 152424 271396
rect 152188 268388 152240 268394
rect 152188 268330 152240 268336
rect 150820 267706 151032 267734
rect 149704 267164 149756 267170
rect 149704 267106 149756 267112
rect 150532 266620 150584 266626
rect 150532 266562 150584 266568
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266562
rect 151004 264330 151032 267706
rect 151004 264302 151386 264330
rect 152200 264316 152228 268330
rect 152384 267734 152412 271390
rect 152752 268394 152780 274722
rect 153304 270230 153332 277780
rect 154316 277766 154514 277794
rect 154316 271182 154344 277766
rect 155696 273698 155724 277780
rect 156604 275732 156656 275738
rect 156604 275674 156656 275680
rect 155684 273692 155736 273698
rect 155684 273634 155736 273640
rect 155960 272808 156012 272814
rect 155960 272750 156012 272756
rect 154304 271176 154356 271182
rect 154304 271118 154356 271124
rect 154028 270768 154080 270774
rect 154028 270710 154080 270716
rect 153292 270224 153344 270230
rect 153292 270166 153344 270172
rect 153844 269204 153896 269210
rect 153844 269146 153896 269152
rect 152740 268388 152792 268394
rect 152740 268330 152792 268336
rect 152384 267706 152688 267734
rect 152660 264330 152688 267706
rect 152660 264302 153042 264330
rect 153856 264316 153884 269146
rect 154040 266626 154068 270710
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 154672 267572 154724 267578
rect 154672 267514 154724 267520
rect 154028 266620 154080 266626
rect 154028 266562 154080 266568
rect 154684 264316 154712 267514
rect 155512 264316 155540 268466
rect 155972 264330 156000 272750
rect 156616 267306 156644 275674
rect 156892 275330 156920 277780
rect 158102 277766 158668 277794
rect 159298 277766 160048 277794
rect 156880 275324 156932 275330
rect 156880 275266 156932 275272
rect 157616 274236 157668 274242
rect 157616 274178 157668 274184
rect 156420 267300 156472 267306
rect 156420 267242 156472 267248
rect 156604 267300 156656 267306
rect 156604 267242 156656 267248
rect 156432 264602 156460 267242
rect 156604 266892 156656 266898
rect 156604 266834 156656 266840
rect 156616 266490 156644 266834
rect 156604 266484 156656 266490
rect 156604 266426 156656 266432
rect 156432 264574 156736 264602
rect 156708 264330 156736 264574
rect 157628 264330 157656 274178
rect 158640 270094 158668 277766
rect 158812 274372 158864 274378
rect 158812 274314 158864 274320
rect 158628 270088 158680 270094
rect 158628 270030 158680 270036
rect 155972 264302 156354 264330
rect 156708 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 274314
rect 160020 268530 160048 277766
rect 160480 275602 160508 277780
rect 160744 276004 160796 276010
rect 160744 275946 160796 275952
rect 160468 275596 160520 275602
rect 160468 275538 160520 275544
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 160008 268524 160060 268530
rect 160008 268466 160060 268472
rect 159640 267300 159692 267306
rect 159640 267242 159692 267248
rect 159652 264316 159680 267242
rect 160480 264316 160508 268602
rect 160756 267306 160784 275946
rect 161584 272678 161612 277780
rect 162124 272944 162176 272950
rect 162124 272886 162176 272892
rect 161572 272672 161624 272678
rect 161572 272614 161624 272620
rect 161294 269784 161350 269793
rect 161294 269719 161350 269728
rect 160744 267300 160796 267306
rect 160744 267242 160796 267248
rect 161308 264316 161336 269719
rect 162136 266626 162164 272886
rect 162780 271454 162808 277780
rect 163976 274786 164004 277780
rect 165186 277766 165568 277794
rect 165540 276026 165568 277766
rect 165540 275998 165660 276026
rect 166368 276010 166396 277780
rect 164148 275460 164200 275466
rect 164148 275402 164200 275408
rect 163964 274780 164016 274786
rect 163964 274722 164016 274728
rect 164160 271726 164188 275402
rect 164976 275188 165028 275194
rect 164976 275130 165028 275136
rect 163320 271720 163372 271726
rect 163320 271662 163372 271668
rect 164148 271720 164200 271726
rect 164148 271662 164200 271668
rect 162768 271448 162820 271454
rect 162768 271390 162820 271396
rect 161940 266620 161992 266626
rect 161940 266562 161992 266568
rect 162124 266620 162176 266626
rect 162124 266562 162176 266568
rect 162952 266620 163004 266626
rect 162952 266562 163004 266568
rect 161952 266354 161980 266562
rect 162124 266484 162176 266490
rect 162124 266426 162176 266432
rect 161940 266348 161992 266354
rect 161940 266290 161992 266296
rect 162136 264316 162164 266426
rect 162964 264316 162992 266562
rect 163332 264330 163360 271662
rect 164792 271584 164844 271590
rect 164792 271526 164844 271532
rect 164804 267734 164832 271526
rect 164988 267734 165016 275130
rect 165632 274242 165660 275998
rect 166356 276004 166408 276010
rect 166356 275946 166408 275952
rect 167564 275466 167592 277780
rect 167552 275460 167604 275466
rect 167552 275402 167604 275408
rect 167644 275052 167696 275058
rect 167644 274994 167696 275000
rect 166264 274916 166316 274922
rect 166264 274858 166316 274864
rect 165620 274236 165672 274242
rect 165620 274178 165672 274184
rect 166276 272270 166304 274858
rect 166080 272264 166132 272270
rect 166080 272206 166132 272212
rect 166264 272264 166316 272270
rect 166264 272206 166316 272212
rect 166092 270042 166120 272206
rect 166092 270014 166488 270042
rect 166264 268932 166316 268938
rect 166264 268874 166316 268880
rect 164804 267706 164924 267734
rect 164988 267706 165108 267734
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 163332 264302 163806 264330
rect 164620 264316 164648 267242
rect 164896 264466 164924 267706
rect 165080 266422 165108 267706
rect 165068 266416 165120 266422
rect 165068 266358 165120 266364
rect 164896 264438 165016 264466
rect 164988 264330 165016 264438
rect 164988 264302 165462 264330
rect 166276 264316 166304 268874
rect 166460 267306 166488 270014
rect 167656 267578 167684 274994
rect 168380 273080 168432 273086
rect 168380 273022 168432 273028
rect 167920 268796 167972 268802
rect 167920 268738 167972 268744
rect 167644 267572 167696 267578
rect 167644 267514 167696 267520
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 166448 267300 166500 267306
rect 166448 267242 166500 267248
rect 167104 264316 167132 267378
rect 167932 264316 167960 268738
rect 168392 264330 168420 273022
rect 168668 268666 168696 277780
rect 169878 277766 170076 277794
rect 170048 270230 170076 277766
rect 171060 275194 171088 277780
rect 171048 275188 171100 275194
rect 171048 275130 171100 275136
rect 172256 274786 172284 277780
rect 173466 277766 173848 277794
rect 172428 275596 172480 275602
rect 172428 275538 172480 275544
rect 170404 274780 170456 274786
rect 170404 274722 170456 274728
rect 172244 274780 172296 274786
rect 172244 274722 172296 274728
rect 169852 270224 169904 270230
rect 169852 270166 169904 270172
rect 170036 270224 170088 270230
rect 170036 270166 170088 270172
rect 168656 268660 168708 268666
rect 168656 268602 168708 268608
rect 169864 266898 169892 270166
rect 170416 267442 170444 274722
rect 171600 274508 171652 274514
rect 171600 274450 171652 274456
rect 171232 269068 171284 269074
rect 171232 269010 171284 269016
rect 170404 267436 170456 267442
rect 170404 267378 170456 267384
rect 169852 266892 169904 266898
rect 169852 266834 169904 266840
rect 170404 266552 170456 266558
rect 170404 266494 170456 266500
rect 169576 266416 169628 266422
rect 169576 266358 169628 266364
rect 168392 264302 168774 264330
rect 169588 264316 169616 266358
rect 170416 264316 170444 266494
rect 171244 264316 171272 269010
rect 171612 264330 171640 274450
rect 172440 268938 172468 275538
rect 173348 269680 173400 269686
rect 173348 269622 173400 269628
rect 172428 268932 172480 268938
rect 172428 268874 172480 268880
rect 172888 267300 172940 267306
rect 172888 267242 172940 267248
rect 171612 264302 172086 264330
rect 172900 264316 172928 267242
rect 173360 264330 173388 269622
rect 173820 268802 173848 277766
rect 174648 275738 174676 277780
rect 174636 275732 174688 275738
rect 174636 275674 174688 275680
rect 174912 274780 174964 274786
rect 174912 274722 174964 274728
rect 174924 269686 174952 274722
rect 175280 274644 175332 274650
rect 175280 274586 175332 274592
rect 174912 269680 174964 269686
rect 174912 269622 174964 269628
rect 173808 268796 173860 268802
rect 173808 268738 173860 268744
rect 174544 268252 174596 268258
rect 174544 268194 174596 268200
rect 173360 264302 173742 264330
rect 174556 264316 174584 268194
rect 175292 264330 175320 274586
rect 175844 270774 175872 277780
rect 176752 271856 176804 271862
rect 176752 271798 176804 271804
rect 175832 270768 175884 270774
rect 175832 270710 175884 270716
rect 176200 270496 176252 270502
rect 176200 270438 176252 270444
rect 175292 264302 175398 264330
rect 176212 264316 176240 270438
rect 176764 264330 176792 271798
rect 176948 270502 176976 277780
rect 178144 271590 178172 277780
rect 179340 274514 179368 277780
rect 179328 274508 179380 274514
rect 179328 274450 179380 274456
rect 180536 274378 180564 277780
rect 181732 275602 181760 277780
rect 182942 277766 183508 277794
rect 184138 277766 184520 277794
rect 182088 276004 182140 276010
rect 182088 275946 182140 275952
rect 181720 275596 181772 275602
rect 181720 275538 181772 275544
rect 180524 274372 180576 274378
rect 180524 274314 180576 274320
rect 181444 273828 181496 273834
rect 181444 273770 181496 273776
rect 181260 273216 181312 273222
rect 181260 273158 181312 273164
rect 179880 272400 179932 272406
rect 179880 272342 179932 272348
rect 178132 271584 178184 271590
rect 178132 271526 178184 271532
rect 177488 271040 177540 271046
rect 177488 270982 177540 270988
rect 176936 270496 176988 270502
rect 176936 270438 176988 270444
rect 177500 264330 177528 270982
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 179524 264316 179552 266698
rect 179892 264330 179920 272342
rect 180892 269408 180944 269414
rect 180892 269350 180944 269356
rect 180904 264330 180932 269350
rect 181272 267734 181300 273158
rect 181456 267734 181484 273770
rect 182100 273086 182128 275946
rect 182088 273080 182140 273086
rect 182088 273022 182140 273028
rect 183480 269550 183508 277766
rect 184492 271590 184520 277766
rect 184204 271584 184256 271590
rect 184204 271526 184256 271532
rect 184480 271584 184532 271590
rect 184480 271526 184532 271532
rect 183652 270360 183704 270366
rect 183652 270302 183704 270308
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 182180 268116 182232 268122
rect 182180 268058 182232 268064
rect 181272 267706 181392 267734
rect 181456 267706 181576 267734
rect 181364 264466 181392 267706
rect 181548 266422 181576 267706
rect 182192 266558 182220 268058
rect 182180 266552 182232 266558
rect 182180 266494 182232 266500
rect 181536 266416 181588 266422
rect 181536 266358 181588 266364
rect 182824 266416 182876 266422
rect 182824 266358 182876 266364
rect 181364 264438 181576 264466
rect 181548 264330 181576 264438
rect 179892 264302 180366 264330
rect 180904 264302 181194 264330
rect 181548 264302 182022 264330
rect 182836 264316 182864 266358
rect 183664 264316 183692 270302
rect 184216 266422 184244 271526
rect 184940 270904 184992 270910
rect 184940 270846 184992 270852
rect 184480 267708 184532 267714
rect 184480 267650 184532 267656
rect 184204 266416 184256 266422
rect 184204 266358 184256 266364
rect 184492 264316 184520 267650
rect 184952 264330 184980 270846
rect 185228 270366 185256 277780
rect 186424 277394 186452 277780
rect 186424 277366 186544 277394
rect 186516 270366 186544 277366
rect 187620 272814 187648 277780
rect 188816 276010 188844 277780
rect 188804 276004 188856 276010
rect 188804 275946 188856 275952
rect 187884 275868 187936 275874
rect 187884 275810 187936 275816
rect 187608 272808 187660 272814
rect 187608 272750 187660 272756
rect 187700 272536 187752 272542
rect 187700 272478 187752 272484
rect 185216 270360 185268 270366
rect 185216 270302 185268 270308
rect 186320 270360 186372 270366
rect 186320 270302 186372 270308
rect 186504 270360 186556 270366
rect 186504 270302 186556 270308
rect 186332 267442 186360 270302
rect 186964 267572 187016 267578
rect 186964 267514 187016 267520
rect 186320 267436 186372 267442
rect 186320 267378 186372 267384
rect 186136 266552 186188 266558
rect 186136 266494 186188 266500
rect 184952 264302 185334 264330
rect 186148 264316 186176 266494
rect 186976 264316 187004 267514
rect 187712 264330 187740 272478
rect 187896 271862 187924 275810
rect 190012 272950 190040 277780
rect 191222 277766 191788 277794
rect 191760 275890 191788 277766
rect 191760 275862 191880 275890
rect 191104 275188 191156 275194
rect 191104 275130 191156 275136
rect 190000 272944 190052 272950
rect 190000 272886 190052 272892
rect 189816 272128 189868 272134
rect 189816 272070 189868 272076
rect 187884 271856 187936 271862
rect 187884 271798 187936 271804
rect 189632 271312 189684 271318
rect 189632 271254 189684 271260
rect 188620 269816 188672 269822
rect 188620 269758 188672 269764
rect 187712 264302 187818 264330
rect 188632 264316 188660 269758
rect 189448 267028 189500 267034
rect 189448 266970 189500 266976
rect 189460 264316 189488 266970
rect 189644 264466 189672 271254
rect 189828 267714 189856 272070
rect 190828 269952 190880 269958
rect 190828 269894 190880 269900
rect 189816 267708 189868 267714
rect 189816 267650 189868 267656
rect 189644 264438 189856 264466
rect 189828 264330 189856 264438
rect 190840 264330 190868 269894
rect 191116 267034 191144 275130
rect 191852 273970 191880 275862
rect 191840 273964 191892 273970
rect 191840 273906 191892 273912
rect 191840 273828 191892 273834
rect 191840 273770 191892 273776
rect 191104 267028 191156 267034
rect 191104 266970 191156 266976
rect 191852 265674 191880 273770
rect 192312 272542 192340 277780
rect 193508 274106 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 195716 277766 195914 277794
rect 193312 274100 193364 274106
rect 193312 274042 193364 274048
rect 193496 274100 193548 274106
rect 193496 274042 193548 274048
rect 192300 272536 192352 272542
rect 192300 272478 192352 272484
rect 192024 272264 192076 272270
rect 192024 272206 192076 272212
rect 191840 265668 191892 265674
rect 191840 265610 191892 265616
rect 192036 265554 192064 272206
rect 192484 265668 192536 265674
rect 192484 265610 192536 265616
rect 191944 265526 192064 265554
rect 189828 264302 190302 264330
rect 190840 264302 191130 264330
rect 191944 264316 191972 265526
rect 192496 264330 192524 265610
rect 193324 264330 193352 274042
rect 194612 269822 194640 277366
rect 194784 271720 194836 271726
rect 194784 271662 194836 271668
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 192496 264302 192786 264330
rect 193324 264302 193614 264330
rect 194428 264316 194456 267106
rect 194796 264330 194824 271662
rect 195716 271318 195744 277766
rect 196440 271856 196492 271862
rect 196440 271798 196492 271804
rect 195704 271312 195756 271318
rect 195704 271254 195756 271260
rect 196072 268388 196124 268394
rect 196072 268330 196124 268336
rect 195244 267572 195296 267578
rect 195244 267514 195296 267520
rect 195256 266626 195284 267514
rect 195244 266620 195296 266626
rect 195244 266562 195296 266568
rect 194796 264302 195270 264330
rect 196084 264316 196112 268330
rect 196452 264330 196480 271798
rect 197096 271726 197124 277780
rect 198096 273692 198148 273698
rect 198096 273634 198148 273640
rect 197084 271720 197136 271726
rect 197084 271662 197136 271668
rect 197912 271176 197964 271182
rect 197912 271118 197964 271124
rect 197924 267734 197952 271118
rect 198108 267734 198136 273634
rect 198292 271182 198320 277780
rect 199292 275324 199344 275330
rect 199292 275266 199344 275272
rect 198280 271176 198332 271182
rect 198280 271118 198332 271124
rect 197728 267708 197780 267714
rect 197924 267706 198044 267734
rect 198108 267706 198228 267734
rect 197728 267650 197780 267656
rect 196452 264302 196926 264330
rect 197740 264316 197768 267650
rect 198016 264330 198044 267706
rect 198200 266898 198228 267706
rect 199304 267170 199332 275266
rect 199488 274854 199516 277780
rect 199476 274848 199528 274854
rect 199476 274790 199528 274796
rect 200396 268524 200448 268530
rect 200396 268466 200448 268472
rect 199292 267164 199344 267170
rect 199292 267106 199344 267112
rect 198188 266892 198240 266898
rect 198188 266834 198240 266840
rect 200212 266892 200264 266898
rect 200212 266834 200264 266840
rect 199384 266756 199436 266762
rect 199384 266698 199436 266704
rect 198016 264302 198582 264330
rect 199396 264316 199424 266698
rect 200224 264316 200252 266834
rect 200408 266422 200436 268466
rect 200592 268394 200620 277780
rect 201788 270094 201816 277780
rect 202998 277766 203288 277794
rect 202788 274848 202840 274854
rect 202788 274790 202840 274796
rect 202800 270366 202828 274790
rect 203260 272678 203288 277766
rect 203064 272672 203116 272678
rect 203064 272614 203116 272620
rect 203248 272672 203300 272678
rect 203248 272614 203300 272620
rect 202328 270360 202380 270366
rect 202328 270302 202380 270308
rect 202788 270360 202840 270366
rect 202788 270302 202840 270308
rect 201040 270088 201092 270094
rect 201040 270030 201092 270036
rect 201776 270088 201828 270094
rect 201776 270030 201828 270036
rect 200580 268388 200632 268394
rect 200580 268330 200632 268336
rect 200396 266416 200448 266422
rect 200396 266358 200448 266364
rect 201052 264316 201080 270030
rect 201868 267164 201920 267170
rect 201868 267106 201920 267112
rect 201880 264316 201908 267106
rect 202340 266898 202368 270302
rect 202328 266892 202380 266898
rect 202328 266834 202380 266840
rect 202696 266416 202748 266422
rect 202696 266358 202748 266364
rect 202708 264316 202736 266358
rect 203076 264330 203104 272614
rect 204180 269958 204208 277780
rect 204720 274644 204772 274650
rect 204720 274586 204772 274592
rect 204732 274106 204760 274586
rect 204720 274100 204772 274106
rect 204720 274042 204772 274048
rect 205376 271454 205404 277780
rect 205732 274236 205784 274242
rect 205732 274178 205784 274184
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 205364 271448 205416 271454
rect 205364 271390 205416 271396
rect 204168 269952 204220 269958
rect 204168 269894 204220 269900
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 204180 267714 204208 269486
rect 204352 268932 204404 268938
rect 204352 268874 204404 268880
rect 204168 267708 204220 267714
rect 204168 267650 204220 267656
rect 203076 264302 203550 264330
rect 204364 264316 204392 268874
rect 204732 264330 204760 271390
rect 205088 269952 205140 269958
rect 205088 269894 205140 269900
rect 205100 269550 205128 269894
rect 205088 269544 205140 269550
rect 205088 269486 205140 269492
rect 205744 264330 205772 274178
rect 206572 274106 206600 277780
rect 207782 277766 208256 277794
rect 206560 274100 206612 274106
rect 206560 274042 206612 274048
rect 207296 273080 207348 273086
rect 207296 273022 207348 273028
rect 206284 270768 206336 270774
rect 206284 270710 206336 270716
rect 205916 270360 205968 270366
rect 205916 270302 205968 270308
rect 205928 270094 205956 270302
rect 205916 270088 205968 270094
rect 205916 270030 205968 270036
rect 206296 267306 206324 270710
rect 206284 267300 206336 267306
rect 206284 267242 206336 267248
rect 206836 267164 206888 267170
rect 206836 267106 206888 267112
rect 207020 267164 207072 267170
rect 207020 267106 207072 267112
rect 204732 264302 205206 264330
rect 205744 264302 206034 264330
rect 206848 264316 206876 267106
rect 207032 266898 207060 267106
rect 207020 266892 207072 266898
rect 207020 266834 207072 266840
rect 207308 264330 207336 273022
rect 208228 268938 208256 277766
rect 208676 275732 208728 275738
rect 208676 275674 208728 275680
rect 208216 268932 208268 268938
rect 208216 268874 208268 268880
rect 208688 268666 208716 275674
rect 208872 274786 208900 277780
rect 209044 275460 209096 275466
rect 209044 275402 209096 275408
rect 208860 274780 208912 274786
rect 208860 274722 208912 274728
rect 208492 268660 208544 268666
rect 208492 268602 208544 268608
rect 208676 268660 208728 268666
rect 208676 268602 208728 268608
rect 207308 264302 207690 264330
rect 208504 264316 208532 268602
rect 209056 264330 209084 275402
rect 210068 274922 210096 277780
rect 211264 275330 211292 277780
rect 212460 275738 212488 277780
rect 212448 275732 212500 275738
rect 212448 275674 212500 275680
rect 211252 275324 211304 275330
rect 211252 275266 211304 275272
rect 210056 274916 210108 274922
rect 210056 274858 210108 274864
rect 212448 274916 212500 274922
rect 212448 274858 212500 274864
rect 210608 274780 210660 274786
rect 210608 274722 210660 274728
rect 210620 270230 210648 274722
rect 210148 270224 210200 270230
rect 210148 270166 210200 270172
rect 210608 270224 210660 270230
rect 210608 270166 210660 270172
rect 209056 264302 209346 264330
rect 210160 264316 210188 270166
rect 210976 269408 211028 269414
rect 210976 269350 211028 269356
rect 210988 264316 211016 269350
rect 212460 268530 212488 274858
rect 213184 274508 213236 274514
rect 213184 274450 213236 274456
rect 212632 268796 212684 268802
rect 212632 268738 212684 268744
rect 212448 268524 212500 268530
rect 212448 268466 212500 268472
rect 211804 267028 211856 267034
rect 211804 266970 211856 266976
rect 211816 264316 211844 266970
rect 212644 264316 212672 268738
rect 213196 266422 213224 274450
rect 213656 274242 213684 277780
rect 214866 277766 215248 277794
rect 215970 277766 216352 277794
rect 213644 274236 213696 274242
rect 213644 274178 213696 274184
rect 214748 270496 214800 270502
rect 214748 270438 214800 270444
rect 214288 268660 214340 268666
rect 214288 268602 214340 268608
rect 213460 267300 213512 267306
rect 213460 267242 213512 267248
rect 213184 266416 213236 266422
rect 213184 266358 213236 266364
rect 213472 264316 213500 267242
rect 214300 264316 214328 268602
rect 214760 264330 214788 270438
rect 215220 268802 215248 277766
rect 216324 271590 216352 277766
rect 216956 274372 217008 274378
rect 216956 274314 217008 274320
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 216312 271584 216364 271590
rect 216312 271526 216364 271532
rect 215208 268796 215260 268802
rect 215208 268738 215260 268744
rect 215956 267170 215984 271526
rect 216968 267734 216996 274314
rect 217152 272950 217180 277780
rect 218348 275466 218376 277780
rect 218612 275596 218664 275602
rect 218612 275538 218664 275544
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217416 273080 217468 273086
rect 217416 273022 217468 273028
rect 217140 272944 217192 272950
rect 217140 272886 217192 272892
rect 216968 267706 217272 267734
rect 216772 267572 216824 267578
rect 216772 267514 216824 267520
rect 215944 267164 215996 267170
rect 215944 267106 215996 267112
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 214760 264302 215142 264330
rect 215956 264316 215984 266358
rect 216784 264316 216812 267514
rect 217244 264330 217272 267706
rect 217428 267306 217456 273022
rect 218428 267708 218480 267714
rect 218428 267650 218480 267656
rect 217416 267300 217468 267306
rect 217416 267242 217468 267248
rect 217244 264302 217626 264330
rect 218440 264316 218468 267650
rect 218624 264330 218652 275538
rect 218796 274644 218848 274650
rect 218796 274586 218848 274592
rect 218808 267578 218836 274586
rect 219544 270366 219572 277780
rect 220544 275732 220596 275738
rect 220544 275674 220596 275680
rect 220556 272814 220584 275674
rect 220740 275670 220768 277780
rect 221936 277394 221964 277780
rect 221936 277366 222056 277394
rect 220728 275664 220780 275670
rect 220728 275606 220780 275612
rect 220084 272808 220136 272814
rect 220084 272750 220136 272756
rect 220544 272808 220596 272814
rect 220544 272750 220596 272756
rect 219532 270360 219584 270366
rect 219532 270302 219584 270308
rect 218796 267572 218848 267578
rect 218796 267514 218848 267520
rect 220096 267306 220124 272750
rect 220820 268796 220872 268802
rect 220820 268738 220872 268744
rect 219900 267300 219952 267306
rect 219900 267242 219952 267248
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 219912 266898 219940 267242
rect 220832 267170 220860 268738
rect 221740 267436 221792 267442
rect 221740 267378 221792 267384
rect 220084 267164 220136 267170
rect 220084 267106 220136 267112
rect 220820 267164 220872 267170
rect 220820 267106 220872 267112
rect 219900 266892 219952 266898
rect 219900 266834 219952 266840
rect 218624 264302 219282 264330
rect 220096 264316 220124 267106
rect 220912 267028 220964 267034
rect 220912 266970 220964 266976
rect 220924 264316 220952 266970
rect 221752 264316 221780 267378
rect 222028 267034 222056 277366
rect 222844 276004 222896 276010
rect 222844 275946 222896 275952
rect 222568 267300 222620 267306
rect 222568 267242 222620 267248
rect 222016 267028 222068 267034
rect 222016 266970 222068 266976
rect 222580 264316 222608 267242
rect 222856 266422 222884 275946
rect 223132 274378 223160 277780
rect 224250 277766 224632 277794
rect 223120 274372 223172 274378
rect 223120 274314 223172 274320
rect 224604 271726 224632 277766
rect 224960 275664 225012 275670
rect 224960 275606 225012 275612
rect 224972 273970 225000 275606
rect 225432 275602 225460 277780
rect 225420 275596 225472 275602
rect 225420 275538 225472 275544
rect 224960 273964 225012 273970
rect 224960 273906 225012 273912
rect 224960 273828 225012 273834
rect 224960 273770 225012 273776
rect 224224 271720 224276 271726
rect 224224 271662 224276 271668
rect 224592 271720 224644 271726
rect 224592 271662 224644 271668
rect 223488 269544 223540 269550
rect 223488 269486 223540 269492
rect 223500 267306 223528 269486
rect 224236 267714 224264 271662
rect 224224 267708 224276 267714
rect 224224 267650 224276 267656
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 223396 266892 223448 266898
rect 223396 266834 223448 266840
rect 222844 266416 222896 266422
rect 222844 266358 222896 266364
rect 223408 264316 223436 266834
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 224236 264316 224264 266358
rect 224972 264330 225000 273770
rect 225512 272536 225564 272542
rect 225512 272478 225564 272484
rect 225524 264330 225552 272478
rect 226628 269686 226656 277780
rect 227838 277766 228128 277794
rect 227904 271312 227956 271318
rect 227904 271254 227956 271260
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 226708 267572 226760 267578
rect 226708 267514 226760 267520
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226720 264316 226748 267514
rect 227272 264330 227300 269758
rect 227720 268932 227772 268938
rect 227720 268874 227772 268880
rect 227732 267442 227760 268874
rect 227720 267436 227772 267442
rect 227720 267378 227772 267384
rect 227916 264330 227944 271254
rect 228100 268666 228128 277766
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 228836 272542 228864 277766
rect 228824 272536 228876 272542
rect 228824 272478 228876 272484
rect 229560 271176 229612 271182
rect 229560 271118 229612 271124
rect 228088 268660 228140 268666
rect 228088 268602 228140 268608
rect 229192 267708 229244 267714
rect 229192 267650 229244 267656
rect 227272 264302 227562 264330
rect 227916 264302 228390 264330
rect 229204 264316 229232 267650
rect 229572 264330 229600 271118
rect 230400 270502 230428 277766
rect 231412 271182 231440 277780
rect 232516 275738 232544 277780
rect 232504 275732 232556 275738
rect 232504 275674 232556 275680
rect 232688 275324 232740 275330
rect 232688 275266 232740 275272
rect 231400 271176 231452 271182
rect 231400 271118 231452 271124
rect 230388 270496 230440 270502
rect 230388 270438 230440 270444
rect 230848 270088 230900 270094
rect 230848 270030 230900 270036
rect 229572 264302 230046 264330
rect 230860 264316 230888 270030
rect 232504 269952 232556 269958
rect 232504 269894 232556 269900
rect 231676 268388 231728 268394
rect 231676 268330 231728 268336
rect 231688 264316 231716 268330
rect 232516 264316 232544 269894
rect 232700 266762 232728 275266
rect 233240 272672 233292 272678
rect 233240 272614 233292 272620
rect 232688 266756 232740 266762
rect 232688 266698 232740 266704
rect 233252 264330 233280 272614
rect 233712 269958 233740 277780
rect 234908 277394 234936 277780
rect 234816 277366 234936 277394
rect 234620 274100 234672 274106
rect 234620 274042 234672 274048
rect 233700 269952 233752 269958
rect 233700 269894 233752 269900
rect 234160 267300 234212 267306
rect 234160 267242 234212 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267242
rect 234632 265674 234660 274042
rect 234816 268394 234844 277366
rect 234988 271448 235040 271454
rect 234988 271390 235040 271396
rect 234804 268388 234856 268394
rect 234804 268330 234856 268336
rect 234620 265668 234672 265674
rect 234620 265610 234672 265616
rect 235000 264316 235028 271390
rect 236104 269686 236132 277780
rect 237300 271318 237328 277780
rect 238496 272542 238524 277780
rect 239404 275460 239456 275466
rect 239404 275402 239456 275408
rect 239220 272808 239272 272814
rect 239220 272750 239272 272756
rect 238024 272536 238076 272542
rect 238024 272478 238076 272484
rect 238484 272536 238536 272542
rect 238484 272478 238536 272484
rect 237288 271312 237340 271318
rect 237288 271254 237340 271260
rect 237472 270224 237524 270230
rect 237472 270166 237524 270172
rect 236092 269680 236144 269686
rect 236092 269622 236144 269628
rect 236644 267436 236696 267442
rect 236644 267378 236696 267384
rect 235540 265668 235592 265674
rect 235540 265610 235592 265616
rect 235552 264330 235580 265610
rect 235552 264302 235842 264330
rect 236656 264316 236684 267378
rect 237484 264316 237512 270166
rect 238036 267306 238064 272478
rect 238300 268524 238352 268530
rect 238300 268466 238352 268472
rect 238024 267300 238076 267306
rect 238024 267242 238076 267248
rect 238312 264316 238340 268466
rect 239232 267734 239260 272750
rect 239416 267734 239444 275402
rect 239600 272678 239628 277780
rect 240810 277766 241376 277794
rect 240416 274236 240468 274242
rect 240416 274178 240468 274184
rect 239588 272672 239640 272678
rect 239588 272614 239640 272620
rect 239232 267706 239352 267734
rect 239416 267706 239536 267734
rect 239128 266756 239180 266762
rect 239128 266698 239180 266704
rect 239140 264316 239168 266698
rect 239324 264466 239352 267706
rect 239508 266422 239536 267706
rect 239496 266416 239548 266422
rect 239496 266358 239548 266364
rect 239324 264438 239536 264466
rect 239508 264330 239536 264438
rect 240428 264330 240456 274178
rect 241348 268530 241376 277766
rect 241992 274990 242020 277780
rect 242256 275596 242308 275602
rect 242256 275538 242308 275544
rect 241980 274984 242032 274990
rect 241980 274926 242032 274932
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241336 268524 241388 268530
rect 241336 268466 241388 268472
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 239508 264302 239982 264330
rect 240428 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271526
rect 242268 266898 242296 275538
rect 243188 274854 243216 277780
rect 244384 275738 244412 277780
rect 245580 277394 245608 277780
rect 245488 277366 245608 277394
rect 244372 275732 244424 275738
rect 244372 275674 244424 275680
rect 244096 274984 244148 274990
rect 244096 274926 244148 274932
rect 243176 274848 243228 274854
rect 243176 274790 243228 274796
rect 242900 272944 242952 272950
rect 242900 272886 242952 272892
rect 242256 266892 242308 266898
rect 242256 266834 242308 266840
rect 242912 264330 242940 272886
rect 244108 270094 244136 274926
rect 244924 270360 244976 270366
rect 244924 270302 244976 270308
rect 244096 270088 244148 270094
rect 244096 270030 244148 270036
rect 243912 269952 243964 269958
rect 243912 269894 243964 269900
rect 243924 267170 243952 269894
rect 243912 267164 243964 267170
rect 243912 267106 243964 267112
rect 244096 266416 244148 266422
rect 244096 266358 244148 266364
rect 242084 264302 242466 264330
rect 242912 264302 243294 264330
rect 244108 264316 244136 266358
rect 244936 264316 244964 270302
rect 245488 269958 245516 277366
rect 245660 275596 245712 275602
rect 245660 275538 245712 275544
rect 245672 274106 245700 275538
rect 246776 275126 246804 277780
rect 247894 277766 248368 277794
rect 247040 275732 247092 275738
rect 247040 275674 247092 275680
rect 246764 275120 246816 275126
rect 246764 275062 246816 275068
rect 245660 274100 245712 274106
rect 245660 274042 245712 274048
rect 247052 273970 247080 275674
rect 248340 274666 248368 277766
rect 249076 275262 249104 277780
rect 249064 275256 249116 275262
rect 249064 275198 249116 275204
rect 249064 274848 249116 274854
rect 249064 274790 249116 274796
rect 248340 274638 248460 274666
rect 247224 274372 247276 274378
rect 247224 274314 247276 274320
rect 245752 273964 245804 273970
rect 245752 273906 245804 273912
rect 247040 273964 247092 273970
rect 247040 273906 247092 273912
rect 245476 269952 245528 269958
rect 245476 269894 245528 269900
rect 245764 264316 245792 273906
rect 246580 267028 246632 267034
rect 246580 266970 246632 266976
rect 246592 264316 246620 266970
rect 247236 264330 247264 274314
rect 247776 271720 247828 271726
rect 247776 271662 247828 271668
rect 247788 264330 247816 271662
rect 248432 271454 248460 274638
rect 248420 271448 248472 271454
rect 248420 271390 248472 271396
rect 249076 267034 249104 274790
rect 250272 269822 250300 277780
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 250260 269816 250312 269822
rect 250260 269758 250312 269764
rect 249064 267028 249116 267034
rect 249064 266970 249116 266976
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 247236 264302 247434 264330
rect 247788 264302 248262 264330
rect 249076 264316 249104 266834
rect 249904 264316 249932 269758
rect 251468 269278 251496 277780
rect 252664 272678 252692 277780
rect 253860 275466 253888 277780
rect 255070 277766 255268 277794
rect 256174 277766 256556 277794
rect 253848 275460 253900 275466
rect 253848 275402 253900 275408
rect 253572 275256 253624 275262
rect 253572 275198 253624 275204
rect 251824 272672 251876 272678
rect 251824 272614 251876 272620
rect 252652 272672 252704 272678
rect 252652 272614 252704 272620
rect 251456 269272 251508 269278
rect 251456 269214 251508 269220
rect 250720 268660 250772 268666
rect 250720 268602 250772 268608
rect 250732 264316 250760 268602
rect 251548 267300 251600 267306
rect 251548 267242 251600 267248
rect 251560 264316 251588 267242
rect 251836 266898 251864 272614
rect 253584 271182 253612 275198
rect 254032 274100 254084 274106
rect 254032 274042 254084 274048
rect 252744 271176 252796 271182
rect 252744 271118 252796 271124
rect 253572 271176 253624 271182
rect 253572 271118 253624 271124
rect 252100 270496 252152 270502
rect 252100 270438 252152 270444
rect 251824 266892 251876 266898
rect 251824 266834 251876 266840
rect 252112 264330 252140 270438
rect 252756 264330 252784 271118
rect 253756 269680 253808 269686
rect 253756 269622 253808 269628
rect 253768 266422 253796 269622
rect 253756 266416 253808 266422
rect 253756 266358 253808 266364
rect 252112 264302 252402 264330
rect 252756 264302 253230 264330
rect 254044 264316 254072 274042
rect 255240 270230 255268 277766
rect 255228 270224 255280 270230
rect 255228 270166 255280 270172
rect 256528 268394 256556 277766
rect 256700 275120 256752 275126
rect 256700 275062 256752 275068
rect 256712 268666 256740 275062
rect 257356 274718 257384 277780
rect 257344 274712 257396 274718
rect 257344 274654 257396 274660
rect 258080 272536 258132 272542
rect 258080 272478 258132 272484
rect 256976 271312 257028 271318
rect 256976 271254 257028 271260
rect 256700 268660 256752 268666
rect 256700 268602 256752 268608
rect 256700 268524 256752 268530
rect 256700 268466 256752 268472
rect 255688 268388 255740 268394
rect 255688 268330 255740 268336
rect 256516 268388 256568 268394
rect 256516 268330 256568 268336
rect 254860 267164 254912 267170
rect 254860 267106 254912 267112
rect 254872 264316 254900 267106
rect 255700 264316 255728 268330
rect 256712 266422 256740 268466
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 256700 266416 256752 266422
rect 256700 266358 256752 266364
rect 256528 264316 256556 266358
rect 256988 264330 257016 271254
rect 258092 264330 258120 272478
rect 258552 272406 258580 277780
rect 259748 275330 259776 277780
rect 260944 275806 260972 277780
rect 262140 277394 262168 277780
rect 262048 277366 262168 277394
rect 260932 275800 260984 275806
rect 260932 275742 260984 275748
rect 261484 275460 261536 275466
rect 261484 275402 261536 275408
rect 259736 275324 259788 275330
rect 259736 275266 259788 275272
rect 260196 274712 260248 274718
rect 260196 274654 260248 274660
rect 258540 272400 258592 272406
rect 258540 272342 258592 272348
rect 260208 271318 260236 274654
rect 260196 271312 260248 271318
rect 260196 271254 260248 271260
rect 260656 270088 260708 270094
rect 260656 270030 260708 270036
rect 258264 269272 258316 269278
rect 258264 269214 258316 269220
rect 258276 266558 258304 269214
rect 259000 266892 259052 266898
rect 259000 266834 259052 266840
rect 258264 266552 258316 266558
rect 258264 266494 258316 266500
rect 256988 264302 257370 264330
rect 258092 264302 258198 264330
rect 259012 264316 259040 266834
rect 259828 266416 259880 266422
rect 259828 266358 259880 266364
rect 259840 264316 259868 266358
rect 260668 264316 260696 270030
rect 261496 267306 261524 275402
rect 262048 270094 262076 277366
rect 263244 274854 263272 277780
rect 264454 277766 264836 277794
rect 265650 277766 266308 277794
rect 263508 275800 263560 275806
rect 263508 275742 263560 275748
rect 263232 274848 263284 274854
rect 263232 274790 263284 274796
rect 263520 273970 263548 275742
rect 262220 273964 262272 273970
rect 262220 273906 262272 273912
rect 263508 273964 263560 273970
rect 263508 273906 263560 273912
rect 262036 270088 262088 270094
rect 262036 270030 262088 270036
rect 261484 267300 261536 267306
rect 261484 267242 261536 267248
rect 261484 267028 261536 267034
rect 261484 266970 261536 266976
rect 261496 264316 261524 266970
rect 262232 264330 262260 273906
rect 264336 271448 264388 271454
rect 264336 271390 264388 271396
rect 263140 269952 263192 269958
rect 263140 269894 263192 269900
rect 262232 264302 262338 264330
rect 263152 264316 263180 269894
rect 263968 268660 264020 268666
rect 263968 268602 264020 268608
rect 263980 264316 264008 268602
rect 264348 264330 264376 271390
rect 264808 267734 264836 277766
rect 265256 271176 265308 271182
rect 265256 271118 265308 271124
rect 264808 267706 265020 267734
rect 264992 266898 265020 267706
rect 264980 266892 265032 266898
rect 264980 266834 265032 266840
rect 265268 264330 265296 271118
rect 266280 269958 266308 277766
rect 266452 274848 266504 274854
rect 266452 274790 266504 274796
rect 266268 269952 266320 269958
rect 266268 269894 266320 269900
rect 266464 268530 266492 274790
rect 266832 269822 266860 277780
rect 268028 275738 268056 277780
rect 269238 277766 269528 277794
rect 268016 275732 268068 275738
rect 268016 275674 268068 275680
rect 269120 275732 269172 275738
rect 269120 275674 269172 275680
rect 268844 275324 268896 275330
rect 268844 275266 268896 275272
rect 268856 273222 268884 275266
rect 269132 274106 269160 275674
rect 269120 274100 269172 274106
rect 269120 274042 269172 274048
rect 268844 273216 268896 273222
rect 268844 273158 268896 273164
rect 267832 272536 267884 272542
rect 267832 272478 267884 272484
rect 266636 269816 266688 269822
rect 266636 269758 266688 269764
rect 266820 269816 266872 269822
rect 266820 269758 266872 269764
rect 266452 268524 266504 268530
rect 266452 268466 266504 268472
rect 266648 264330 266676 269758
rect 267280 266552 267332 266558
rect 267280 266494 267332 266500
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266478 264302 266676 264330
rect 267292 264316 267320 266494
rect 267844 264330 267872 272478
rect 269500 271182 269528 277766
rect 270420 275126 270448 277780
rect 270408 275120 270460 275126
rect 270408 275062 270460 275068
rect 269764 272400 269816 272406
rect 269764 272342 269816 272348
rect 269488 271176 269540 271182
rect 269488 271118 269540 271124
rect 269396 270224 269448 270230
rect 269396 270166 269448 270172
rect 268936 267300 268988 267306
rect 268936 267242 268988 267248
rect 267844 264302 268134 264330
rect 268948 264316 268976 267242
rect 269408 264330 269436 270166
rect 269776 266422 269804 272342
rect 271524 271318 271552 277780
rect 272734 277766 273116 277794
rect 272616 273216 272668 273222
rect 272616 273158 272668 273164
rect 270960 271312 271012 271318
rect 270960 271254 271012 271260
rect 271512 271312 271564 271318
rect 271512 271254 271564 271260
rect 270592 268388 270644 268394
rect 270592 268330 270644 268336
rect 269764 266416 269816 266422
rect 269764 266358 269816 266364
rect 269408 264302 269790 264330
rect 270604 264316 270632 268330
rect 270972 264330 271000 271254
rect 272248 266416 272300 266422
rect 272248 266358 272300 266364
rect 270972 264302 271446 264330
rect 272260 264316 272288 266358
rect 272628 264330 272656 273158
rect 272892 269952 272944 269958
rect 272892 269894 272944 269900
rect 272904 266422 272932 269894
rect 273088 269414 273116 277766
rect 273536 273964 273588 273970
rect 273536 273906 273588 273912
rect 273076 269408 273128 269414
rect 273076 269350 273128 269356
rect 272892 266416 272944 266422
rect 272892 266358 272944 266364
rect 273548 264330 273576 273906
rect 273916 272542 273944 277780
rect 273904 272536 273956 272542
rect 273904 272478 273956 272484
rect 275112 270502 275140 277780
rect 276308 275330 276336 277780
rect 276296 275324 276348 275330
rect 276296 275266 276348 275272
rect 276204 275120 276256 275126
rect 276204 275062 276256 275068
rect 275100 270496 275152 270502
rect 275100 270438 275152 270444
rect 276020 270496 276072 270502
rect 276020 270438 276072 270444
rect 274732 270088 274784 270094
rect 274732 270030 274784 270036
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274744 264316 274772 270030
rect 275560 268524 275612 268530
rect 275560 268466 275612 268472
rect 275572 264316 275600 268466
rect 276032 267034 276060 270438
rect 276216 268394 276244 275062
rect 277504 274854 277532 277780
rect 278700 277394 278728 277780
rect 278608 277366 278728 277394
rect 277492 274848 277544 274854
rect 277492 274790 277544 274796
rect 278608 270366 278636 277366
rect 278780 274100 278832 274106
rect 278780 274042 278832 274048
rect 278596 270360 278648 270366
rect 278596 270302 278648 270308
rect 278044 269816 278096 269822
rect 278044 269758 278096 269764
rect 277400 269408 277452 269414
rect 277400 269350 277452 269356
rect 276204 268388 276256 268394
rect 276204 268330 276256 268336
rect 276020 267028 276072 267034
rect 276020 266970 276072 266976
rect 276388 266892 276440 266898
rect 276388 266834 276440 266840
rect 276400 264316 276428 266834
rect 277412 266422 277440 269350
rect 277216 266416 277268 266422
rect 277216 266358 277268 266364
rect 277400 266416 277452 266422
rect 277400 266358 277452 266364
rect 277228 264316 277256 266358
rect 278056 264316 278084 269758
rect 278792 264330 278820 274042
rect 279804 273970 279832 277780
rect 281014 277766 281488 277794
rect 282210 277766 282868 277794
rect 279792 273964 279844 273970
rect 279792 273906 279844 273912
rect 280896 271312 280948 271318
rect 280896 271254 280948 271260
rect 279240 271176 279292 271182
rect 279240 271118 279292 271124
rect 279252 264330 279280 271118
rect 280528 268388 280580 268394
rect 280528 268330 280580 268336
rect 278792 264302 278898 264330
rect 279252 264302 279726 264330
rect 280540 264316 280568 268330
rect 280908 264330 280936 271254
rect 281460 270502 281488 277766
rect 281448 270496 281500 270502
rect 281448 270438 281500 270444
rect 282840 267170 282868 277766
rect 283196 274848 283248 274854
rect 283196 274790 283248 274796
rect 283012 272536 283064 272542
rect 283012 272478 283064 272484
rect 282828 267164 282880 267170
rect 282828 267106 282880 267112
rect 282184 266416 282236 266422
rect 282184 266358 282236 266364
rect 280908 264302 281382 264330
rect 282196 264316 282224 266358
rect 283024 264316 283052 272478
rect 283208 271862 283236 274790
rect 283392 274718 283420 277780
rect 284588 275330 284616 277780
rect 284300 275324 284352 275330
rect 284300 275266 284352 275272
rect 284576 275324 284628 275330
rect 284576 275266 284628 275272
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283196 271856 283248 271862
rect 283196 271798 283248 271804
rect 283840 267028 283892 267034
rect 283840 266970 283892 266976
rect 283852 264316 283880 266970
rect 284312 264330 284340 275266
rect 285128 271856 285180 271862
rect 285128 271798 285180 271804
rect 285140 264330 285168 271798
rect 285784 271182 285812 277780
rect 286888 277394 286916 277780
rect 288098 277766 288296 277794
rect 286888 277366 287008 277394
rect 285772 271176 285824 271182
rect 285772 271118 285824 271124
rect 285680 270496 285732 270502
rect 285680 270438 285732 270444
rect 285692 266898 285720 270438
rect 286324 270360 286376 270366
rect 286324 270302 286376 270308
rect 285680 266892 285732 266898
rect 285680 266834 285732 266840
rect 284312 264302 284694 264330
rect 285140 264302 285522 264330
rect 286336 264316 286364 270302
rect 286980 269958 287008 277366
rect 287152 273964 287204 273970
rect 287152 273906 287204 273912
rect 286968 269952 287020 269958
rect 286968 269894 287020 269900
rect 287164 264316 287192 273906
rect 288268 270230 288296 277766
rect 289280 274854 289308 277780
rect 290096 275324 290148 275330
rect 290096 275266 290148 275272
rect 289268 274848 289320 274854
rect 289268 274790 289320 274796
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 288256 270224 288308 270230
rect 288256 270166 288308 270172
rect 288808 267164 288860 267170
rect 288808 267106 288860 267112
rect 287980 266892 288032 266898
rect 287980 266834 288032 266840
rect 287992 264316 288020 266834
rect 288820 264316 288848 267106
rect 289188 264330 289216 274654
rect 290108 264330 290136 275266
rect 290476 274718 290504 277780
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 291200 271176 291252 271182
rect 291200 271118 291252 271124
rect 291212 264330 291240 271118
rect 291672 270366 291700 277780
rect 292868 270502 292896 277780
rect 294064 277394 294092 277780
rect 294064 277366 294184 277394
rect 293408 274848 293460 274854
rect 293408 274790 293460 274796
rect 292856 270496 292908 270502
rect 292856 270438 292908 270444
rect 291660 270360 291712 270366
rect 291660 270302 291712 270308
rect 292948 270224 293000 270230
rect 292948 270166 293000 270172
rect 292120 269952 292172 269958
rect 292120 269894 292172 269900
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291212 264302 291318 264330
rect 292132 264316 292160 269894
rect 292960 264316 292988 270166
rect 293420 264330 293448 274790
rect 293960 270496 294012 270502
rect 293960 270438 294012 270444
rect 293972 266422 294000 270438
rect 294156 269142 294184 277366
rect 294328 274712 294380 274718
rect 294328 274654 294380 274660
rect 295168 274666 295196 277780
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 294144 269136 294196 269142
rect 294144 269078 294196 269084
rect 293960 266416 294012 266422
rect 293960 266358 294012 266364
rect 294340 264330 294368 274654
rect 295168 274638 295380 274666
rect 296352 274654 296404 274660
rect 295352 269278 295380 274638
rect 297928 270502 297956 277766
rect 298756 274718 298784 277780
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298744 274712 298796 274718
rect 298744 274654 298796 274660
rect 297916 270496 297968 270502
rect 297916 270438 297968 270444
rect 295524 270360 295576 270366
rect 295524 270302 295576 270308
rect 295340 269272 295392 269278
rect 295340 269214 295392 269220
rect 295536 267734 295564 270302
rect 297916 269272 297968 269278
rect 297916 269214 297968 269220
rect 297088 269136 297140 269142
rect 297088 269078 297140 269084
rect 295444 267706 295564 267734
rect 293420 264302 293802 264330
rect 294340 264302 294630 264330
rect 295444 264316 295472 267706
rect 296260 266416 296312 266422
rect 296260 266358 296312 266364
rect 296272 264316 296300 266358
rect 297100 264316 297128 269078
rect 297928 264316 297956 269214
rect 298388 264330 298416 274654
rect 299952 270502 299980 277780
rect 301148 277394 301176 277780
rect 301056 277366 301176 277394
rect 302344 277394 302372 277780
rect 302344 277366 302464 277394
rect 300124 274712 300176 274718
rect 300124 274654 300176 274660
rect 299572 270496 299624 270502
rect 299572 270438 299624 270444
rect 299940 270496 299992 270502
rect 299940 270438 299992 270444
rect 298388 264302 298770 264330
rect 299584 264316 299612 270438
rect 300136 264330 300164 274654
rect 300860 270496 300912 270502
rect 300860 270438 300912 270444
rect 300872 264330 300900 270438
rect 301056 266422 301084 277366
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300136 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303448 270450 303476 277780
rect 304092 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 303448 270422 303660 270450
rect 303632 264330 303660 270422
rect 304092 264330 304120 277766
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 266892 312872 266898
rect 312820 266834 312872 266840
rect 312360 266688 312412 266694
rect 312360 266630 312412 266636
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312372 264330 312400 266630
rect 312018 264302 312400 264330
rect 312832 264316 312860 266834
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313648 266484 313700 266490
rect 313648 266426 313700 266432
rect 313660 264316 313688 266426
rect 314488 264316 314516 269758
rect 314672 266694 314700 277766
rect 316512 277394 316540 277780
rect 316420 277366 316540 277394
rect 317432 277766 317722 277794
rect 318826 277766 319024 277794
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266688 314712 266694
rect 314660 266630 314712 266636
rect 315776 264330 315804 271254
rect 316420 266898 316448 277366
rect 316960 270088 317012 270094
rect 316960 270030 317012 270036
rect 316408 266892 316460 266898
rect 316408 266834 316460 266840
rect 316132 266620 316184 266626
rect 316132 266562 316184 266568
rect 315330 264302 315804 264330
rect 316144 264316 316172 266562
rect 316972 264316 317000 270030
rect 317432 266490 317460 277766
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317788 266756 317840 266762
rect 317788 266698 317840 266704
rect 317420 266484 317472 266490
rect 317420 266426 317472 266432
rect 317800 264316 317828 266698
rect 318628 264316 318656 271730
rect 318996 269822 319024 277766
rect 320008 271318 320036 277780
rect 320560 277766 321218 277794
rect 321572 277766 322414 277794
rect 322952 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318984 269816 319036 269822
rect 318984 269758 319036 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320560 266626 320588 277766
rect 321100 270224 321152 270230
rect 321100 270166 321152 270172
rect 320548 266620 320600 266626
rect 320548 266562 320600 266568
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 270166
rect 321572 270094 321600 277766
rect 322756 272536 322808 272542
rect 322756 272478 322808 272484
rect 321560 270088 321612 270094
rect 321560 270030 321612 270036
rect 321928 266892 321980 266898
rect 321928 266834 321980 266840
rect 321940 264316 321968 266834
rect 322768 264316 322796 272478
rect 322952 266762 322980 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 324964 274712 325016 274718
rect 324964 274654 325016 274660
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 323584 269952 323636 269958
rect 323584 269894 323636 269900
rect 322940 266756 322992 266762
rect 322940 266698 322992 266704
rect 323596 264316 323624 269894
rect 324412 267164 324464 267170
rect 324412 267106 324464 267112
rect 324424 264316 324452 267106
rect 324976 266422 325004 274654
rect 325516 271312 325568 271318
rect 325516 271254 325568 271260
rect 324964 266416 325016 266422
rect 324964 266358 325016 266364
rect 325528 264330 325556 271254
rect 325712 269142 325740 277766
rect 327092 274718 327120 277780
rect 327460 277766 328302 277794
rect 328472 277766 329498 277794
rect 327080 274712 327132 274718
rect 327080 274654 327132 274660
rect 327080 270496 327132 270502
rect 327080 270438 327132 270444
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326068 268524 326120 268530
rect 326068 268466 326120 268472
rect 325266 264302 325556 264330
rect 326080 264316 326108 268466
rect 326908 264316 326936 269758
rect 327092 266898 327120 270438
rect 327460 270230 327488 277766
rect 328092 271176 328144 271182
rect 328092 271118 328144 271124
rect 327448 270224 327500 270230
rect 327448 270166 327500 270172
rect 327080 266892 327132 266898
rect 327080 266834 327132 266840
rect 328104 264330 328132 271118
rect 328472 270502 328500 277766
rect 330484 273284 330536 273290
rect 330484 273226 330536 273232
rect 328460 270496 328512 270502
rect 328460 270438 328512 270444
rect 329380 270224 329432 270230
rect 329380 270166 329432 270172
rect 328552 267776 328604 267782
rect 328552 267718 328604 267724
rect 327750 264302 328132 264330
rect 328564 264316 328592 267718
rect 329392 264316 329420 270166
rect 330496 267170 330524 273226
rect 330680 272542 330708 277780
rect 331232 277766 331890 277794
rect 330668 272536 330720 272542
rect 330668 272478 330720 272484
rect 331036 272536 331088 272542
rect 331036 272478 331088 272484
rect 330484 267164 330536 267170
rect 330484 267106 330536 267112
rect 330208 266552 330260 266558
rect 330208 266494 330260 266500
rect 330220 264316 330248 266494
rect 331048 264316 331076 272478
rect 331232 269958 331260 277766
rect 331404 274712 331456 274718
rect 331404 274654 331456 274660
rect 331220 269952 331272 269958
rect 331220 269894 331272 269900
rect 331416 268530 331444 274654
rect 333072 273290 333100 277780
rect 333796 273964 333848 273970
rect 333796 273906 333848 273912
rect 333060 273284 333112 273290
rect 333060 273226 333112 273232
rect 332232 270088 332284 270094
rect 332232 270030 332284 270036
rect 331404 268524 331456 268530
rect 331404 268466 331456 268472
rect 332244 264330 332272 270030
rect 333520 267164 333572 267170
rect 333520 267106 333572 267112
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 331890 264302 332272 264330
rect 332704 264316 332732 266358
rect 333532 264316 333560 267106
rect 333808 266422 333836 273906
rect 334176 271318 334204 277780
rect 335372 274718 335400 277780
rect 335556 277766 336582 277794
rect 335360 274712 335412 274718
rect 335360 274654 335412 274660
rect 334164 271312 334216 271318
rect 334164 271254 334216 271260
rect 334624 271312 334676 271318
rect 334624 271254 334676 271260
rect 334348 267300 334400 267306
rect 334348 267242 334400 267248
rect 333796 266416 333848 266422
rect 333796 266358 333848 266364
rect 334360 264316 334388 267242
rect 334636 266558 334664 271254
rect 335556 269822 335584 277766
rect 336648 274848 336700 274854
rect 336648 274790 336700 274796
rect 336660 270094 336688 274790
rect 337108 274712 337160 274718
rect 337108 274654 337160 274660
rect 336648 270088 336700 270094
rect 336648 270030 336700 270036
rect 336004 269952 336056 269958
rect 336004 269894 336056 269900
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 335176 268524 335228 268530
rect 335176 268466 335228 268472
rect 334624 266552 334676 266558
rect 334624 266494 334676 266500
rect 335188 264316 335216 268466
rect 336016 264316 336044 269894
rect 336832 269816 336884 269822
rect 336832 269758 336884 269764
rect 336844 264316 336872 269758
rect 337120 267782 337148 274654
rect 337764 271182 337792 277780
rect 338960 274718 338988 277780
rect 339512 277766 340170 277794
rect 339132 275324 339184 275330
rect 339132 275266 339184 275272
rect 338948 274712 339000 274718
rect 338948 274654 339000 274660
rect 337752 271176 337804 271182
rect 337752 271118 337804 271124
rect 337660 268388 337712 268394
rect 337660 268330 337712 268336
rect 337108 267776 337160 267782
rect 337108 267718 337160 267724
rect 337672 264316 337700 268330
rect 339144 267734 339172 275266
rect 339316 271176 339368 271182
rect 339316 271118 339368 271124
rect 338960 267706 339172 267734
rect 338960 264330 338988 267706
rect 338514 264302 338988 264330
rect 339328 264316 339356 271118
rect 339512 270230 339540 277766
rect 340604 271584 340656 271590
rect 340604 271526 340656 271532
rect 339500 270224 339552 270230
rect 339500 270166 339552 270172
rect 340616 264330 340644 271526
rect 341352 271318 341380 277780
rect 342456 272542 342484 277780
rect 343652 274854 343680 277780
rect 344480 277766 344862 277794
rect 345124 277766 346058 277794
rect 343640 274848 343692 274854
rect 343640 274790 343692 274796
rect 344284 274712 344336 274718
rect 344284 274654 344336 274660
rect 343548 272808 343600 272814
rect 343548 272750 343600 272756
rect 342444 272536 342496 272542
rect 342444 272478 342496 272484
rect 341340 271312 341392 271318
rect 341340 271254 341392 271260
rect 341800 269680 341852 269686
rect 341800 269622 341852 269628
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341812 264316 341840 269622
rect 342260 269136 342312 269142
rect 342260 269078 342312 269084
rect 342272 267170 342300 269078
rect 342260 267164 342312 267170
rect 342260 267106 342312 267112
rect 343364 267028 343416 267034
rect 343364 266970 343416 266976
rect 342628 266416 342680 266422
rect 342628 266358 342680 266364
rect 342640 264316 342668 266358
rect 343376 264330 343404 266970
rect 343560 266422 343588 272750
rect 344296 267306 344324 274654
rect 344480 273970 344508 277766
rect 344468 273964 344520 273970
rect 344468 273906 344520 273912
rect 344652 273964 344704 273970
rect 344652 273906 344704 273912
rect 344284 267300 344336 267306
rect 344284 267242 344336 267248
rect 343548 266416 343600 266422
rect 343548 266358 343600 266364
rect 344664 264330 344692 273906
rect 345124 269142 345152 277766
rect 347240 274718 347268 277780
rect 347792 277766 348450 277794
rect 347412 275596 347464 275602
rect 347412 275538 347464 275544
rect 347228 274712 347280 274718
rect 347228 274654 347280 274660
rect 345940 270224 345992 270230
rect 345940 270166 345992 270172
rect 345112 269136 345164 269142
rect 345112 269078 345164 269084
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 343376 264302 343482 264330
rect 344310 264302 344692 264330
rect 345124 264316 345152 266358
rect 345952 264316 345980 270166
rect 347424 270094 347452 275538
rect 347596 272672 347648 272678
rect 347596 272614 347648 272620
rect 347412 270088 347464 270094
rect 347412 270030 347464 270036
rect 346768 269952 346820 269958
rect 346768 269894 346820 269900
rect 346780 264316 346808 269894
rect 347608 264316 347636 272614
rect 347792 268530 347820 277766
rect 349632 275602 349660 277780
rect 350552 277766 350750 277794
rect 349620 275596 349672 275602
rect 349620 275538 349672 275544
rect 349712 275460 349764 275466
rect 349712 275402 349764 275408
rect 349724 273970 349752 275402
rect 349896 274100 349948 274106
rect 349896 274042 349948 274048
rect 349712 273964 349764 273970
rect 349712 273906 349764 273912
rect 348884 271448 348936 271454
rect 348884 271390 348936 271396
rect 347780 268524 347832 268530
rect 347780 268466 347832 268472
rect 348896 264330 348924 271390
rect 349712 270088 349764 270094
rect 349712 270030 349764 270036
rect 349724 269686 349752 270030
rect 349712 269680 349764 269686
rect 349712 269622 349764 269628
rect 349252 266892 349304 266898
rect 349252 266834 349304 266840
rect 348450 264302 348924 264330
rect 349264 264316 349292 266834
rect 349908 266422 349936 274042
rect 350356 273828 350408 273834
rect 350356 273770 350408 273776
rect 349896 266416 349948 266422
rect 349896 266358 349948 266364
rect 350368 264330 350396 273770
rect 350552 269822 350580 277766
rect 350540 269816 350592 269822
rect 350540 269758 350592 269764
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 350908 267164 350960 267170
rect 350908 267106 350960 267112
rect 350106 264302 350396 264330
rect 350920 264316 350948 267106
rect 351748 264316 351776 269758
rect 351932 268394 351960 277780
rect 352380 275596 352432 275602
rect 352380 275538 352432 275544
rect 351920 268388 351972 268394
rect 351920 268330 351972 268336
rect 352392 267034 352420 275538
rect 353128 275330 353156 277780
rect 353116 275324 353168 275330
rect 353116 275266 353168 275272
rect 354324 271182 354352 277780
rect 355152 277766 355534 277794
rect 356072 277766 356730 277794
rect 357452 277766 357926 277794
rect 355152 271590 355180 277766
rect 355140 271584 355192 271590
rect 355140 271526 355192 271532
rect 355324 271584 355376 271590
rect 355324 271526 355376 271532
rect 354588 271312 354640 271318
rect 354588 271254 354640 271260
rect 354312 271176 354364 271182
rect 354312 271118 354364 271124
rect 352564 268388 352616 268394
rect 352564 268330 352616 268336
rect 352380 267028 352432 267034
rect 352380 266970 352432 266976
rect 352576 264316 352604 268330
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 353404 264316 353432 266970
rect 354600 264330 354628 271254
rect 355336 266898 355364 271526
rect 355876 268660 355928 268666
rect 355876 268602 355928 268608
rect 355324 266892 355376 266898
rect 355324 266834 355376 266840
rect 355048 266416 355100 266422
rect 355048 266358 355100 266364
rect 354246 264302 354628 264330
rect 355060 264316 355088 266358
rect 355888 264316 355916 268602
rect 356072 267782 356100 277766
rect 356704 272536 356756 272542
rect 356704 272478 356756 272484
rect 356060 267776 356112 267782
rect 356060 267718 356112 267724
rect 356716 266422 356744 272478
rect 357452 270094 357480 277766
rect 359016 272814 359044 277780
rect 360212 275602 360240 277780
rect 360200 275596 360252 275602
rect 360200 275538 360252 275544
rect 361408 275466 361436 277780
rect 361396 275460 361448 275466
rect 361396 275402 361448 275408
rect 359464 275324 359516 275330
rect 359464 275266 359516 275272
rect 359004 272808 359056 272814
rect 359004 272750 359056 272756
rect 359188 270360 359240 270366
rect 359188 270302 359240 270308
rect 357440 270088 357492 270094
rect 357440 270030 357492 270036
rect 357532 268524 357584 268530
rect 357532 268466 357584 268472
rect 357072 267572 357124 267578
rect 357072 267514 357124 267520
rect 356704 266416 356756 266422
rect 356704 266358 356756 266364
rect 357084 264330 357112 267514
rect 356730 264302 357112 264330
rect 357544 264316 357572 268466
rect 358360 267436 358412 267442
rect 358360 267378 358412 267384
rect 358372 264316 358400 267378
rect 359200 264316 359228 270302
rect 359476 267170 359504 275266
rect 360200 274712 360252 274718
rect 360200 274654 360252 274660
rect 360212 270502 360240 274654
rect 362604 274106 362632 277780
rect 362960 275460 363012 275466
rect 362960 275402 363012 275408
rect 362776 274236 362828 274242
rect 362776 274178 362828 274184
rect 362592 274100 362644 274106
rect 362592 274042 362644 274048
rect 360844 272808 360896 272814
rect 360844 272750 360896 272756
rect 360200 270496 360252 270502
rect 360200 270438 360252 270444
rect 360200 270224 360252 270230
rect 360200 270166 360252 270172
rect 360212 267734 360240 270166
rect 360028 267706 360240 267734
rect 359464 267164 359516 267170
rect 359464 267106 359516 267112
rect 360028 264316 360056 267706
rect 360856 267442 360884 272750
rect 362788 271266 362816 274178
rect 362972 271454 363000 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 363604 271720 363656 271726
rect 363604 271662 363656 271668
rect 362960 271448 363012 271454
rect 362960 271390 363012 271396
rect 362788 271238 362908 271266
rect 362684 271176 362736 271182
rect 362684 271118 362736 271124
rect 360844 267436 360896 267442
rect 360844 267378 360896 267384
rect 360844 267300 360896 267306
rect 360844 267242 360896 267248
rect 360856 264316 360884 267242
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 361684 264316 361712 266358
rect 362696 264330 362724 271118
rect 362880 266422 362908 271238
rect 363328 267164 363380 267170
rect 363328 267106 363380 267112
rect 362868 266416 362920 266422
rect 362868 266358 362920 266364
rect 362526 264302 362724 264330
rect 363340 264316 363368 267106
rect 363616 267034 363644 271662
rect 364156 270088 364208 270094
rect 364156 270030 364208 270036
rect 363604 267028 363656 267034
rect 363604 266970 363656 266976
rect 364168 264316 364196 270030
rect 364352 269958 364380 277766
rect 365904 275732 365956 275738
rect 365904 275674 365956 275680
rect 365916 273970 365944 275674
rect 365904 273964 365956 273970
rect 365904 273906 365956 273912
rect 366100 272678 366128 277780
rect 367296 275466 367324 277780
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 367836 275460 367888 275466
rect 367836 275402 367888 275408
rect 367008 273964 367060 273970
rect 367008 273906 367060 273912
rect 366088 272672 366140 272678
rect 366088 272614 366140 272620
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 364340 269952 364392 269958
rect 364340 269894 364392 269900
rect 364984 269952 365036 269958
rect 364984 269894 365036 269900
rect 364996 264316 365024 269894
rect 366376 267442 366404 271390
rect 366364 267436 366416 267442
rect 366364 267378 366416 267384
rect 365812 267028 365864 267034
rect 365812 266970 365864 266976
rect 365824 264316 365852 266970
rect 367020 264330 367048 273906
rect 367848 268666 367876 275402
rect 368296 274100 368348 274106
rect 368296 274042 368348 274048
rect 367836 268660 367888 268666
rect 367836 268602 367888 268608
rect 368112 267708 368164 267714
rect 368112 267650 368164 267656
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 367048 264330
rect 367480 264316 367508 266358
rect 368124 264330 368152 267650
rect 368308 266422 368336 274042
rect 368492 271590 368520 277780
rect 369688 275738 369716 277780
rect 369676 275732 369728 275738
rect 369676 275674 369728 275680
rect 370884 275330 370912 277780
rect 371252 277766 372094 277794
rect 370872 275324 370924 275330
rect 370872 275266 370924 275272
rect 369860 274848 369912 274854
rect 369860 274790 369912 274796
rect 368756 274712 368808 274718
rect 368756 274654 368808 274660
rect 368480 271584 368532 271590
rect 368480 271526 368532 271532
rect 368768 268394 368796 274654
rect 369492 271584 369544 271590
rect 369492 271526 369544 271532
rect 368756 268388 368808 268394
rect 368756 268330 368808 268336
rect 368296 266416 368348 266422
rect 368296 266358 368348 266364
rect 369504 264330 369532 271526
rect 369872 271318 369900 274790
rect 370964 272672 371016 272678
rect 370964 272614 371016 272620
rect 369860 271312 369912 271318
rect 369860 271254 369912 271260
rect 369952 268388 370004 268394
rect 369952 268330 370004 268336
rect 368124 264302 368322 264330
rect 369150 264302 369532 264330
rect 369964 264316 369992 268330
rect 370976 264330 371004 272614
rect 371252 269822 371280 277766
rect 373080 275732 373132 275738
rect 373080 275674 373132 275680
rect 372528 271312 372580 271318
rect 372528 271254 372580 271260
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 372344 268660 372396 268666
rect 372344 268602 372396 268608
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 370806 264302 371004 264330
rect 371620 264316 371648 266358
rect 372356 264330 372384 268602
rect 372540 266422 372568 271254
rect 373092 267306 373120 275674
rect 373276 274718 373304 277780
rect 373264 274712 373316 274718
rect 373264 274654 373316 274660
rect 374380 271726 374408 277780
rect 375576 274854 375604 277780
rect 376576 275596 376628 275602
rect 376576 275538 376628 275544
rect 375564 274848 375616 274854
rect 375564 274790 375616 274796
rect 376588 273970 376616 275538
rect 376576 273964 376628 273970
rect 376576 273906 376628 273912
rect 376576 273828 376628 273834
rect 376576 273770 376628 273776
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374368 271720 374420 271726
rect 374368 271662 374420 271668
rect 374920 269816 374972 269822
rect 374920 269758 374972 269764
rect 373264 267572 373316 267578
rect 373264 267514 373316 267520
rect 373080 267300 373132 267306
rect 373080 267242 373132 267248
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267514
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 269758
rect 375300 266422 375328 271798
rect 375748 267436 375800 267442
rect 375748 267378 375800 267384
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 375760 264316 375788 267378
rect 376588 264316 376616 273770
rect 376772 272542 376800 277780
rect 377968 275466 377996 277780
rect 377956 275460 378008 275466
rect 377956 275402 378008 275408
rect 377404 275324 377456 275330
rect 377404 275266 377456 275272
rect 376760 272536 376812 272542
rect 376760 272478 376812 272484
rect 377416 271590 377444 275266
rect 378784 274508 378836 274514
rect 378784 274450 378836 274456
rect 377404 271584 377456 271590
rect 377404 271526 377456 271532
rect 377956 270360 378008 270366
rect 377956 270302 378008 270308
rect 377404 268796 377456 268802
rect 377404 268738 377456 268744
rect 377416 264316 377444 268738
rect 377968 267170 377996 270302
rect 378796 267714 378824 274450
rect 379164 271454 379192 277780
rect 379532 277766 380374 277794
rect 379336 271584 379388 271590
rect 379336 271526 379388 271532
rect 379152 271448 379204 271454
rect 379152 271390 379204 271396
rect 378784 267708 378836 267714
rect 378784 267650 378836 267656
rect 378232 267300 378284 267306
rect 378232 267242 378284 267248
rect 377956 267164 378008 267170
rect 377956 267106 378008 267112
rect 378244 264316 378272 267242
rect 379348 264330 379376 271526
rect 379532 268530 379560 277766
rect 381556 272814 381584 277780
rect 382292 277766 382674 277794
rect 383672 277766 383870 277794
rect 382004 273080 382056 273086
rect 382004 273022 382056 273028
rect 381544 272808 381596 272814
rect 381544 272750 381596 272756
rect 380808 272536 380860 272542
rect 380808 272478 380860 272484
rect 379520 268524 379572 268530
rect 379520 268466 379572 268472
rect 380624 267708 380676 267714
rect 380624 267650 380676 267656
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379376 264330
rect 379900 264316 379928 266358
rect 380636 264330 380664 267650
rect 380820 266422 380848 272478
rect 380808 266416 380860 266422
rect 380808 266358 380860 266364
rect 382016 264330 382044 273022
rect 382292 270502 382320 277766
rect 382464 275460 382516 275466
rect 382464 275402 382516 275408
rect 382476 271318 382504 275402
rect 383384 271448 383436 271454
rect 383384 271390 383436 271396
rect 382464 271312 382516 271318
rect 382464 271254 382516 271260
rect 382280 270496 382332 270502
rect 382280 270438 382332 270444
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 380636 264302 380742 264330
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 383396 264330 383424 271390
rect 383672 270230 383700 277766
rect 385052 275738 385080 277780
rect 385960 276004 386012 276010
rect 385960 275946 386012 275952
rect 385040 275732 385092 275738
rect 385040 275674 385092 275680
rect 384948 274372 385000 274378
rect 384948 274314 385000 274320
rect 384764 271720 384816 271726
rect 384764 271662 384816 271668
rect 383844 270496 383896 270502
rect 383844 270438 383896 270444
rect 383660 270224 383712 270230
rect 383660 270166 383712 270172
rect 383856 267170 383884 270438
rect 383844 267164 383896 267170
rect 383844 267106 383896 267112
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 383226 264302 383424 264330
rect 384040 264316 384068 266358
rect 384776 264330 384804 271662
rect 384960 266422 384988 274314
rect 385972 268666 386000 275946
rect 386248 274242 386276 277780
rect 387168 277766 387458 277794
rect 387812 277766 388654 277794
rect 389192 277766 389758 277794
rect 390572 277766 390954 277794
rect 391952 277766 392150 277794
rect 386236 274236 386288 274242
rect 386236 274178 386288 274184
rect 387168 271182 387196 277766
rect 387524 271312 387576 271318
rect 387524 271254 387576 271260
rect 387156 271176 387208 271182
rect 387156 271118 387208 271124
rect 385960 268660 386012 268666
rect 385960 268602 386012 268608
rect 387340 268660 387392 268666
rect 387340 268602 387392 268608
rect 385684 267164 385736 267170
rect 385684 267106 385736 267112
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 384776 264302 384882 264330
rect 385696 264316 385724 267106
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387352 264316 387380 268602
rect 387536 266422 387564 271254
rect 387812 270366 387840 277766
rect 388812 272944 388864 272950
rect 388812 272886 388864 272892
rect 387800 270360 387852 270366
rect 387800 270302 387852 270308
rect 387708 270224 387760 270230
rect 387708 270166 387760 270172
rect 387720 267578 387748 270166
rect 388168 269544 388220 269550
rect 388168 269486 388220 269492
rect 387708 267572 387760 267578
rect 387708 267514 387760 267520
rect 387524 266416 387576 266422
rect 387524 266358 387576 266364
rect 388180 264316 388208 269486
rect 388824 264330 388852 272886
rect 389192 270094 389220 277766
rect 389180 270088 389232 270094
rect 389180 270030 389232 270036
rect 389640 270088 389692 270094
rect 389640 270030 389692 270036
rect 389652 267442 389680 270030
rect 390572 269958 390600 277766
rect 391756 271176 391808 271182
rect 391756 271118 391808 271124
rect 390560 269952 390612 269958
rect 390560 269894 390612 269900
rect 389640 267436 389692 267442
rect 389640 267378 389692 267384
rect 389824 267300 389876 267306
rect 389824 267242 389876 267248
rect 388824 264302 389022 264330
rect 389836 264316 389864 267242
rect 390652 266756 390704 266762
rect 390652 266698 390704 266704
rect 390664 264316 390692 266698
rect 391768 264330 391796 271118
rect 391952 270502 391980 277766
rect 393332 275602 393360 277780
rect 393872 275868 393924 275874
rect 393872 275810 393924 275816
rect 393320 275596 393372 275602
rect 393320 275538 393372 275544
rect 393884 271590 393912 275810
rect 394528 274106 394556 277780
rect 395068 275596 395120 275602
rect 395068 275538 395120 275544
rect 394516 274100 394568 274106
rect 394516 274042 394568 274048
rect 394332 272808 394384 272814
rect 394332 272750 394384 272756
rect 393872 271584 393924 271590
rect 393872 271526 393924 271532
rect 391940 270496 391992 270502
rect 391940 270438 391992 270444
rect 391940 269952 391992 269958
rect 391940 269894 391992 269900
rect 391952 267034 391980 269894
rect 393320 269680 393372 269686
rect 393320 269622 393372 269628
rect 393332 267714 393360 269622
rect 393320 267708 393372 267714
rect 393320 267650 393372 267656
rect 391940 267028 391992 267034
rect 391940 266970 391992 266976
rect 392308 267028 392360 267034
rect 392308 266970 392360 266976
rect 391506 264302 391796 264330
rect 392320 264316 392348 266970
rect 393136 266892 393188 266898
rect 393136 266834 393188 266840
rect 393148 264316 393176 266834
rect 394344 264330 394372 272750
rect 395080 271862 395108 275538
rect 395724 274514 395752 277780
rect 396920 275330 396948 277780
rect 397472 277766 398038 277794
rect 396908 275324 396960 275330
rect 396908 275266 396960 275272
rect 395712 274508 395764 274514
rect 395712 274450 395764 274456
rect 395344 274100 395396 274106
rect 395344 274042 395396 274048
rect 395068 271856 395120 271862
rect 395068 271798 395120 271804
rect 394792 267436 394844 267442
rect 394792 267378 394844 267384
rect 393990 264302 394372 264330
rect 394804 264316 394832 267378
rect 395356 267306 395384 274042
rect 397276 273828 397328 273834
rect 397276 273770 397328 273776
rect 395528 271584 395580 271590
rect 395528 271526 395580 271532
rect 395344 267300 395396 267306
rect 395344 267242 395396 267248
rect 395540 266762 395568 271526
rect 397092 267300 397144 267306
rect 397092 267242 397144 267248
rect 395528 266756 395580 266762
rect 395528 266698 395580 266704
rect 395620 266552 395672 266558
rect 395620 266494 395672 266500
rect 395632 264316 395660 266494
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 396460 264316 396488 266358
rect 397104 264330 397132 267242
rect 397288 266422 397316 273770
rect 397472 268394 397500 277766
rect 399220 272678 399248 277780
rect 400220 275732 400272 275738
rect 400220 275674 400272 275680
rect 400232 274378 400260 275674
rect 400416 275466 400444 277780
rect 401612 276010 401640 277780
rect 401796 277766 402822 277794
rect 401600 276004 401652 276010
rect 401600 275946 401652 275952
rect 400404 275460 400456 275466
rect 400404 275402 400456 275408
rect 400404 275324 400456 275330
rect 400404 275266 400456 275272
rect 400220 274372 400272 274378
rect 400220 274314 400272 274320
rect 400128 274236 400180 274242
rect 400128 274178 400180 274184
rect 399208 272672 399260 272678
rect 399208 272614 399260 272620
rect 398748 268524 398800 268530
rect 398748 268466 398800 268472
rect 397460 268388 397512 268394
rect 397460 268330 397512 268336
rect 398760 266898 398788 268466
rect 399760 268388 399812 268394
rect 399760 268330 399812 268336
rect 398748 266892 398800 266898
rect 398748 266834 398800 266840
rect 398104 266756 398156 266762
rect 398104 266698 398156 266704
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 266698
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 268330
rect 400140 266422 400168 274178
rect 400416 272950 400444 275266
rect 401508 273216 401560 273222
rect 401508 273158 401560 273164
rect 400404 272944 400456 272950
rect 400404 272886 400456 272892
rect 400588 270496 400640 270502
rect 400588 270438 400640 270444
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 270438
rect 401520 267734 401548 273158
rect 401796 270230 401824 277766
rect 404004 275602 404032 277780
rect 404372 277766 405214 277794
rect 405752 277766 406318 277794
rect 403992 275596 404044 275602
rect 403992 275538 404044 275544
rect 403624 275460 403676 275466
rect 403624 275402 403676 275408
rect 403636 271182 403664 275402
rect 403992 274644 404044 274650
rect 403992 274586 404044 274592
rect 403624 271176 403676 271182
rect 403624 271118 403676 271124
rect 401784 270224 401836 270230
rect 401784 270166 401836 270172
rect 401692 269408 401744 269414
rect 401692 269350 401744 269356
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401704 267170 401732 269350
rect 404004 267734 404032 274586
rect 404176 271176 404228 271182
rect 404176 271118 404228 271124
rect 402244 267708 402296 267714
rect 402244 267650 402296 267656
rect 403912 267706 404032 267734
rect 401692 267164 401744 267170
rect 401692 267106 401744 267112
rect 402256 264316 402284 267650
rect 403072 266892 403124 266898
rect 403072 266834 403124 266840
rect 403084 264316 403112 266834
rect 403912 264316 403940 267706
rect 404188 266898 404216 271118
rect 404372 269822 404400 277766
rect 405004 270904 405056 270910
rect 405004 270846 405056 270852
rect 404360 269816 404412 269822
rect 404360 269758 404412 269764
rect 404728 267572 404780 267578
rect 404728 267514 404780 267520
rect 404176 266892 404228 266898
rect 404176 266834 404228 266840
rect 404740 264316 404768 267514
rect 405016 266558 405044 270846
rect 405752 270094 405780 277766
rect 407500 273970 407528 277780
rect 408512 277766 408710 277794
rect 407672 275596 407724 275602
rect 407672 275538 407724 275544
rect 407488 273964 407540 273970
rect 407488 273906 407540 273912
rect 406844 272944 406896 272950
rect 406844 272886 406896 272892
rect 405740 270088 405792 270094
rect 405740 270030 405792 270036
rect 405556 266892 405608 266898
rect 405556 266834 405608 266840
rect 405004 266552 405056 266558
rect 405004 266494 405056 266500
rect 405568 264316 405596 266834
rect 406856 264330 406884 272886
rect 407684 272814 407712 275538
rect 407672 272808 407724 272814
rect 407672 272750 407724 272756
rect 408132 272808 408184 272814
rect 408132 272750 408184 272756
rect 407212 270360 407264 270366
rect 407212 270302 407264 270308
rect 406410 264302 406884 264330
rect 407224 264316 407252 270302
rect 408144 267734 408172 272750
rect 408512 268802 408540 277766
rect 409236 274508 409288 274514
rect 409236 274450 409288 274456
rect 408500 268796 408552 268802
rect 408500 268738 408552 268744
rect 408052 267706 408172 267734
rect 408052 264316 408080 267706
rect 409248 264330 409276 274450
rect 409696 270088 409748 270094
rect 409696 270030 409748 270036
rect 408894 264302 409276 264330
rect 409708 264316 409736 270030
rect 409892 269958 409920 277780
rect 411088 275874 411116 277780
rect 412008 277766 412298 277794
rect 412652 277766 413402 277794
rect 411076 275868 411128 275874
rect 411076 275810 411128 275816
rect 411260 275868 411312 275874
rect 411260 275810 411312 275816
rect 410524 270224 410576 270230
rect 410524 270166 410576 270172
rect 409880 269952 409932 269958
rect 409880 269894 409932 269900
rect 410536 264316 410564 270166
rect 411272 268938 411300 275810
rect 412008 272542 412036 277766
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411996 272536 412048 272542
rect 411996 272478 412048 272484
rect 411260 268932 411312 268938
rect 411260 268874 411312 268880
rect 412284 266422 412312 272614
rect 412456 269952 412508 269958
rect 412456 269894 412508 269900
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 411364 264316 411392 266358
rect 412468 264330 412496 269894
rect 412652 269686 412680 277766
rect 414584 273086 414612 277780
rect 415780 275874 415808 277780
rect 415768 275868 415820 275874
rect 415768 275810 415820 275816
rect 415308 274780 415360 274786
rect 415308 274722 415360 274728
rect 414572 273080 414624 273086
rect 414572 273022 414624 273028
rect 413836 272536 413888 272542
rect 413836 272478 413888 272484
rect 412640 269680 412692 269686
rect 412640 269622 412692 269628
rect 413008 268252 413060 268258
rect 413008 268194 413060 268200
rect 412206 264302 412496 264330
rect 413020 264316 413048 268194
rect 413848 264316 413876 272478
rect 415320 271726 415348 274722
rect 416596 274372 416648 274378
rect 416596 274314 416648 274320
rect 415308 271720 415360 271726
rect 415308 271662 415360 271668
rect 414480 270632 414532 270638
rect 414480 270574 414532 270580
rect 414492 266762 414520 270574
rect 416412 268796 416464 268802
rect 416412 268738 416464 268744
rect 416424 267442 416452 268738
rect 416412 267436 416464 267442
rect 416412 267378 416464 267384
rect 414664 267164 414716 267170
rect 414664 267106 414716 267112
rect 414480 266756 414532 266762
rect 414480 266698 414532 266704
rect 414676 264316 414704 267106
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 415504 264316 415532 266358
rect 416608 264330 416636 274314
rect 416976 271454 417004 277780
rect 418172 275738 418200 277780
rect 418160 275732 418212 275738
rect 418160 275674 418212 275680
rect 418344 275732 418396 275738
rect 418344 275674 418396 275680
rect 418356 273834 418384 275674
rect 418528 274916 418580 274922
rect 418528 274858 418580 274864
rect 418344 273828 418396 273834
rect 418344 273770 418396 273776
rect 416964 271448 417016 271454
rect 416964 271390 417016 271396
rect 418068 271040 418120 271046
rect 418068 270982 418120 270988
rect 417148 269816 417200 269822
rect 417148 269758 417200 269764
rect 416346 264302 416636 264330
rect 417160 264316 417188 269758
rect 418080 267734 418108 270982
rect 418540 268666 418568 274858
rect 419368 274786 419396 277780
rect 419552 277766 420578 277794
rect 421392 277766 421682 277794
rect 419356 274780 419408 274786
rect 419356 274722 419408 274728
rect 418988 271448 419040 271454
rect 418988 271390 419040 271396
rect 418528 268660 418580 268666
rect 418528 268602 418580 268608
rect 417988 267706 418108 267734
rect 417988 264316 418016 267706
rect 419000 267034 419028 271390
rect 419552 269414 419580 277766
rect 420736 273964 420788 273970
rect 420736 273906 420788 273912
rect 419540 269408 419592 269414
rect 419540 269350 419592 269356
rect 419816 269408 419868 269414
rect 419816 269350 419868 269356
rect 419632 267436 419684 267442
rect 419632 267378 419684 267384
rect 418988 267028 419040 267034
rect 418988 266970 419040 266976
rect 418804 266620 418856 266626
rect 418804 266562 418856 266568
rect 418816 264316 418844 266562
rect 419644 264316 419672 267378
rect 419828 266422 419856 269350
rect 419816 266416 419868 266422
rect 419816 266358 419868 266364
rect 420748 264330 420776 273906
rect 421392 271318 421420 277766
rect 422864 274922 422892 277780
rect 423588 275868 423640 275874
rect 423588 275810 423640 275816
rect 422852 274916 422904 274922
rect 422852 274858 422904 274864
rect 423036 274780 423088 274786
rect 423036 274722 423088 274728
rect 421380 271312 421432 271318
rect 421380 271254 421432 271260
rect 421564 271312 421616 271318
rect 421564 271254 421616 271260
rect 421576 267306 421604 271254
rect 422116 269680 422168 269686
rect 422116 269622 422168 269628
rect 421564 267300 421616 267306
rect 421564 267242 421616 267248
rect 421288 266484 421340 266490
rect 421288 266426 421340 266432
rect 420486 264302 420776 264330
rect 421300 264316 421328 266426
rect 422128 264316 422156 269622
rect 423048 269550 423076 274722
rect 423600 274242 423628 275810
rect 424060 274786 424088 277780
rect 425256 275330 425284 277780
rect 425244 275324 425296 275330
rect 425244 275266 425296 275272
rect 426256 275052 426308 275058
rect 426256 274994 426308 275000
rect 424048 274780 424100 274786
rect 424048 274722 424100 274728
rect 423588 274236 423640 274242
rect 423588 274178 423640 274184
rect 424968 273080 425020 273086
rect 424968 273022 425020 273028
rect 423036 269544 423088 269550
rect 423036 269486 423088 269492
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267714 422340 268058
rect 422300 267708 422352 267714
rect 422300 267650 422352 267656
rect 422944 267028 422996 267034
rect 422944 266970 422996 266976
rect 422956 264316 422984 266970
rect 423772 266756 423824 266762
rect 423772 266698 423824 266704
rect 423784 264316 423812 266698
rect 424612 264316 424640 269486
rect 424980 266762 425008 273022
rect 425704 270768 425756 270774
rect 425704 270710 425756 270716
rect 425716 266898 425744 270710
rect 426072 267300 426124 267306
rect 426072 267242 426124 267248
rect 425704 266892 425756 266898
rect 425704 266834 425756 266840
rect 424968 266756 425020 266762
rect 424968 266698 425020 266704
rect 425428 266756 425480 266762
rect 425428 266698 425480 266704
rect 425440 264316 425468 266698
rect 426084 264330 426112 267242
rect 426268 266762 426296 274994
rect 426452 274106 426480 277780
rect 427452 274236 427504 274242
rect 427452 274178 427504 274184
rect 426440 274100 426492 274106
rect 426440 274042 426492 274048
rect 426256 266756 426308 266762
rect 426256 266698 426308 266704
rect 427464 264330 427492 274178
rect 427648 271590 427676 277780
rect 428844 275466 428872 277780
rect 429672 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275460 428884 275466
rect 428832 275402 428884 275408
rect 427820 275324 427872 275330
rect 427820 275266 427872 275272
rect 427832 273222 427860 275266
rect 429200 275188 429252 275194
rect 429200 275130 429252 275136
rect 429212 273306 429240 275130
rect 428936 273278 429240 273306
rect 427820 273216 427872 273222
rect 427820 273158 427872 273164
rect 427636 271584 427688 271590
rect 427636 271526 427688 271532
rect 428740 269068 428792 269074
rect 428740 269010 428792 269016
rect 427912 266756 427964 266762
rect 427912 266698 427964 266704
rect 426084 264302 426282 264330
rect 427110 264302 427492 264330
rect 427924 264316 427952 266698
rect 428752 264316 428780 269010
rect 428936 266762 428964 273278
rect 429672 271454 429700 277766
rect 429844 272400 429896 272406
rect 429844 272342 429896 272348
rect 429660 271448 429712 271454
rect 429660 271390 429712 271396
rect 429568 268932 429620 268938
rect 429568 268874 429620 268880
rect 428924 266756 428976 266762
rect 428924 266698 428976 266704
rect 429580 264316 429608 268874
rect 429856 267578 429884 272342
rect 430592 268530 430620 277766
rect 432340 275602 432368 277780
rect 433352 277766 433550 277794
rect 432972 276004 433024 276010
rect 432972 275946 433024 275952
rect 432328 275596 432380 275602
rect 432328 275538 432380 275544
rect 431684 274100 431736 274106
rect 431684 274042 431736 274048
rect 430580 268524 430632 268530
rect 430580 268466 430632 268472
rect 430396 267708 430448 267714
rect 430396 267650 430448 267656
rect 429844 267572 429896 267578
rect 429844 267514 429896 267520
rect 430408 264316 430436 267650
rect 431696 264330 431724 274042
rect 432984 267734 433012 275946
rect 433156 271856 433208 271862
rect 433156 271798 433208 271804
rect 432892 267706 433012 267734
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267706
rect 433168 266422 433196 271798
rect 433352 268802 433380 277766
rect 434444 271584 434496 271590
rect 434444 271526 434496 271532
rect 433340 268796 433392 268802
rect 433340 268738 433392 268744
rect 433708 268524 433760 268530
rect 433708 268466 433760 268472
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433720 264316 433748 268466
rect 434456 264330 434484 271526
rect 434732 270910 434760 277780
rect 435928 275738 435956 277780
rect 435916 275732 435968 275738
rect 435916 275674 435968 275680
rect 435732 275460 435784 275466
rect 435732 275402 435784 275408
rect 434720 270904 434772 270910
rect 434720 270846 434772 270852
rect 435744 264330 435772 275402
rect 437032 271318 437060 277780
rect 437952 277766 438242 277794
rect 437204 271720 437256 271726
rect 437204 271662 437256 271668
rect 437020 271312 437072 271318
rect 437020 271254 437072 271260
rect 436192 267844 436244 267850
rect 436192 267786 436244 267792
rect 434456 264302 434562 264330
rect 435390 264302 435772 264330
rect 436204 264316 436232 267786
rect 436744 267572 436796 267578
rect 436744 267514 436796 267520
rect 436756 267170 436784 267514
rect 436744 267164 436796 267170
rect 436744 267106 436796 267112
rect 437216 264330 437244 271662
rect 437952 270638 437980 277766
rect 439424 275874 439452 277780
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439412 275868 439464 275874
rect 439412 275810 439464 275816
rect 438860 275596 438912 275602
rect 438860 275538 438912 275544
rect 438872 274650 438900 275538
rect 438860 274644 438912 274650
rect 438860 274586 438912 274592
rect 439320 273828 439372 273834
rect 439320 273770 439372 273776
rect 438124 273692 438176 273698
rect 438124 273634 438176 273640
rect 437940 270632 437992 270638
rect 437940 270574 437992 270580
rect 438136 266898 438164 273634
rect 438768 273216 438820 273222
rect 438768 273158 438820 273164
rect 438780 267734 438808 273158
rect 438688 267706 438808 267734
rect 438124 266892 438176 266898
rect 438124 266834 438176 266840
rect 437848 266756 437900 266762
rect 437848 266698 437900 266704
rect 437046 264302 437244 264330
rect 437860 264316 437888 266698
rect 438688 264316 438716 267706
rect 439332 266422 439360 273770
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 439320 266416 439372 266422
rect 439320 266358 439372 266364
rect 439976 264330 440004 271390
rect 440252 268394 440280 277766
rect 441632 270502 441660 277766
rect 443012 275330 443040 277780
rect 443288 277766 444222 277794
rect 443000 275324 443052 275330
rect 443000 275266 443052 275272
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269272 441672 269278
rect 441620 269214 441672 269220
rect 441160 268796 441212 268802
rect 441160 268738 441212 268744
rect 440240 268388 440292 268394
rect 440240 268330 440292 268336
rect 440332 267164 440384 267170
rect 440332 267106 440384 267112
rect 439530 264302 440004 264330
rect 440344 264316 440372 267106
rect 441172 264316 441200 268738
rect 441632 267578 441660 269214
rect 443288 268122 443316 277766
rect 443644 275868 443696 275874
rect 443644 275810 443696 275816
rect 443276 268116 443328 268122
rect 443276 268058 443328 268064
rect 441620 267572 441672 267578
rect 441620 267514 441672 267520
rect 442816 267572 442868 267578
rect 442816 267514 442868 267520
rect 441988 266552 442040 266558
rect 441988 266494 442040 266500
rect 442000 264316 442028 266494
rect 442828 264316 442856 267514
rect 443656 267170 443684 275810
rect 445312 271182 445340 277780
rect 446508 275602 446536 277780
rect 446496 275596 446548 275602
rect 446496 275538 446548 275544
rect 446404 273556 446456 273562
rect 446404 273498 446456 273504
rect 445668 271312 445720 271318
rect 445668 271254 445720 271260
rect 445300 271176 445352 271182
rect 445300 271118 445352 271124
rect 445024 270632 445076 270638
rect 445024 270574 445076 270580
rect 443920 268660 443972 268666
rect 443920 268602 443972 268608
rect 443644 267164 443696 267170
rect 443644 267106 443696 267112
rect 443932 264330 443960 268602
rect 445036 266558 445064 270574
rect 445300 267164 445352 267170
rect 445300 267106 445352 267112
rect 445024 266552 445076 266558
rect 445024 266494 445076 266500
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 443670 264302 443960 264330
rect 444484 264316 444512 266358
rect 445312 264316 445340 267106
rect 445680 266422 445708 271254
rect 446416 267442 446444 273498
rect 447704 272406 447732 277780
rect 448244 275324 448296 275330
rect 448244 275266 448296 275272
rect 447692 272400 447744 272406
rect 447692 272342 447744 272348
rect 447784 272128 447836 272134
rect 447784 272070 447836 272076
rect 446404 267436 446456 267442
rect 446404 267378 446456 267384
rect 446956 266892 447008 266898
rect 446956 266834 447008 266840
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446128 266416 446180 266422
rect 446128 266358 446180 266364
rect 446140 264316 446168 266358
rect 446968 264316 446996 266834
rect 447796 266422 447824 272070
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 448256 264330 448284 275266
rect 448900 270774 448928 277780
rect 450096 272950 450124 277780
rect 451306 277766 451504 277794
rect 450084 272944 450136 272950
rect 450084 272886 450136 272892
rect 451096 272944 451148 272950
rect 451096 272886 451148 272892
rect 449808 271176 449860 271182
rect 449808 271118 449860 271124
rect 448888 270768 448940 270774
rect 448888 270710 448940 270716
rect 448612 267980 448664 267986
rect 448612 267922 448664 267928
rect 447810 264302 448284 264330
rect 448624 264316 448652 267922
rect 449820 264330 449848 271118
rect 450268 267436 450320 267442
rect 450268 267378 450320 267384
rect 449466 264302 449848 264330
rect 450280 264316 450308 267378
rect 451108 264316 451136 272886
rect 451476 270366 451504 277766
rect 452120 277766 452502 277794
rect 452120 272814 452148 277766
rect 453592 274718 453620 277780
rect 454144 277766 454802 277794
rect 455432 277766 455998 277794
rect 453948 275596 454000 275602
rect 453948 275538 454000 275544
rect 453580 274712 453632 274718
rect 453580 274654 453632 274660
rect 453304 274508 453356 274514
rect 453304 274450 453356 274456
rect 452108 272808 452160 272814
rect 452108 272750 452160 272756
rect 452292 272808 452344 272814
rect 452292 272750 452344 272756
rect 451464 270360 451516 270366
rect 451464 270302 451516 270308
rect 452304 264330 452332 272750
rect 453316 267306 453344 274450
rect 453960 274378 453988 275538
rect 453948 274372 454000 274378
rect 453948 274314 454000 274320
rect 453580 270496 453632 270502
rect 453580 270438 453632 270444
rect 453304 267300 453356 267306
rect 453304 267242 453356 267248
rect 452752 266756 452804 266762
rect 452752 266698 452804 266704
rect 451950 264302 452332 264330
rect 452764 264316 452792 266698
rect 453592 264316 453620 270438
rect 454144 270094 454172 277766
rect 455432 270230 455460 277766
rect 457180 272678 457208 277780
rect 458192 277766 458390 277794
rect 459586 277766 459784 277794
rect 457444 275732 457496 275738
rect 457444 275674 457496 275680
rect 457168 272672 457220 272678
rect 457168 272614 457220 272620
rect 455788 271312 455840 271318
rect 455840 271260 456380 271266
rect 455788 271254 456380 271260
rect 455800 271238 456380 271254
rect 456352 271182 456380 271238
rect 456340 271176 456392 271182
rect 456340 271118 456392 271124
rect 456064 270904 456116 270910
rect 456064 270846 456116 270852
rect 455420 270224 455472 270230
rect 455420 270166 455472 270172
rect 454132 270088 454184 270094
rect 454132 270030 454184 270036
rect 454500 270088 454552 270094
rect 454500 270030 454552 270036
rect 454512 267034 454540 270030
rect 455236 267300 455288 267306
rect 455236 267242 455288 267248
rect 454500 267028 454552 267034
rect 454500 266970 454552 266976
rect 454776 267028 454828 267034
rect 454776 266970 454828 266976
rect 454788 264330 454816 266970
rect 454434 264302 454816 264330
rect 455248 264316 455276 267242
rect 456076 266898 456104 270846
rect 456432 270360 456484 270366
rect 456432 270302 456484 270308
rect 456064 266892 456116 266898
rect 456064 266834 456116 266840
rect 456444 264330 456472 270302
rect 457456 266762 457484 275674
rect 457996 272672 458048 272678
rect 457996 272614 458048 272620
rect 457720 266892 457772 266898
rect 457720 266834 457772 266840
rect 457444 266756 457496 266762
rect 457444 266698 457496 266704
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456090 264302 456472 264330
rect 456904 264316 456932 266358
rect 457732 264316 457760 266834
rect 458008 266422 458036 272614
rect 458192 269958 458220 277766
rect 458824 274644 458876 274650
rect 458824 274586 458876 274592
rect 458180 269952 458232 269958
rect 458180 269894 458232 269900
rect 458548 269952 458600 269958
rect 458548 269894 458600 269900
rect 457996 266416 458048 266422
rect 457996 266358 458048 266364
rect 458560 264316 458588 269894
rect 458836 267714 458864 274586
rect 459560 268388 459612 268394
rect 459560 268330 459612 268336
rect 458824 267708 458876 267714
rect 458824 267650 458876 267656
rect 459572 267186 459600 268330
rect 459756 268258 459784 277766
rect 460676 272542 460704 277780
rect 460952 277766 461886 277794
rect 462332 277766 463082 277794
rect 460664 272536 460716 272542
rect 460664 272478 460716 272484
rect 460952 269278 460980 277766
rect 461952 272536 462004 272542
rect 461952 272478 462004 272484
rect 461400 270224 461452 270230
rect 461400 270166 461452 270172
rect 460940 269272 460992 269278
rect 460940 269214 460992 269220
rect 459744 268252 459796 268258
rect 459744 268194 459796 268200
rect 460204 267708 460256 267714
rect 460204 267650 460256 267656
rect 459204 267158 459600 267186
rect 459204 267034 459232 267158
rect 459192 267028 459244 267034
rect 459192 266970 459244 266976
rect 459376 267028 459428 267034
rect 459376 266970 459428 266976
rect 459388 264316 459416 266970
rect 460216 264316 460244 267650
rect 461412 264330 461440 270166
rect 461964 267734 461992 272478
rect 462332 269414 462360 277766
rect 464264 275602 464292 277780
rect 465092 277766 465474 277794
rect 464804 276820 464856 276826
rect 464804 276762 464856 276768
rect 464252 275596 464304 275602
rect 464252 275538 464304 275544
rect 464436 275596 464488 275602
rect 464436 275538 464488 275544
rect 463792 271040 463844 271046
rect 463792 270982 463844 270988
rect 463804 270774 463832 270982
rect 463792 270768 463844 270774
rect 463792 270710 463844 270716
rect 462320 269408 462372 269414
rect 462320 269350 462372 269356
rect 463516 269272 463568 269278
rect 463516 269214 463568 269220
rect 461058 264302 461440 264330
rect 461872 267706 461992 267734
rect 461872 264316 461900 267706
rect 462688 266756 462740 266762
rect 462688 266698 462740 266704
rect 462700 264316 462728 266698
rect 463528 264316 463556 269214
rect 464448 266898 464476 275538
rect 464436 266892 464488 266898
rect 464436 266834 464488 266840
rect 464816 264330 464844 276762
rect 465092 269822 465120 277766
rect 465724 271312 465776 271318
rect 465724 271254 465776 271260
rect 465908 271312 465960 271318
rect 465908 271254 465960 271260
rect 465736 271046 465764 271254
rect 465724 271040 465776 271046
rect 465724 270982 465776 270988
rect 465920 270910 465948 271254
rect 465908 270904 465960 270910
rect 465908 270846 465960 270852
rect 466656 270774 466684 277780
rect 467852 273698 467880 277780
rect 467840 273692 467892 273698
rect 467840 273634 467892 273640
rect 468956 273562 468984 277780
rect 470152 273970 470180 277780
rect 470140 273964 470192 273970
rect 470140 273906 470192 273912
rect 470416 273964 470468 273970
rect 470416 273906 470468 273912
rect 468944 273556 468996 273562
rect 468944 273498 468996 273504
rect 467748 272264 467800 272270
rect 467748 272206 467800 272212
rect 466644 270768 466696 270774
rect 466644 270710 466696 270716
rect 467104 270768 467156 270774
rect 467104 270710 467156 270716
rect 465080 269816 465132 269822
rect 465080 269758 465132 269764
rect 466000 269816 466052 269822
rect 466000 269758 466052 269764
rect 465172 266756 465224 266762
rect 465172 266698 465224 266704
rect 464370 264302 464844 264330
rect 465184 264316 465212 266698
rect 466012 264316 466040 269758
rect 467116 267034 467144 270710
rect 467104 267028 467156 267034
rect 467104 266970 467156 266976
rect 467288 267028 467340 267034
rect 467288 266970 467340 266976
rect 467300 266626 467328 266970
rect 467288 266620 467340 266626
rect 467288 266562 467340 266568
rect 467564 266620 467616 266626
rect 467564 266562 467616 266568
rect 466828 266416 466880 266422
rect 466828 266358 466880 266364
rect 466840 264316 466868 266358
rect 467576 264330 467604 266562
rect 467760 266422 467788 272206
rect 468482 269784 468538 269793
rect 468482 269719 468538 269728
rect 467748 266416 467800 266422
rect 467748 266358 467800 266364
rect 467576 264302 467682 264330
rect 468496 264316 468524 269719
rect 469496 268252 469548 268258
rect 469496 268194 469548 268200
rect 469508 267034 469536 268194
rect 469496 267028 469548 267034
rect 469496 266970 469548 266976
rect 469956 266892 470008 266898
rect 469956 266834 470008 266840
rect 470140 266892 470192 266898
rect 470140 266834 470192 266840
rect 469312 266416 469364 266422
rect 469312 266358 469364 266364
rect 469324 264316 469352 266358
rect 469968 266286 469996 266834
rect 469956 266280 470008 266286
rect 469956 266222 470008 266228
rect 470152 264316 470180 266834
rect 470428 266422 470456 273906
rect 471348 273834 471376 277780
rect 472084 277766 472558 277794
rect 473372 277766 473754 277794
rect 471888 274780 471940 274786
rect 471888 274722 471940 274728
rect 471336 273828 471388 273834
rect 471336 273770 471388 273776
rect 471900 273222 471928 274722
rect 471888 273216 471940 273222
rect 471888 273158 471940 273164
rect 471612 272400 471664 272406
rect 471612 272342 471664 272348
rect 470966 269240 471022 269249
rect 470966 269175 471022 269184
rect 470416 266416 470468 266422
rect 470416 266358 470468 266364
rect 470980 264316 471008 269175
rect 471624 264330 471652 272342
rect 472084 269686 472112 277766
rect 473084 273828 473136 273834
rect 473084 273770 473136 273776
rect 472072 269680 472124 269686
rect 472072 269622 472124 269628
rect 473096 264330 473124 273770
rect 473372 270094 473400 277766
rect 474372 274372 474424 274378
rect 474372 274314 474424 274320
rect 473360 270088 473412 270094
rect 473360 270030 473412 270036
rect 474384 266898 474412 274314
rect 474936 273086 474964 277780
rect 475752 273420 475804 273426
rect 475752 273362 475804 273368
rect 474924 273080 474976 273086
rect 474924 273022 474976 273028
rect 474648 269680 474700 269686
rect 474648 269622 474700 269628
rect 473452 266892 473504 266898
rect 473452 266834 473504 266840
rect 474372 266892 474424 266898
rect 474372 266834 474424 266840
rect 471624 264302 471822 264330
rect 472650 264302 473124 264330
rect 473464 264316 473492 266834
rect 474660 264330 474688 269622
rect 475200 269068 475252 269074
rect 475200 269010 475252 269016
rect 475384 269068 475436 269074
rect 475384 269010 475436 269016
rect 475212 268122 475240 269010
rect 475396 268258 475424 269010
rect 475384 268252 475436 268258
rect 475384 268194 475436 268200
rect 475200 268116 475252 268122
rect 475200 268058 475252 268064
rect 475108 266892 475160 266898
rect 475108 266834 475160 266840
rect 474306 264302 474688 264330
rect 475120 264316 475148 266834
rect 475764 264330 475792 273362
rect 475936 273216 475988 273222
rect 475936 273158 475988 273164
rect 475948 266898 475976 273158
rect 476132 269550 476160 277780
rect 477236 275058 477264 277780
rect 477224 275052 477276 275058
rect 477224 274994 477276 275000
rect 478432 274514 478460 277780
rect 479352 277766 479642 277794
rect 478972 274916 479024 274922
rect 478972 274858 479024 274864
rect 478420 274508 478472 274514
rect 478420 274450 478472 274456
rect 478788 273556 478840 273562
rect 478788 273498 478840 273504
rect 476120 269544 476172 269550
rect 476120 269486 476172 269492
rect 476764 269544 476816 269550
rect 476764 269486 476816 269492
rect 475936 266892 475988 266898
rect 475936 266834 475988 266840
rect 475764 264302 475962 264330
rect 476776 264316 476804 269486
rect 477590 266384 477646 266393
rect 477590 266319 477646 266328
rect 477604 264316 477632 266319
rect 478800 264330 478828 273498
rect 478984 268122 479012 274858
rect 479352 274242 479380 277766
rect 480824 275194 480852 277780
rect 480812 275188 480864 275194
rect 480812 275130 480864 275136
rect 482020 274922 482048 277780
rect 483216 277394 483244 277780
rect 483124 277366 483244 277394
rect 482836 276684 482888 276690
rect 482836 276626 482888 276632
rect 482008 274916 482060 274922
rect 482008 274858 482060 274864
rect 481364 274508 481416 274514
rect 481364 274450 481416 274456
rect 479340 274236 479392 274242
rect 479340 274178 479392 274184
rect 479706 271416 479762 271425
rect 479706 271351 479762 271360
rect 478972 268116 479024 268122
rect 478972 268058 479024 268064
rect 479720 266393 479748 271351
rect 479706 266384 479762 266393
rect 479706 266319 479762 266328
rect 480076 266348 480128 266354
rect 480076 266290 480128 266296
rect 479248 265396 479300 265402
rect 479248 265338 479300 265344
rect 478446 264302 478828 264330
rect 479260 264316 479288 265338
rect 480088 264316 480116 266290
rect 481376 264330 481404 274450
rect 481732 265532 481784 265538
rect 481732 265474 481784 265480
rect 480930 264302 481404 264330
rect 481744 264316 481772 265474
rect 482848 264330 482876 276626
rect 483124 268938 483152 277366
rect 484320 274650 484348 277780
rect 485044 275052 485096 275058
rect 485044 274994 485096 275000
rect 484308 274644 484360 274650
rect 484308 274586 484360 274592
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483112 268932 483164 268938
rect 483112 268874 483164 268880
rect 484122 267064 484178 267073
rect 484122 266999 484178 267008
rect 483204 266756 483256 266762
rect 483204 266698 483256 266704
rect 483216 266490 483244 266698
rect 483204 266484 483256 266490
rect 483204 266426 483256 266432
rect 483388 266484 483440 266490
rect 483388 266426 483440 266432
rect 482586 264302 482876 264330
rect 483400 264316 483428 266426
rect 484136 264330 484164 266999
rect 484320 266490 484348 273634
rect 485056 267578 485084 274994
rect 485516 274106 485544 277780
rect 485504 274100 485556 274106
rect 485504 274042 485556 274048
rect 486712 271862 486740 277780
rect 487908 276010 487936 277780
rect 488552 277766 489118 277794
rect 487896 276004 487948 276010
rect 487896 275946 487948 275952
rect 487160 275188 487212 275194
rect 487160 275130 487212 275136
rect 486976 274236 487028 274242
rect 486976 274178 487028 274184
rect 486700 271856 486752 271862
rect 486700 271798 486752 271804
rect 485044 267572 485096 267578
rect 485044 267514 485096 267520
rect 486988 266490 487016 274178
rect 487172 273834 487200 275130
rect 487804 274916 487856 274922
rect 487804 274858 487856 274864
rect 487160 273828 487212 273834
rect 487160 273770 487212 273776
rect 487816 267578 487844 274858
rect 488356 273828 488408 273834
rect 488356 273770 488408 273776
rect 487160 267572 487212 267578
rect 487160 267514 487212 267520
rect 487804 267572 487856 267578
rect 487804 267514 487856 267520
rect 487172 266762 487200 267514
rect 487160 266756 487212 266762
rect 487160 266698 487212 266704
rect 487528 266756 487580 266762
rect 487528 266698 487580 266704
rect 484308 266484 484360 266490
rect 484308 266426 484360 266432
rect 485872 266484 485924 266490
rect 485872 266426 485924 266432
rect 486976 266484 487028 266490
rect 486976 266426 487028 266432
rect 485044 266212 485096 266218
rect 485044 266154 485096 266160
rect 484136 264302 484242 264330
rect 485056 264316 485084 266154
rect 485884 264316 485912 266426
rect 486700 266076 486752 266082
rect 486700 266018 486752 266024
rect 486712 264316 486740 266018
rect 487540 264316 487568 266698
rect 488368 264316 488396 273770
rect 488552 268530 488580 277766
rect 490300 271590 490328 277780
rect 491496 275466 491524 277780
rect 491864 277766 492614 277794
rect 491484 275460 491536 275466
rect 491484 275402 491536 275408
rect 490288 271584 490340 271590
rect 490288 271526 490340 271532
rect 488540 268524 488592 268530
rect 488540 268466 488592 268472
rect 490840 268252 490892 268258
rect 490840 268194 490892 268200
rect 489184 268116 489236 268122
rect 489184 268058 489236 268064
rect 489196 264316 489224 268058
rect 490012 266484 490064 266490
rect 490012 266426 490064 266432
rect 490024 264316 490052 266426
rect 490852 264316 490880 268194
rect 491864 267850 491892 277766
rect 493140 274644 493192 274650
rect 493140 274586 493192 274592
rect 492036 270904 492088 270910
rect 492036 270846 492088 270852
rect 491852 267844 491904 267850
rect 491852 267786 491904 267792
rect 492048 264330 492076 270846
rect 493152 266626 493180 274586
rect 493796 271726 493824 277780
rect 494256 277766 495006 277794
rect 494060 275460 494112 275466
rect 494060 275402 494112 275408
rect 494072 275058 494100 275402
rect 494060 275052 494112 275058
rect 494060 274994 494112 275000
rect 493784 271720 493836 271726
rect 493784 271662 493836 271668
rect 494256 269074 494284 277766
rect 494428 275052 494480 275058
rect 494428 274994 494480 275000
rect 494440 274650 494468 274994
rect 496188 274786 496216 277780
rect 496176 274780 496228 274786
rect 496176 274722 496228 274728
rect 494428 274644 494480 274650
rect 494428 274586 494480 274592
rect 496544 271856 496596 271862
rect 496544 271798 496596 271804
rect 494704 271584 494756 271590
rect 494704 271526 494756 271532
rect 494716 270638 494744 271526
rect 494704 270632 494756 270638
rect 494704 270574 494756 270580
rect 495348 270632 495400 270638
rect 495348 270574 495400 270580
rect 494244 269068 494296 269074
rect 494244 269010 494296 269016
rect 493324 267844 493376 267850
rect 493324 267786 493376 267792
rect 493140 266620 493192 266626
rect 493140 266562 493192 266568
rect 492496 265940 492548 265946
rect 492496 265882 492548 265888
rect 491694 264302 492076 264330
rect 492508 264316 492536 265882
rect 493336 264316 493364 267786
rect 494704 267572 494756 267578
rect 494704 267514 494756 267520
rect 494716 267170 494744 267514
rect 494704 267164 494756 267170
rect 494704 267106 494756 267112
rect 494888 267164 494940 267170
rect 494888 267106 494940 267112
rect 494704 266756 494756 266762
rect 494900 266744 494928 267106
rect 494756 266716 494928 266744
rect 494704 266698 494756 266704
rect 495164 266620 495216 266626
rect 495164 266562 495216 266568
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 494164 264316 494192 266426
rect 495176 264330 495204 266562
rect 495360 266490 495388 270574
rect 495808 269068 495860 269074
rect 495808 269010 495860 269016
rect 495348 266484 495400 266490
rect 495348 266426 495400 266432
rect 495006 264302 495204 264330
rect 495820 264316 495848 269010
rect 496556 264330 496584 271798
rect 497384 271454 497412 277780
rect 498580 275874 498608 277780
rect 498568 275868 498620 275874
rect 498568 275810 498620 275816
rect 499776 274718 499804 277780
rect 500512 277766 500894 277794
rect 498476 274712 498528 274718
rect 498476 274654 498528 274660
rect 499764 274712 499816 274718
rect 499764 274654 499816 274660
rect 497372 271448 497424 271454
rect 497372 271390 497424 271396
rect 497462 269512 497518 269521
rect 497462 269447 497518 269456
rect 497476 266762 497504 269447
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 497464 266756 497516 266762
rect 497464 266698 497516 266704
rect 497464 266620 497516 266626
rect 497464 266562 497516 266568
rect 496556 264302 496662 264330
rect 497476 264316 497504 266562
rect 498304 264316 498332 268874
rect 498488 268802 498516 274654
rect 499488 271720 499540 271726
rect 499488 271662 499540 271668
rect 498476 268796 498528 268802
rect 498476 268738 498528 268744
rect 499500 264330 499528 271662
rect 500512 271590 500540 277766
rect 502076 275466 502104 277780
rect 502352 277766 503286 277794
rect 504192 277766 504482 277794
rect 502064 275460 502116 275466
rect 502064 275402 502116 275408
rect 501604 274712 501656 274718
rect 501604 274654 501656 274660
rect 500868 273080 500920 273086
rect 500868 273022 500920 273028
rect 500500 271584 500552 271590
rect 500500 271526 500552 271532
rect 500684 268796 500736 268802
rect 500684 268738 500736 268744
rect 499948 266756 500000 266762
rect 499948 266698 500000 266704
rect 499146 264302 499528 264330
rect 499960 264316 499988 266698
rect 500696 264330 500724 268738
rect 500880 266762 500908 273022
rect 501616 267578 501644 274654
rect 501972 271584 502024 271590
rect 501972 271526 502024 271532
rect 501604 267572 501656 267578
rect 501604 267514 501656 267520
rect 500868 266756 500920 266762
rect 500868 266698 500920 266704
rect 501984 264330 502012 271526
rect 502352 268666 502380 277766
rect 504192 271182 504220 277766
rect 504732 275868 504784 275874
rect 504732 275810 504784 275816
rect 504180 271176 504232 271182
rect 504180 271118 504232 271124
rect 504548 271040 504600 271046
rect 504548 270982 504600 270988
rect 504560 270638 504588 270982
rect 504548 270632 504600 270638
rect 504548 270574 504600 270580
rect 502340 268660 502392 268666
rect 502340 268602 502392 268608
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 267572 502484 267578
rect 502432 267514 502484 267520
rect 500696 264302 500802 264330
rect 501630 264302 502012 264330
rect 502444 264316 502472 267514
rect 503272 264316 503300 268602
rect 504088 266756 504140 266762
rect 504088 266698 504140 266704
rect 504100 264316 504128 266698
rect 504744 264330 504772 275810
rect 505664 274718 505692 277780
rect 505836 275460 505888 275466
rect 505836 275402 505888 275408
rect 505652 274712 505704 274718
rect 505652 274654 505704 274660
rect 504916 271448 504968 271454
rect 504916 271390 504968 271396
rect 504928 266762 504956 271390
rect 505848 267442 505876 275402
rect 506480 274712 506532 274718
rect 506480 274654 506532 274660
rect 506110 268424 506166 268433
rect 506110 268359 506166 268368
rect 505836 267436 505888 267442
rect 505836 267378 505888 267384
rect 504916 266756 504968 266762
rect 504916 266698 504968 266704
rect 506124 264330 506152 268359
rect 506492 267986 506520 274654
rect 506860 272134 506888 277780
rect 506848 272128 506900 272134
rect 506848 272070 506900 272076
rect 507308 272128 507360 272134
rect 507308 272070 507360 272076
rect 506480 267980 506532 267986
rect 506480 267922 506532 267928
rect 507320 267170 507348 272070
rect 507964 271318 507992 277780
rect 509160 275330 509188 277780
rect 509148 275324 509200 275330
rect 509148 275266 509200 275272
rect 510356 274718 510384 277780
rect 510528 274780 510580 274786
rect 510528 274722 510580 274728
rect 510344 274712 510396 274718
rect 510344 274654 510396 274660
rect 507952 271312 508004 271318
rect 507952 271254 508004 271260
rect 509148 271312 509200 271318
rect 509148 271254 509200 271260
rect 507766 271144 507822 271153
rect 507766 271079 507822 271088
rect 507584 267572 507636 267578
rect 507584 267514 507636 267520
rect 507308 267164 507360 267170
rect 507308 267106 507360 267112
rect 506572 266756 506624 266762
rect 506572 266698 506624 266704
rect 504744 264302 504942 264330
rect 505770 264302 506152 264330
rect 506584 264316 506612 266698
rect 507596 264330 507624 267514
rect 507780 266762 507808 271079
rect 507952 269408 508004 269414
rect 507952 269350 508004 269356
rect 507964 267073 507992 269350
rect 509160 267734 509188 271254
rect 509068 267706 509188 267734
rect 508412 267436 508464 267442
rect 508412 267378 508464 267384
rect 508228 267164 508280 267170
rect 508228 267106 508280 267112
rect 507950 267064 508006 267073
rect 507950 266999 508006 267008
rect 507768 266756 507820 266762
rect 507768 266698 507820 266704
rect 507426 264302 507624 264330
rect 508240 264316 508268 267106
rect 508424 266762 508452 267378
rect 508412 266756 508464 266762
rect 508412 266698 508464 266704
rect 509068 264316 509096 267706
rect 509884 267436 509936 267442
rect 509884 267378 509936 267384
rect 509896 264316 509924 267378
rect 510540 267306 510568 274722
rect 511552 271182 511580 277780
rect 512552 276004 512604 276010
rect 512552 275946 512604 275952
rect 511540 271176 511592 271182
rect 511540 271118 511592 271124
rect 511908 271176 511960 271182
rect 511908 271118 511960 271124
rect 510712 268524 510764 268530
rect 510712 268466 510764 268472
rect 510528 267300 510580 267306
rect 510528 267242 510580 267248
rect 510724 264316 510752 268466
rect 511920 264330 511948 271118
rect 512564 267714 512592 275946
rect 512748 275466 512776 277780
rect 512736 275460 512788 275466
rect 512736 275402 512788 275408
rect 513748 275324 513800 275330
rect 513748 275266 513800 275272
rect 513194 274136 513250 274145
rect 513194 274071 513250 274080
rect 512552 267708 512604 267714
rect 512552 267650 512604 267656
rect 512368 267300 512420 267306
rect 512368 267242 512420 267248
rect 511566 264302 511948 264330
rect 512380 264316 512408 267242
rect 513208 264316 513236 274071
rect 513760 266898 513788 275266
rect 513944 272950 513972 277780
rect 513932 272944 513984 272950
rect 513932 272886 513984 272892
rect 515140 272814 515168 277780
rect 516244 275738 516272 277780
rect 516520 277766 517454 277794
rect 517624 277766 518650 277794
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 515128 272808 515180 272814
rect 515128 272750 515180 272756
rect 516048 271992 516100 271998
rect 516048 271934 516100 271940
rect 514392 267708 514444 267714
rect 514392 267650 514444 267656
rect 513748 266892 513800 266898
rect 513748 266834 513800 266840
rect 514024 266892 514076 266898
rect 514024 266834 514076 266840
rect 514036 266490 514064 266834
rect 514024 266484 514076 266490
rect 514024 266426 514076 266432
rect 514404 264330 514432 267650
rect 516060 266490 516088 271934
rect 516520 270502 516548 277766
rect 516692 275732 516744 275738
rect 516692 275674 516744 275680
rect 516704 271998 516732 275674
rect 516692 271992 516744 271998
rect 516692 271934 516744 271940
rect 517336 271992 517388 271998
rect 517336 271934 517388 271940
rect 516508 270496 516560 270502
rect 516508 270438 516560 270444
rect 517150 267064 517206 267073
rect 517150 266999 517206 267008
rect 514852 266484 514904 266490
rect 514852 266426 514904 266432
rect 516048 266484 516100 266490
rect 516048 266426 516100 266432
rect 516508 266484 516560 266490
rect 516508 266426 516560 266432
rect 514050 264302 514432 264330
rect 514864 264316 514892 266426
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266426
rect 517164 264330 517192 266999
rect 517348 266490 517376 271934
rect 517624 268394 517652 277766
rect 519832 274786 519860 277780
rect 520292 277766 521042 277794
rect 519820 274780 519872 274786
rect 519820 274722 519872 274728
rect 520096 272944 520148 272950
rect 520096 272886 520148 272892
rect 517796 270496 517848 270502
rect 517796 270438 517848 270444
rect 517612 268388 517664 268394
rect 517612 268330 517664 268336
rect 517808 267442 517836 270438
rect 517796 267436 517848 267442
rect 517796 267378 517848 267384
rect 519818 267336 519874 267345
rect 519818 267271 519874 267280
rect 518716 266892 518768 266898
rect 518716 266834 518768 266840
rect 518900 266892 518952 266898
rect 518900 266834 518952 266840
rect 518728 266642 518756 266834
rect 518912 266642 518940 266834
rect 518728 266614 518940 266642
rect 517336 266484 517388 266490
rect 517336 266426 517388 266432
rect 518992 266484 519044 266490
rect 518992 266426 519044 266432
rect 518164 265668 518216 265674
rect 518164 265610 518216 265616
rect 517164 264302 517362 264330
rect 518176 264316 518204 265610
rect 519004 264316 519032 266426
rect 519832 264316 519860 267271
rect 520108 266490 520136 272886
rect 520292 270366 520320 277766
rect 521474 273048 521530 273057
rect 521474 272983 521530 272992
rect 520280 270360 520332 270366
rect 520280 270302 520332 270308
rect 520648 267300 520700 267306
rect 520648 267242 520700 267248
rect 520096 266484 520148 266490
rect 520096 266426 520148 266432
rect 520660 264316 520688 267242
rect 521488 264316 521516 272983
rect 522224 272678 522252 277780
rect 523420 275602 523448 277780
rect 524524 277394 524552 277780
rect 524432 277366 524552 277394
rect 525352 277766 525734 277794
rect 523408 275596 523460 275602
rect 523408 275538 523460 275544
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 522396 274644 522448 274650
rect 522396 274586 522448 274592
rect 522212 272672 522264 272678
rect 522212 272614 522264 272620
rect 522408 267170 522436 274586
rect 523696 274378 523724 274722
rect 523684 274372 523736 274378
rect 523684 274314 523736 274320
rect 524052 272808 524104 272814
rect 524052 272750 524104 272756
rect 523132 270360 523184 270366
rect 523132 270302 523184 270308
rect 522396 267164 522448 267170
rect 522396 267106 522448 267112
rect 522672 267164 522724 267170
rect 522672 267106 522724 267112
rect 522684 264330 522712 267106
rect 522330 264302 522712 264330
rect 523144 264316 523172 270302
rect 524064 267734 524092 272750
rect 524432 269958 524460 277366
rect 525352 270774 525380 277766
rect 526916 276010 526944 277780
rect 527192 277766 528126 277794
rect 526904 276004 526956 276010
rect 526904 275946 526956 275952
rect 525800 275596 525852 275602
rect 525800 275538 525852 275544
rect 525616 275460 525668 275466
rect 525616 275402 525668 275408
rect 525340 270768 525392 270774
rect 525340 270710 525392 270716
rect 525628 270178 525656 275402
rect 525812 271998 525840 275538
rect 526812 272672 526864 272678
rect 526812 272614 526864 272620
rect 525800 271992 525852 271998
rect 525800 271934 525852 271940
rect 526444 270768 526496 270774
rect 526444 270710 526496 270716
rect 525628 270150 525748 270178
rect 525524 270088 525576 270094
rect 525524 270030 525576 270036
rect 524420 269952 524472 269958
rect 524420 269894 524472 269900
rect 523972 267706 524092 267734
rect 523972 264316 524000 267706
rect 524788 266484 524840 266490
rect 524788 266426 524840 266432
rect 524800 264316 524828 266426
rect 525536 264330 525564 270030
rect 525720 266490 525748 270150
rect 526456 266898 526484 270710
rect 526628 267164 526680 267170
rect 526628 267106 526680 267112
rect 526640 266898 526668 267106
rect 526444 266892 526496 266898
rect 526444 266834 526496 266840
rect 526628 266892 526680 266898
rect 526628 266834 526680 266840
rect 525708 266484 525760 266490
rect 525708 266426 525760 266432
rect 526824 264330 526852 272614
rect 527192 270230 527220 277766
rect 527364 276004 527416 276010
rect 527364 275946 527416 275952
rect 527376 275602 527404 275946
rect 527364 275596 527416 275602
rect 527364 275538 527416 275544
rect 529308 272542 529336 277780
rect 530504 274922 530532 277780
rect 531332 277766 531622 277794
rect 530492 274916 530544 274922
rect 530492 274858 530544 274864
rect 530676 274916 530728 274922
rect 530676 274858 530728 274864
rect 529848 274100 529900 274106
rect 529848 274042 529900 274048
rect 529296 272536 529348 272542
rect 529296 272478 529348 272484
rect 529480 272536 529532 272542
rect 529480 272478 529532 272484
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 528100 270224 528152 270230
rect 528100 270166 528152 270172
rect 527272 266484 527324 266490
rect 527272 266426 527324 266432
rect 525536 264302 525642 264330
rect 526470 264302 526852 264330
rect 527284 264316 527312 266426
rect 528112 264316 528140 270166
rect 529492 267734 529520 272478
rect 529860 267734 529888 274042
rect 529400 267706 529520 267734
rect 529768 267706 529888 267734
rect 529400 264330 529428 267706
rect 528954 264302 529428 264330
rect 529768 264316 529796 267706
rect 530688 267034 530716 274858
rect 530950 270328 531006 270337
rect 530950 270263 531006 270272
rect 530676 267028 530728 267034
rect 530676 266970 530728 266976
rect 530964 264330 530992 270263
rect 531332 269278 531360 277766
rect 532804 276826 532832 277780
rect 532792 276820 532844 276826
rect 532792 276762 532844 276768
rect 532700 275596 532752 275602
rect 532700 275538 532752 275544
rect 532712 274106 532740 275538
rect 534000 275330 534028 277780
rect 534368 277766 535210 277794
rect 533988 275324 534040 275330
rect 533988 275266 534040 275272
rect 532700 274100 532752 274106
rect 532700 274042 532752 274048
rect 533434 273864 533490 273873
rect 533434 273799 533490 273808
rect 531688 269952 531740 269958
rect 531688 269894 531740 269900
rect 531320 269272 531372 269278
rect 531320 269214 531372 269220
rect 531700 264330 531728 269894
rect 532240 267164 532292 267170
rect 532240 267106 532292 267112
rect 530610 264302 530992 264330
rect 531438 264302 531728 264330
rect 532252 264316 532280 267106
rect 533448 264330 533476 273799
rect 533894 272776 533950 272785
rect 533894 272711 533950 272720
rect 533094 264302 533476 264330
rect 533908 264316 533936 272711
rect 534368 269822 534396 277766
rect 535734 275224 535790 275233
rect 535734 275159 535790 275168
rect 534356 269816 534408 269822
rect 534356 269758 534408 269764
rect 535552 269816 535604 269822
rect 535552 269758 535604 269764
rect 534724 268388 534776 268394
rect 534724 268330 534776 268336
rect 534736 264316 534764 268330
rect 535564 264316 535592 269758
rect 535748 268394 535776 275159
rect 536392 272270 536420 277780
rect 537312 277766 537602 277794
rect 537312 275058 537340 277766
rect 538784 275058 538812 277780
rect 539508 275324 539560 275330
rect 539508 275266 539560 275272
rect 537300 275052 537352 275058
rect 537300 274994 537352 275000
rect 537668 275052 537720 275058
rect 537668 274994 537720 275000
rect 538772 275052 538824 275058
rect 538772 274994 538824 275000
rect 537484 274372 537536 274378
rect 537484 274314 537536 274320
rect 536380 272264 536432 272270
rect 536380 272206 536432 272212
rect 535736 268388 535788 268394
rect 535736 268330 535788 268336
rect 536380 268388 536432 268394
rect 536380 268330 536432 268336
rect 536392 264316 536420 268330
rect 537496 267306 537524 274314
rect 537680 269793 537708 274994
rect 539322 272504 539378 272513
rect 539322 272439 539378 272448
rect 538034 270056 538090 270065
rect 538034 269991 538090 270000
rect 537666 269784 537722 269793
rect 537666 269719 537722 269728
rect 537484 267300 537536 267306
rect 537484 267242 537536 267248
rect 537208 267028 537260 267034
rect 537208 266970 537260 266976
rect 537220 264316 537248 266970
rect 538048 264316 538076 269991
rect 539336 264330 539364 272439
rect 539520 269249 539548 275266
rect 539888 273970 539916 277780
rect 541084 274922 541112 277780
rect 542280 275330 542308 277780
rect 542268 275324 542320 275330
rect 542268 275266 542320 275272
rect 543280 275324 543332 275330
rect 543280 275266 543332 275272
rect 541992 275052 542044 275058
rect 541992 274994 542044 275000
rect 541072 274916 541124 274922
rect 541072 274858 541124 274864
rect 540888 274100 540940 274106
rect 540888 274042 540940 274048
rect 539876 273964 539928 273970
rect 539876 273906 539928 273912
rect 540518 269784 540574 269793
rect 540518 269719 540574 269728
rect 539506 269240 539562 269249
rect 539506 269175 539562 269184
rect 539692 267300 539744 267306
rect 539692 267242 539744 267248
rect 538890 264302 539364 264330
rect 539704 264316 539732 267242
rect 540532 264316 540560 269719
rect 540900 267306 540928 274042
rect 542004 273426 542032 274994
rect 542176 273964 542228 273970
rect 542176 273906 542228 273912
rect 541992 273420 542044 273426
rect 541992 273362 542044 273368
rect 541624 272264 541676 272270
rect 541624 272206 541676 272212
rect 541636 267714 541664 272206
rect 541624 267708 541676 267714
rect 541624 267650 541676 267656
rect 542188 267306 542216 273906
rect 540888 267300 540940 267306
rect 540888 267242 540940 267248
rect 541348 267300 541400 267306
rect 541348 267242 541400 267248
rect 542176 267300 542228 267306
rect 542176 267242 542228 267248
rect 542360 267300 542412 267306
rect 542360 267242 542412 267248
rect 541360 264316 541388 267242
rect 542372 267186 542400 267242
rect 542188 267158 542400 267186
rect 542188 264316 542216 267158
rect 543292 264330 543320 275266
rect 543476 272406 543504 277780
rect 544672 275194 544700 277780
rect 544660 275188 544712 275194
rect 544660 275130 544712 275136
rect 545120 274916 545172 274922
rect 545120 274858 545172 274864
rect 545132 273562 545160 274858
rect 545868 274786 545896 277780
rect 546512 277766 547078 277794
rect 545856 274780 545908 274786
rect 545856 274722 545908 274728
rect 545120 273556 545172 273562
rect 545120 273498 545172 273504
rect 543464 272400 543516 272406
rect 543464 272342 543516 272348
rect 546512 269686 546540 277766
rect 548168 273222 548196 277780
rect 549364 275058 549392 277780
rect 549916 277766 550574 277794
rect 549352 275052 549404 275058
rect 549352 274994 549404 275000
rect 548156 273216 548208 273222
rect 548156 273158 548208 273164
rect 546500 269680 546552 269686
rect 546500 269622 546552 269628
rect 549916 269550 549944 277766
rect 551284 274780 551336 274786
rect 551284 274722 551336 274728
rect 549904 269544 549956 269550
rect 549904 269486 549956 269492
rect 551296 267850 551324 274722
rect 551756 271425 551784 277780
rect 552572 275188 552624 275194
rect 552572 275130 552624 275136
rect 552584 273698 552612 275130
rect 552952 274922 552980 277780
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552940 274916 552992 274922
rect 552940 274858 552992 274864
rect 552572 273692 552624 273698
rect 552572 273634 552624 273640
rect 552664 273556 552716 273562
rect 552664 273498 552716 273504
rect 551742 271416 551798 271425
rect 551742 271351 551798 271360
rect 551284 267844 551336 267850
rect 551284 267786 551336 267792
rect 552676 266626 552704 273498
rect 552664 266620 552716 266626
rect 552664 266562 552716 266568
rect 553412 265402 553440 277766
rect 554792 266354 554820 277766
rect 556448 274514 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 274508 556488 274514
rect 556436 274450 556488 274456
rect 554780 266348 554832 266354
rect 554780 266290 554832 266296
rect 557552 265538 557580 277366
rect 558840 276690 558868 277780
rect 558828 276684 558880 276690
rect 558828 276626 558880 276632
rect 560036 275194 560064 277780
rect 560312 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 275188 560076 275194
rect 560024 275130 560076 275136
rect 559196 274916 559248 274922
rect 559196 274858 559248 274864
rect 559208 273834 559236 274858
rect 559564 274508 559616 274514
rect 559564 274450 559616 274456
rect 559196 273828 559248 273834
rect 559196 273770 559248 273776
rect 559576 266762 559604 274450
rect 560312 269414 560340 277766
rect 560300 269408 560352 269414
rect 560300 269350 560352 269356
rect 559564 266756 559616 266762
rect 559564 266698 559616 266704
rect 561692 266218 561720 277766
rect 563532 274242 563560 277780
rect 564452 277766 564742 277794
rect 563520 274236 563572 274242
rect 563520 274178 563572 274184
rect 563704 274236 563756 274242
rect 563704 274178 563756 274184
rect 563716 267345 563744 274178
rect 563702 267336 563758 267345
rect 563702 267271 563758 267280
rect 561680 266212 561732 266218
rect 561680 266154 561732 266160
rect 564452 266082 564480 277766
rect 565924 272134 565952 277780
rect 567120 277394 567148 277780
rect 567028 277366 567148 277394
rect 567304 277766 568330 277794
rect 568592 277766 569526 277794
rect 569972 277766 570722 277794
rect 567028 274922 567056 277366
rect 567016 274916 567068 274922
rect 567016 274858 567068 274864
rect 565912 272128 565964 272134
rect 565912 272070 565964 272076
rect 567304 268122 567332 277766
rect 568592 269521 568620 277766
rect 568578 269512 568634 269521
rect 568578 269447 568634 269456
rect 569972 268258 570000 277766
rect 571812 270910 571840 277780
rect 572732 277766 573022 277794
rect 571800 270904 571852 270910
rect 571800 270846 571852 270852
rect 569960 268252 570012 268258
rect 569960 268194 570012 268200
rect 567292 268116 567344 268122
rect 567292 268058 567344 268064
rect 564440 266076 564492 266082
rect 564440 266018 564492 266024
rect 572732 265946 572760 277766
rect 574204 274786 574232 277780
rect 574192 274780 574244 274786
rect 574192 274722 574244 274728
rect 575400 271046 575428 277780
rect 575388 271040 575440 271046
rect 575388 270982 575440 270988
rect 576124 271040 576176 271046
rect 576124 270982 576176 270988
rect 576136 267578 576164 270982
rect 576596 270774 576624 277780
rect 576872 277766 577806 277794
rect 576584 270768 576636 270774
rect 576584 270710 576636 270716
rect 576872 269074 576900 277766
rect 578896 271862 578924 277780
rect 580092 273562 580120 277780
rect 581012 277766 581302 277794
rect 580264 275120 580316 275126
rect 580264 275062 580316 275068
rect 580080 273556 580132 273562
rect 580080 273498 580132 273504
rect 580276 273086 580304 275062
rect 580264 273080 580316 273086
rect 580264 273022 580316 273028
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 269068 576912 269074
rect 576860 269010 576912 269016
rect 581012 268938 581040 277766
rect 582484 271726 582512 277780
rect 583680 275126 583708 277780
rect 583864 277766 584890 277794
rect 585612 277766 586086 277794
rect 583668 275120 583720 275126
rect 583668 275062 583720 275068
rect 582472 271720 582524 271726
rect 582472 271662 582524 271668
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 582288 268932 582340 268938
rect 582288 268874 582340 268880
rect 576124 267572 576176 267578
rect 576124 267514 576176 267520
rect 582300 267442 582328 268874
rect 583864 268802 583892 277766
rect 585612 271590 585640 277766
rect 587176 274514 587204 277780
rect 587912 277766 588386 277794
rect 587164 274508 587216 274514
rect 587164 274450 587216 274456
rect 585600 271584 585652 271590
rect 585600 271526 585652 271532
rect 585784 271584 585836 271590
rect 585784 271526 585836 271532
rect 583852 268796 583904 268802
rect 583852 268738 583904 268744
rect 582288 267436 582340 267442
rect 582288 267378 582340 267384
rect 585796 267073 585824 271526
rect 587912 268666 587940 277766
rect 589568 271454 589596 277780
rect 590764 275874 590792 277780
rect 591132 277766 591974 277794
rect 590752 275868 590804 275874
rect 590752 275810 590804 275816
rect 589556 271448 589608 271454
rect 589556 271390 589608 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 591132 268433 591160 277766
rect 592684 271448 592736 271454
rect 592684 271390 592736 271396
rect 591118 268424 591174 268433
rect 591118 268359 591174 268368
rect 585782 267064 585838 267073
rect 585782 266999 585838 267008
rect 592696 266490 592724 271390
rect 593156 271153 593184 277780
rect 593142 271144 593198 271153
rect 593142 271079 593198 271088
rect 594352 271046 594380 277780
rect 595456 274650 595484 277780
rect 595444 274644 595496 274650
rect 595444 274586 595496 274592
rect 596652 271318 596680 277780
rect 597572 277766 597862 277794
rect 596640 271312 596692 271318
rect 596640 271254 596692 271260
rect 596824 271312 596876 271318
rect 596824 271254 596876 271260
rect 594340 271040 594392 271046
rect 594340 270982 594392 270988
rect 596836 267170 596864 271254
rect 597572 270502 597600 277766
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597560 270496 597612 270502
rect 597560 270438 597612 270444
rect 598952 268530 598980 277366
rect 600240 271182 600268 277780
rect 600608 277766 601450 277794
rect 600228 271176 600280 271182
rect 600228 271118 600280 271124
rect 600608 268938 600636 277766
rect 602540 274145 602568 277780
rect 602526 274136 602582 274145
rect 602526 274071 602582 274080
rect 603736 272270 603764 277780
rect 604932 275738 604960 277780
rect 605852 277766 606142 277794
rect 604920 275732 604972 275738
rect 604920 275674 604972 275680
rect 605104 275732 605156 275738
rect 605104 275674 605156 275680
rect 603724 272264 603776 272270
rect 603724 272206 603776 272212
rect 605116 270366 605144 275674
rect 605104 270360 605156 270366
rect 605104 270302 605156 270308
rect 600596 268932 600648 268938
rect 600596 268874 600648 268880
rect 598940 268524 598992 268530
rect 598940 268466 598992 268472
rect 596824 267164 596876 267170
rect 596824 267106 596876 267112
rect 592684 266484 592736 266490
rect 592684 266426 592736 266432
rect 572720 265940 572772 265946
rect 572720 265882 572772 265888
rect 605852 265810 605880 277766
rect 607324 276010 607352 277780
rect 607312 276004 607364 276010
rect 607312 275946 607364 275952
rect 608520 271590 608548 277780
rect 608704 277766 609730 277794
rect 608508 271584 608560 271590
rect 608508 271526 608560 271532
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 608704 265674 608732 277766
rect 610820 272950 610848 277780
rect 612016 274242 612044 277780
rect 613212 274378 613240 277780
rect 613200 274372 613252 274378
rect 613200 274314 613252 274320
rect 612004 274236 612056 274242
rect 612004 274178 612056 274184
rect 614408 273057 614436 277780
rect 615604 277394 615632 277780
rect 615512 277366 615632 277394
rect 614394 273048 614450 273057
rect 614394 272983 614450 272992
rect 610808 272944 610860 272950
rect 610808 272886 610860 272892
rect 615512 266898 615540 277366
rect 616800 275738 616828 277780
rect 616788 275732 616840 275738
rect 616788 275674 616840 275680
rect 617996 272814 618024 277780
rect 619100 275466 619128 277780
rect 619652 277766 620310 277794
rect 619088 275460 619140 275466
rect 619088 275402 619140 275408
rect 619180 274712 619232 274718
rect 619180 274654 619232 274660
rect 617984 272808 618036 272814
rect 617984 272750 618036 272756
rect 619192 270230 619220 274654
rect 619180 270224 619232 270230
rect 619180 270166 619232 270172
rect 619652 270094 619680 277766
rect 621492 272678 621520 277780
rect 621480 272672 621532 272678
rect 621480 272614 621532 272620
rect 622688 271454 622716 277780
rect 623884 274718 623912 277780
rect 624712 277766 625094 277794
rect 623872 274712 623924 274718
rect 623872 274654 623924 274660
rect 624712 272542 624740 277766
rect 626184 275602 626212 277780
rect 626644 277766 627394 277794
rect 627932 277766 628590 277794
rect 626172 275596 626224 275602
rect 626172 275538 626224 275544
rect 626448 275460 626500 275466
rect 626448 275402 626500 275408
rect 626460 274106 626488 275402
rect 626448 274100 626500 274106
rect 626448 274042 626500 274048
rect 624700 272536 624752 272542
rect 624700 272478 624752 272484
rect 622676 271448 622728 271454
rect 622676 271390 622728 271396
rect 623044 271176 623096 271182
rect 623044 271118 623096 271124
rect 619640 270088 619692 270094
rect 619640 270030 619692 270036
rect 623056 267306 623084 271118
rect 626644 270337 626672 277766
rect 626630 270328 626686 270337
rect 626630 270263 626686 270272
rect 627932 269958 627960 277766
rect 629772 271318 629800 277780
rect 630968 273873 630996 277780
rect 630954 273864 631010 273873
rect 630954 273799 631010 273808
rect 632164 272785 632192 277780
rect 633360 275233 633388 277780
rect 633544 277766 634478 277794
rect 634832 277766 635674 277794
rect 636212 277766 636870 277794
rect 637592 277766 638066 277794
rect 633346 275224 633402 275233
rect 633346 275159 633402 275168
rect 632150 272776 632206 272785
rect 632150 272711 632206 272720
rect 629760 271312 629812 271318
rect 629760 271254 629812 271260
rect 627920 269952 627972 269958
rect 627920 269894 627972 269900
rect 633544 269822 633572 277766
rect 633532 269816 633584 269822
rect 633532 269758 633584 269764
rect 634832 268394 634860 277766
rect 634820 268388 634872 268394
rect 634820 268330 634872 268336
rect 623044 267300 623096 267306
rect 623044 267242 623096 267248
rect 636212 267034 636240 277766
rect 637592 270065 637620 277766
rect 639248 272513 639276 277780
rect 640444 275466 640472 277780
rect 640720 277766 641654 277794
rect 640432 275460 640484 275466
rect 640432 275402 640484 275408
rect 639234 272504 639290 272513
rect 639234 272439 639290 272448
rect 637578 270056 637634 270065
rect 637578 269991 637634 270000
rect 640720 269793 640748 277766
rect 642744 273970 642772 277780
rect 642732 273964 642784 273970
rect 642732 273906 642784 273912
rect 643940 271182 643968 277780
rect 645136 275330 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645124 275324 645176 275330
rect 645124 275266 645176 275272
rect 643928 271176 643980 271182
rect 643928 271118 643980 271124
rect 640706 269784 640762 269793
rect 640706 269719 640762 269728
rect 636200 267028 636252 267034
rect 636200 266970 636252 266976
rect 615500 266892 615552 266898
rect 615500 266834 615552 266840
rect 608692 265668 608744 265674
rect 608692 265610 608744 265616
rect 557540 265532 557592 265538
rect 557540 265474 557592 265480
rect 553400 265396 553452 265402
rect 553400 265338 553452 265344
rect 543030 264302 543320 264330
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 645872 261526 645900 277766
rect 571984 261520 572036 261526
rect 571984 261462 572036 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 563704 259480 563756 259486
rect 563704 259422 563756 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 560944 256760 560996 256766
rect 560944 256702 560996 256708
rect 553766 255640 553822 255649
rect 553766 255575 553822 255584
rect 553780 255338 553808 255575
rect 553768 255332 553820 255338
rect 553768 255274 553820 255280
rect 556804 255332 556856 255338
rect 556804 255274 556856 255280
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 553490 251288 553546 251297
rect 553490 251223 553492 251232
rect 553544 251223 553546 251232
rect 555424 251252 555476 251258
rect 553492 251194 553544 251200
rect 555424 251194 555476 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 124128 230784 124180 230790
rect 124128 230726 124180 230732
rect 97908 230648 97960 230654
rect 97908 230590 97960 230596
rect 91008 230512 91060 230518
rect 91008 230454 91060 230460
rect 71042 230072 71098 230081
rect 71042 230007 71098 230016
rect 86224 230036 86276 230042
rect 65522 229800 65578 229809
rect 65522 229735 65578 229744
rect 64144 228540 64196 228546
rect 64144 228482 64196 228488
rect 62946 224496 63002 224505
rect 62946 224431 63002 224440
rect 63408 224256 63460 224262
rect 63408 224198 63460 224204
rect 63132 218680 63184 218686
rect 63132 218622 63184 218628
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 62028 218068 62080 218074
rect 62028 218010 62080 218016
rect 62304 218068 62356 218074
rect 62304 218010 62356 218016
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218010
rect 63144 217138 63172 218622
rect 63420 218074 63448 224198
rect 63960 219292 64012 219298
rect 63960 219234 64012 219240
rect 63408 218068 63460 218074
rect 63408 218010 63460 218016
rect 63972 217138 64000 219234
rect 64156 218210 64184 228482
rect 64786 222864 64842 222873
rect 64786 222799 64842 222808
rect 64144 218204 64196 218210
rect 64144 218146 64196 218152
rect 64800 217274 64828 222799
rect 65536 219298 65564 229735
rect 68284 227180 68336 227186
rect 68284 227122 68336 227128
rect 66902 224496 66958 224505
rect 66902 224431 66958 224440
rect 66444 220652 66496 220658
rect 66444 220594 66496 220600
rect 65524 219292 65576 219298
rect 65524 219234 65576 219240
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 64754 217246 64828 217274
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217274 66484 220594
rect 66916 218074 66944 224431
rect 68296 218686 68324 227122
rect 70308 225888 70360 225894
rect 70308 225830 70360 225836
rect 68928 222896 68980 222902
rect 68928 222838 68980 222844
rect 68284 218680 68336 218686
rect 68284 218622 68336 218628
rect 68744 218340 68796 218346
rect 68744 218282 68796 218288
rect 67272 218204 67324 218210
rect 67272 218146 67324 218152
rect 66904 218068 66956 218074
rect 66904 218010 66956 218016
rect 65582 217110 65656 217138
rect 66410 217246 66484 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217246
rect 67284 217138 67312 218146
rect 68100 218068 68152 218074
rect 68100 218010 68152 218016
rect 68112 217138 68140 218010
rect 68756 217274 68784 218282
rect 68940 218074 68968 222838
rect 70320 218074 70348 225830
rect 70584 219428 70636 219434
rect 70584 219370 70636 219376
rect 68928 218068 68980 218074
rect 68928 218010 68980 218016
rect 69756 218068 69808 218074
rect 69756 218010 69808 218016
rect 70308 218068 70360 218074
rect 70308 218010 70360 218016
rect 68756 217246 68922 217274
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69768 217138 69796 218010
rect 70596 217138 70624 219370
rect 71056 218210 71084 230007
rect 86224 229978 86276 229984
rect 73710 228304 73766 228313
rect 73710 228239 73766 228248
rect 72422 224768 72478 224777
rect 72422 224703 72478 224712
rect 71410 223136 71466 223145
rect 71410 223071 71466 223080
rect 71044 218204 71096 218210
rect 71044 218146 71096 218152
rect 71424 217274 71452 223071
rect 72436 218346 72464 224703
rect 73068 220108 73120 220114
rect 73068 220050 73120 220056
rect 72424 218340 72476 218346
rect 72424 218282 72476 218288
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 69722 217110 69796 217138
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 69722 216988 69750 217110
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220050
rect 73724 218074 73752 228239
rect 81348 227316 81400 227322
rect 81348 227258 81400 227264
rect 79966 226944 80022 226953
rect 79966 226879 80022 226888
rect 76564 224392 76616 224398
rect 76564 224334 76616 224340
rect 75828 223032 75880 223038
rect 75828 222974 75880 222980
rect 73896 221604 73948 221610
rect 73896 221546 73948 221552
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221546
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 222974
rect 76380 220380 76432 220386
rect 76380 220322 76432 220328
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220322
rect 76576 218210 76604 224334
rect 78588 223304 78640 223310
rect 78588 223246 78640 223252
rect 77206 218648 77262 218657
rect 77206 218583 77262 218592
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218583
rect 78600 218074 78628 223246
rect 79692 220244 79744 220250
rect 79692 220186 79744 220192
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220186
rect 79980 218074 80008 226879
rect 81164 223168 81216 223174
rect 81164 223110 81216 223116
rect 81176 219434 81204 223110
rect 81176 219406 81296 219434
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80520 218068 80572 218074
rect 80520 218010 80572 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80532 217138 80560 218010
rect 81268 217274 81296 219406
rect 81360 218090 81388 227258
rect 84108 226024 84160 226030
rect 84108 225966 84160 225972
rect 82726 225584 82782 225593
rect 82726 225519 82782 225528
rect 81360 218074 81480 218090
rect 82740 218074 82768 225519
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 81360 218068 81492 218074
rect 81360 218062 81440 218068
rect 81440 218010 81492 218016
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 82728 218068 82780 218074
rect 82728 218010 82780 218016
rect 83004 218068 83056 218074
rect 83004 218010 83056 218016
rect 81268 217246 81342 217274
rect 80486 217110 80560 217138
rect 80486 216988 80514 217110
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217138 83044 218010
rect 83844 217138 83872 218826
rect 84120 218074 84148 225966
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 84660 221468 84712 221474
rect 84660 221410 84712 221416
rect 84108 218068 84160 218074
rect 84108 218010 84160 218016
rect 84672 217274 84700 221410
rect 85500 217274 85528 224470
rect 86236 221610 86264 229978
rect 89626 227216 89682 227225
rect 89626 227151 89682 227160
rect 89442 225856 89498 225865
rect 89442 225791 89498 225800
rect 87972 223576 88024 223582
rect 87972 223518 88024 223524
rect 86224 221604 86276 221610
rect 86224 221546 86276 221552
rect 86316 220516 86368 220522
rect 86316 220458 86368 220464
rect 86328 217274 86356 220458
rect 87144 219156 87196 219162
rect 87144 219098 87196 219104
rect 87156 217274 87184 219098
rect 87984 217274 88012 223518
rect 89456 218074 89484 225791
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 82142 217110 82216 217138
rect 82970 217110 83044 217138
rect 83798 217110 83872 217138
rect 84626 217246 84700 217274
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 87110 217246 87184 217274
rect 87938 217246 88012 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217110
rect 83798 216988 83826 217110
rect 84626 216988 84654 217246
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87110 216988 87138 217246
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227151
rect 91020 218074 91048 230454
rect 95240 229628 95292 229634
rect 95240 229570 95292 229576
rect 94504 229492 94556 229498
rect 94504 229434 94556 229440
rect 94516 229094 94544 229434
rect 94424 229066 94544 229094
rect 93768 228676 93820 228682
rect 93768 228618 93820 228624
rect 92110 223408 92166 223417
rect 92110 223343 92166 223352
rect 91284 221604 91336 221610
rect 91284 221546 91336 221552
rect 90456 218068 90508 218074
rect 90456 218010 90508 218016
rect 91008 218068 91060 218074
rect 91008 218010 91060 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 218010
rect 91296 217274 91324 221546
rect 92124 217274 92152 223343
rect 93780 218754 93808 228618
rect 94424 221746 94452 229066
rect 95252 227322 95280 229570
rect 95240 227316 95292 227322
rect 95240 227258 95292 227264
rect 96252 227316 96304 227322
rect 96252 227258 96304 227264
rect 94412 221740 94464 221746
rect 94412 221682 94464 221688
rect 94596 221740 94648 221746
rect 94596 221682 94648 221688
rect 92940 218748 92992 218754
rect 92940 218690 92992 218696
rect 93768 218748 93820 218754
rect 93768 218690 93820 218696
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218690
rect 93768 218612 93820 218618
rect 93768 218554 93820 218560
rect 93780 217138 93808 218554
rect 94608 217308 94636 221682
rect 95422 221504 95478 221513
rect 95422 221439 95478 221448
rect 95436 217308 95464 221439
rect 96264 217308 96292 227258
rect 97722 221776 97778 221785
rect 97722 221711 97778 221720
rect 97736 219434 97764 221711
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217280 94636 217308
rect 95390 217280 95464 217308
rect 96218 217280 96292 217308
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217280
rect 95390 216988 95418 217280
rect 96218 216988 96246 217280
rect 97092 217138 97120 218010
rect 97828 217308 97856 219406
rect 97920 218090 97948 230590
rect 117228 229900 117280 229906
rect 117228 229842 117280 229848
rect 110328 229764 110380 229770
rect 110328 229706 110380 229712
rect 106924 229220 106976 229226
rect 106924 229162 106976 229168
rect 100668 228948 100720 228954
rect 100668 228890 100720 228896
rect 99288 226160 99340 226166
rect 99288 226102 99340 226108
rect 97920 218074 98040 218090
rect 99300 218074 99328 226102
rect 100392 218748 100444 218754
rect 100392 218690 100444 218696
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217280 97902 217308
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217280
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218690
rect 100680 218074 100708 228890
rect 106188 228812 106240 228818
rect 106188 228754 106240 228760
rect 103428 227452 103480 227458
rect 103428 227394 103480 227400
rect 102048 223440 102100 223446
rect 102048 223382 102100 223388
rect 101220 221876 101272 221882
rect 101220 221818 101272 221824
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217308 101260 221818
rect 102060 217308 102088 223382
rect 103440 218074 103468 227394
rect 106004 224664 106056 224670
rect 106004 224606 106056 224612
rect 104532 222012 104584 222018
rect 104532 221954 104584 221960
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217280 101260 217308
rect 102014 217280 102088 217308
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217280
rect 102014 216988 102042 217280
rect 102888 217138 102916 218010
rect 104544 217274 104572 221954
rect 106016 218074 106044 224606
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 103658 217252 103710 217258
rect 103658 217194 103710 217200
rect 104498 217246 104572 217274
rect 102842 217110 102916 217138
rect 102842 216988 102870 217110
rect 103670 216988 103698 217194
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 228754
rect 106936 219162 106964 229162
rect 110144 227588 110196 227594
rect 110144 227530 110196 227536
rect 108670 222048 108726 222057
rect 108670 221983 108726 221992
rect 107844 220788 107896 220794
rect 107844 220730 107896 220736
rect 106924 219156 106976 219162
rect 106924 219098 106976 219104
rect 107108 219156 107160 219162
rect 107108 219098 107160 219104
rect 107120 217274 107148 219098
rect 107856 217274 107884 220730
rect 108684 217274 108712 221983
rect 110156 218074 110184 227530
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 106982 217246 107148 217274
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 106982 216988 107010 217246
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217274 110368 229706
rect 112994 228576 113050 228585
rect 112994 228511 113050 228520
rect 112812 224800 112864 224806
rect 112812 224742 112864 224748
rect 111156 222148 111208 222154
rect 111156 222090 111208 222096
rect 111168 217274 111196 222090
rect 112824 218074 112852 224742
rect 111984 218068 112036 218074
rect 111984 218010 112036 218016
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 109466 217110 109540 217138
rect 110294 217246 110368 217274
rect 111122 217246 111196 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 216988 111150 217246
rect 111996 217138 112024 218010
rect 113008 217274 113036 228511
rect 116952 227724 117004 227730
rect 116952 227666 117004 227672
rect 115848 224120 115900 224126
rect 115848 224062 115900 224068
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113640 219292 113692 219298
rect 113640 219234 113692 219240
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 219234
rect 114480 217274 114508 219914
rect 115860 218074 115888 224062
rect 116964 218074 116992 227666
rect 117240 219434 117268 229842
rect 119988 229084 120040 229090
rect 119988 229026 120040 229032
rect 118608 224936 118660 224942
rect 118608 224878 118660 224884
rect 117778 220144 117834 220153
rect 117778 220079 117834 220088
rect 117148 219406 117268 219434
rect 115296 218068 115348 218074
rect 115296 218010 115348 218016
rect 115848 218068 115900 218074
rect 115848 218010 115900 218016
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 116952 218068 117004 218074
rect 116952 218010 117004 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 218010
rect 116136 217138 116164 218010
rect 117148 217274 117176 219406
rect 117792 217274 117820 220079
rect 118620 217274 118648 224878
rect 120000 218074 120028 229026
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 223984 122616 223990
rect 122564 223926 122616 223932
rect 121092 221332 121144 221338
rect 121092 221274 121144 221280
rect 120264 218340 120316 218346
rect 120264 218282 120316 218288
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217246 117176 217274
rect 117746 217246 117820 217274
rect 118574 217246 118648 217274
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217246
rect 117746 216988 117774 217246
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217274 120304 218282
rect 121104 217274 121132 221274
rect 122576 218074 122604 223926
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217246 120304 217274
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217246
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 226850
rect 124140 218074 124168 230726
rect 133788 230308 133840 230314
rect 133788 230250 133840 230256
rect 126888 230172 126940 230178
rect 126888 230114 126940 230120
rect 126704 228268 126756 228274
rect 126704 228210 126756 228216
rect 125230 226128 125286 226137
rect 125230 226063 125286 226072
rect 124402 220416 124458 220425
rect 124402 220351 124458 220360
rect 123576 218068 123628 218074
rect 123576 218010 123628 218016
rect 124128 218068 124180 218074
rect 124128 218010 124180 218016
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 218010
rect 124416 217274 124444 220351
rect 125244 217274 125272 226063
rect 126716 218074 126744 228210
rect 126060 218068 126112 218074
rect 126060 218010 126112 218016
rect 126704 218068 126756 218074
rect 126704 218010 126756 218016
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218010
rect 126900 217274 126928 230114
rect 133512 228132 133564 228138
rect 133512 228074 133564 228080
rect 129372 226772 129424 226778
rect 129372 226714 129424 226720
rect 127716 219836 127768 219842
rect 127716 219778 127768 219784
rect 127728 217274 127756 219778
rect 128544 217456 128596 217462
rect 128544 217398 128596 217404
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 127682 217246 127756 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127682 216988 127710 217246
rect 128556 217138 128584 217398
rect 129384 217274 129412 226714
rect 132408 225480 132460 225486
rect 132408 225422 132460 225428
rect 131028 222760 131080 222766
rect 131028 222702 131080 222708
rect 130200 218204 130252 218210
rect 130200 218146 130252 218152
rect 128510 217110 128584 217138
rect 129338 217246 129412 217274
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218146
rect 131040 217274 131068 222702
rect 132420 218074 132448 225422
rect 133524 218074 133552 228074
rect 133800 219434 133828 230250
rect 137284 229356 137336 229362
rect 137284 229298 137336 229304
rect 136546 227488 136602 227497
rect 136546 227423 136602 227432
rect 135168 226296 135220 226302
rect 135168 226238 135220 226244
rect 134984 222488 135036 222494
rect 134984 222430 135036 222436
rect 133708 219406 133828 219434
rect 131856 218068 131908 218074
rect 131856 218010 131908 218016
rect 132408 218068 132460 218074
rect 132408 218010 132460 218016
rect 132684 218068 132736 218074
rect 132684 218010 132736 218016
rect 133512 218068 133564 218074
rect 133512 218010 133564 218016
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 218010
rect 132696 217138 132724 218010
rect 133708 217274 133736 219406
rect 134996 218074 135024 222430
rect 134340 218068 134392 218074
rect 134340 218010 134392 218016
rect 134984 218068 135036 218074
rect 134984 218010 135036 218016
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134352 217138 134380 218010
rect 135180 217274 135208 226238
rect 136560 218074 136588 227423
rect 137296 219026 137324 229298
rect 141160 228410 141188 231676
rect 141148 228404 141200 228410
rect 141148 228346 141200 228352
rect 139308 227996 139360 228002
rect 139308 227938 139360 227944
rect 139124 225344 139176 225350
rect 139124 225286 139176 225292
rect 137652 219700 137704 219706
rect 137652 219642 137704 219648
rect 137284 219020 137336 219026
rect 137284 218962 137336 218968
rect 136824 218340 136876 218346
rect 136824 218282 136876 218288
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 136548 218068 136600 218074
rect 136548 218010 136600 218016
rect 134306 217110 134380 217138
rect 135134 217246 135208 217274
rect 134306 216988 134334 217110
rect 135134 216988 135162 217246
rect 136008 217138 136036 218010
rect 136836 217138 136864 218282
rect 137664 217274 137692 219642
rect 139136 218074 139164 225286
rect 138480 218068 138532 218074
rect 138480 218010 138532 218016
rect 139124 218068 139176 218074
rect 139124 218010 139176 218016
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 218010
rect 139320 217274 139348 227938
rect 141804 225758 141832 231676
rect 142448 227050 142476 231676
rect 143092 228546 143120 231676
rect 143736 229362 143764 231676
rect 143724 229356 143776 229362
rect 143724 229298 143776 229304
rect 144184 229356 144236 229362
rect 144184 229298 144236 229304
rect 144196 229094 144224 229298
rect 144104 229066 144224 229094
rect 143080 228540 143132 228546
rect 143080 228482 143132 228488
rect 143448 227860 143500 227866
rect 143448 227802 143500 227808
rect 142436 227044 142488 227050
rect 142436 226986 142488 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141792 225752 141844 225758
rect 141792 225694 141844 225700
rect 141976 225752 142028 225758
rect 141976 225694 142028 225700
rect 139952 223848 140004 223854
rect 139952 223790 140004 223796
rect 139964 218618 139992 223790
rect 140964 221060 141016 221066
rect 140964 221002 141016 221008
rect 139952 218612 140004 218618
rect 139952 218554 140004 218560
rect 140136 218612 140188 218618
rect 140136 218554 140188 218560
rect 139492 218340 139544 218346
rect 139492 218282 139544 218288
rect 139504 218074 139532 218282
rect 139492 218068 139544 218074
rect 139492 218010 139544 218016
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218554
rect 140976 217274 141004 221002
rect 141988 219434 142016 225694
rect 141804 219406 142016 219434
rect 141804 217274 141832 219406
rect 143276 218210 143304 226986
rect 142620 218204 142672 218210
rect 142620 218146 142672 218152
rect 143264 218204 143316 218210
rect 143264 218146 143316 218152
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218146
rect 143460 217274 143488 227802
rect 144104 220658 144132 229066
rect 144380 225622 144408 231676
rect 144368 225616 144420 225622
rect 144368 225558 144420 225564
rect 145024 224233 145052 231676
rect 145668 229498 145696 231676
rect 146312 230330 146340 231676
rect 146680 231662 146970 231690
rect 146312 230302 146432 230330
rect 145656 229492 145708 229498
rect 145656 229434 145708 229440
rect 146208 229492 146260 229498
rect 146208 229434 146260 229440
rect 145932 228404 145984 228410
rect 145932 228346 145984 228352
rect 145010 224224 145066 224233
rect 145010 224159 145066 224168
rect 144092 220652 144144 220658
rect 144092 220594 144144 220600
rect 144276 220652 144328 220658
rect 144276 220594 144328 220600
rect 143724 219020 143776 219026
rect 143724 218962 143776 218968
rect 143736 218618 143764 218962
rect 143724 218612 143776 218618
rect 143724 218554 143776 218560
rect 144288 217274 144316 220594
rect 145104 218204 145156 218210
rect 145104 218146 145156 218152
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 144242 217246 144316 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144242 216988 144270 217246
rect 145116 217138 145144 218146
rect 145944 217274 145972 228346
rect 146220 227866 146248 229434
rect 146208 227860 146260 227866
rect 146208 227802 146260 227808
rect 146404 227186 146432 230302
rect 146392 227180 146444 227186
rect 146392 227122 146444 227128
rect 146680 222873 146708 231662
rect 147600 224262 147628 231676
rect 148244 229809 148272 231676
rect 148230 229800 148286 229809
rect 148230 229735 148286 229744
rect 148888 229362 148916 231676
rect 148876 229356 148928 229362
rect 148876 229298 148928 229304
rect 147588 224256 147640 224262
rect 146942 224224 146998 224233
rect 147588 224198 147640 224204
rect 146942 224159 146998 224168
rect 146666 222864 146722 222873
rect 146666 222799 146722 222808
rect 146116 222624 146168 222630
rect 146116 222566 146168 222572
rect 146128 218210 146156 222566
rect 146956 218754 146984 224159
rect 149532 222902 149560 231676
rect 149808 231662 150190 231690
rect 149808 224505 149836 231662
rect 150820 230081 150848 231676
rect 150806 230072 150862 230081
rect 150806 230007 150862 230016
rect 150072 229356 150124 229362
rect 150072 229298 150124 229304
rect 149794 224496 149850 224505
rect 149794 224431 149850 224440
rect 149520 222896 149572 222902
rect 149520 222838 149572 222844
rect 148416 221196 148468 221202
rect 148416 221138 148468 221144
rect 147586 220688 147642 220697
rect 147586 220623 147642 220632
rect 146944 218748 146996 218754
rect 146944 218690 146996 218696
rect 146760 218612 146812 218618
rect 146760 218554 146812 218560
rect 146116 218204 146168 218210
rect 146116 218146 146168 218152
rect 146772 217274 146800 218554
rect 147600 217274 147628 220623
rect 145070 217110 145144 217138
rect 145898 217246 145972 217274
rect 146726 217246 146800 217274
rect 147554 217246 147628 217274
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146726 216988 146754 217246
rect 147554 216988 147582 217246
rect 148428 217138 148456 221138
rect 149060 219428 149112 219434
rect 149060 219370 149112 219376
rect 149244 219428 149296 219434
rect 149244 219370 149296 219376
rect 149072 218754 149100 219370
rect 149060 218748 149112 218754
rect 149060 218690 149112 218696
rect 149256 217138 149284 219370
rect 150084 217274 150112 229298
rect 150256 226636 150308 226642
rect 150256 226578 150308 226584
rect 150268 219434 150296 226578
rect 151464 225894 151492 231676
rect 151452 225888 151504 225894
rect 151452 225830 151504 225836
rect 151728 224256 151780 224262
rect 151728 224198 151780 224204
rect 150898 222864 150954 222873
rect 150898 222799 150954 222808
rect 150256 219428 150308 219434
rect 150256 219370 150308 219376
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150112 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150912 217138 150940 222799
rect 151740 217138 151768 224198
rect 152108 223145 152136 231676
rect 152752 224777 152780 231676
rect 153410 231662 153608 231690
rect 153108 228540 153160 228546
rect 153108 228482 153160 228488
rect 152924 227180 152976 227186
rect 152924 227122 152976 227128
rect 152936 226642 152964 227122
rect 152924 226636 152976 226642
rect 152924 226578 152976 226584
rect 152738 224768 152794 224777
rect 152738 224703 152794 224712
rect 152094 223136 152150 223145
rect 152094 223071 152150 223080
rect 153120 219434 153148 228482
rect 153580 224954 153608 231662
rect 153304 224926 153608 224954
rect 153764 231662 154054 231690
rect 152556 219428 152608 219434
rect 152556 219370 152608 219376
rect 153108 219428 153160 219434
rect 153108 219370 153160 219376
rect 152568 217138 152596 219370
rect 153304 218906 153332 224926
rect 153764 220114 153792 231662
rect 154684 223038 154712 231676
rect 155328 228313 155356 231676
rect 155972 230042 156000 231676
rect 156156 231662 156630 231690
rect 155960 230036 156012 230042
rect 155960 229978 156012 229984
rect 155314 228304 155370 228313
rect 155314 228239 155370 228248
rect 155868 225616 155920 225622
rect 155868 225558 155920 225564
rect 155684 225208 155736 225214
rect 155684 225150 155736 225156
rect 155696 224954 155724 225150
rect 155696 224926 155816 224954
rect 154672 223032 154724 223038
rect 154672 222974 154724 222980
rect 154212 222896 154264 222902
rect 154212 222838 154264 222844
rect 153752 220108 153804 220114
rect 153752 220050 153804 220056
rect 153212 218878 153332 218906
rect 153212 218754 153240 218878
rect 153200 218748 153252 218754
rect 153200 218690 153252 218696
rect 153384 218748 153436 218754
rect 153384 218690 153436 218696
rect 153396 217138 153424 218690
rect 154224 217138 154252 222838
rect 155040 219428 155092 219434
rect 155040 219370 155092 219376
rect 155052 217138 155080 219370
rect 155788 217274 155816 224926
rect 155880 219434 155908 225558
rect 156156 220386 156184 231662
rect 157064 230036 157116 230042
rect 157064 229978 157116 229984
rect 157076 224954 157104 229978
rect 156708 224926 157104 224954
rect 156144 220380 156196 220386
rect 156144 220322 156196 220328
rect 155880 219428 156012 219434
rect 155880 219406 155960 219428
rect 155960 219370 156012 219376
rect 156144 219428 156196 219434
rect 156144 219370 156196 219376
rect 156156 218890 156184 219370
rect 156144 218884 156196 218890
rect 156144 218826 156196 218832
rect 156708 217274 156736 224926
rect 157260 223310 157288 231676
rect 157904 224398 157932 231676
rect 158088 231662 158562 231690
rect 158916 231662 159206 231690
rect 157892 224392 157944 224398
rect 157892 224334 157944 224340
rect 157248 223304 157300 223310
rect 157248 223246 157300 223252
rect 157524 220108 157576 220114
rect 157524 220050 157576 220056
rect 157536 217274 157564 220050
rect 158088 219434 158116 231662
rect 158352 225888 158404 225894
rect 158352 225830 158404 225836
rect 157720 219406 158116 219434
rect 157720 218657 157748 219406
rect 157706 218648 157762 218657
rect 157706 218583 157762 218592
rect 158364 217274 158392 225830
rect 158916 220250 158944 231662
rect 159364 223304 159416 223310
rect 159364 223246 159416 223252
rect 158904 220244 158956 220250
rect 158904 220186 158956 220192
rect 159376 219162 159404 223246
rect 159836 223174 159864 231676
rect 160480 226953 160508 231676
rect 161124 229634 161152 231676
rect 161112 229628 161164 229634
rect 161112 229570 161164 229576
rect 161296 229628 161348 229634
rect 161296 229570 161348 229576
rect 160466 226944 160522 226953
rect 160466 226879 160522 226888
rect 160008 226636 160060 226642
rect 160008 226578 160060 226584
rect 159824 223168 159876 223174
rect 159824 223110 159876 223116
rect 159364 219156 159416 219162
rect 159364 219098 159416 219104
rect 159822 218648 159878 218657
rect 159822 218583 159878 218592
rect 159180 218204 159232 218210
rect 159180 218146 159232 218152
rect 155788 217246 155862 217274
rect 150866 217110 150940 217138
rect 151694 217110 151768 217138
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217110 154252 217138
rect 155006 217110 155080 217138
rect 150866 216988 150894 217110
rect 151694 216988 151722 217110
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217110
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156662 217246 156736 217274
rect 157490 217246 157564 217274
rect 158318 217246 158392 217274
rect 156662 216988 156690 217246
rect 157490 216988 157518 217246
rect 158318 216988 158346 217246
rect 159192 217138 159220 218146
rect 159836 217274 159864 218583
rect 160020 218210 160048 226578
rect 161308 219434 161336 229570
rect 161768 226030 161796 231676
rect 162044 231662 162426 231690
rect 162044 229094 162072 231662
rect 161952 229066 162072 229094
rect 161756 226024 161808 226030
rect 161756 225966 161808 225972
rect 161952 221898 161980 229066
rect 163056 225593 163084 231676
rect 163332 231662 163714 231690
rect 163042 225584 163098 225593
rect 163042 225519 163098 225528
rect 161584 221870 161980 221898
rect 161584 221626 161612 221870
rect 161492 221598 161612 221626
rect 161492 221474 161520 221598
rect 161480 221468 161532 221474
rect 161480 221410 161532 221416
rect 161664 221468 161716 221474
rect 161664 221410 161716 221416
rect 160756 219406 161336 219434
rect 160756 219026 160784 219406
rect 160744 219020 160796 219026
rect 160744 218962 160796 218968
rect 160008 218204 160060 218210
rect 160008 218146 160060 218152
rect 160836 218204 160888 218210
rect 160836 218146 160888 218152
rect 159836 217246 160002 217274
rect 159146 217110 159220 217138
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160848 217138 160876 218146
rect 161676 217274 161704 221410
rect 161940 220244 161992 220250
rect 161940 220186 161992 220192
rect 161952 218210 161980 220186
rect 163332 219434 163360 231662
rect 164056 223032 164108 223038
rect 164056 222974 164108 222980
rect 162860 219428 163360 219434
rect 162912 219406 163360 219428
rect 162860 219370 162912 219376
rect 163320 219156 163372 219162
rect 163320 219098 163372 219104
rect 162492 219020 162544 219026
rect 162492 218962 162544 218968
rect 161940 218204 161992 218210
rect 161940 218146 161992 218152
rect 160802 217110 160876 217138
rect 161630 217246 161704 217274
rect 160802 216988 160830 217110
rect 161630 216988 161658 217246
rect 162504 217138 162532 218962
rect 163332 217138 163360 219098
rect 164068 217274 164096 222974
rect 164344 220522 164372 231676
rect 164988 223582 165016 231676
rect 165632 224534 165660 231676
rect 166276 229226 166304 231676
rect 166264 229220 166316 229226
rect 166264 229162 166316 229168
rect 166920 227225 166948 231676
rect 167104 231662 167578 231690
rect 166906 227216 166962 227225
rect 166906 227151 166962 227160
rect 166264 225072 166316 225078
rect 166264 225014 166316 225020
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165528 224392 165580 224398
rect 165528 224334 165580 224340
rect 164976 223576 165028 223582
rect 164976 223518 165028 223524
rect 164332 220516 164384 220522
rect 164332 220458 164384 220464
rect 165540 218210 165568 224334
rect 165804 219428 165856 219434
rect 165804 219370 165856 219376
rect 164976 218204 165028 218210
rect 164976 218146 165028 218152
rect 165528 218204 165580 218210
rect 165528 218146 165580 218152
rect 164068 217246 164142 217274
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217246
rect 164988 217138 165016 218146
rect 165816 217138 165844 219370
rect 166276 219298 166304 225014
rect 166448 223576 166500 223582
rect 166448 223518 166500 223524
rect 166264 219292 166316 219298
rect 166264 219234 166316 219240
rect 166460 218482 166488 223518
rect 167104 221610 167132 231662
rect 167644 229220 167696 229226
rect 167644 229162 167696 229168
rect 167092 221604 167144 221610
rect 167092 221546 167144 221552
rect 167656 218890 167684 229162
rect 168208 225865 168236 231676
rect 168852 230518 168880 231676
rect 168840 230512 168892 230518
rect 168840 230454 168892 230460
rect 169496 228682 169524 231676
rect 169772 231662 170154 231690
rect 169484 228676 169536 228682
rect 169484 228618 169536 228624
rect 168930 228304 168986 228313
rect 168930 228239 168986 228248
rect 168194 225856 168250 225865
rect 168194 225791 168250 225800
rect 168288 223168 168340 223174
rect 168288 223110 168340 223116
rect 167644 218884 167696 218890
rect 167644 218826 167696 218832
rect 166632 218748 166684 218754
rect 166632 218690 166684 218696
rect 166448 218476 166500 218482
rect 166448 218418 166500 218424
rect 166644 217138 166672 218690
rect 168104 218476 168156 218482
rect 168104 218418 168156 218424
rect 167460 218204 167512 218210
rect 167460 218146 167512 218152
rect 167472 217138 167500 218146
rect 168116 217274 168144 218418
rect 168300 218210 168328 223110
rect 168944 219026 168972 228239
rect 169576 227860 169628 227866
rect 169576 227802 169628 227808
rect 168932 219020 168984 219026
rect 168932 218962 168984 218968
rect 169588 218210 169616 227802
rect 169772 221746 169800 231662
rect 169944 228676 169996 228682
rect 169944 228618 169996 228624
rect 169956 227866 169984 228618
rect 169944 227860 169996 227866
rect 169944 227802 169996 227808
rect 170784 223417 170812 231676
rect 171428 223854 171456 231676
rect 172072 227322 172100 231676
rect 172060 227316 172112 227322
rect 172060 227258 172112 227264
rect 172336 224528 172388 224534
rect 172336 224470 172388 224476
rect 171416 223848 171468 223854
rect 171416 223790 171468 223796
rect 170770 223408 170826 223417
rect 170770 223343 170826 223352
rect 169760 221740 169812 221746
rect 169760 221682 169812 221688
rect 171046 221232 171102 221241
rect 171046 221167 171102 221176
rect 170772 220380 170824 220386
rect 170772 220322 170824 220328
rect 169944 219156 169996 219162
rect 169944 219098 169996 219104
rect 169760 218748 169812 218754
rect 169760 218690 169812 218696
rect 169772 218210 169800 218690
rect 168288 218204 168340 218210
rect 168288 218146 168340 218152
rect 169116 218204 169168 218210
rect 169116 218146 169168 218152
rect 169576 218204 169628 218210
rect 169576 218146 169628 218152
rect 169760 218204 169812 218210
rect 169760 218146 169812 218152
rect 168116 217246 168282 217274
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 218146
rect 169956 217138 169984 219098
rect 170784 217274 170812 220322
rect 171060 218482 171088 221167
rect 171416 218748 171468 218754
rect 171416 218690 171468 218696
rect 171048 218476 171100 218482
rect 171048 218418 171100 218424
rect 171428 218074 171456 218690
rect 172152 218476 172204 218482
rect 172152 218418 172204 218424
rect 171416 218068 171468 218074
rect 171416 218010 171468 218016
rect 171600 218068 171652 218074
rect 171600 218010 171652 218016
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217246 170812 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217246
rect 171612 217138 171640 218010
rect 172164 217274 172192 218418
rect 172348 218074 172376 224470
rect 172716 221785 172744 231676
rect 172992 231662 173374 231690
rect 172702 221776 172758 221785
rect 172702 221711 172758 221720
rect 172992 221513 173020 231662
rect 174004 230654 174032 231676
rect 173992 230648 174044 230654
rect 173992 230590 174044 230596
rect 174648 228954 174676 231676
rect 175306 231662 175504 231690
rect 175096 229628 175148 229634
rect 175096 229570 175148 229576
rect 175280 229628 175332 229634
rect 175280 229570 175332 229576
rect 175108 229226 175136 229570
rect 174912 229220 174964 229226
rect 174912 229162 174964 229168
rect 175096 229220 175148 229226
rect 175096 229162 175148 229168
rect 174924 229106 174952 229162
rect 175292 229106 175320 229570
rect 174924 229078 175320 229106
rect 174636 228948 174688 228954
rect 174636 228890 174688 228896
rect 173164 227316 173216 227322
rect 173164 227258 173216 227264
rect 172978 221504 173034 221513
rect 172978 221439 173034 221448
rect 172612 220924 172664 220930
rect 172612 220866 172664 220872
rect 172624 218346 172652 220866
rect 173176 219434 173204 227258
rect 174912 223848 174964 223854
rect 174912 223790 174964 223796
rect 173164 219428 173216 219434
rect 173164 219370 173216 219376
rect 173256 218884 173308 218890
rect 173256 218826 173308 218832
rect 172612 218340 172664 218346
rect 172612 218282 172664 218288
rect 172336 218068 172388 218074
rect 172336 218010 172388 218016
rect 172164 217246 172422 217274
rect 171566 217110 171640 217138
rect 171566 216988 171594 217110
rect 172394 216988 172422 217246
rect 173268 217138 173296 218826
rect 174084 218340 174136 218346
rect 174084 218282 174136 218288
rect 174096 217138 174124 218282
rect 174924 217274 174952 223790
rect 175476 221882 175504 231662
rect 175936 226166 175964 231676
rect 176384 228948 176436 228954
rect 176384 228890 176436 228896
rect 175924 226160 175976 226166
rect 175924 226102 175976 226108
rect 175922 224224 175978 224233
rect 175922 224159 175978 224168
rect 175464 221876 175516 221882
rect 175464 221818 175516 221824
rect 175936 218754 175964 224159
rect 176396 219434 176424 228890
rect 176580 224505 176608 231676
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 177212 226500 177264 226506
rect 177212 226442 177264 226448
rect 176566 224496 176622 224505
rect 176566 224431 176622 224440
rect 176396 219406 176516 219434
rect 175924 218748 175976 218754
rect 175924 218690 175976 218696
rect 176292 218748 176344 218754
rect 176292 218690 176344 218696
rect 175740 218068 175792 218074
rect 175740 218010 175792 218016
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217246 174952 217274
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217246
rect 175752 217138 175780 218010
rect 176304 217274 176332 218690
rect 176488 218074 176516 219406
rect 177224 218482 177252 226442
rect 177408 222018 177436 231662
rect 178512 223446 178540 231676
rect 178788 231662 179170 231690
rect 178500 223440 178552 223446
rect 178500 223382 178552 223388
rect 177396 222012 177448 222018
rect 177396 221954 177448 221960
rect 177396 221740 177448 221746
rect 177396 221682 177448 221688
rect 177212 218476 177264 218482
rect 177212 218418 177264 218424
rect 176476 218068 176528 218074
rect 176476 218010 176528 218016
rect 177408 217274 177436 221682
rect 178224 221604 178276 221610
rect 178224 221546 178276 221552
rect 178236 217274 178264 221546
rect 178788 219434 178816 231662
rect 179800 228818 179828 231676
rect 179984 231662 180458 231690
rect 179788 228812 179840 228818
rect 179788 228754 179840 228760
rect 179984 220794 180012 231662
rect 181088 224670 181116 231676
rect 181076 224664 181128 224670
rect 181076 224606 181128 224612
rect 181732 223310 181760 231676
rect 182376 227594 182404 231676
rect 182560 231662 183034 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181996 224664 182048 224670
rect 181996 224606 182048 224612
rect 181720 223304 181772 223310
rect 181720 223246 181772 223252
rect 179972 220788 180024 220794
rect 179972 220730 180024 220736
rect 180708 220516 180760 220522
rect 180708 220458 180760 220464
rect 179420 219564 179472 219570
rect 179420 219506 179472 219512
rect 178420 219406 178816 219434
rect 179052 219428 179104 219434
rect 178420 217326 178448 219406
rect 179052 219370 179104 219376
rect 176304 217246 176562 217274
rect 175706 217110 175780 217138
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 217246 177436 217274
rect 178190 217246 178264 217274
rect 178408 217320 178460 217326
rect 178408 217262 178460 217268
rect 177362 216988 177390 217246
rect 178190 216988 178218 217246
rect 179064 217138 179092 219370
rect 179432 218346 179460 219506
rect 179880 218476 179932 218482
rect 179880 218418 179932 218424
rect 179420 218340 179472 218346
rect 179420 218282 179472 218288
rect 179892 217138 179920 218418
rect 180720 217274 180748 220458
rect 182008 218074 182036 224606
rect 182560 222154 182588 231662
rect 183468 228812 183520 228818
rect 183468 228754 183520 228760
rect 182824 227588 182876 227594
rect 182824 227530 182876 227536
rect 182548 222148 182600 222154
rect 182548 222090 182600 222096
rect 182836 219434 182864 227530
rect 182824 219428 182876 219434
rect 182824 219370 182876 219376
rect 183192 219428 183244 219434
rect 183192 219370 183244 219376
rect 181536 218068 181588 218074
rect 181536 218010 181588 218016
rect 181996 218068 182048 218074
rect 181996 218010 182048 218016
rect 182364 218068 182416 218074
rect 182364 218010 182416 218016
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181548 217138 181576 218010
rect 182376 217138 182404 218010
rect 183204 217138 183232 219370
rect 183480 218074 183508 228754
rect 183664 222057 183692 231676
rect 184112 230444 184164 230450
rect 184112 230386 184164 230392
rect 184124 229906 184152 230386
rect 184112 229900 184164 229906
rect 184112 229842 184164 229848
rect 184308 229770 184336 231676
rect 184480 229900 184532 229906
rect 184480 229842 184532 229848
rect 184296 229764 184348 229770
rect 184296 229706 184348 229712
rect 184020 222148 184072 222154
rect 184020 222090 184072 222096
rect 183650 222048 183706 222057
rect 183650 221983 183706 221992
rect 183468 218068 183520 218074
rect 183468 218010 183520 218016
rect 184032 217274 184060 222090
rect 184492 219434 184520 229842
rect 184952 228585 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184938 228576 184994 228585
rect 184938 228511 184994 228520
rect 184940 227316 184992 227322
rect 184940 227258 184992 227264
rect 184952 226914 184980 227258
rect 184940 226908 184992 226914
rect 184940 226850 184992 226856
rect 185136 224754 185164 231662
rect 185584 229764 185636 229770
rect 185584 229706 185636 229712
rect 185596 229226 185624 229706
rect 185584 229220 185636 229226
rect 185584 229162 185636 229168
rect 185584 227452 185636 227458
rect 185584 227394 185636 227400
rect 185596 226914 185624 227394
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185044 224726 185164 224754
rect 185044 219978 185072 224726
rect 185216 224664 185268 224670
rect 185214 224632 185216 224641
rect 185400 224664 185452 224670
rect 185268 224632 185270 224641
rect 185400 224606 185452 224612
rect 185214 224567 185270 224576
rect 185032 219972 185084 219978
rect 185032 219914 185084 219920
rect 184216 219406 184520 219434
rect 185412 219434 185440 224606
rect 185596 223718 185624 224878
rect 185872 224806 185900 231662
rect 186044 226024 186096 226030
rect 186044 225966 186096 225972
rect 185860 224800 185912 224806
rect 185860 224742 185912 224748
rect 185584 223712 185636 223718
rect 185584 223654 185636 223660
rect 186056 219434 186084 225966
rect 186884 225078 186912 231676
rect 187528 227730 187556 231676
rect 187896 231662 188186 231690
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 186872 225072 186924 225078
rect 186872 225014 186924 225020
rect 186228 224664 186280 224670
rect 186226 224632 186228 224641
rect 186280 224632 186282 224641
rect 186226 224567 186282 224576
rect 187332 220788 187384 220794
rect 187332 220730 187384 220736
rect 185412 219406 185532 219434
rect 186056 219406 186176 219434
rect 184216 219026 184244 219406
rect 184204 219020 184256 219026
rect 184204 218962 184256 218968
rect 185504 218074 185532 219406
rect 186148 218074 186176 219406
rect 186504 219020 186556 219026
rect 186504 218962 186556 218968
rect 184848 218068 184900 218074
rect 184848 218010 184900 218016
rect 185492 218068 185544 218074
rect 185492 218010 185544 218016
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 181502 217110 181576 217138
rect 182330 217110 182404 217138
rect 183158 217110 183232 217138
rect 183986 217246 184060 217274
rect 181502 216988 181530 217110
rect 182330 216988 182358 217110
rect 183158 216988 183186 217110
rect 183986 216988 184014 217246
rect 184860 217138 184888 218010
rect 185688 217138 185716 218010
rect 186516 217138 186544 218962
rect 187344 217274 187372 220730
rect 187896 220153 187924 231662
rect 188816 224126 188844 231676
rect 189460 230450 189488 231676
rect 189448 230444 189500 230450
rect 189448 230386 189500 230392
rect 189724 229220 189776 229226
rect 189724 229162 189776 229168
rect 188988 227452 189040 227458
rect 188988 227394 189040 227400
rect 188804 224120 188856 224126
rect 188804 224062 188856 224068
rect 187882 220144 187938 220153
rect 187882 220079 187938 220088
rect 188160 218068 188212 218074
rect 188160 218010 188212 218016
rect 184814 217110 184888 217138
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 184814 216988 184842 217110
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188172 217138 188200 218010
rect 189000 217274 189028 227394
rect 189172 221876 189224 221882
rect 189172 221818 189224 221824
rect 189184 218074 189212 221818
rect 189736 218754 189764 229162
rect 190104 229090 190132 231676
rect 190656 231662 190762 231690
rect 191024 231662 191406 231690
rect 190092 229084 190144 229090
rect 190092 229026 190144 229032
rect 189908 224120 189960 224126
rect 189908 224062 189960 224068
rect 189724 218748 189776 218754
rect 189724 218690 189776 218696
rect 189920 218618 189948 224062
rect 190656 221338 190684 231662
rect 191024 223718 191052 231662
rect 191472 224936 191524 224942
rect 191472 224878 191524 224884
rect 191012 223712 191064 223718
rect 191012 223654 191064 223660
rect 190644 221332 190696 221338
rect 190644 221274 190696 221280
rect 189908 218612 189960 218618
rect 189908 218554 189960 218560
rect 190644 218340 190696 218346
rect 190644 218282 190696 218288
rect 189172 218068 189224 218074
rect 189172 218010 189224 218016
rect 189816 218068 189868 218074
rect 189816 218010 189868 218016
rect 188126 217110 188200 217138
rect 188954 217246 189028 217274
rect 188126 216988 188154 217110
rect 188954 216988 188982 217246
rect 189828 217138 189856 218010
rect 190656 217138 190684 218282
rect 191484 217274 191512 224878
rect 192036 223582 192064 231676
rect 192680 227322 192708 231676
rect 193128 229084 193180 229090
rect 193128 229026 193180 229032
rect 192668 227316 192720 227322
rect 192668 227258 192720 227264
rect 192024 223576 192076 223582
rect 192024 223518 192076 223524
rect 191656 223304 191708 223310
rect 191656 223246 191708 223252
rect 191668 218346 191696 223246
rect 192944 219292 192996 219298
rect 192944 219234 192996 219240
rect 191656 218340 191708 218346
rect 191656 218282 191708 218288
rect 192300 218340 192352 218346
rect 192300 218282 192352 218288
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 218282
rect 192956 217274 192984 219234
rect 193140 218346 193168 229026
rect 193324 220425 193352 231676
rect 193968 223990 193996 231676
rect 194612 230790 194640 231676
rect 194600 230784 194652 230790
rect 194600 230726 194652 230732
rect 195256 228274 195284 231676
rect 195440 231662 195914 231690
rect 195244 228268 195296 228274
rect 195244 228210 195296 228216
rect 193956 223984 194008 223990
rect 193956 223926 194008 223932
rect 194508 223576 194560 223582
rect 194508 223518 194560 223524
rect 193310 220416 193366 220425
rect 193310 220351 193366 220360
rect 194520 218346 194548 223518
rect 194784 222012 194836 222018
rect 194784 221954 194836 221960
rect 193128 218340 193180 218346
rect 193128 218282 193180 218288
rect 193956 218340 194008 218346
rect 193956 218282 194008 218288
rect 194508 218340 194560 218346
rect 194508 218282 194560 218288
rect 192956 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218282
rect 194796 217274 194824 221954
rect 195440 219842 195468 231662
rect 196072 230444 196124 230450
rect 196072 230386 196124 230392
rect 195612 225072 195664 225078
rect 195612 225014 195664 225020
rect 195428 219836 195480 219842
rect 195428 219778 195480 219784
rect 195624 217274 195652 225014
rect 196084 222766 196112 230386
rect 196544 226137 196572 231676
rect 197188 230178 197216 231676
rect 197176 230172 197228 230178
rect 197176 230114 197228 230120
rect 197452 230172 197504 230178
rect 197452 230114 197504 230120
rect 196716 227860 196768 227866
rect 196716 227802 196768 227808
rect 196530 226128 196586 226137
rect 196530 226063 196586 226072
rect 196072 222760 196124 222766
rect 196072 222702 196124 222708
rect 196728 219434 196756 227802
rect 197268 223440 197320 223446
rect 197268 223382 197320 223388
rect 196636 219406 196756 219434
rect 196636 219162 196664 219406
rect 196624 219156 196676 219162
rect 196624 219098 196676 219104
rect 196440 218476 196492 218482
rect 196440 218418 196492 218424
rect 196452 217274 196480 218418
rect 197280 217274 197308 223382
rect 197464 222494 197492 230114
rect 197832 226778 197860 231676
rect 198476 230450 198504 231676
rect 198464 230444 198516 230450
rect 198464 230386 198516 230392
rect 198648 227316 198700 227322
rect 198648 227258 198700 227264
rect 197820 226772 197872 226778
rect 197820 226714 197872 226720
rect 197452 222488 197504 222494
rect 197452 222430 197504 222436
rect 198660 218346 198688 227258
rect 198924 218612 198976 218618
rect 198924 218554 198976 218560
rect 198096 218340 198148 218346
rect 198096 218282 198148 218288
rect 198648 218340 198700 218346
rect 198648 218282 198700 218288
rect 193922 217110 193996 217138
rect 194750 217246 194824 217274
rect 195578 217246 195652 217274
rect 196406 217246 196480 217274
rect 197234 217246 197308 217274
rect 193922 216988 193950 217110
rect 194750 216988 194778 217246
rect 195578 216988 195606 217246
rect 196406 216988 196434 217246
rect 197234 216988 197262 217246
rect 198108 217138 198136 218282
rect 198936 217138 198964 218554
rect 199120 217462 199148 231676
rect 199488 231662 199778 231690
rect 199488 220930 199516 231662
rect 200408 228138 200436 231676
rect 201052 230178 201080 231676
rect 201040 230172 201092 230178
rect 201040 230114 201092 230120
rect 200396 228132 200448 228138
rect 200396 228074 200448 228080
rect 200028 227724 200080 227730
rect 200028 227666 200080 227672
rect 199476 220924 199528 220930
rect 199476 220866 199528 220872
rect 199292 219428 199344 219434
rect 199292 219370 199344 219376
rect 199752 219428 199804 219434
rect 199752 219370 199804 219376
rect 199304 218346 199332 219370
rect 199292 218340 199344 218346
rect 199292 218282 199344 218288
rect 199108 217456 199160 217462
rect 199108 217398 199160 217404
rect 199764 217138 199792 219370
rect 200040 218618 200068 227666
rect 201696 225486 201724 231676
rect 202340 230314 202368 231676
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202144 230172 202196 230178
rect 202144 230114 202196 230120
rect 201684 225480 201736 225486
rect 201684 225422 201736 225428
rect 200764 223984 200816 223990
rect 200764 223926 200816 223932
rect 200580 219972 200632 219978
rect 200580 219914 200632 219920
rect 200028 218612 200080 218618
rect 200028 218554 200080 218560
rect 200592 217274 200620 219914
rect 200776 218657 200804 223926
rect 201408 221332 201460 221338
rect 201408 221274 201460 221280
rect 200762 218648 200818 218657
rect 200762 218583 200818 218592
rect 201420 217274 201448 221274
rect 202156 219434 202184 230114
rect 202984 227497 203012 231676
rect 203168 231662 203642 231690
rect 202970 227488 203026 227497
rect 202970 227423 203026 227432
rect 202696 226160 202748 226166
rect 202696 226102 202748 226108
rect 202064 219406 202184 219434
rect 201868 218612 201920 218618
rect 201868 218554 201920 218560
rect 201880 218210 201908 218554
rect 202064 218346 202092 219406
rect 202052 218340 202104 218346
rect 202052 218282 202104 218288
rect 202708 218210 202736 226102
rect 203168 219706 203196 231662
rect 204272 226302 204300 231676
rect 204260 226296 204312 226302
rect 204260 226238 204312 226244
rect 204916 224233 204944 231676
rect 205364 228268 205416 228274
rect 205364 228210 205416 228216
rect 204902 224224 204958 224233
rect 204902 224159 204958 224168
rect 203892 222488 203944 222494
rect 203892 222430 203944 222436
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 203064 219428 203116 219434
rect 203064 219370 203116 219376
rect 203076 219162 203104 219370
rect 203064 219156 203116 219162
rect 203064 219098 203116 219104
rect 203064 218340 203116 218346
rect 203064 218282 203116 218288
rect 201868 218204 201920 218210
rect 201868 218146 201920 218152
rect 202236 218204 202288 218210
rect 202236 218146 202288 218152
rect 202696 218204 202748 218210
rect 202696 218146 202748 218152
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217246 200620 217274
rect 201374 217246 201448 217274
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217246
rect 201374 216988 201402 217246
rect 202248 217138 202276 218146
rect 203076 217138 203104 218282
rect 203904 217274 203932 222430
rect 205376 219434 205404 228210
rect 205560 228002 205588 231676
rect 205836 231662 206218 231690
rect 206388 231662 206862 231690
rect 205548 227996 205600 228002
rect 205548 227938 205600 227944
rect 205548 226296 205600 226302
rect 205548 226238 205600 226244
rect 205560 219434 205588 226238
rect 205836 221066 205864 231662
rect 206192 225480 206244 225486
rect 206192 225422 206244 225428
rect 205824 221060 205876 221066
rect 205824 221002 205876 221008
rect 204720 219428 204772 219434
rect 205376 219406 205496 219434
rect 205560 219428 205692 219434
rect 205560 219406 205640 219428
rect 204720 219370 204772 219376
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 219370
rect 205468 217274 205496 219406
rect 205640 219370 205692 219376
rect 205652 219339 205680 219370
rect 206204 218618 206232 225422
rect 206388 225350 206416 231662
rect 207492 229770 207520 231676
rect 207664 230444 207716 230450
rect 207664 230386 207716 230392
rect 207480 229764 207532 229770
rect 207480 229706 207532 229712
rect 206744 226160 206796 226166
rect 206744 226102 206796 226108
rect 206756 225486 206784 226102
rect 206744 225480 206796 225486
rect 206744 225422 206796 225428
rect 206376 225344 206428 225350
rect 206376 225286 206428 225292
rect 207204 219836 207256 219842
rect 207204 219778 207256 219784
rect 206192 218612 206244 218618
rect 206192 218554 206244 218560
rect 206376 218612 206428 218618
rect 206376 218554 206428 218560
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218554
rect 207216 217274 207244 219778
rect 207676 218482 207704 230386
rect 208136 227050 208164 231676
rect 208596 231662 208794 231690
rect 208124 227044 208176 227050
rect 208124 226986 208176 226992
rect 208032 222760 208084 222766
rect 208032 222702 208084 222708
rect 207664 218476 207716 218482
rect 207664 218418 207716 218424
rect 208044 217274 208072 222702
rect 208596 220658 208624 231662
rect 209424 225758 209452 231676
rect 210068 229498 210096 231676
rect 210424 229764 210476 229770
rect 210424 229706 210476 229712
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 209412 225752 209464 225758
rect 209412 225694 209464 225700
rect 209596 225752 209648 225758
rect 209596 225694 209648 225700
rect 208584 220652 208636 220658
rect 208584 220594 208636 220600
rect 209608 219586 209636 225694
rect 209516 219558 209636 219586
rect 209516 218210 209544 219558
rect 210436 219434 210464 229706
rect 210712 228410 210740 231676
rect 210700 228404 210752 228410
rect 210700 228346 210752 228352
rect 211068 228132 211120 228138
rect 211068 228074 211120 228080
rect 209688 219428 209740 219434
rect 209688 219370 209740 219376
rect 210332 219428 210464 219434
rect 210384 219406 210464 219428
rect 210332 219370 210384 219376
rect 208860 218204 208912 218210
rect 208860 218146 208912 218152
rect 209504 218204 209556 218210
rect 209504 218146 209556 218152
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 207998 217246 208072 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 207998 216988 208026 217246
rect 208872 217138 208900 218146
rect 209700 217138 209728 219370
rect 210884 218884 210936 218890
rect 210884 218826 210936 218832
rect 210896 218482 210924 218826
rect 210884 218476 210936 218482
rect 210884 218418 210936 218424
rect 211080 218210 211108 228074
rect 211356 220697 211384 231676
rect 212000 222630 212028 231676
rect 212172 226908 212224 226914
rect 212172 226850 212224 226856
rect 211988 222624 212040 222630
rect 211988 222566 212040 222572
rect 211342 220688 211398 220697
rect 211342 220623 211398 220632
rect 210516 218204 210568 218210
rect 210516 218146 210568 218152
rect 211068 218204 211120 218210
rect 211068 218146 211120 218152
rect 211344 218204 211396 218210
rect 211344 218146 211396 218152
rect 210528 217138 210556 218146
rect 211356 217138 211384 218146
rect 212184 217274 212212 226850
rect 212644 224126 212672 231676
rect 213092 229356 213144 229362
rect 213092 229298 213144 229304
rect 213104 229094 213132 229298
rect 213288 229094 213316 231676
rect 213104 229066 213224 229094
rect 213288 229066 213408 229094
rect 212632 224120 212684 224126
rect 212632 224062 212684 224068
rect 212816 219428 212868 219434
rect 212816 219370 212868 219376
rect 212828 218618 212856 219370
rect 212816 218612 212868 218618
rect 212816 218554 212868 218560
rect 213000 218612 213052 218618
rect 213000 218554 213052 218560
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217110 210556 217138
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217110
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 218554
rect 213196 218346 213224 229066
rect 213380 227186 213408 229066
rect 213368 227180 213420 227186
rect 213368 227122 213420 227128
rect 213932 222873 213960 231676
rect 214116 231662 214590 231690
rect 213918 222864 213974 222873
rect 213918 222799 213974 222808
rect 213828 222624 213880 222630
rect 213828 222566 213880 222572
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 222566
rect 214116 221202 214144 231662
rect 214380 230172 214432 230178
rect 214380 230114 214432 230120
rect 214392 229906 214420 230114
rect 214380 229900 214432 229906
rect 214380 229842 214432 229848
rect 215220 229498 215248 231676
rect 215208 229492 215260 229498
rect 215208 229434 215260 229440
rect 215864 228546 215892 231676
rect 216232 231662 216522 231690
rect 215852 228540 215904 228546
rect 215852 228482 215904 228488
rect 215208 228404 215260 228410
rect 215208 228346 215260 228352
rect 214104 221196 214156 221202
rect 214104 221138 214156 221144
rect 214288 221196 214340 221202
rect 214288 221138 214340 221144
rect 214300 218210 214328 221138
rect 215220 218210 215248 228346
rect 216232 222902 216260 231662
rect 217152 224262 217180 231676
rect 217796 229634 217824 231676
rect 217784 229628 217836 229634
rect 217784 229570 217836 229576
rect 217324 229492 217376 229498
rect 217324 229434 217376 229440
rect 217140 224256 217192 224262
rect 217140 224198 217192 224204
rect 216588 224120 216640 224126
rect 216588 224062 216640 224068
rect 216220 222896 216272 222902
rect 216220 222838 216272 222844
rect 216312 220652 216364 220658
rect 216312 220594 216364 220600
rect 214288 218204 214340 218210
rect 214288 218146 214340 218152
rect 214656 218204 214708 218210
rect 214656 218146 214708 218152
rect 215208 218204 215260 218210
rect 215208 218146 215260 218152
rect 215484 218204 215536 218210
rect 215484 218146 215536 218152
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218146
rect 215496 217138 215524 218146
rect 216324 217274 216352 220594
rect 216600 218210 216628 224062
rect 217336 220658 217364 229434
rect 218440 225214 218468 231676
rect 218716 231662 219098 231690
rect 218428 225208 218480 225214
rect 218428 225150 218480 225156
rect 217876 222896 217928 222902
rect 217876 222838 217928 222844
rect 217324 220652 217376 220658
rect 217324 220594 217376 220600
rect 217508 220652 217560 220658
rect 217508 220594 217560 220600
rect 217520 219434 217548 220594
rect 217152 219406 217548 219434
rect 216588 218204 216640 218210
rect 216588 218146 216640 218152
rect 217152 217274 217180 219406
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217246 216352 217274
rect 217106 217246 217180 217274
rect 217888 217274 217916 222838
rect 218716 220114 218744 231662
rect 219348 226296 219400 226302
rect 219348 226238 219400 226244
rect 218704 220108 218756 220114
rect 218704 220050 218756 220056
rect 219360 218210 219388 226238
rect 219728 225622 219756 231676
rect 220372 229906 220400 231676
rect 220360 229900 220412 229906
rect 220360 229842 220412 229848
rect 221016 226642 221044 231676
rect 221292 231662 221674 231690
rect 221004 226636 221056 226642
rect 221004 226578 221056 226584
rect 219716 225616 219768 225622
rect 219716 225558 219768 225564
rect 220452 225616 220504 225622
rect 220452 225558 220504 225564
rect 219624 218340 219676 218346
rect 219624 218282 219676 218288
rect 218796 218204 218848 218210
rect 218796 218146 218848 218152
rect 219348 218204 219400 218210
rect 219348 218146 219400 218152
rect 217888 217246 217962 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217246
rect 217106 216988 217134 217246
rect 217934 216988 217962 217246
rect 218808 217138 218836 218146
rect 219636 217138 219664 218282
rect 220464 217274 220492 225558
rect 220820 220244 220872 220250
rect 220820 220186 220872 220192
rect 220832 218482 220860 220186
rect 221292 220114 221320 231662
rect 222016 228540 222068 228546
rect 222016 228482 222068 228488
rect 221280 220108 221332 220114
rect 221280 220050 221332 220056
rect 220820 218476 220872 218482
rect 220820 218418 220872 218424
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 228482
rect 222304 225894 222332 231676
rect 222292 225888 222344 225894
rect 222292 225830 222344 225836
rect 222948 223990 222976 231676
rect 223592 228313 223620 231676
rect 224040 229900 224092 229906
rect 224040 229842 224092 229848
rect 224052 229498 224080 229842
rect 224040 229492 224092 229498
rect 224040 229434 224092 229440
rect 223578 228304 223634 228313
rect 223578 228239 223634 228248
rect 223488 224256 223540 224262
rect 223488 224198 223540 224204
rect 222936 223984 222988 223990
rect 222936 223926 222988 223932
rect 222568 221060 222620 221066
rect 222568 221002 222620 221008
rect 222580 218074 222608 221002
rect 223500 218074 223528 224198
rect 224236 223038 224264 231676
rect 224512 231662 224894 231690
rect 224512 229094 224540 231662
rect 225524 230178 225552 231676
rect 225512 230172 225564 230178
rect 225512 230114 225564 230120
rect 225788 230036 225840 230042
rect 225788 229978 225840 229984
rect 224420 229066 224540 229094
rect 224224 223032 224276 223038
rect 224224 222974 224276 222980
rect 224420 221474 224448 229066
rect 224776 227180 224828 227186
rect 224776 227122 224828 227128
rect 224592 226772 224644 226778
rect 224592 226714 224644 226720
rect 224408 221468 224460 221474
rect 224408 221410 224460 221416
rect 224604 218074 224632 226714
rect 222568 218068 222620 218074
rect 222568 218010 222620 218016
rect 222936 218068 222988 218074
rect 222936 218010 222988 218016
rect 223488 218068 223540 218074
rect 223488 218010 223540 218016
rect 223764 218068 223816 218074
rect 223764 218010 223816 218016
rect 224592 218068 224644 218074
rect 224592 218010 224644 218016
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218010
rect 223776 217138 223804 218010
rect 224788 217274 224816 227122
rect 225604 225208 225656 225214
rect 225604 225150 225656 225156
rect 225616 218210 225644 225150
rect 225800 224262 225828 229978
rect 226168 227050 226196 231676
rect 226156 227044 226208 227050
rect 226156 226986 226208 226992
rect 225788 224256 225840 224262
rect 225788 224198 225840 224204
rect 226156 223984 226208 223990
rect 226156 223926 226208 223932
rect 225972 218476 226024 218482
rect 225972 218418 226024 218424
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217246 224816 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218418
rect 226168 218074 226196 223926
rect 226812 223174 226840 231676
rect 227456 224398 227484 231676
rect 228100 225350 228128 231676
rect 228744 228682 228772 231676
rect 229112 231662 229402 231690
rect 229572 231662 230046 231690
rect 228732 228676 228784 228682
rect 228732 228618 228784 228624
rect 228732 227044 228784 227050
rect 228732 226986 228784 226992
rect 228088 225344 228140 225350
rect 228088 225286 228140 225292
rect 227444 224392 227496 224398
rect 227444 224334 227496 224340
rect 227628 223712 227680 223718
rect 227628 223654 227680 223660
rect 226800 223168 226852 223174
rect 226800 223110 226852 223116
rect 227640 218074 227668 223654
rect 227904 220924 227956 220930
rect 227904 220866 227956 220872
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227076 218068 227128 218074
rect 227076 218010 227128 218016
rect 227628 218068 227680 218074
rect 227628 218010 227680 218016
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227088 217138 227116 218010
rect 227916 217274 227944 220866
rect 228744 217274 228772 226986
rect 229112 220386 229140 231662
rect 229572 221241 229600 231662
rect 230480 230172 230532 230178
rect 230480 230114 230532 230120
rect 230492 223530 230520 230114
rect 230676 227866 230704 231676
rect 230664 227860 230716 227866
rect 230664 227802 230716 227808
rect 231320 226506 231348 231676
rect 231308 226500 231360 226506
rect 231308 226442 231360 226448
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 230400 223502 230520 223530
rect 229558 221232 229614 221241
rect 229558 221167 229614 221176
rect 229100 220380 229152 220386
rect 229100 220322 229152 220328
rect 230204 220108 230256 220114
rect 230204 220050 230256 220056
rect 230216 219434 230244 220050
rect 230216 219406 230336 219434
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 227042 217110 227116 217138
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217110
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230308 217274 230336 219406
rect 230400 218090 230428 223502
rect 230400 218074 230520 218090
rect 231688 218074 231716 224198
rect 231964 219570 231992 231676
rect 232608 224534 232636 231676
rect 233266 231662 233464 231690
rect 232596 224528 232648 224534
rect 232596 224470 232648 224476
rect 233148 224528 233200 224534
rect 233148 224470 233200 224476
rect 232688 220516 232740 220522
rect 232688 220458 232740 220464
rect 231952 219564 232004 219570
rect 231952 219506 232004 219512
rect 232700 218754 232728 220458
rect 232872 218884 232924 218890
rect 232872 218826 232924 218832
rect 232688 218748 232740 218754
rect 232688 218690 232740 218696
rect 230400 218068 230532 218074
rect 230400 218062 230480 218068
rect 230480 218010 230532 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217138 232912 218826
rect 233160 218074 233188 224470
rect 233436 220250 233464 231662
rect 233896 228954 233924 231676
rect 234172 231662 234554 231690
rect 233884 228948 233936 228954
rect 233884 228890 233936 228896
rect 234172 221746 234200 231662
rect 234528 228948 234580 228954
rect 234528 228890 234580 228896
rect 234160 221740 234212 221746
rect 234160 221682 234212 221688
rect 234344 221468 234396 221474
rect 234344 221410 234396 221416
rect 233424 220244 233476 220250
rect 233424 220186 233476 220192
rect 234356 219434 234384 221410
rect 234356 219406 234476 219434
rect 233884 219292 233936 219298
rect 233884 219234 233936 219240
rect 233896 218754 233924 219234
rect 233884 218748 233936 218754
rect 233884 218690 233936 218696
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233700 218068 233752 218074
rect 233700 218010 233752 218016
rect 233712 217138 233740 218010
rect 234448 217274 234476 219406
rect 234540 218090 234568 228890
rect 235184 223854 235212 231676
rect 235828 229226 235856 231676
rect 235816 229220 235868 229226
rect 235816 229162 235868 229168
rect 235816 228676 235868 228682
rect 235816 228618 235868 228624
rect 235172 223848 235224 223854
rect 235172 223790 235224 223796
rect 235632 220380 235684 220386
rect 235632 220322 235684 220328
rect 235644 219026 235672 220322
rect 235632 219020 235684 219026
rect 235632 218962 235684 218968
rect 234540 218074 234660 218090
rect 235828 218074 235856 228618
rect 236472 227594 236500 231676
rect 236656 231662 237130 231690
rect 237392 231662 237774 231690
rect 238036 231662 238418 231690
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 236656 220250 236684 231662
rect 237392 221610 237420 231662
rect 237380 221604 237432 221610
rect 237380 221546 237432 221552
rect 238036 220522 238064 231662
rect 239048 228818 239076 231676
rect 239232 231662 239706 231690
rect 239036 228812 239088 228818
rect 239036 228754 239088 228760
rect 238668 223032 238720 223038
rect 238668 222974 238720 222980
rect 238024 220516 238076 220522
rect 238024 220458 238076 220464
rect 236644 220244 236696 220250
rect 236644 220186 236696 220192
rect 237012 220244 237064 220250
rect 237012 220186 237064 220192
rect 236184 219700 236236 219706
rect 236184 219642 236236 219648
rect 234540 218068 234672 218074
rect 234540 218062 234620 218068
rect 234620 218010 234672 218016
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 234448 217246 234522 217274
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217110 233740 217138
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217110
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217274 236224 219642
rect 237024 217274 237052 220186
rect 237840 219292 237892 219298
rect 237840 219234 237892 219240
rect 235322 217110 235396 217138
rect 236150 217246 236224 217274
rect 236978 217246 237052 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217246
rect 236978 216988 237006 217246
rect 237852 217138 237880 219234
rect 238680 217274 238708 222974
rect 239232 222154 239260 231662
rect 239404 225888 239456 225894
rect 239404 225830 239456 225836
rect 239220 222148 239272 222154
rect 239220 222090 239272 222096
rect 238852 221604 238904 221610
rect 238852 221546 238904 221552
rect 238864 218754 238892 221546
rect 239416 219298 239444 225830
rect 240336 224670 240364 231676
rect 240980 230314 241008 231676
rect 240968 230308 241020 230314
rect 240968 230250 241020 230256
rect 241624 226030 241652 231676
rect 241808 231662 242282 231690
rect 241612 226024 241664 226030
rect 241612 225966 241664 225972
rect 240324 224664 240376 224670
rect 240324 224606 240376 224612
rect 241152 224392 241204 224398
rect 241152 224334 241204 224340
rect 240324 220516 240376 220522
rect 240324 220458 240376 220464
rect 239404 219292 239456 219298
rect 239404 219234 239456 219240
rect 238852 218748 238904 218754
rect 238852 218690 238904 218696
rect 239496 218748 239548 218754
rect 239496 218690 239548 218696
rect 237806 217110 237880 217138
rect 238634 217246 238708 217274
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 218690
rect 240336 217274 240364 220458
rect 241164 217274 241192 224334
rect 241808 220794 241836 231662
rect 242532 230308 242584 230314
rect 242532 230250 242584 230256
rect 242544 229094 242572 230250
rect 242544 229066 242756 229094
rect 241980 227588 242032 227594
rect 241980 227530 242032 227536
rect 241796 220788 241848 220794
rect 241796 220730 241848 220736
rect 241992 217274 242020 227530
rect 239462 217110 239536 217138
rect 240290 217246 240364 217274
rect 241118 217246 241192 217274
rect 241946 217246 242020 217274
rect 242728 217274 242756 229066
rect 242912 224806 242940 231676
rect 243096 231662 243570 231690
rect 242900 224800 242952 224806
rect 242900 224742 242952 224748
rect 243096 220386 243124 231662
rect 244200 227458 244228 231676
rect 244188 227452 244240 227458
rect 244188 227394 244240 227400
rect 244844 223310 244872 231676
rect 245028 231662 245502 231690
rect 244832 223304 244884 223310
rect 244832 223246 244884 223252
rect 244096 222352 244148 222358
rect 244096 222294 244148 222300
rect 243084 220380 243136 220386
rect 243084 220322 243136 220328
rect 244108 218074 244136 222294
rect 245028 221882 245056 231662
rect 245292 226024 245344 226030
rect 245292 225966 245344 225972
rect 245016 221876 245068 221882
rect 245016 221818 245068 221824
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 242728 217246 242802 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217246
rect 241118 216988 241146 217246
rect 241946 216988 241974 217246
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217138 244504 218010
rect 245304 217274 245332 225966
rect 246132 225214 246160 231676
rect 246776 229090 246804 231676
rect 246764 229084 246816 229090
rect 246764 229026 246816 229032
rect 246304 228812 246356 228818
rect 246304 228754 246356 228760
rect 246120 225208 246172 225214
rect 246120 225150 246172 225156
rect 246120 219020 246172 219026
rect 246120 218962 246172 218968
rect 246132 217274 246160 218962
rect 246316 218074 246344 228754
rect 247420 223582 247448 231676
rect 248064 224942 248092 231676
rect 248616 231662 248722 231690
rect 248052 224936 248104 224942
rect 248052 224878 248104 224884
rect 247408 223576 247460 223582
rect 247408 223518 247460 223524
rect 248236 223168 248288 223174
rect 248236 223110 248288 223116
rect 247132 221740 247184 221746
rect 247132 221682 247184 221688
rect 246948 220380 247000 220386
rect 246948 220322 247000 220328
rect 246304 218068 246356 218074
rect 246304 218010 246356 218016
rect 246960 217274 246988 220322
rect 247144 219162 247172 221682
rect 247132 219156 247184 219162
rect 247132 219098 247184 219104
rect 248248 218074 248276 223110
rect 248616 221610 248644 231662
rect 249352 225078 249380 231676
rect 249340 225072 249392 225078
rect 249340 225014 249392 225020
rect 249616 224664 249668 224670
rect 249616 224606 249668 224612
rect 248604 221604 248656 221610
rect 248604 221546 248656 221552
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 243602 217110 243676 217138
rect 244430 217110 244504 217138
rect 245258 217246 245332 217274
rect 246086 217246 246160 217274
rect 246914 217246 246988 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246086 216988 246114 217246
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218146
rect 249628 218074 249656 224606
rect 249996 223446 250024 231676
rect 250180 231662 250654 231690
rect 249984 223440 250036 223446
rect 249984 223382 250036 223388
rect 250180 222018 250208 231662
rect 251284 230450 251312 231676
rect 251272 230444 251324 230450
rect 251272 230386 251324 230392
rect 251732 229628 251784 229634
rect 251732 229570 251784 229576
rect 251088 227452 251140 227458
rect 251088 227394 251140 227400
rect 250168 222012 250220 222018
rect 250168 221954 250220 221960
rect 250260 221604 250312 221610
rect 250260 221546 250312 221552
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250272 217274 250300 221546
rect 251100 217274 251128 227394
rect 251744 218210 251772 229570
rect 251928 227730 251956 231676
rect 252586 231662 252784 231690
rect 252376 227996 252428 228002
rect 252376 227938 252428 227944
rect 251916 227724 251968 227730
rect 251916 227666 251968 227672
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 252388 218074 252416 227938
rect 252560 221876 252612 221882
rect 252560 221818 252612 221824
rect 252572 219434 252600 221818
rect 252756 219978 252784 231662
rect 253216 227322 253244 231676
rect 253400 231662 253874 231690
rect 253204 227316 253256 227322
rect 253204 227258 253256 227264
rect 253400 221746 253428 231662
rect 254504 225486 254532 231676
rect 254872 231662 255162 231690
rect 255424 231662 255806 231690
rect 254492 225480 254544 225486
rect 254492 225422 254544 225428
rect 253572 223576 253624 223582
rect 253572 223518 253624 223524
rect 253388 221740 253440 221746
rect 253388 221682 253440 221688
rect 252744 219972 252796 219978
rect 252744 219914 252796 219920
rect 252560 219428 252612 219434
rect 252560 219370 252612 219376
rect 252744 219292 252796 219298
rect 252744 219234 252796 219240
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252376 218068 252428 218074
rect 252376 218010 252428 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217246 250300 217274
rect 251054 217246 251128 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217246
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217274 252784 219234
rect 253584 217274 253612 223518
rect 254872 222494 254900 231662
rect 255228 225480 255280 225486
rect 255228 225422 255280 225428
rect 255044 225344 255096 225350
rect 255044 225286 255096 225292
rect 254860 222488 254912 222494
rect 254860 222430 254912 222436
rect 255056 219434 255084 225286
rect 255240 219434 255268 225422
rect 255424 221338 255452 231662
rect 256436 229498 256464 231676
rect 256608 230444 256660 230450
rect 256608 230386 256660 230392
rect 256424 229492 256476 229498
rect 256424 229434 256476 229440
rect 255412 221332 255464 221338
rect 255412 221274 255464 221280
rect 256620 219434 256648 230386
rect 257080 228274 257108 231676
rect 257264 231662 257738 231690
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 256884 219972 256936 219978
rect 256884 219914 256936 219920
rect 254400 219428 254452 219434
rect 255056 219406 255176 219434
rect 255240 219428 255372 219434
rect 255240 219406 255320 219428
rect 254400 219370 254452 219376
rect 251882 217110 251956 217138
rect 252710 217246 252784 217274
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217246
rect 253538 216988 253566 217246
rect 254412 217138 254440 219370
rect 255148 217274 255176 219406
rect 255320 219370 255372 219376
rect 256528 219406 256648 219434
rect 256528 218074 256556 219406
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 255148 217246 255222 217274
rect 254366 217110 254440 217138
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217274 256924 219914
rect 257264 219842 257292 231662
rect 257712 229084 257764 229090
rect 257712 229026 257764 229032
rect 257252 219836 257304 219842
rect 257252 219778 257304 219784
rect 257724 217274 257752 229026
rect 258368 226166 258396 231676
rect 258644 231662 259026 231690
rect 258356 226160 258408 226166
rect 258356 226102 258408 226108
rect 258080 222012 258132 222018
rect 258080 221954 258132 221960
rect 258092 218346 258120 221954
rect 258644 221882 258672 231662
rect 259368 227316 259420 227322
rect 259368 227258 259420 227264
rect 258632 221876 258684 221882
rect 258632 221818 258684 221824
rect 259184 219292 259236 219298
rect 259184 219234 259236 219240
rect 258080 218340 258132 218346
rect 258080 218282 258132 218288
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217246 256924 217274
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217246
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259196 217274 259224 219234
rect 259380 218074 259408 227258
rect 259656 225758 259684 231676
rect 260300 228138 260328 231676
rect 260288 228132 260340 228138
rect 260288 228074 260340 228080
rect 259644 225752 259696 225758
rect 259644 225694 259696 225700
rect 260012 225004 260064 225010
rect 260012 224946 260064 224952
rect 260024 218618 260052 224946
rect 260944 222766 260972 231676
rect 261588 229770 261616 231676
rect 261576 229764 261628 229770
rect 261576 229706 261628 229712
rect 261484 229356 261536 229362
rect 261484 229298 261536 229304
rect 260932 222760 260984 222766
rect 260932 222702 260984 222708
rect 260196 221740 260248 221746
rect 260196 221682 260248 221688
rect 260012 218612 260064 218618
rect 260012 218554 260064 218560
rect 259368 218068 259420 218074
rect 259368 218010 259420 218016
rect 260208 217274 260236 221682
rect 261024 220788 261076 220794
rect 261024 220730 261076 220736
rect 261036 217274 261064 220730
rect 261496 219706 261524 229298
rect 262232 226914 262260 231676
rect 262220 226908 262272 226914
rect 262220 226850 262272 226856
rect 261852 223304 261904 223310
rect 261852 223246 261904 223252
rect 261484 219700 261536 219706
rect 261484 219642 261536 219648
rect 261864 217274 261892 223246
rect 262876 222630 262904 231676
rect 263152 231662 263534 231690
rect 262864 222624 262916 222630
rect 262864 222566 262916 222572
rect 263152 221202 263180 231662
rect 263416 227724 263468 227730
rect 263416 227666 263468 227672
rect 263140 221196 263192 221202
rect 263140 221138 263192 221144
rect 262680 218612 262732 218618
rect 262680 218554 262732 218560
rect 259196 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260162 217246 260236 217274
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 260162 216988 260190 217246
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262692 217138 262720 218554
rect 263428 217274 263456 227666
rect 264164 225010 264192 231676
rect 264440 231662 264822 231690
rect 265084 231662 265466 231690
rect 264152 225004 264204 225010
rect 264152 224946 264204 224952
rect 264440 224126 264468 231662
rect 264888 225752 264940 225758
rect 264888 225694 264940 225700
rect 264428 224120 264480 224126
rect 264428 224062 264480 224068
rect 264900 218074 264928 225694
rect 265084 220658 265112 231662
rect 266096 228410 266124 231676
rect 266740 229906 266768 231676
rect 266728 229900 266780 229906
rect 266728 229842 266780 229848
rect 266084 228404 266136 228410
rect 266084 228346 266136 228352
rect 265624 228268 265676 228274
rect 265624 228210 265676 228216
rect 265072 220652 265124 220658
rect 265072 220594 265124 220600
rect 265636 218482 265664 228210
rect 267384 226302 267412 231676
rect 267372 226296 267424 226302
rect 267372 226238 267424 226244
rect 268028 225622 268056 231676
rect 268016 225616 268068 225622
rect 268016 225558 268068 225564
rect 266268 224936 266320 224942
rect 266268 224878 266320 224884
rect 265624 218476 265676 218482
rect 265624 218418 265676 218424
rect 265992 218476 266044 218482
rect 265992 218418 266044 218424
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264888 218068 264940 218074
rect 264888 218010 264940 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263428 217246 263502 217274
rect 262646 217110 262720 217138
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 218418
rect 266280 218074 266308 224878
rect 267556 223440 267608 223446
rect 267556 223382 267608 223388
rect 266820 221876 266872 221882
rect 266820 221818 266872 221824
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266832 217274 266860 221818
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267568 217274 267596 223382
rect 268672 222902 268700 231676
rect 269224 231662 269330 231690
rect 269028 225616 269080 225622
rect 269028 225558 269080 225564
rect 268660 222896 268712 222902
rect 268660 222838 268712 222844
rect 269040 218074 269068 225558
rect 269224 222018 269252 231662
rect 269960 228546 269988 231676
rect 270132 229764 270184 229770
rect 270132 229706 270184 229712
rect 270144 229094 270172 229706
rect 270144 229066 270264 229094
rect 269948 228540 270000 228546
rect 269948 228482 270000 228488
rect 269212 222012 269264 222018
rect 269212 221954 269264 221960
rect 270040 222012 270092 222018
rect 270040 221954 270092 221960
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 269028 218068 269080 218074
rect 269028 218010 269080 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 267568 217246 267642 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270052 217274 270080 221954
rect 270236 218074 270264 229066
rect 270604 226778 270632 231676
rect 270880 231662 271262 231690
rect 270592 226772 270644 226778
rect 270592 226714 270644 226720
rect 270880 221066 270908 231662
rect 271892 230042 271920 231676
rect 271880 230036 271932 230042
rect 271880 229978 271932 229984
rect 271788 228404 271840 228410
rect 271788 228346 271840 228352
rect 271604 224800 271656 224806
rect 271604 224742 271656 224748
rect 270868 221060 270920 221066
rect 270868 221002 270920 221008
rect 270776 219564 270828 219570
rect 270776 219506 270828 219512
rect 270788 218890 270816 219506
rect 270776 218884 270828 218890
rect 270776 218826 270828 218832
rect 271616 218074 271644 224742
rect 270224 218068 270276 218074
rect 270224 218010 270276 218016
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 271604 218068 271656 218074
rect 271604 218010 271656 218016
rect 270052 217246 270126 217274
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 228346
rect 272536 223990 272564 231676
rect 272524 223984 272576 223990
rect 272524 223926 272576 223932
rect 273180 223718 273208 231676
rect 273824 227186 273852 231676
rect 274088 228540 274140 228546
rect 274088 228482 274140 228488
rect 273812 227180 273864 227186
rect 273812 227122 273864 227128
rect 273168 223712 273220 223718
rect 273168 223654 273220 223660
rect 272432 219428 272484 219434
rect 272432 219370 272484 219376
rect 272444 218482 272472 219370
rect 272432 218476 272484 218482
rect 272432 218418 272484 218424
rect 272616 218476 272668 218482
rect 272616 218418 272668 218424
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272628 217138 272656 218418
rect 274100 218074 274128 228482
rect 274468 228274 274496 231676
rect 274456 228268 274508 228274
rect 274456 228210 274508 228216
rect 274272 227180 274324 227186
rect 274272 227122 274324 227128
rect 273444 218068 273496 218074
rect 273444 218010 273496 218016
rect 274088 218068 274140 218074
rect 274088 218010 274140 218016
rect 273456 217138 273484 218010
rect 274284 217274 274312 227122
rect 275112 227050 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 227044 275152 227050
rect 275100 226986 275152 226992
rect 275296 220114 275324 231662
rect 275652 226908 275704 226914
rect 275652 226850 275704 226856
rect 275284 220108 275336 220114
rect 275284 220050 275336 220056
rect 275664 218074 275692 226850
rect 275836 224120 275888 224126
rect 275836 224062 275888 224068
rect 275100 218068 275152 218074
rect 275100 218010 275152 218016
rect 275652 218068 275704 218074
rect 275652 218010 275704 218016
rect 272582 217110 272656 217138
rect 273410 217110 273484 217138
rect 274238 217246 274312 217274
rect 272582 216988 272610 217110
rect 273410 216988 273438 217110
rect 274238 216988 274266 217246
rect 275112 217138 275140 218010
rect 275848 217274 275876 224062
rect 276124 220930 276152 231662
rect 277044 230178 277072 231676
rect 277032 230172 277084 230178
rect 277032 230114 277084 230120
rect 276664 229492 276716 229498
rect 276664 229434 276716 229440
rect 276112 220924 276164 220930
rect 276112 220866 276164 220872
rect 276676 219434 276704 229434
rect 277688 224534 277716 231676
rect 278332 228954 278360 231676
rect 278320 228948 278372 228954
rect 278320 228890 278372 228896
rect 277676 224528 277728 224534
rect 277676 224470 277728 224476
rect 278976 224262 279004 231676
rect 279252 231662 279634 231690
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 278412 222896 278464 222902
rect 278412 222838 278464 222844
rect 277584 221468 277636 221474
rect 277584 221410 277636 221416
rect 276848 220108 276900 220114
rect 276848 220050 276900 220056
rect 276860 219434 276888 220050
rect 276584 219406 276704 219434
rect 276768 219406 276888 219434
rect 276584 218618 276612 219406
rect 276572 218612 276624 218618
rect 276572 218554 276624 218560
rect 276768 217274 276796 219406
rect 277596 217274 277624 221410
rect 278424 217274 278452 222838
rect 279252 219570 279280 231662
rect 280264 228682 280292 231676
rect 280448 231662 280922 231690
rect 281566 231662 281764 231690
rect 280252 228676 280304 228682
rect 280252 228618 280304 228624
rect 280068 220652 280120 220658
rect 280068 220594 280120 220600
rect 279240 219564 279292 219570
rect 279240 219506 279292 219512
rect 279240 218612 279292 218618
rect 279240 218554 279292 218560
rect 275848 217246 275922 217274
rect 275066 217110 275140 217138
rect 275066 216988 275094 217110
rect 275894 216988 275922 217246
rect 276722 217246 276796 217274
rect 277550 217246 277624 217274
rect 278378 217246 278452 217274
rect 276722 216988 276750 217246
rect 277550 216988 277578 217246
rect 278378 216988 278406 217246
rect 279252 217138 279280 218554
rect 280080 217274 280108 220594
rect 280448 220250 280476 231662
rect 280712 227860 280764 227866
rect 280712 227802 280764 227808
rect 280436 220244 280488 220250
rect 280436 220186 280488 220192
rect 280724 218754 280752 227802
rect 281448 224256 281500 224262
rect 281448 224198 281500 224204
rect 280712 218748 280764 218754
rect 280712 218690 280764 218696
rect 281460 218074 281488 224198
rect 281736 221338 281764 231662
rect 282196 229362 282224 231676
rect 282184 229356 282236 229362
rect 282184 229298 282236 229304
rect 282460 224528 282512 224534
rect 282460 224470 282512 224476
rect 281724 221332 281776 221338
rect 281724 221274 281776 221280
rect 282472 218074 282500 224470
rect 282840 223038 282868 231676
rect 283116 231662 283498 231690
rect 282828 223032 282880 223038
rect 282828 222974 282880 222980
rect 282644 222148 282696 222154
rect 282644 222090 282696 222096
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282460 218068 282512 218074
rect 282460 218010 282512 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282656 217274 282684 222090
rect 283116 220522 283144 231662
rect 283564 229900 283616 229906
rect 283564 229842 283616 229848
rect 283576 222154 283604 229842
rect 284128 225894 284156 231676
rect 284772 227866 284800 231676
rect 284760 227860 284812 227866
rect 284760 227802 284812 227808
rect 285416 227594 285444 231676
rect 285588 228676 285640 228682
rect 285588 228618 285640 228624
rect 285404 227588 285456 227594
rect 285404 227530 285456 227536
rect 284852 227044 284904 227050
rect 284852 226986 284904 226992
rect 284116 225888 284168 225894
rect 284116 225830 284168 225836
rect 283564 222148 283616 222154
rect 283564 222090 283616 222096
rect 283748 222148 283800 222154
rect 283748 222090 283800 222096
rect 283760 221474 283788 222090
rect 283748 221468 283800 221474
rect 283748 221410 283800 221416
rect 284024 221468 284076 221474
rect 284024 221410 284076 221416
rect 283104 220516 283156 220522
rect 283104 220458 283156 220464
rect 283380 220516 283432 220522
rect 283380 220458 283432 220464
rect 283392 217274 283420 220458
rect 284036 219026 284064 221410
rect 284024 219020 284076 219026
rect 284024 218962 284076 218968
rect 284864 218074 284892 226986
rect 285600 219434 285628 228618
rect 286060 222358 286088 231676
rect 286704 229094 286732 231676
rect 287348 230314 287376 231676
rect 287624 231662 288006 231690
rect 288544 231662 288650 231690
rect 287336 230308 287388 230314
rect 287336 230250 287388 230256
rect 286520 229066 286732 229094
rect 286520 224398 286548 229066
rect 286692 226160 286744 226166
rect 286692 226102 286744 226108
rect 286508 224392 286560 224398
rect 286508 224334 286560 224340
rect 286048 222352 286100 222358
rect 286048 222294 286100 222300
rect 285508 219406 285628 219434
rect 285508 218074 285536 219406
rect 285864 218884 285916 218890
rect 285864 218826 285916 218832
rect 284208 218068 284260 218074
rect 284208 218010 284260 218016
rect 284852 218068 284904 218074
rect 284852 218010 284904 218016
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282684 217274
rect 283346 217246 283420 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284220 217138 284248 218010
rect 285048 217138 285076 218010
rect 285876 217138 285904 218826
rect 286704 217274 286732 226102
rect 287624 226030 287652 231662
rect 288072 228948 288124 228954
rect 288072 228890 288124 228896
rect 287612 226024 287664 226030
rect 287612 225966 287664 225972
rect 288084 218074 288112 228890
rect 288256 225888 288308 225894
rect 288256 225830 288308 225836
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 288072 218068 288124 218074
rect 288072 218010 288124 218016
rect 284174 217110 284248 217138
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 284174 216988 284202 217110
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 225830
rect 288544 220386 288572 231662
rect 288716 229356 288768 229362
rect 288716 229298 288768 229304
rect 288728 224126 288756 229298
rect 289280 228818 289308 231676
rect 289268 228812 289320 228818
rect 289268 228754 289320 228760
rect 288716 224120 288768 224126
rect 288716 224062 288768 224068
rect 289084 223916 289136 223922
rect 289084 223858 289136 223864
rect 288532 220380 288584 220386
rect 288532 220322 288584 220328
rect 288440 219836 288492 219842
rect 288440 219778 288492 219784
rect 288452 218482 288480 219778
rect 289096 219026 289124 223858
rect 289924 221474 289952 231676
rect 290568 224670 290596 231676
rect 291226 231662 291424 231690
rect 290556 224664 290608 224670
rect 290556 224606 290608 224612
rect 291016 224392 291068 224398
rect 291016 224334 291068 224340
rect 290832 222760 290884 222766
rect 290832 222702 290884 222708
rect 289912 221468 289964 221474
rect 289912 221410 289964 221416
rect 289084 219020 289136 219026
rect 289084 218962 289136 218968
rect 288440 218476 288492 218482
rect 288440 218418 288492 218424
rect 289176 218204 289228 218210
rect 289176 218146 289228 218152
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218146
rect 290844 218074 290872 222702
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 290832 218068 290884 218074
rect 290832 218010 290884 218016
rect 290016 217138 290044 218010
rect 291028 217274 291056 224334
rect 291396 221610 291424 231662
rect 291856 223174 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 293144 228002 293172 231676
rect 293512 231662 293802 231690
rect 293132 227996 293184 228002
rect 293132 227938 293184 227944
rect 293512 223582 293540 231662
rect 293776 227588 293828 227594
rect 293776 227530 293828 227536
rect 293500 223576 293552 223582
rect 293500 223518 293552 223524
rect 291844 223168 291896 223174
rect 291844 223110 291896 223116
rect 292488 223032 292540 223038
rect 292488 222974 292540 222980
rect 291384 221604 291436 221610
rect 291384 221546 291436 221552
rect 292304 221332 292356 221338
rect 292304 221274 292356 221280
rect 292316 219298 292344 221274
rect 292304 219292 292356 219298
rect 292304 219234 292356 219240
rect 291660 218748 291712 218754
rect 291660 218690 291712 218696
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 291056 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291672 217138 291700 218690
rect 292500 217274 292528 222974
rect 293788 218074 293816 227530
rect 294432 227458 294460 231676
rect 294800 231662 295090 231690
rect 294604 230172 294656 230178
rect 294604 230114 294656 230120
rect 294420 227452 294472 227458
rect 294420 227394 294472 227400
rect 294144 219020 294196 219026
rect 294144 218962 294196 218968
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 291626 217110 291700 217138
rect 292454 217246 292528 217274
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218962
rect 294616 218210 294644 230114
rect 294800 223922 294828 231662
rect 295720 225350 295748 231676
rect 295996 231662 296378 231690
rect 295708 225344 295760 225350
rect 295708 225286 295760 225292
rect 294972 224664 295024 224670
rect 294972 224606 295024 224612
rect 294788 223916 294840 223922
rect 294788 223858 294840 223864
rect 294604 218204 294656 218210
rect 294604 218146 294656 218152
rect 294984 217274 295012 224606
rect 295996 219978 296024 231662
rect 296628 226024 296680 226030
rect 296628 225966 296680 225972
rect 296444 221468 296496 221474
rect 296444 221410 296496 221416
rect 295984 219972 296036 219978
rect 295984 219914 296036 219920
rect 296456 219434 296484 221410
rect 296456 219406 296576 219434
rect 295800 218068 295852 218074
rect 295800 218010 295852 218016
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 218010
rect 296548 217274 296576 219406
rect 296640 218090 296668 225966
rect 297008 225486 297036 231676
rect 297652 230450 297680 231676
rect 297640 230444 297692 230450
rect 297640 230386 297692 230392
rect 297364 227860 297416 227866
rect 297364 227802 297416 227808
rect 296996 225480 297048 225486
rect 296996 225422 297048 225428
rect 297180 221876 297232 221882
rect 297180 221818 297232 221824
rect 297192 221474 297220 221818
rect 297180 221468 297232 221474
rect 297180 221410 297232 221416
rect 297376 219434 297404 227802
rect 298296 227322 298324 231676
rect 298572 231662 298954 231690
rect 298284 227316 298336 227322
rect 298284 227258 298336 227264
rect 298572 221882 298600 231662
rect 299584 229090 299612 231676
rect 299952 231662 300242 231690
rect 299572 229084 299624 229090
rect 299572 229026 299624 229032
rect 298560 221876 298612 221882
rect 298560 221818 298612 221824
rect 298284 221740 298336 221746
rect 298284 221682 298336 221688
rect 297364 219428 297416 219434
rect 297364 219370 297416 219376
rect 297456 218204 297508 218210
rect 297456 218146 297508 218152
rect 296640 218074 296760 218090
rect 296640 218068 296772 218074
rect 296640 218062 296720 218068
rect 296720 218010 296772 218016
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218146
rect 298296 217274 298324 221682
rect 299952 221338 299980 231662
rect 300124 230036 300176 230042
rect 300124 229978 300176 229984
rect 299940 221332 299992 221338
rect 299940 221274 299992 221280
rect 299112 220244 299164 220250
rect 299112 220186 299164 220192
rect 299124 217274 299152 220186
rect 300136 218210 300164 229978
rect 300872 223310 300900 231676
rect 301516 227730 301544 231676
rect 301700 231662 302174 231690
rect 301504 227724 301556 227730
rect 301504 227666 301556 227672
rect 300860 223304 300912 223310
rect 300860 223246 300912 223252
rect 300768 223168 300820 223174
rect 300768 223110 300820 223116
rect 300584 219156 300636 219162
rect 300584 219098 300636 219104
rect 300124 218204 300176 218210
rect 300124 218146 300176 218152
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217246 298324 217274
rect 299078 217246 299152 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217246
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300596 217274 300624 219098
rect 300780 218074 300808 223110
rect 301700 220794 301728 231662
rect 302804 229498 302832 231676
rect 302792 229492 302844 229498
rect 302792 229434 302844 229440
rect 302148 227452 302200 227458
rect 302148 227394 302200 227400
rect 301688 220788 301740 220794
rect 301688 220730 301740 220736
rect 302160 218074 302188 227394
rect 303252 226296 303304 226302
rect 303252 226238 303304 226244
rect 302424 221468 302476 221474
rect 302424 221410 302476 221416
rect 300768 218068 300820 218074
rect 300768 218010 300820 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300596 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 221410
rect 303264 217274 303292 226238
rect 303448 224942 303476 231676
rect 303816 231662 304106 231690
rect 303436 224936 303488 224942
rect 303436 224878 303488 224884
rect 303816 221338 303844 231662
rect 304736 225758 304764 231676
rect 304908 228812 304960 228818
rect 304908 228754 304960 228760
rect 304724 225752 304776 225758
rect 304724 225694 304776 225700
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304920 219434 304948 228754
rect 305380 227866 305408 231676
rect 305644 230308 305696 230314
rect 305644 230250 305696 230256
rect 305368 227860 305420 227866
rect 305368 227802 305420 227808
rect 304828 219406 304948 219434
rect 304080 218204 304132 218210
rect 304080 218146 304132 218152
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 218146
rect 304828 217274 304856 219406
rect 305656 218210 305684 230250
rect 306024 225622 306052 231676
rect 306576 231662 306682 231690
rect 306012 225616 306064 225622
rect 306012 225558 306064 225564
rect 306196 225616 306248 225622
rect 306196 225558 306248 225564
rect 305644 218204 305696 218210
rect 305644 218146 305696 218152
rect 306208 218074 306236 225558
rect 306576 222018 306604 231662
rect 307024 223576 307076 223582
rect 307024 223518 307076 223524
rect 306564 222012 306616 222018
rect 306564 221954 306616 221960
rect 306564 221876 306616 221882
rect 306564 221818 306616 221824
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 304828 217246 304902 217274
rect 304046 217110 304120 217138
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217274 306604 221818
rect 307036 218618 307064 223518
rect 307312 223446 307340 231676
rect 307956 229770 307984 231676
rect 307944 229764 307996 229770
rect 307944 229706 307996 229712
rect 308600 228410 308628 231676
rect 308772 229084 308824 229090
rect 308772 229026 308824 229032
rect 308588 228404 308640 228410
rect 308588 228346 308640 228352
rect 307300 223440 307352 223446
rect 307300 223382 307352 223388
rect 307392 219292 307444 219298
rect 307392 219234 307444 219240
rect 307024 218612 307076 218618
rect 307024 218554 307076 218560
rect 305702 217110 305776 217138
rect 306530 217246 306604 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217246
rect 307404 217138 307432 219234
rect 308784 218074 308812 229026
rect 309244 228546 309272 231676
rect 309232 228540 309284 228546
rect 309232 228482 309284 228488
rect 309692 228268 309744 228274
rect 309692 228210 309744 228216
rect 308956 227316 309008 227322
rect 308956 227258 309008 227264
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308772 218068 308824 218074
rect 308772 218010 308824 218016
rect 308232 217138 308260 218010
rect 308968 217274 308996 227258
rect 309704 219026 309732 228210
rect 309888 224806 309916 231676
rect 310546 231662 310744 231690
rect 309876 224800 309928 224806
rect 309876 224742 309928 224748
rect 309876 220380 309928 220386
rect 309876 220322 309928 220328
rect 309692 219020 309744 219026
rect 309692 218962 309744 218968
rect 309888 217274 309916 220322
rect 310716 219842 310744 231662
rect 311176 226914 311204 231676
rect 311452 231662 311834 231690
rect 311452 229094 311480 231662
rect 311900 229628 311952 229634
rect 311900 229570 311952 229576
rect 311360 229066 311480 229094
rect 311164 226908 311216 226914
rect 311164 226850 311216 226856
rect 311360 220114 311388 229066
rect 311912 223802 311940 229570
rect 312464 227186 312492 231676
rect 313108 229362 313136 231676
rect 313096 229356 313148 229362
rect 313096 229298 313148 229304
rect 313004 228404 313056 228410
rect 313004 228346 313056 228352
rect 312452 227180 312504 227186
rect 312452 227122 312504 227128
rect 311820 223774 311940 223802
rect 311348 220108 311400 220114
rect 311348 220050 311400 220056
rect 311532 220108 311584 220114
rect 311532 220050 311584 220056
rect 310704 219836 310756 219842
rect 310704 219778 310756 219784
rect 310704 218068 310756 218074
rect 310704 218010 310756 218016
rect 308968 217246 309042 217274
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309842 217246 309916 217274
rect 309842 216988 309870 217246
rect 310716 217138 310744 218010
rect 311544 217274 311572 220050
rect 311820 218074 311848 223774
rect 313016 219434 313044 228346
rect 313188 224800 313240 224806
rect 313188 224742 313240 224748
rect 313200 219434 313228 224742
rect 313752 222902 313780 231676
rect 313936 231662 314410 231690
rect 314856 231662 315054 231690
rect 313936 229094 313964 231662
rect 313936 229066 314056 229094
rect 313740 222896 313792 222902
rect 313740 222838 313792 222844
rect 313832 220788 313884 220794
rect 313832 220730 313884 220736
rect 312360 219428 312412 219434
rect 313016 219406 313136 219434
rect 313200 219428 313332 219434
rect 313200 219406 313280 219428
rect 312360 219370 312412 219376
rect 311808 218068 311860 218074
rect 311808 218010 311860 218016
rect 310670 217110 310744 217138
rect 311498 217246 311572 217274
rect 310670 216988 310698 217110
rect 311498 216988 311526 217246
rect 312372 217138 312400 219370
rect 313108 217274 313136 219406
rect 313280 219370 313332 219376
rect 313292 219339 313320 219370
rect 313844 218890 313872 220730
rect 314028 220658 314056 229066
rect 314856 222154 314884 231662
rect 315684 223582 315712 231676
rect 316328 224534 316356 231676
rect 316604 231662 316986 231690
rect 316316 224528 316368 224534
rect 316316 224470 316368 224476
rect 315672 223576 315724 223582
rect 315672 223518 315724 223524
rect 315856 223304 315908 223310
rect 315856 223246 315908 223252
rect 315672 222896 315724 222902
rect 315672 222838 315724 222844
rect 314844 222148 314896 222154
rect 314844 222090 314896 222096
rect 314016 220652 314068 220658
rect 314016 220594 314068 220600
rect 314016 219020 314068 219026
rect 314016 218962 314068 218968
rect 313832 218884 313884 218890
rect 313832 218826 313884 218832
rect 313108 217246 313182 217274
rect 312326 217110 312400 217138
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218962
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 314856 217138 314884 218010
rect 315684 217274 315712 222838
rect 315868 218074 315896 223246
rect 316604 220522 316632 231662
rect 317144 224528 317196 224534
rect 317144 224470 317196 224476
rect 316592 220516 316644 220522
rect 316592 220458 316644 220464
rect 317156 218074 317184 224470
rect 317616 224262 317644 231676
rect 318260 229906 318288 231676
rect 318248 229900 318300 229906
rect 318248 229842 318300 229848
rect 318432 229900 318484 229906
rect 318432 229842 318484 229848
rect 318444 229094 318472 229842
rect 317984 229066 318472 229094
rect 317604 224256 317656 224262
rect 317604 224198 317656 224204
rect 317984 218074 318012 229066
rect 318904 228682 318932 231676
rect 318892 228676 318944 228682
rect 318892 228618 318944 228624
rect 319548 226166 319576 231676
rect 319812 227180 319864 227186
rect 319812 227122 319864 227128
rect 319536 226160 319588 226166
rect 319536 226102 319588 226108
rect 318156 220652 318208 220658
rect 318156 220594 318208 220600
rect 315856 218068 315908 218074
rect 315856 218010 315908 218016
rect 316500 218068 316552 218074
rect 316500 218010 316552 218016
rect 317144 218068 317196 218074
rect 317144 218010 317196 218016
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217246 315712 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217246
rect 316512 217138 316540 218010
rect 317340 217138 317368 218010
rect 318168 217274 318196 220594
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 316466 217110 316540 217138
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 316466 216988 316494 217110
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 227122
rect 320192 227050 320220 231676
rect 320376 231662 320850 231690
rect 320180 227044 320232 227050
rect 320180 226986 320232 226992
rect 319996 225752 320048 225758
rect 319996 225694 320048 225700
rect 320008 218074 320036 225694
rect 320376 220794 320404 231662
rect 321480 225894 321508 231676
rect 321848 231662 322138 231690
rect 321468 225888 321520 225894
rect 321468 225830 321520 225836
rect 321468 224936 321520 224942
rect 321468 224878 321520 224884
rect 320364 220788 320416 220794
rect 320364 220730 320416 220736
rect 320640 218612 320692 218618
rect 320640 218554 320692 218560
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 218554
rect 321480 217274 321508 224878
rect 321848 222766 321876 231662
rect 322768 228954 322796 231676
rect 323412 230178 323440 231676
rect 323584 230444 323636 230450
rect 323584 230386 323636 230392
rect 323400 230172 323452 230178
rect 323400 230114 323452 230120
rect 322756 228948 322808 228954
rect 322756 228890 322808 228896
rect 322296 224256 322348 224262
rect 322296 224198 322348 224204
rect 321836 222760 321888 222766
rect 321836 222702 321888 222708
rect 320606 217110 320680 217138
rect 321434 217246 321508 217274
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 224198
rect 322848 223440 322900 223446
rect 322848 223382 322900 223388
rect 322860 219162 322888 223382
rect 323124 219428 323176 219434
rect 323124 219370 323176 219376
rect 322848 219156 322900 219162
rect 322848 219098 322900 219104
rect 323136 217138 323164 219370
rect 323596 218754 323624 230386
rect 324056 224398 324084 231676
rect 324700 230450 324728 231676
rect 324688 230444 324740 230450
rect 324688 230386 324740 230392
rect 324964 230172 325016 230178
rect 324964 230114 325016 230120
rect 324228 225888 324280 225894
rect 324228 225830 324280 225836
rect 324044 224392 324096 224398
rect 324044 224334 324096 224340
rect 324240 219434 324268 225830
rect 324228 219428 324280 219434
rect 324228 219370 324280 219376
rect 324780 219428 324832 219434
rect 324780 219370 324832 219376
rect 323952 219292 324004 219298
rect 323952 219234 324004 219240
rect 323584 218748 323636 218754
rect 323584 218690 323636 218696
rect 323964 217138 323992 219234
rect 324792 217138 324820 219370
rect 324976 219298 325004 230114
rect 325344 227594 325372 231676
rect 325332 227588 325384 227594
rect 325332 227530 325384 227536
rect 325516 227044 325568 227050
rect 325516 226986 325568 226992
rect 325528 219434 325556 226986
rect 325988 224670 326016 231676
rect 325976 224664 326028 224670
rect 325976 224606 326028 224612
rect 326632 223038 326660 231676
rect 326896 228540 326948 228546
rect 326896 228482 326948 228488
rect 326620 223032 326672 223038
rect 326620 222974 326672 222980
rect 326908 219434 326936 228482
rect 327276 228274 327304 231676
rect 327552 231662 327934 231690
rect 327264 228268 327316 228274
rect 327264 228210 327316 228216
rect 327552 221610 327580 231662
rect 327724 228948 327776 228954
rect 327724 228890 327776 228896
rect 327540 221604 327592 221610
rect 327540 221546 327592 221552
rect 327736 219434 327764 228890
rect 328564 221746 328592 231676
rect 329208 226030 329236 231676
rect 329852 230042 329880 231676
rect 330128 231662 330510 231690
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 329196 226024 329248 226030
rect 329196 225966 329248 225972
rect 330128 223174 330156 231662
rect 331140 227458 331168 231676
rect 331416 231662 331798 231690
rect 331416 229094 331444 231662
rect 331324 229066 331444 229094
rect 331128 227452 331180 227458
rect 331128 227394 331180 227400
rect 330392 226024 330444 226030
rect 330392 225966 330444 225972
rect 330116 223168 330168 223174
rect 330116 223110 330168 223116
rect 329748 223032 329800 223038
rect 329748 222974 329800 222980
rect 328552 221740 328604 221746
rect 328552 221682 328604 221688
rect 328092 221604 328144 221610
rect 328092 221546 328144 221552
rect 325516 219428 325568 219434
rect 325516 219370 325568 219376
rect 326436 219428 326488 219434
rect 326436 219370 326488 219376
rect 326896 219428 326948 219434
rect 326896 219370 326948 219376
rect 327724 219428 327776 219434
rect 327724 219370 327776 219376
rect 324964 219292 325016 219298
rect 324964 219234 325016 219240
rect 325608 219156 325660 219162
rect 325608 219098 325660 219104
rect 325620 217138 325648 219098
rect 326448 217138 326476 219370
rect 327264 219292 327316 219298
rect 327264 219234 327316 219240
rect 327276 217274 327304 219234
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217110 323992 217138
rect 324746 217110 324820 217138
rect 325574 217110 325648 217138
rect 326402 217110 326476 217138
rect 327230 217246 327304 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217110
rect 324746 216988 324774 217110
rect 325574 216988 325602 217110
rect 326402 216988 326430 217110
rect 327230 216988 327258 217246
rect 328104 217138 328132 221546
rect 328920 220516 328972 220522
rect 328920 220458 328972 220464
rect 328932 217138 328960 220458
rect 329760 217138 329788 222974
rect 330404 219162 330432 225966
rect 330576 222012 330628 222018
rect 330576 221954 330628 221960
rect 330392 219156 330444 219162
rect 330392 219098 330444 219104
rect 330588 217138 330616 221954
rect 331324 221864 331352 229066
rect 332428 223446 332456 231676
rect 333072 226302 333100 231676
rect 333716 228818 333744 231676
rect 334084 231662 334374 231690
rect 333704 228812 333756 228818
rect 333704 228754 333756 228760
rect 333888 227452 333940 227458
rect 333888 227394 333940 227400
rect 333060 226296 333112 226302
rect 333060 226238 333112 226244
rect 332416 223440 332468 223446
rect 332416 223382 332468 223388
rect 331232 221836 331352 221864
rect 331232 220250 331260 221836
rect 331404 221740 331456 221746
rect 331404 221682 331456 221688
rect 331220 220244 331272 220250
rect 331220 220186 331272 220192
rect 331416 217274 331444 221682
rect 333704 218748 333756 218754
rect 333704 218690 333756 218696
rect 332232 218204 332284 218210
rect 332232 218146 332284 218152
rect 328058 217110 328132 217138
rect 328886 217110 328960 217138
rect 329714 217110 329788 217138
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 328058 216988 328086 217110
rect 328886 216988 328914 217110
rect 329714 216988 329742 217110
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332244 217138 332272 218146
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 333072 217138 333100 218010
rect 333716 217274 333744 218690
rect 333900 218074 333928 227394
rect 334084 221474 334112 231662
rect 335004 230314 335032 231676
rect 335464 231662 335662 231690
rect 334992 230308 335044 230314
rect 334992 230250 335044 230256
rect 335268 228812 335320 228818
rect 335268 228754 335320 228760
rect 334072 221468 334124 221474
rect 334072 221410 334124 221416
rect 334992 221468 335044 221474
rect 334992 221410 335044 221416
rect 335004 218210 335032 221410
rect 334992 218204 335044 218210
rect 334992 218146 335044 218152
rect 335280 218074 335308 228754
rect 335464 221882 335492 231662
rect 336292 229090 336320 231676
rect 336280 229084 336332 229090
rect 336280 229026 336332 229032
rect 336556 228676 336608 228682
rect 336556 228618 336608 228624
rect 336372 223168 336424 223174
rect 336372 223110 336424 223116
rect 335452 221876 335504 221882
rect 335452 221818 335504 221824
rect 336384 218074 336412 223110
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335268 218068 335320 218074
rect 335268 218010 335320 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 336372 218068 336424 218074
rect 336372 218010 336424 218016
rect 333716 217246 333882 217274
rect 332198 217110 332272 217138
rect 333026 217110 333100 217138
rect 332198 216988 332226 217110
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336568 217274 336596 228618
rect 336936 225622 336964 231676
rect 337580 228954 337608 231676
rect 338132 231662 338238 231690
rect 338408 231662 338882 231690
rect 337844 230036 337896 230042
rect 337844 229978 337896 229984
rect 337568 228948 337620 228954
rect 337568 228890 337620 228896
rect 336924 225616 336976 225622
rect 336924 225558 336976 225564
rect 337856 218074 337884 229978
rect 338132 220386 338160 231662
rect 338120 220380 338172 220386
rect 338120 220322 338172 220328
rect 338028 220244 338080 220250
rect 338028 220186 338080 220192
rect 337200 218068 337252 218074
rect 337200 218010 337252 218016
rect 337844 218068 337896 218074
rect 337844 218010 337896 218016
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336596 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218010
rect 338040 217274 338068 220186
rect 338408 220114 338436 231662
rect 339512 227322 339540 231676
rect 340156 229770 340184 231676
rect 340144 229764 340196 229770
rect 340144 229706 340196 229712
rect 340800 228410 340828 231676
rect 340788 228404 340840 228410
rect 340788 228346 340840 228352
rect 340144 228268 340196 228274
rect 340144 228210 340196 228216
rect 339500 227316 339552 227322
rect 339500 227258 339552 227264
rect 339224 220788 339276 220794
rect 339224 220730 339276 220736
rect 338396 220108 338448 220114
rect 338396 220050 338448 220056
rect 339236 219026 339264 220730
rect 339224 219020 339276 219026
rect 339224 218962 339276 218968
rect 340156 218210 340184 228210
rect 340696 225616 340748 225622
rect 340696 225558 340748 225564
rect 340512 219020 340564 219026
rect 340512 218962 340564 218968
rect 338856 218204 338908 218210
rect 338856 218146 338908 218152
rect 340144 218204 340196 218210
rect 340144 218146 340196 218152
rect 337166 217110 337240 217138
rect 337994 217246 338068 217274
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218146
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 339696 217138 339724 218010
rect 340524 217274 340552 218962
rect 340708 218074 340736 225558
rect 341444 223310 341472 231676
rect 342088 224806 342116 231676
rect 342456 231662 342746 231690
rect 343008 231662 343390 231690
rect 343836 231662 344034 231690
rect 342076 224800 342128 224806
rect 342076 224742 342128 224748
rect 341984 224392 342036 224398
rect 341984 224334 342036 224340
rect 341432 223304 341484 223310
rect 341432 223246 341484 223252
rect 341996 219434 342024 224334
rect 342168 223304 342220 223310
rect 342168 223246 342220 223252
rect 342180 219434 342208 223246
rect 342456 220794 342484 231662
rect 343008 224534 343036 231662
rect 342996 224528 343048 224534
rect 342996 224470 343048 224476
rect 343456 224528 343508 224534
rect 343456 224470 343508 224476
rect 342444 220788 342496 220794
rect 342444 220730 342496 220736
rect 342720 220108 342772 220114
rect 342720 220050 342772 220056
rect 341340 219428 341392 219434
rect 341996 219406 342116 219434
rect 342180 219428 342312 219434
rect 342180 219406 342260 219428
rect 341340 219370 341392 219376
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217246 340552 217274
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217246
rect 341352 217138 341380 219370
rect 342088 217274 342116 219406
rect 342260 219370 342312 219376
rect 342732 219298 342760 220050
rect 342720 219292 342772 219298
rect 342720 219234 342772 219240
rect 343468 218074 343496 224470
rect 343836 220658 343864 231662
rect 344664 222902 344692 231676
rect 345308 229906 345336 231676
rect 345860 231662 345966 231690
rect 345296 229900 345348 229906
rect 345296 229842 345348 229848
rect 345664 229764 345716 229770
rect 345664 229706 345716 229712
rect 344652 222896 344704 222902
rect 344652 222838 344704 222844
rect 345676 222018 345704 229706
rect 345860 227186 345888 231662
rect 345848 227180 345900 227186
rect 345848 227122 345900 227128
rect 346124 227180 346176 227186
rect 346124 227122 346176 227128
rect 345664 222012 345716 222018
rect 345664 221954 345716 221960
rect 344652 221876 344704 221882
rect 344652 221818 344704 221824
rect 343824 220652 343876 220658
rect 343824 220594 343876 220600
rect 343640 220380 343692 220386
rect 343640 220322 343692 220328
rect 343652 218890 343680 220322
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 343640 218884 343692 218890
rect 343640 218826 343692 218832
rect 342996 218068 343048 218074
rect 342996 218010 343048 218016
rect 343456 218068 343508 218074
rect 343456 218010 343508 218016
rect 342088 217246 342162 217274
rect 341306 217110 341380 217138
rect 341306 216988 341334 217110
rect 342134 216988 342162 217246
rect 343008 217138 343036 218010
rect 343836 217138 343864 219370
rect 344664 217274 344692 221818
rect 346136 219434 346164 227122
rect 346596 224942 346624 231676
rect 347240 225758 347268 231676
rect 347228 225752 347280 225758
rect 347228 225694 347280 225700
rect 346584 224936 346636 224942
rect 346584 224878 346636 224884
rect 347044 224664 347096 224670
rect 347044 224606 347096 224612
rect 346308 222896 346360 222902
rect 346308 222838 346360 222844
rect 346136 219406 346256 219434
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 342962 217110 343036 217138
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 342962 216988 342990 217110
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346228 217274 346256 219406
rect 346320 218090 346348 222838
rect 347056 219434 347084 224606
rect 347884 220386 347912 231676
rect 348528 225894 348556 231676
rect 349172 227050 349200 231676
rect 349160 227044 349212 227050
rect 349160 226986 349212 226992
rect 348516 225888 348568 225894
rect 348516 225830 348568 225836
rect 349068 225752 349120 225758
rect 349068 225694 349120 225700
rect 347872 220380 347924 220386
rect 347872 220322 347924 220328
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347136 218884 347188 218890
rect 347136 218826 347188 218832
rect 346320 218074 346440 218090
rect 346320 218068 346452 218074
rect 346320 218062 346400 218068
rect 346400 218010 346452 218016
rect 346228 217246 346302 217274
rect 345446 217110 345520 217138
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347148 217138 347176 218826
rect 348792 218204 348844 218210
rect 348792 218146 348844 218152
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 347976 217138 348004 218010
rect 348804 217138 348832 218146
rect 349080 218074 349108 225694
rect 349816 224262 349844 231676
rect 350460 230178 350488 231676
rect 350448 230172 350500 230178
rect 350448 230114 350500 230120
rect 350172 228948 350224 228954
rect 350172 228890 350224 228896
rect 349804 224256 349856 224262
rect 349804 224198 349856 224204
rect 350184 218074 350212 228890
rect 351104 228546 351132 231676
rect 351288 231662 351762 231690
rect 351932 231662 352406 231690
rect 352576 231662 353050 231690
rect 351092 228540 351144 228546
rect 351092 228482 351144 228488
rect 351092 227316 351144 227322
rect 351092 227258 351144 227264
rect 350356 226160 350408 226166
rect 350356 226102 350408 226108
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 349632 217138 349660 218010
rect 350368 217274 350396 226102
rect 351104 219026 351132 227258
rect 351288 221610 351316 231662
rect 351932 226030 351960 231662
rect 352576 229094 352604 231662
rect 352392 229066 352604 229094
rect 351920 226024 351972 226030
rect 351920 225966 351972 225972
rect 351736 224256 351788 224262
rect 351736 224198 351788 224204
rect 351276 221604 351328 221610
rect 351276 221546 351328 221552
rect 351092 219020 351144 219026
rect 351092 218962 351144 218968
rect 351748 218074 351776 224198
rect 352392 220114 352420 229066
rect 352564 226024 352616 226030
rect 352564 225966 352616 225972
rect 352380 220108 352432 220114
rect 352380 220050 352432 220056
rect 352576 218754 352604 225966
rect 353680 223038 353708 231676
rect 353864 231662 354338 231690
rect 354692 231662 354982 231690
rect 353668 223032 353720 223038
rect 353668 222974 353720 222980
rect 353864 221746 353892 231662
rect 353852 221740 353904 221746
rect 353852 221682 353904 221688
rect 353300 221604 353352 221610
rect 353300 221546 353352 221552
rect 352932 220380 352984 220386
rect 352932 220322 352984 220328
rect 352564 218748 352616 218754
rect 352564 218690 352616 218696
rect 351276 218068 351328 218074
rect 351276 218010 351328 218016
rect 351736 218068 351788 218074
rect 351736 218010 351788 218016
rect 352104 218068 352156 218074
rect 352104 218010 352156 218016
rect 350368 217246 350442 217274
rect 347102 217110 347176 217138
rect 347930 217110 348004 217138
rect 348758 217110 348832 217138
rect 349586 217110 349660 217138
rect 347102 216988 347130 217110
rect 347930 216988 347958 217110
rect 348758 216988 348786 217110
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351288 217138 351316 218010
rect 352116 217138 352144 218010
rect 352944 217274 352972 220322
rect 353312 218210 353340 221546
rect 354692 220522 354720 231662
rect 354864 230172 354916 230178
rect 354864 230114 354916 230120
rect 354876 226166 354904 230114
rect 355612 229770 355640 231676
rect 355600 229764 355652 229770
rect 355600 229706 355652 229712
rect 356256 227458 356284 231676
rect 356900 228818 356928 231676
rect 357072 229764 357124 229770
rect 357072 229706 357124 229712
rect 356888 228812 356940 228818
rect 356888 228754 356940 228760
rect 356244 227452 356296 227458
rect 356244 227394 356296 227400
rect 354864 226160 354916 226166
rect 354864 226102 354916 226108
rect 355324 225888 355376 225894
rect 355324 225830 355376 225836
rect 354680 220516 354732 220522
rect 354680 220458 354732 220464
rect 354404 220108 354456 220114
rect 354404 220050 354456 220056
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 353300 218204 353352 218210
rect 353300 218146 353352 218152
rect 351242 217110 351316 217138
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 351242 216988 351270 217110
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354416 218074 354444 220050
rect 355336 219434 355364 225830
rect 355968 223032 356020 223038
rect 355968 222974 356020 222980
rect 354588 219428 354640 219434
rect 354588 219370 354640 219376
rect 355324 219428 355376 219434
rect 355324 219370 355376 219376
rect 354404 218068 354456 218074
rect 354404 218010 354456 218016
rect 354600 217138 354628 219370
rect 355980 218074 356008 222974
rect 355416 218068 355468 218074
rect 355416 218010 355468 218016
rect 355968 218068 356020 218074
rect 355968 218010 356020 218016
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 355428 217138 355456 218010
rect 356256 217138 356284 218010
rect 357084 217274 357112 229706
rect 357256 227044 357308 227050
rect 357256 226986 357308 226992
rect 357268 218074 357296 226986
rect 357544 221474 357572 231676
rect 358188 226030 358216 231676
rect 358832 228682 358860 231676
rect 359016 231662 359490 231690
rect 359752 231662 360134 231690
rect 358820 228676 358872 228682
rect 358820 228618 358872 228624
rect 358176 226024 358228 226030
rect 358176 225966 358228 225972
rect 357532 221468 357584 221474
rect 357532 221410 357584 221416
rect 357900 221468 357952 221474
rect 357900 221410 357952 221416
rect 357256 218068 357308 218074
rect 357256 218010 357308 218016
rect 357912 217274 357940 221410
rect 359016 220250 359044 231662
rect 359752 223174 359780 231662
rect 360764 230042 360792 231676
rect 360752 230036 360804 230042
rect 360752 229978 360804 229984
rect 361212 229900 361264 229906
rect 361212 229842 361264 229848
rect 361224 229094 361252 229842
rect 361408 229094 361436 231676
rect 361224 229066 361344 229094
rect 361408 229066 361528 229094
rect 360108 228540 360160 228546
rect 360108 228482 360160 228488
rect 359740 223168 359792 223174
rect 359740 223110 359792 223116
rect 359004 220244 359056 220250
rect 359004 220186 359056 220192
rect 358728 219292 358780 219298
rect 358728 219234 358780 219240
rect 353726 217110 353800 217138
rect 354554 217110 354628 217138
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357112 217274
rect 357866 217246 357940 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217110
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357866 216988 357894 217246
rect 358740 217138 358768 219234
rect 360120 218074 360148 228482
rect 361120 220244 361172 220250
rect 361120 220186 361172 220192
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361132 217274 361160 220186
rect 361316 218074 361344 229066
rect 361500 225622 361528 229066
rect 361488 225616 361540 225622
rect 361488 225558 361540 225564
rect 362052 223310 362080 231676
rect 362696 228410 362724 231676
rect 362684 228404 362736 228410
rect 362684 228346 362736 228352
rect 362868 228404 362920 228410
rect 362868 228346 362920 228352
rect 362040 223304 362092 223310
rect 362040 223246 362092 223252
rect 362040 221740 362092 221746
rect 362040 221682 362092 221688
rect 361304 218068 361356 218074
rect 361304 218010 361356 218016
rect 362052 217274 362080 221682
rect 362880 219434 362908 228346
rect 363340 227322 363368 231676
rect 363328 227316 363380 227322
rect 363328 227258 363380 227264
rect 363512 227316 363564 227322
rect 363512 227258 363564 227264
rect 361132 217246 361206 217274
rect 358694 217110 358768 217138
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 358694 216988 358722 217110
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362006 217246 362080 217274
rect 362788 219406 362908 219434
rect 362788 217274 362816 219406
rect 363524 218890 363552 227258
rect 363984 224670 364012 231676
rect 364536 231662 364642 231690
rect 363972 224664 364024 224670
rect 363972 224606 364024 224612
rect 363788 224528 363840 224534
rect 363788 224470 363840 224476
rect 363800 219298 363828 224470
rect 364536 221882 364564 231662
rect 365272 224398 365300 231676
rect 365536 225616 365588 225622
rect 365536 225558 365588 225564
rect 365260 224392 365312 224398
rect 365260 224334 365312 224340
rect 364524 221876 364576 221882
rect 364524 221818 364576 221824
rect 363788 219292 363840 219298
rect 363788 219234 363840 219240
rect 363696 219156 363748 219162
rect 363696 219098 363748 219104
rect 363512 218884 363564 218890
rect 363512 218826 363564 218832
rect 362788 217246 362862 217274
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363708 217138 363736 219098
rect 365352 218340 365404 218346
rect 365352 218282 365404 218288
rect 364524 218068 364576 218074
rect 364524 218010 364576 218016
rect 364536 217138 364564 218010
rect 365364 217138 365392 218282
rect 365548 218074 365576 225558
rect 365916 224806 365944 231676
rect 366560 227186 366588 231676
rect 366548 227180 366600 227186
rect 366548 227122 366600 227128
rect 367204 225758 367232 231676
rect 367480 231662 367862 231690
rect 367192 225752 367244 225758
rect 367192 225694 367244 225700
rect 365904 224800 365956 224806
rect 365904 224742 365956 224748
rect 366732 223304 366784 223310
rect 366732 223246 366784 223252
rect 366744 218074 366772 223246
rect 366916 223168 366968 223174
rect 366916 223110 366968 223116
rect 365536 218068 365588 218074
rect 365536 218010 365588 218016
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366732 218068 366784 218074
rect 366732 218010 366784 218016
rect 366192 217138 366220 218010
rect 366928 217274 366956 223110
rect 367480 222902 367508 231662
rect 368492 227322 368520 231676
rect 369136 228954 369164 231676
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 368480 227316 368532 227322
rect 368480 227258 368532 227264
rect 369492 227180 369544 227186
rect 369492 227122 369544 227128
rect 367652 225004 367704 225010
rect 367652 224946 367704 224952
rect 367468 222896 367520 222902
rect 367468 222838 367520 222844
rect 367664 218754 367692 224946
rect 368388 224392 368440 224398
rect 368388 224334 368440 224340
rect 367652 218748 367704 218754
rect 367652 218690 367704 218696
rect 368400 218074 368428 224334
rect 368664 218204 368716 218210
rect 368664 218146 368716 218152
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218146
rect 369504 217274 369532 227122
rect 369780 224262 369808 231676
rect 369964 231662 370438 231690
rect 369768 224256 369820 224262
rect 369768 224198 369820 224204
rect 369964 221610 369992 231662
rect 371068 230178 371096 231676
rect 371436 231662 371726 231690
rect 371056 230172 371108 230178
rect 371056 230114 371108 230120
rect 371056 228676 371108 228682
rect 371056 228618 371108 228624
rect 369952 221604 370004 221610
rect 369952 221546 370004 221552
rect 370504 221604 370556 221610
rect 370504 221546 370556 221552
rect 370320 219020 370372 219026
rect 370320 218962 370372 218968
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370332 217138 370360 218962
rect 370516 218346 370544 221546
rect 370504 218340 370556 218346
rect 370504 218282 370556 218288
rect 371068 217274 371096 228618
rect 371436 220386 371464 231662
rect 372356 225894 372384 231676
rect 372816 231662 373014 231690
rect 372344 225888 372396 225894
rect 372344 225830 372396 225836
rect 372436 224256 372488 224262
rect 372436 224198 372488 224204
rect 371424 220380 371476 220386
rect 371424 220322 371476 220328
rect 372252 220380 372304 220386
rect 372252 220322 372304 220328
rect 372264 218210 372292 220322
rect 372252 218204 372304 218210
rect 372252 218146 372304 218152
rect 372448 218074 372476 224198
rect 372816 220114 372844 231662
rect 373644 225010 373672 231676
rect 373816 228812 373868 228818
rect 373816 228754 373868 228760
rect 373632 225004 373684 225010
rect 373632 224946 373684 224952
rect 372804 220108 372856 220114
rect 372804 220050 372856 220056
rect 373632 219428 373684 219434
rect 373632 219370 373684 219376
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372436 218068 372488 218074
rect 372436 218010 372488 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 371068 217246 371142 217274
rect 370286 217110 370360 217138
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217138 373672 219370
rect 373828 218074 373856 228754
rect 374288 227050 374316 231676
rect 374564 231662 374946 231690
rect 374276 227044 374328 227050
rect 374276 226986 374328 226992
rect 374564 221474 374592 231662
rect 375288 225752 375340 225758
rect 375288 225694 375340 225700
rect 374552 221468 374604 221474
rect 374552 221410 374604 221416
rect 374000 221196 374052 221202
rect 374000 221138 374052 221144
rect 374012 219162 374040 221138
rect 374000 219156 374052 219162
rect 374000 219098 374052 219104
rect 375104 218204 375156 218210
rect 375104 218146 375156 218152
rect 373816 218068 373868 218074
rect 373816 218010 373868 218016
rect 374460 218068 374512 218074
rect 374460 218010 374512 218016
rect 374472 217138 374500 218010
rect 375116 217274 375144 218146
rect 375300 218074 375328 225694
rect 375576 223038 375604 231676
rect 376024 230376 376076 230382
rect 376024 230318 376076 230324
rect 375564 223032 375616 223038
rect 375564 222974 375616 222980
rect 376036 221746 376064 230318
rect 376220 229770 376248 231676
rect 376208 229764 376260 229770
rect 376208 229706 376260 229712
rect 376864 228546 376892 231676
rect 377048 231662 377522 231690
rect 376852 228540 376904 228546
rect 376852 228482 376904 228488
rect 376668 227044 376720 227050
rect 376668 226986 376720 226992
rect 376024 221740 376076 221746
rect 376024 221682 376076 221688
rect 375472 221468 375524 221474
rect 375472 221410 375524 221416
rect 375484 219026 375512 221410
rect 375472 219020 375524 219026
rect 375472 218962 375524 218968
rect 376680 218074 376708 226986
rect 377048 220250 377076 231662
rect 377772 228540 377824 228546
rect 377772 228482 377824 228488
rect 377036 220244 377088 220250
rect 377036 220186 377088 220192
rect 376944 218748 376996 218754
rect 376944 218690 376996 218696
rect 375288 218068 375340 218074
rect 375288 218010 375340 218016
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 375116 217246 375282 217274
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217110 373672 217138
rect 374426 217110 374500 217138
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217110
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218690
rect 377784 217274 377812 228482
rect 378152 224534 378180 231676
rect 378796 229906 378824 231676
rect 378784 229900 378836 229906
rect 378784 229842 378836 229848
rect 379440 228410 379468 231676
rect 379808 231662 380098 231690
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 379244 228268 379296 228274
rect 379244 228210 379296 228216
rect 378140 224528 378192 224534
rect 378140 224470 378192 224476
rect 378048 220244 378100 220250
rect 378048 220186 378100 220192
rect 378060 219434 378088 220186
rect 378048 219428 378100 219434
rect 378048 219370 378100 219376
rect 379256 218074 379284 228210
rect 379808 225622 379836 231662
rect 380728 230382 380756 231676
rect 381096 231662 381386 231690
rect 380716 230376 380768 230382
rect 380716 230318 380768 230324
rect 380716 229764 380768 229770
rect 380716 229706 380768 229712
rect 379796 225616 379848 225622
rect 379796 225558 379848 225564
rect 380072 225616 380124 225622
rect 380072 225558 380124 225564
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 218210 380112 225558
rect 380072 218204 380124 218210
rect 380072 218146 380124 218152
rect 380728 218074 380756 229706
rect 381096 221202 381124 231662
rect 382016 223310 382044 231676
rect 382660 229094 382688 231676
rect 382844 231662 383318 231690
rect 382844 229094 382872 231662
rect 382568 229066 382688 229094
rect 382752 229066 382872 229094
rect 382568 224398 382596 229066
rect 382556 224392 382608 224398
rect 382556 224334 382608 224340
rect 382004 223304 382056 223310
rect 382004 223246 382056 223252
rect 382096 223032 382148 223038
rect 382096 222974 382148 222980
rect 381084 221196 381136 221202
rect 381084 221138 381136 221144
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 380256 218068 380308 218074
rect 380256 218010 380308 218016
rect 380716 218068 380768 218074
rect 380716 218010 380768 218016
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 218010
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 222974
rect 382752 221746 382780 229066
rect 382924 224392 382976 224398
rect 382924 224334 382976 224340
rect 382740 221740 382792 221746
rect 382740 221682 382792 221688
rect 382740 221604 382792 221610
rect 382740 221546 382792 221552
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217274 382780 221546
rect 382936 218210 382964 224334
rect 383948 223174 383976 231676
rect 384592 227186 384620 231676
rect 385236 228682 385264 231676
rect 385420 231662 385894 231690
rect 385224 228676 385276 228682
rect 385224 228618 385276 228624
rect 384580 227180 384632 227186
rect 384580 227122 384632 227128
rect 384948 226908 385000 226914
rect 384948 226850 385000 226856
rect 383936 223168 383988 223174
rect 383936 223110 383988 223116
rect 383568 219020 383620 219026
rect 383568 218962 383620 218968
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217246 382780 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217246
rect 383580 217138 383608 218962
rect 384960 218074 384988 226850
rect 385420 220522 385448 231662
rect 385684 227316 385736 227322
rect 385684 227258 385736 227264
rect 385408 220516 385460 220522
rect 385408 220458 385460 220464
rect 385696 218754 385724 227258
rect 386328 222896 386380 222902
rect 386328 222838 386380 222844
rect 385684 218748 385736 218754
rect 385684 218690 385736 218696
rect 386052 218748 386104 218754
rect 386052 218690 386104 218696
rect 384396 218068 384448 218074
rect 384396 218010 384448 218016
rect 384948 218068 385000 218074
rect 384948 218010 385000 218016
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 384408 217138 384436 218010
rect 385236 217138 385264 218010
rect 386064 217138 386092 218690
rect 386340 218074 386368 222838
rect 386524 221474 386552 231676
rect 387168 228818 387196 231676
rect 387340 230240 387392 230246
rect 387340 230182 387392 230188
rect 387156 228812 387208 228818
rect 387156 228754 387208 228760
rect 387352 224262 387380 230182
rect 387812 225758 387840 231676
rect 388456 230246 388484 231676
rect 388640 231662 389114 231690
rect 388444 230240 388496 230246
rect 388444 230182 388496 230188
rect 387800 225752 387852 225758
rect 387800 225694 387852 225700
rect 388444 225752 388496 225758
rect 388444 225694 388496 225700
rect 387708 224528 387760 224534
rect 387708 224470 387760 224476
rect 387340 224256 387392 224262
rect 387340 224198 387392 224204
rect 386880 222148 386932 222154
rect 386880 222090 386932 222096
rect 386512 221468 386564 221474
rect 386512 221410 386564 221416
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 386892 217274 386920 222090
rect 387720 217274 387748 224470
rect 388456 219026 388484 225694
rect 388640 220250 388668 231662
rect 389744 227050 389772 231676
rect 389916 229900 389968 229906
rect 389916 229842 389968 229848
rect 389732 227044 389784 227050
rect 389732 226986 389784 226992
rect 389928 222154 389956 229842
rect 390388 228546 390416 231676
rect 390376 228540 390428 228546
rect 390376 228482 390428 228488
rect 390100 228268 390152 228274
rect 390100 228210 390152 228216
rect 389916 222148 389968 222154
rect 389916 222090 389968 222096
rect 388628 220244 388680 220250
rect 388628 220186 388680 220192
rect 388444 219020 388496 219026
rect 388444 218962 388496 218968
rect 388536 218612 388588 218618
rect 388536 218554 388588 218560
rect 383534 217110 383608 217138
rect 384362 217110 384436 217138
rect 385190 217110 385264 217138
rect 386018 217110 386092 217138
rect 386846 217246 386920 217274
rect 387674 217246 387748 217274
rect 383534 216988 383562 217110
rect 384362 216988 384390 217110
rect 385190 216988 385218 217110
rect 386018 216988 386046 217110
rect 386846 216988 386874 217246
rect 387674 216988 387702 217246
rect 388548 217138 388576 218554
rect 390112 218074 390140 228210
rect 391032 225622 391060 231676
rect 391676 227322 391704 231676
rect 392136 231662 392334 231690
rect 391664 227316 391716 227322
rect 391664 227258 391716 227264
rect 391572 227180 391624 227186
rect 391572 227122 391624 227128
rect 391020 225616 391072 225622
rect 391020 225558 391072 225564
rect 390284 221468 390336 221474
rect 390284 221410 390336 221416
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 390100 218068 390152 218074
rect 390100 218010 390152 218016
rect 389376 217138 389404 218010
rect 390296 217274 390324 221410
rect 391584 218074 391612 227122
rect 391756 225616 391808 225622
rect 391756 225558 391808 225564
rect 391020 218068 391072 218074
rect 391020 218010 391072 218016
rect 391572 218068 391624 218074
rect 391572 218010 391624 218016
rect 388502 217110 388576 217138
rect 389330 217110 389404 217138
rect 390158 217246 390324 217274
rect 388502 216988 388530 217110
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 391032 217138 391060 218010
rect 391768 217274 391796 225558
rect 392136 220114 392164 231662
rect 392964 223038 392992 231676
rect 393608 228410 393636 231676
rect 394252 229770 394280 231676
rect 394240 229764 394292 229770
rect 394240 229706 394292 229712
rect 393596 228404 393648 228410
rect 393596 228346 393648 228352
rect 393964 227928 394016 227934
rect 393964 227870 394016 227876
rect 392952 223032 393004 223038
rect 392952 222974 393004 222980
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 392676 218884 392728 218890
rect 392676 218826 392728 218832
rect 391768 217246 391842 217274
rect 390986 217110 391060 217138
rect 390986 216988 391014 217110
rect 391814 216988 391842 217246
rect 392688 217138 392716 218826
rect 393976 218618 394004 227870
rect 394516 224256 394568 224262
rect 394516 224198 394568 224204
rect 393964 218612 394016 218618
rect 393964 218554 394016 218560
rect 394332 218204 394384 218210
rect 394332 218146 394384 218152
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 393516 217138 393544 218010
rect 394344 217138 394372 218146
rect 394528 218074 394556 224198
rect 394896 221610 394924 231676
rect 395540 226914 395568 231676
rect 395804 227044 395856 227050
rect 395804 226986 395856 226992
rect 395528 226908 395580 226914
rect 395528 226850 395580 226856
rect 394884 221604 394936 221610
rect 394884 221546 394936 221552
rect 395816 218074 395844 226986
rect 396184 224398 396212 231676
rect 396552 231662 396842 231690
rect 396552 229094 396580 231662
rect 396460 229066 396580 229094
rect 396460 225758 396488 229066
rect 397472 227798 397500 231676
rect 396632 227792 396684 227798
rect 396632 227734 396684 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396448 225752 396500 225758
rect 396448 225694 396500 225700
rect 396172 224392 396224 224398
rect 396172 224334 396224 224340
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396644 218754 396672 227734
rect 398116 224534 398144 231676
rect 398392 231662 398774 231690
rect 398392 229094 398420 231662
rect 399404 229906 399432 231676
rect 399392 229900 399444 229906
rect 399392 229842 399444 229848
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 398300 229066 398420 229094
rect 398104 224528 398156 224534
rect 398104 224470 398156 224476
rect 398300 222902 398328 229066
rect 398656 228132 398708 228138
rect 398656 228074 398708 228080
rect 398288 222896 398340 222902
rect 398288 222838 398340 222844
rect 398472 222896 398524 222902
rect 398472 222838 398524 222844
rect 396816 221604 396868 221610
rect 396816 221546 396868 221552
rect 396632 218748 396684 218754
rect 396632 218690 396684 218696
rect 396828 217274 396856 221546
rect 398484 218074 398512 222838
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 398472 218068 398524 218074
rect 398472 218010 398524 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217110 394372 217138
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217110
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397656 217138 397684 218010
rect 398668 217274 398696 228074
rect 399864 219434 399892 229706
rect 400048 228274 400076 231676
rect 400692 229094 400720 231676
rect 400600 229066 400720 229094
rect 400220 228540 400272 228546
rect 400220 228482 400272 228488
rect 400036 228268 400088 228274
rect 400036 228210 400088 228216
rect 400232 228154 400260 228482
rect 400140 228126 400260 228154
rect 400140 219434 400168 228126
rect 400600 227186 400628 229066
rect 401336 227934 401364 231676
rect 401704 231662 401994 231690
rect 401324 227928 401376 227934
rect 401324 227870 401376 227876
rect 400772 227792 400824 227798
rect 400772 227734 400824 227740
rect 400588 227180 400640 227186
rect 400588 227122 400640 227128
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 397610 217110 397684 217138
rect 398438 217246 398696 217274
rect 397610 216988 397638 217110
rect 398438 216988 398466 217246
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400784 218890 400812 227734
rect 401508 227180 401560 227186
rect 401508 227122 401560 227128
rect 400772 218884 400824 218890
rect 400772 218826 400824 218832
rect 401520 218074 401548 227122
rect 401704 221474 401732 231662
rect 402244 227928 402296 227934
rect 402244 227870 402296 227876
rect 401692 221468 401744 221474
rect 401692 221410 401744 221416
rect 401784 218884 401836 218890
rect 401784 218826 401836 218832
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 401508 218068 401560 218074
rect 401508 218010 401560 218016
rect 400048 217246 400122 217274
rect 399266 217110 399340 217138
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218826
rect 402256 218210 402284 227870
rect 402624 227798 402652 231676
rect 403268 227798 403296 231676
rect 403544 231662 403926 231690
rect 402612 227792 402664 227798
rect 402612 227734 402664 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 403544 225622 403572 231662
rect 404176 228676 404228 228682
rect 404176 228618 404228 228624
rect 403532 225616 403584 225622
rect 403532 225558 403584 225564
rect 403440 219428 403492 219434
rect 403440 219370 403492 219376
rect 402612 218748 402664 218754
rect 402612 218690 402664 218696
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402624 217138 402652 218690
rect 403452 217138 403480 219370
rect 404188 217274 404216 228618
rect 404360 225072 404412 225078
rect 404280 225020 404360 225026
rect 404280 225014 404412 225020
rect 404280 224998 404400 225014
rect 404280 219434 404308 224998
rect 404556 224262 404584 231676
rect 404740 231662 405214 231690
rect 404544 224256 404596 224262
rect 404544 224198 404596 224204
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 404280 219428 404412 219434
rect 404280 219406 404360 219428
rect 404360 219370 404412 219376
rect 405568 218074 405596 224198
rect 405844 222902 405872 231676
rect 406488 227050 406516 231676
rect 407146 231662 407344 231690
rect 406476 227044 406528 227050
rect 406476 226986 406528 226992
rect 406752 223304 406804 223310
rect 406752 223246 406804 223252
rect 405832 222896 405884 222902
rect 405832 222838 405884 222844
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223246
rect 407316 221610 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 409064 228274 409092 231676
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228404 409840 228410
rect 409788 228346 409840 228352
rect 409052 228268 409104 228274
rect 409052 228210 409104 228216
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 407304 221604 407356 221610
rect 407304 221546 407356 221552
rect 407776 218890 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218884 407816 218890
rect 407764 218826 407816 218832
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218754 409092 227734
rect 409052 218748 409104 218754
rect 409052 218690 409104 218696
rect 409800 218074 409828 228346
rect 410352 227798 410380 231676
rect 410800 229900 410852 229906
rect 410800 229842 410852 229848
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410812 219434 410840 229842
rect 410996 228682 411024 231676
rect 410984 228676 411036 228682
rect 410984 228618 411036 228624
rect 410984 228540 411036 228546
rect 410984 228482 411036 228488
rect 410996 219434 411024 228482
rect 411640 226370 411668 231676
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411628 226364 411680 226370
rect 411628 226306 411680 226312
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 225078 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 225072 412324 225078
rect 412272 225014 412324 225020
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 230240 413888 230246
rect 413836 230182 413888 230188
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 230182
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223310 414888 231676
rect 415504 228410 415532 231676
rect 416148 228546 416176 231676
rect 416792 229094 416820 231676
rect 417436 229906 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229900 417476 229906
rect 417424 229842 417476 229848
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416136 228540 416188 228546
rect 416136 228482 416188 228488
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416688 227792 416740 227798
rect 416688 227734 416740 227740
rect 415032 224052 415084 224058
rect 415032 223994 415084 224000
rect 414848 223304 414900 223310
rect 414848 223246 414900 223252
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 223994
rect 416504 223576 416556 223582
rect 416504 223518 416556 223524
rect 416516 219434 416544 223518
rect 416700 219434 416728 227734
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 220794 418384 231662
rect 419368 227050 419396 231676
rect 420012 230246 420040 231676
rect 420000 230240 420052 230246
rect 420000 230182 420052 230188
rect 419632 229152 419684 229158
rect 419632 229094 419684 229100
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 419448 226908 419500 226914
rect 419448 226850 419500 226856
rect 418344 220788 418396 220794
rect 418344 220730 418396 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 419172 219156 419224 219162
rect 419172 219098 419224 219104
rect 418344 218068 418396 218074
rect 418344 218010 418396 218016
rect 418356 217138 418384 218010
rect 419184 217138 419212 219098
rect 419460 218074 419488 226850
rect 419644 224058 419672 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 224256 420880 224262
rect 420828 224198 420880 224204
rect 419632 224052 419684 224058
rect 419632 223994 419684 224000
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 420656 219434 420684 220798
rect 420656 219406 420776 219434
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 224198
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 223582 422248 229066
rect 422208 223576 422260 223582
rect 422208 223518 422260 223524
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 220862 423904 231676
rect 424520 226914 424548 231676
rect 424508 226908 424560 226914
rect 424508 226850 424560 226856
rect 425164 224262 425192 231676
rect 425440 231662 425822 231690
rect 425152 224256 425204 224262
rect 425152 224198 425204 224204
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 423864 220856 423916 220862
rect 423864 220798 423916 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219162 422708 219406
rect 422668 219156 422720 219162
rect 422668 219098 422720 219104
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 417482 217110 417556 217138
rect 418310 217110 418384 217138
rect 419138 217110 419212 217138
rect 419966 217110 420040 217138
rect 417482 216988 417510 217110
rect 418310 216988 418338 217110
rect 419138 216988 419166 217110
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 224942 426480 231676
rect 426820 231662 427110 231690
rect 426440 224936 426492 224942
rect 426440 224878 426492 224884
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 426992 224936 427044 224942
rect 426992 224878 427044 224884
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 224878
rect 427912 220176 427964 220182
rect 427912 220118 427964 220124
rect 427924 218074 427952 220118
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 219370
rect 428476 218210 428504 229066
rect 428752 220182 428780 231662
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 428740 220176 428792 220182
rect 428740 220118 428792 220124
rect 429948 219434 429976 231662
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220244 432288 220250
rect 432236 220186 432288 220192
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220186
rect 429580 219406 429976 219434
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 431972 219406 432276 219434
rect 429580 218346 429608 219406
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217138 429148 218010
rect 429948 217138 429976 218690
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 219406
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220250 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436416 231690
rect 434812 220244 434864 220250
rect 434812 220186 434864 220192
rect 435284 218210 435312 231662
rect 436388 224398 436416 231662
rect 436572 231662 436770 231690
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436572 229094 436600 231662
rect 436572 229066 436692 229094
rect 436376 224392 436428 224398
rect 436376 224334 436428 224340
rect 436284 224256 436336 224262
rect 436284 224198 436336 224204
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218204 435784 218210
rect 435732 218146 435784 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434904 218068 434956 218074
rect 434904 218010 434956 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218010
rect 435744 217138 435772 218146
rect 436296 218074 436324 224198
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436468 218068 436520 218074
rect 436468 218010 436520 218016
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436480 217138 436508 218010
rect 436664 217546 436692 229066
rect 436836 224392 436888 224398
rect 436836 224334 436888 224340
rect 436848 218210 436876 224334
rect 437032 224262 437060 231662
rect 437020 224256 437072 224262
rect 437020 224198 437072 224204
rect 436836 218204 436888 218210
rect 436836 218146 436888 218152
rect 437768 218074 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 224954 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 224954 439360 230318
rect 438872 224926 438992 224954
rect 439056 224926 439360 224954
rect 438872 219434 438900 224926
rect 438216 219428 438268 219434
rect 438216 219370 438268 219376
rect 438860 219428 438912 219434
rect 438860 219370 438912 219376
rect 437756 218068 437808 218074
rect 437756 218010 437808 218016
rect 436664 217518 437336 217546
rect 437308 217274 437336 217518
rect 437308 217246 437382 217274
rect 436480 217110 436554 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217246
rect 438228 217138 438256 219370
rect 439056 217274 439084 224926
rect 440344 219434 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 219428 439924 219434
rect 439872 219370 439924 219376
rect 440332 219428 440384 219434
rect 440332 219370 440384 219376
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 219370
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443210 231662 443408 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 224954 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 224926 441752 224954
rect 441632 218090 441660 224926
rect 441540 218062 441660 218090
rect 441540 217274 441568 218062
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441494 217246 441568 217274
rect 442276 217274 442304 229066
rect 443380 224954 443408 231662
rect 443552 230444 443604 230450
rect 443552 230386 443604 230392
rect 443564 229094 443592 230386
rect 443840 230246 443868 231676
rect 444484 230450 444512 231676
rect 444668 231662 445142 231690
rect 444472 230444 444524 230450
rect 444472 230386 444524 230392
rect 444668 230330 444696 231662
rect 444484 230302 444696 230330
rect 443828 230240 443880 230246
rect 443828 230182 443880 230188
rect 443564 229066 443960 229094
rect 443196 224926 443408 224954
rect 443196 217274 443224 224926
rect 442276 217246 442350 217274
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441494 216988 441522 217246
rect 442322 216988 442350 217246
rect 443150 217246 443224 217274
rect 443932 217274 443960 229066
rect 444484 224954 444512 230302
rect 444656 230240 444708 230246
rect 444656 230182 444708 230188
rect 444668 224954 444696 230182
rect 445772 224954 445800 231676
rect 446416 229158 446444 231676
rect 446404 229152 446456 229158
rect 446404 229094 446456 229100
rect 447060 227934 447088 231676
rect 447244 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 444484 224926 444604 224954
rect 444668 224926 445616 224954
rect 445772 224926 446444 224954
rect 444576 217274 444604 224926
rect 445588 217274 445616 224926
rect 446416 217274 446444 224926
rect 447244 219434 447272 231662
rect 447600 230444 447652 230450
rect 447600 230386 447652 230392
rect 447612 219434 447640 230386
rect 448348 229294 448376 231676
rect 448992 229566 449020 231676
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448336 229288 448388 229294
rect 448336 229230 448388 229236
rect 449636 229158 449664 231676
rect 450280 229294 450308 231676
rect 450924 229430 450952 231676
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 449808 229288 449860 229294
rect 449808 229230 449860 229236
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 448520 229152 448572 229158
rect 448520 229094 448572 229100
rect 449624 229152 449676 229158
rect 449624 229094 449676 229100
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 448532 219434 448560 229094
rect 449820 224954 449848 229230
rect 451568 229158 451596 231676
rect 452226 231662 452608 231690
rect 452200 229560 452252 229566
rect 452200 229502 452252 229508
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 450728 229152 450780 229158
rect 450728 229094 450780 229100
rect 451556 229152 451608 229158
rect 451556 229094 451608 229100
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 449728 224926 449848 224954
rect 448532 219406 448652 219434
rect 443932 217246 444006 217274
rect 444576 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448624 217274 448652 219406
rect 449728 217274 449756 224926
rect 450556 217274 450584 227870
rect 450740 218346 450768 229094
rect 451752 219434 451780 229230
rect 451476 219406 451780 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448624 217246 448974 217274
rect 449728 217246 449802 217274
rect 450556 217246 450630 217274
rect 448106 217194 448158 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449774 216988 449802 217246
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229502
rect 452580 222154 452608 231662
rect 452856 229294 452884 231676
rect 453500 229430 453528 231676
rect 453028 229424 453080 229430
rect 453028 229366 453080 229372
rect 453488 229424 453540 229430
rect 453488 229366 453540 229372
rect 452844 229288 452896 229294
rect 452844 229230 452896 229236
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229366
rect 454144 229158 454172 231676
rect 454788 229378 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455788 229424 455840 229430
rect 454788 229350 454908 229378
rect 455788 229366 455840 229372
rect 454684 229288 454736 229294
rect 454684 229230 454736 229236
rect 453304 229152 453356 229158
rect 453304 229094 453356 229100
rect 454132 229152 454184 229158
rect 454132 229094 454184 229100
rect 453316 218074 453344 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229230
rect 454880 223582 454908 229350
rect 455328 229152 455380 229158
rect 455328 229094 455380 229100
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220726 455368 229094
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220720 455380 220726
rect 455328 220662 455380 220668
rect 455616 218074 455644 222090
rect 455800 219434 455828 229366
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220862 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220856 456760 220862
rect 456708 220798 456760 220804
rect 457180 219434 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 458824 220720 458876 220726
rect 458824 220662 458876 220668
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220662
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 224942 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224936 460624 224942
rect 460572 224878 460624 224884
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224398 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224392 462556 224398
rect 462504 224334 462556 224340
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 225762
rect 463160 225078 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225072 463200 225078
rect 463148 225014 463200 225020
rect 463148 224936 463200 224942
rect 463148 224878 463200 224884
rect 463160 218074 463188 224878
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 230042 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 230036 465500 230042
rect 465448 229978 465500 229984
rect 465736 220794 465764 230318
rect 465920 226506 465948 231662
rect 466104 231662 466394 231690
rect 467038 231662 467328 231690
rect 465908 226500 465960 226506
rect 465908 226442 465960 226448
rect 465724 220788 465776 220794
rect 465724 220730 465776 220736
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466104 219162 466132 231662
rect 467300 222902 467328 231662
rect 467668 225622 467696 231676
rect 468312 230450 468340 231676
rect 468864 231662 468970 231690
rect 468300 230444 468352 230450
rect 468300 230386 468352 230392
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 225072 467524 225078
rect 467472 225014 467524 225020
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 467288 222896 467340 222902
rect 467288 222838 467340 222844
rect 466092 219156 466144 219162
rect 466092 219098 466144 219104
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467484 219434 467512 225014
rect 468668 222148 468720 222154
rect 468668 222090 468720 222096
rect 467300 219406 467512 219434
rect 468680 219434 468708 222090
rect 468864 220250 468892 231662
rect 469036 230444 469088 230450
rect 469036 230386 469088 230392
rect 469048 221610 469076 230386
rect 469312 224392 469364 224398
rect 469312 224334 469364 224340
rect 469036 221604 469088 221610
rect 469036 221546 469088 221552
rect 468852 220244 468904 220250
rect 468852 220186 468904 220192
rect 468680 219406 468800 219434
rect 467300 218074 467328 219406
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 219406
rect 468772 217246 468846 217274
rect 469324 217258 469352 224334
rect 469600 224262 469628 231676
rect 470244 228410 470272 231676
rect 470888 230246 470916 231676
rect 470876 230240 470928 230246
rect 470876 230182 470928 230188
rect 470232 228404 470284 228410
rect 470232 228346 470284 228352
rect 471532 226982 471560 231676
rect 472176 230450 472204 231676
rect 472834 231662 473308 231690
rect 472164 230444 472216 230450
rect 472164 230386 472216 230392
rect 473084 230444 473136 230450
rect 473084 230386 473136 230392
rect 471888 230240 471940 230246
rect 471888 230182 471940 230188
rect 471520 226976 471572 226982
rect 471520 226918 471572 226924
rect 469864 226500 469916 226506
rect 469864 226442 469916 226448
rect 469588 224256 469640 224262
rect 469588 224198 469640 224204
rect 469588 220788 469640 220794
rect 469588 220730 469640 220736
rect 469600 217274 469628 220730
rect 469876 218618 469904 226442
rect 471900 220794 471928 230182
rect 473096 221474 473124 230386
rect 473084 221468 473136 221474
rect 473084 221410 473136 221416
rect 471888 220788 471940 220794
rect 471888 220730 471940 220736
rect 473280 220114 473308 231662
rect 473464 230382 473492 231676
rect 473452 230376 473504 230382
rect 473452 230318 473504 230324
rect 474108 230246 474136 231676
rect 474556 230376 474608 230382
rect 474556 230318 474608 230324
rect 474096 230240 474148 230246
rect 474096 230182 474148 230188
rect 473728 230036 473780 230042
rect 473728 229978 473780 229984
rect 473268 220108 473320 220114
rect 473268 220050 473320 220056
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 472084 217274 472112 219574
rect 472900 219156 472952 219162
rect 472900 219098 472952 219104
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 219098
rect 473740 217274 473768 229978
rect 474568 222170 474596 230318
rect 474752 227798 474780 231676
rect 475410 231662 475792 231690
rect 474740 227792 474792 227798
rect 474740 227734 474792 227740
rect 475384 222896 475436 222902
rect 475384 222838 475436 222844
rect 474568 222142 474780 222170
rect 474556 221604 474608 221610
rect 474556 221546 474608 221552
rect 474568 217274 474596 221546
rect 474752 218618 474780 222142
rect 474740 218612 474792 218618
rect 474740 218554 474792 218560
rect 475396 217274 475424 222838
rect 475764 221746 475792 231662
rect 476040 225758 476068 231676
rect 476028 225752 476080 225758
rect 476028 225694 476080 225700
rect 476684 222902 476712 231676
rect 477328 230382 477356 231676
rect 477316 230376 477368 230382
rect 477316 230318 477368 230324
rect 477408 230240 477460 230246
rect 477408 230182 477460 230188
rect 477420 227322 477448 230182
rect 477408 227316 477460 227322
rect 477408 227258 477460 227264
rect 477040 225616 477092 225622
rect 477040 225558 477092 225564
rect 476672 222896 476724 222902
rect 476672 222838 476724 222844
rect 475752 221740 475804 221746
rect 475752 221682 475804 221688
rect 476212 220244 476264 220250
rect 476212 220186 476264 220192
rect 476224 217274 476252 220186
rect 477052 217274 477080 225558
rect 477592 224256 477644 224262
rect 477592 224198 477644 224204
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 477052 217246 477126 217274
rect 477604 217258 477632 224198
rect 477972 223174 478000 231676
rect 478616 224398 478644 231676
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 479708 228404 479760 228410
rect 479708 228346 479760 228352
rect 479524 226976 479576 226982
rect 479524 226918 479576 226924
rect 478604 224392 478656 224398
rect 478604 224334 478656 224340
rect 477960 223168 478012 223174
rect 477960 223110 478012 223116
rect 477868 220788 477920 220794
rect 477868 220730 477920 220736
rect 477880 217274 477908 220730
rect 479536 217274 479564 226918
rect 479720 219298 479748 228346
rect 479904 226914 479932 231676
rect 480548 230382 480576 231676
rect 480076 230376 480128 230382
rect 480076 230318 480128 230324
rect 480536 230376 480588 230382
rect 480536 230318 480588 230324
rect 480088 228546 480116 230318
rect 480076 228540 480128 228546
rect 480076 228482 480128 228488
rect 479892 226908 479944 226914
rect 479892 226850 479944 226856
rect 481192 225622 481220 231676
rect 481548 230376 481600 230382
rect 481548 230318 481600 230324
rect 481180 225616 481232 225622
rect 481180 225558 481232 225564
rect 481180 221468 481232 221474
rect 481180 221410 481232 221416
rect 479708 219292 479760 219298
rect 479708 219234 479760 219240
rect 480352 219292 480404 219298
rect 480352 219234 480404 219240
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477592 217252 477644 217258
rect 477880 217246 477954 217274
rect 477592 217194 477644 217200
rect 477926 216988 477954 217246
rect 478742 217252 478794 217258
rect 479536 217246 479610 217274
rect 478742 217194 478794 217200
rect 478754 216988 478782 217194
rect 479582 216988 479610 217246
rect 480364 217138 480392 219234
rect 481192 217274 481220 221410
rect 481560 220250 481588 230318
rect 481836 228410 481864 231676
rect 482494 231662 482784 231690
rect 481824 228404 481876 228410
rect 481824 228346 481876 228352
rect 481548 220244 481600 220250
rect 481548 220186 481600 220192
rect 482756 220114 482784 231662
rect 482928 227792 482980 227798
rect 482928 227734 482980 227740
rect 482940 222494 482968 227734
rect 483124 223038 483152 231676
rect 483768 227186 483796 231676
rect 484412 229974 484440 231676
rect 484400 229968 484452 229974
rect 484400 229910 484452 229916
rect 485056 228818 485084 231676
rect 485516 231662 485714 231690
rect 485044 228812 485096 228818
rect 485044 228754 485096 228760
rect 485044 227316 485096 227322
rect 485044 227258 485096 227264
rect 483756 227180 483808 227186
rect 483756 227122 483808 227128
rect 483572 225752 483624 225758
rect 483572 225694 483624 225700
rect 483112 223032 483164 223038
rect 483112 222974 483164 222980
rect 482928 222488 482980 222494
rect 482928 222430 482980 222436
rect 482008 220108 482060 220114
rect 482008 220050 482060 220056
rect 482744 220108 482796 220114
rect 482744 220050 482796 220056
rect 482020 217274 482048 220050
rect 482940 218754 482968 222430
rect 482928 218748 482980 218754
rect 482928 218690 482980 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480364 217110 480438 217138
rect 480410 216988 480438 217110
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483584 218074 483612 225694
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 483572 218068 483624 218074
rect 483572 218010 483624 218016
rect 483768 217274 483796 221410
rect 485056 218113 485084 227258
rect 485516 221610 485544 231662
rect 486344 230110 486372 231676
rect 486896 231662 487002 231690
rect 487646 231662 488212 231690
rect 486332 230104 486384 230110
rect 486332 230046 486384 230052
rect 486896 228682 486924 231662
rect 487068 230104 487120 230110
rect 487068 230046 487120 230052
rect 486884 228676 486936 228682
rect 486884 228618 486936 228624
rect 487080 221746 487108 230046
rect 488184 229094 488212 231662
rect 488092 229066 488212 229094
rect 487804 222896 487856 222902
rect 487804 222838 487856 222844
rect 486148 221740 486200 221746
rect 486148 221682 486200 221688
rect 487068 221740 487120 221746
rect 487068 221682 487120 221688
rect 485504 221604 485556 221610
rect 485504 221546 485556 221552
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 484582 218104 484638 218113
rect 484582 218039 484638 218048
rect 485042 218104 485098 218113
rect 485042 218039 485098 218048
rect 483722 217246 483796 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484596 217138 484624 218039
rect 484550 217110 484624 217138
rect 485332 217138 485360 218690
rect 486160 217138 486188 221682
rect 487816 218385 487844 222838
rect 488092 220522 488120 229066
rect 488276 222902 488304 231676
rect 488920 224262 488948 231676
rect 489184 228540 489236 228546
rect 489184 228482 489236 228488
rect 489196 224954 489224 228482
rect 489564 225758 489592 231676
rect 490208 230110 490236 231676
rect 490196 230104 490248 230110
rect 490196 230046 490248 230052
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 489552 225752 489604 225758
rect 489552 225694 489604 225700
rect 489104 224926 489224 224954
rect 488908 224256 488960 224262
rect 488908 224198 488960 224204
rect 488264 222896 488316 222902
rect 488264 222838 488316 222844
rect 488080 220516 488132 220522
rect 488080 220458 488132 220464
rect 487802 218376 487858 218385
rect 487802 218311 487858 218320
rect 486976 218068 487028 218074
rect 486976 218010 487028 218016
rect 486988 217138 487016 218010
rect 487816 217138 487844 218311
rect 489104 217274 489132 224926
rect 489932 224058 489960 229706
rect 490852 227322 490880 231676
rect 490840 227316 490892 227322
rect 490840 227258 490892 227264
rect 491496 227050 491524 231676
rect 491484 227044 491536 227050
rect 491484 226986 491536 226992
rect 491944 226908 491996 226914
rect 491944 226850 491996 226856
rect 490288 224392 490340 224398
rect 490288 224334 490340 224340
rect 489920 224052 489972 224058
rect 489920 223994 489972 224000
rect 489460 223168 489512 223174
rect 489460 223110 489512 223116
rect 488690 217246 489132 217274
rect 485332 217110 485406 217138
rect 486160 217110 486234 217138
rect 486988 217110 487062 217138
rect 487816 217110 487890 217138
rect 484550 216988 484578 217110
rect 485378 216988 485406 217110
rect 486206 216988 486234 217110
rect 487034 216988 487062 217110
rect 487862 216988 487890 217110
rect 488690 216988 488718 217246
rect 489104 217161 489132 217246
rect 489090 217152 489146 217161
rect 489472 217138 489500 223110
rect 490300 218657 490328 224334
rect 491116 224052 491168 224058
rect 491116 223994 491168 224000
rect 491128 223650 491156 223994
rect 491116 223644 491168 223650
rect 491116 223586 491168 223592
rect 490286 218648 490342 218657
rect 490286 218583 490342 218592
rect 490300 217138 490328 218583
rect 491128 217274 491156 223586
rect 491956 219473 491984 226850
rect 492140 224398 492168 231676
rect 492784 225486 492812 231676
rect 493442 231662 494008 231690
rect 494086 231662 494376 231690
rect 494730 231662 495204 231690
rect 493692 225616 493744 225622
rect 493692 225558 493744 225564
rect 492772 225480 492824 225486
rect 492772 225422 492824 225428
rect 492128 224392 492180 224398
rect 492128 224334 492180 224340
rect 492772 220244 492824 220250
rect 492772 220186 492824 220192
rect 491942 219464 491998 219473
rect 491942 219399 491998 219408
rect 491956 217274 491984 219399
rect 491128 217246 491202 217274
rect 491956 217246 492030 217274
rect 489472 217110 489546 217138
rect 490300 217110 490374 217138
rect 489090 217087 489146 217096
rect 489518 216988 489546 217110
rect 490346 216988 490374 217110
rect 491174 216988 491202 217246
rect 492002 216988 492030 217246
rect 492784 217138 492812 220186
rect 493704 218929 493732 225558
rect 493980 220386 494008 231662
rect 494348 229770 494376 231662
rect 494336 229764 494388 229770
rect 494336 229706 494388 229712
rect 494704 228404 494756 228410
rect 494704 228346 494756 228352
rect 493968 220380 494020 220386
rect 493968 220322 494020 220328
rect 494716 219201 494744 228346
rect 495176 220250 495204 231662
rect 495360 228546 495388 231676
rect 495348 228540 495400 228546
rect 495348 228482 495400 228488
rect 496004 225894 496032 231676
rect 495992 225888 496044 225894
rect 495992 225830 496044 225836
rect 496648 223174 496676 231676
rect 496820 229968 496872 229974
rect 496820 229910 496872 229916
rect 496832 223786 496860 229910
rect 497292 228410 497320 231676
rect 497936 229294 497964 231676
rect 497924 229288 497976 229294
rect 497924 229230 497976 229236
rect 497280 228404 497332 228410
rect 497280 228346 497332 228352
rect 498580 227186 498608 231676
rect 498752 228812 498804 228818
rect 498752 228754 498804 228760
rect 497556 227180 497608 227186
rect 497556 227122 497608 227128
rect 498568 227180 498620 227186
rect 498568 227122 498620 227128
rect 496820 223780 496872 223786
rect 496820 223722 496872 223728
rect 497372 223780 497424 223786
rect 497372 223722 497424 223728
rect 496636 223168 496688 223174
rect 496636 223110 496688 223116
rect 496084 223032 496136 223038
rect 496084 222974 496136 222980
rect 495164 220244 495216 220250
rect 495164 220186 495216 220192
rect 495256 220108 495308 220114
rect 495256 220050 495308 220056
rect 494702 219192 494758 219201
rect 494532 219150 494702 219178
rect 493690 218920 493746 218929
rect 493690 218855 493746 218864
rect 493704 217274 493732 218855
rect 494532 217274 494560 219150
rect 494702 219127 494758 219136
rect 495268 217297 495296 220050
rect 493658 217246 493732 217274
rect 494486 217246 494560 217274
rect 495254 217288 495310 217297
rect 492784 217110 492858 217138
rect 492830 216988 492858 217110
rect 493658 216988 493686 217246
rect 494486 216988 494514 217246
rect 496096 217274 496124 222974
rect 497002 218648 497058 218657
rect 497002 218583 497058 218592
rect 497016 217274 497044 218583
rect 497384 217546 497412 223722
rect 497568 218657 497596 227122
rect 498764 219434 498792 228754
rect 499224 224670 499252 231676
rect 499868 230382 499896 231676
rect 500052 231662 500526 231690
rect 499856 230376 499908 230382
rect 499856 230318 499908 230324
rect 500052 225298 500080 231662
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 500236 229094 500264 229230
rect 500236 229066 500448 229094
rect 500052 225270 500264 225298
rect 499212 224664 499264 224670
rect 499212 224606 499264 224612
rect 500040 221740 500092 221746
rect 500040 221682 500092 221688
rect 499396 221604 499448 221610
rect 499396 221546 499448 221552
rect 498672 219406 498792 219434
rect 497554 218648 497610 218657
rect 497554 218583 497610 218592
rect 498672 218210 498700 219406
rect 499210 218920 499266 218929
rect 499210 218855 499266 218864
rect 498660 218204 498712 218210
rect 498660 218146 498712 218152
rect 497384 217518 497780 217546
rect 496096 217246 496170 217274
rect 495254 217223 495310 217232
rect 495268 217138 495296 217223
rect 495268 217110 495342 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217246
rect 496970 217246 497044 217274
rect 497752 217274 497780 217518
rect 498672 217274 498700 218146
rect 499224 217841 499252 218855
rect 499210 217832 499266 217841
rect 499210 217767 499266 217776
rect 497752 217246 497826 217274
rect 496970 216988 496998 217246
rect 497798 216988 497826 217246
rect 498626 217246 498700 217274
rect 499408 217274 499436 221546
rect 499580 218884 499632 218890
rect 499580 218826 499632 218832
rect 499592 218385 499620 218826
rect 500052 218482 500080 221682
rect 500236 221610 500264 225270
rect 500224 221604 500276 221610
rect 500224 221546 500276 221552
rect 500420 220386 500448 229066
rect 500960 228676 501012 228682
rect 500960 228618 501012 228624
rect 500408 220380 500460 220386
rect 500408 220322 500460 220328
rect 500972 219434 501000 228618
rect 501156 226166 501184 231676
rect 501800 230382 501828 231676
rect 501604 230376 501656 230382
rect 501604 230318 501656 230324
rect 501788 230376 501840 230382
rect 501788 230318 501840 230324
rect 501144 226160 501196 226166
rect 501144 226102 501196 226108
rect 501616 221746 501644 230318
rect 502444 223038 502472 231676
rect 503102 231662 503392 231690
rect 502984 224256 503036 224262
rect 502984 224198 503036 224204
rect 502432 223032 502484 223038
rect 502432 222974 502484 222980
rect 501604 221740 501656 221746
rect 501604 221682 501656 221688
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 500972 219406 501092 219434
rect 500040 218476 500092 218482
rect 500040 218418 500092 218424
rect 500224 218476 500276 218482
rect 500224 218418 500276 218424
rect 499578 218376 499634 218385
rect 499578 218311 499634 218320
rect 499762 218376 499818 218385
rect 499762 218311 499818 218320
rect 499776 217841 499804 218311
rect 499762 217832 499818 217841
rect 499762 217767 499818 217776
rect 499408 217246 499482 217274
rect 498626 216988 498654 217246
rect 499454 216988 499482 217246
rect 500236 217138 500264 218418
rect 501064 217569 501092 219406
rect 501050 217560 501106 217569
rect 501050 217495 501106 217504
rect 501064 217138 501092 217495
rect 501892 217274 501920 220458
rect 502800 218748 502852 218754
rect 502800 218690 502852 218696
rect 501892 217246 501966 217274
rect 500236 217110 500310 217138
rect 501064 217110 501138 217138
rect 500282 216988 500310 217110
rect 501110 216988 501138 217110
rect 501938 216988 501966 217246
rect 502812 217138 502840 218690
rect 502996 217569 503024 224198
rect 503168 222896 503220 222902
rect 503168 222838 503220 222844
rect 503180 218754 503208 222838
rect 503364 222766 503392 231662
rect 503732 230178 503760 231676
rect 503720 230172 503772 230178
rect 503720 230114 503772 230120
rect 504180 225752 504232 225758
rect 504180 225694 504232 225700
rect 503352 222760 503404 222766
rect 503352 222702 503404 222708
rect 504192 219434 504220 225694
rect 504376 224262 504404 231676
rect 505020 224534 505048 231676
rect 505664 230042 505692 231676
rect 505652 230036 505704 230042
rect 505652 229978 505704 229984
rect 505744 229900 505796 229906
rect 505744 229842 505796 229848
rect 505468 227316 505520 227322
rect 505468 227258 505520 227264
rect 505008 224528 505060 224534
rect 505008 224470 505060 224476
rect 504364 224256 504416 224262
rect 504364 224198 504416 224204
rect 504192 219406 504404 219434
rect 503168 218748 503220 218754
rect 503168 218690 503220 218696
rect 503628 218204 503680 218210
rect 503628 218146 503680 218152
rect 503640 217569 503668 218146
rect 502982 217560 503038 217569
rect 502982 217495 503038 217504
rect 503350 217560 503406 217569
rect 503350 217495 503406 217504
rect 503626 217560 503682 217569
rect 503626 217495 503682 217504
rect 503364 217274 503392 217495
rect 504376 217274 504404 219406
rect 505098 219192 505154 219201
rect 505098 219127 505154 219136
rect 505282 219192 505338 219201
rect 505282 219127 505338 219136
rect 505112 219026 505140 219127
rect 505100 219020 505152 219026
rect 505100 218962 505152 218968
rect 505296 218890 505324 219127
rect 505284 218884 505336 218890
rect 505284 218826 505336 218832
rect 505284 218748 505336 218754
rect 505284 218690 505336 218696
rect 505296 218210 505324 218690
rect 505284 218204 505336 218210
rect 505284 218146 505336 218152
rect 503364 217246 503622 217274
rect 504376 217246 504450 217274
rect 502766 217110 502840 217138
rect 502766 216988 502794 217110
rect 503594 216988 503622 217246
rect 504422 216988 504450 217246
rect 505296 217138 505324 218146
rect 505480 217569 505508 227258
rect 505756 218754 505784 229842
rect 506308 228682 506336 231676
rect 506296 228676 506348 228682
rect 506296 228618 506348 228624
rect 506952 227322 506980 231676
rect 506940 227316 506992 227322
rect 506940 227258 506992 227264
rect 506848 227044 506900 227050
rect 506848 226986 506900 226992
rect 505744 218748 505796 218754
rect 505744 218690 505796 218696
rect 505466 217560 505522 217569
rect 505466 217495 505522 217504
rect 506110 217560 506166 217569
rect 506110 217495 506166 217504
rect 506124 217138 506152 217495
rect 506860 217308 506888 226986
rect 507596 222902 507624 231676
rect 508240 229022 508268 231676
rect 508504 230376 508556 230382
rect 508504 230318 508556 230324
rect 508228 229016 508280 229022
rect 508228 228958 508280 228964
rect 507768 224392 507820 224398
rect 507768 224334 507820 224340
rect 507584 222896 507636 222902
rect 507584 222838 507636 222844
rect 507780 217841 507808 224334
rect 508516 220658 508544 230318
rect 508884 225622 508912 231676
rect 509528 230382 509556 231676
rect 509516 230376 509568 230382
rect 509516 230318 509568 230324
rect 509884 229764 509936 229770
rect 509884 229706 509936 229712
rect 508872 225616 508924 225622
rect 508872 225558 508924 225564
rect 508688 225480 508740 225486
rect 508688 225422 508740 225428
rect 508504 220652 508556 220658
rect 508504 220594 508556 220600
rect 507766 217832 507822 217841
rect 507766 217767 507822 217776
rect 506860 217280 506934 217308
rect 505250 217110 505324 217138
rect 506078 217110 506152 217138
rect 505250 216988 505278 217110
rect 506078 216988 506106 217110
rect 506906 216988 506934 217280
rect 507780 217138 507808 217767
rect 508700 217569 508728 225422
rect 509896 224954 509924 229706
rect 510172 225758 510200 231676
rect 510816 229974 510844 231676
rect 510804 229968 510856 229974
rect 510804 229910 510856 229916
rect 511460 228546 511488 231676
rect 511816 229968 511868 229974
rect 511816 229910 511868 229916
rect 510620 228540 510672 228546
rect 510620 228482 510672 228488
rect 511448 228540 511500 228546
rect 511448 228482 511500 228488
rect 510160 225752 510212 225758
rect 510160 225694 510212 225700
rect 509896 224926 510200 224954
rect 509332 220244 509384 220250
rect 509332 220186 509384 220192
rect 508686 217560 508742 217569
rect 508686 217495 508742 217504
rect 508700 217308 508728 217495
rect 507734 217110 507808 217138
rect 508562 217280 508728 217308
rect 507734 216988 507762 217110
rect 508562 216988 508590 217280
rect 509344 217138 509372 220186
rect 510172 218346 510200 224926
rect 510160 218340 510212 218346
rect 510160 218282 510212 218288
rect 510172 217308 510200 218282
rect 510172 217280 510246 217308
rect 509344 217110 509418 217138
rect 509390 216988 509418 217110
rect 510218 216988 510246 217280
rect 510632 217258 510660 228482
rect 511828 220114 511856 229910
rect 512104 227050 512132 231676
rect 512762 231662 513144 231690
rect 512644 230172 512696 230178
rect 512644 230114 512696 230120
rect 512092 227044 512144 227050
rect 512092 226986 512144 226992
rect 512460 225888 512512 225894
rect 512460 225830 512512 225836
rect 512472 223922 512500 225830
rect 512460 223916 512512 223922
rect 512460 223858 512512 223864
rect 510988 220108 511040 220114
rect 510988 220050 511040 220056
rect 511816 220108 511868 220114
rect 511816 220050 511868 220056
rect 511000 217841 511028 220050
rect 510986 217832 511042 217841
rect 510986 217767 511042 217776
rect 510620 217252 510672 217258
rect 510620 217194 510672 217200
rect 511000 217138 511028 217767
rect 512472 217308 512500 223858
rect 512656 221882 512684 230114
rect 513116 223310 513144 231662
rect 513392 229226 513420 231676
rect 513380 229220 513432 229226
rect 513380 229162 513432 229168
rect 514036 227458 514064 231676
rect 514300 228404 514352 228410
rect 514300 228346 514352 228352
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 513104 223304 513156 223310
rect 513104 223246 513156 223252
rect 513564 223168 513616 223174
rect 513564 223110 513616 223116
rect 513576 222057 513604 223110
rect 513562 222048 513618 222057
rect 513562 221983 513618 221992
rect 512644 221876 512696 221882
rect 512644 221818 512696 221824
rect 513576 217308 513604 221983
rect 512472 217280 512730 217308
rect 511862 217252 511914 217258
rect 511862 217194 511914 217200
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217194
rect 512702 216988 512730 217280
rect 513530 217280 513604 217308
rect 514312 217308 514340 228346
rect 514680 224398 514708 231676
rect 515324 230178 515352 231676
rect 515312 230172 515364 230178
rect 515312 230114 515364 230120
rect 515404 229832 515456 229838
rect 515404 229774 515456 229780
rect 515416 227594 515444 229774
rect 515404 227588 515456 227594
rect 515404 227530 515456 227536
rect 515772 227180 515824 227186
rect 515772 227122 515824 227128
rect 514668 224392 514720 224398
rect 514668 224334 514720 224340
rect 515784 221241 515812 227122
rect 515968 226030 515996 231676
rect 516626 231662 517192 231690
rect 517270 231662 517468 231690
rect 515956 226024 516008 226030
rect 515956 225966 516008 225972
rect 516784 224664 516836 224670
rect 516784 224606 516836 224612
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 515128 220380 515180 220386
rect 515128 220322 515180 220328
rect 515140 217841 515168 220322
rect 515784 219434 515812 221167
rect 515784 219406 516088 219434
rect 514942 217832 514998 217841
rect 514942 217767 514944 217776
rect 514996 217767 514998 217776
rect 515126 217832 515182 217841
rect 515126 217767 515182 217776
rect 514944 217738 514996 217744
rect 515140 217308 515168 217767
rect 516060 217308 516088 219406
rect 514312 217280 514386 217308
rect 515140 217280 515214 217308
rect 513530 216988 513558 217280
rect 514358 216988 514386 217280
rect 515186 216988 515214 217280
rect 516014 217280 516088 217308
rect 516796 217308 516824 224606
rect 517164 220386 517192 231662
rect 517440 229362 517468 231662
rect 517428 229356 517480 229362
rect 517428 229298 517480 229304
rect 517900 228954 517928 231676
rect 518164 230376 518216 230382
rect 518164 230318 518216 230324
rect 517888 228948 517940 228954
rect 517888 228890 517940 228896
rect 517704 221740 517756 221746
rect 517704 221682 517756 221688
rect 517520 221604 517572 221610
rect 517520 221546 517572 221552
rect 517532 220969 517560 221546
rect 517518 220960 517574 220969
rect 517518 220895 517574 220904
rect 517152 220380 517204 220386
rect 517152 220322 517204 220328
rect 517716 217666 517744 221682
rect 518176 221610 518204 230318
rect 518544 224670 518572 231676
rect 519188 229906 519216 231676
rect 519176 229900 519228 229906
rect 519176 229842 519228 229848
rect 519544 229220 519596 229226
rect 519544 229162 519596 229168
rect 519268 226160 519320 226166
rect 519268 226102 519320 226108
rect 518532 224664 518584 224670
rect 518532 224606 518584 224612
rect 518164 221604 518216 221610
rect 518164 221546 518216 221552
rect 518530 220960 518586 220969
rect 518530 220895 518586 220904
rect 518346 217832 518402 217841
rect 518346 217767 518402 217776
rect 517704 217660 517756 217666
rect 517704 217602 517756 217608
rect 517716 217308 517744 217602
rect 518360 217530 518388 217767
rect 518348 217524 518400 217530
rect 518348 217466 518400 217472
rect 518544 217308 518572 220895
rect 518898 219736 518954 219745
rect 518898 219671 518954 219680
rect 518912 218958 518940 219671
rect 518900 218952 518952 218958
rect 518900 218894 518952 218900
rect 519084 218816 519136 218822
rect 519084 218758 519136 218764
rect 519096 218113 519124 218758
rect 518898 218104 518954 218113
rect 518898 218039 518954 218048
rect 519082 218104 519138 218113
rect 519082 218039 519138 218048
rect 518912 217938 518940 218039
rect 518900 217932 518952 217938
rect 518900 217874 518952 217880
rect 518714 217832 518770 217841
rect 518714 217767 518716 217776
rect 518768 217767 518770 217776
rect 518900 217796 518952 217802
rect 518716 217738 518768 217744
rect 518900 217738 518952 217744
rect 518912 217569 518940 217738
rect 518898 217560 518954 217569
rect 518898 217495 518954 217504
rect 519082 217560 519138 217569
rect 519082 217495 519084 217504
rect 519136 217495 519138 217504
rect 519084 217466 519136 217472
rect 516796 217280 516870 217308
rect 516014 216988 516042 217280
rect 516842 216988 516870 217280
rect 517670 217280 517744 217308
rect 518498 217280 518572 217308
rect 519280 217308 519308 226102
rect 519556 220522 519584 229162
rect 519832 223174 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 520280 229356 520332 229362
rect 520280 229298 520332 229304
rect 520292 223446 520320 229298
rect 521120 229294 521148 231676
rect 521476 230376 521528 230382
rect 521476 230318 521528 230324
rect 521108 229288 521160 229294
rect 521108 229230 521160 229236
rect 520280 223440 520332 223446
rect 520280 223382 520332 223388
rect 519820 223168 519872 223174
rect 519820 223110 519872 223116
rect 521016 223032 521068 223038
rect 521016 222974 521068 222980
rect 521028 221513 521056 222974
rect 521014 221504 521070 221513
rect 521014 221439 521070 221448
rect 520188 220652 520240 220658
rect 520188 220594 520240 220600
rect 519544 220516 519596 220522
rect 519544 220458 519596 220464
rect 519452 218952 519504 218958
rect 519452 218894 519504 218900
rect 519464 218074 519492 218894
rect 520200 218074 520228 220594
rect 519452 218068 519504 218074
rect 519452 218010 519504 218016
rect 520188 218068 520240 218074
rect 520188 218010 520240 218016
rect 519280 217280 519354 217308
rect 517670 216988 517698 217280
rect 518498 216988 518526 217280
rect 519326 216988 519354 217280
rect 520200 217138 520228 218010
rect 521028 217308 521056 221439
rect 521488 220658 521516 230318
rect 521764 228410 521792 231676
rect 522422 231662 522896 231690
rect 521752 228404 521804 228410
rect 521752 228346 521804 228352
rect 521844 222760 521896 222766
rect 521844 222702 521896 222708
rect 521476 220652 521528 220658
rect 521476 220594 521528 220600
rect 521856 217308 521884 222702
rect 522580 221876 522632 221882
rect 522580 221818 522632 221824
rect 522592 220561 522620 221818
rect 522868 221746 522896 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523316 229084 523368 229090
rect 523316 229026 523368 229032
rect 523328 228274 523356 229026
rect 523316 228268 523368 228274
rect 523316 228210 523368 228216
rect 523696 224534 523724 231676
rect 524340 225894 524368 231676
rect 524984 229158 525012 231676
rect 525156 230172 525208 230178
rect 525156 230114 525208 230120
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524972 227588 525024 227594
rect 524972 227530 525024 227536
rect 524328 225888 524380 225894
rect 524328 225830 524380 225836
rect 523040 224528 523092 224534
rect 523040 224470 523092 224476
rect 523684 224528 523736 224534
rect 523684 224470 523736 224476
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 522578 220552 522634 220561
rect 522578 220487 522634 220496
rect 520154 217110 520228 217138
rect 520982 217280 521056 217308
rect 521810 217280 521884 217308
rect 522592 217308 522620 220487
rect 522592 217280 522666 217308
rect 520154 216988 520182 217110
rect 520982 216988 521010 217280
rect 521810 216988 521838 217280
rect 522638 216988 522666 217280
rect 523052 217258 523080 224470
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 217308 523540 224198
rect 524984 220017 525012 227530
rect 525168 221882 525196 230114
rect 525628 227186 525656 231676
rect 526272 228818 526300 231676
rect 526916 229634 526944 231676
rect 526904 229628 526956 229634
rect 526904 229570 526956 229576
rect 526444 229288 526496 229294
rect 526444 229230 526496 229236
rect 526260 228812 526312 228818
rect 526260 228754 526312 228760
rect 526456 227594 526484 229230
rect 526628 228676 526680 228682
rect 526628 228618 526680 228624
rect 526444 227588 526496 227594
rect 526444 227530 526496 227536
rect 526352 227316 526404 227322
rect 526352 227258 526404 227264
rect 525616 227180 525668 227186
rect 525616 227122 525668 227128
rect 526364 224954 526392 227258
rect 526640 224954 526668 228618
rect 526364 224926 526576 224954
rect 526640 224926 526760 224954
rect 525156 221876 525208 221882
rect 525156 221818 525208 221824
rect 524970 220008 525026 220017
rect 524970 219943 525026 219952
rect 524788 218952 524840 218958
rect 524788 218894 524840 218900
rect 524420 218816 524472 218822
rect 524420 218758 524472 218764
rect 524432 218113 524460 218758
rect 524418 218104 524474 218113
rect 524418 218039 524474 218048
rect 524602 218104 524658 218113
rect 524800 218074 524828 218894
rect 524602 218039 524658 218048
rect 524788 218068 524840 218074
rect 524616 217938 524644 218039
rect 524788 218010 524840 218016
rect 524604 217932 524656 217938
rect 524604 217874 524656 217880
rect 523466 217280 523540 217308
rect 523040 217252 523092 217258
rect 523040 217194 523092 217200
rect 523466 217122 523494 217280
rect 524984 217274 525012 219943
rect 525984 217864 526036 217870
rect 525984 217806 526036 217812
rect 524282 217252 524334 217258
rect 524984 217246 525150 217274
rect 524282 217194 524334 217200
rect 523454 217116 523506 217122
rect 523454 217058 523506 217064
rect 523466 216988 523494 217058
rect 524294 216988 524322 217194
rect 525122 216988 525150 217246
rect 525996 217138 526024 217806
rect 526548 217274 526576 224926
rect 526732 217870 526760 224926
rect 527560 223038 527588 231676
rect 527732 228268 527784 228274
rect 527732 228210 527784 228216
rect 527548 223032 527600 223038
rect 527548 222974 527600 222980
rect 527548 222896 527600 222902
rect 527548 222838 527600 222844
rect 527560 220289 527588 222838
rect 527546 220280 527602 220289
rect 527546 220215 527602 220224
rect 526720 217864 526772 217870
rect 526720 217806 526772 217812
rect 526732 217598 526760 217806
rect 526720 217592 526772 217598
rect 526720 217534 526772 217540
rect 526548 217246 526806 217274
rect 525950 217110 526024 217138
rect 525950 216988 525978 217110
rect 526778 216988 526806 217246
rect 527560 217138 527588 220215
rect 527744 219434 527772 228210
rect 528204 227322 528232 231676
rect 528848 230042 528876 231676
rect 528836 230036 528888 230042
rect 528836 229978 528888 229984
rect 529204 229900 529256 229906
rect 529204 229842 529256 229848
rect 529216 229094 529244 229842
rect 529032 229066 529244 229094
rect 528192 227316 528244 227322
rect 528192 227258 528244 227264
rect 529032 219910 529060 229066
rect 529492 225622 529520 231676
rect 530136 230382 530164 231676
rect 530124 230376 530176 230382
rect 530124 230318 530176 230324
rect 530780 230246 530808 231676
rect 531228 230376 531280 230382
rect 531228 230318 531280 230324
rect 530768 230240 530820 230246
rect 530768 230182 530820 230188
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 226166 529980 229094
rect 529940 226160 529992 226166
rect 529940 226102 529992 226108
rect 530860 225752 530912 225758
rect 530860 225694 530912 225700
rect 529204 225616 529256 225622
rect 529204 225558 529256 225564
rect 529480 225616 529532 225622
rect 529480 225558 529532 225564
rect 529020 219904 529072 219910
rect 529020 219846 529072 219852
rect 528466 219736 528522 219745
rect 528466 219671 528522 219680
rect 527732 219428 527784 219434
rect 527732 219370 527784 219376
rect 528284 219428 528336 219434
rect 528284 219370 528336 219376
rect 528296 217734 528324 219370
rect 528480 218958 528508 219671
rect 528468 218952 528520 218958
rect 528468 218894 528520 218900
rect 528284 217728 528336 217734
rect 528284 217670 528336 217676
rect 528296 217274 528324 217670
rect 529216 217274 529244 225558
rect 530872 221785 530900 225694
rect 530858 221776 530914 221785
rect 530858 221711 530914 221720
rect 530032 221604 530084 221610
rect 530032 221546 530084 221552
rect 530044 220017 530072 221546
rect 530030 220008 530086 220017
rect 530030 219943 530086 219952
rect 528296 217246 528462 217274
rect 529216 217246 529290 217274
rect 527560 217110 527634 217138
rect 527606 216988 527634 217110
rect 528434 216988 528462 217246
rect 529262 216988 529290 217246
rect 530044 217138 530072 219943
rect 530872 217274 530900 221711
rect 531240 221610 531268 230318
rect 531424 228682 531452 231676
rect 532082 231662 532464 231690
rect 531412 228676 531464 228682
rect 531412 228618 531464 228624
rect 531964 228540 532016 228546
rect 531964 228482 532016 228488
rect 531228 221604 531280 221610
rect 531228 221546 531280 221552
rect 531688 220108 531740 220114
rect 531688 220050 531740 220056
rect 531700 217274 531728 220050
rect 531976 219162 532004 228482
rect 532436 222902 532464 231662
rect 532712 230178 532740 231676
rect 533370 231662 533752 231690
rect 533528 230308 533580 230314
rect 533528 230250 533580 230256
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 533540 230042 533568 230250
rect 533528 230036 533580 230042
rect 533528 229978 533580 229984
rect 533436 227044 533488 227050
rect 533436 226986 533488 226992
rect 533448 224954 533476 226986
rect 533356 224926 533476 224954
rect 532424 222896 532476 222902
rect 532424 222838 532476 222844
rect 531964 219156 532016 219162
rect 531964 219098 532016 219104
rect 532516 219156 532568 219162
rect 532516 219098 532568 219104
rect 530872 217246 530946 217274
rect 531700 217246 531774 217274
rect 530044 217110 530118 217138
rect 530090 216988 530118 217110
rect 530918 216988 530946 217246
rect 531746 216988 531774 217246
rect 532528 217138 532556 219098
rect 533356 217258 533384 224926
rect 533724 224262 533752 231662
rect 534000 225758 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534908 229764 534960 229770
rect 534908 229706 534960 229712
rect 534724 229628 534776 229634
rect 534724 229570 534776 229576
rect 533988 225752 534040 225758
rect 533988 225694 534040 225700
rect 533712 224256 533764 224262
rect 533712 224198 533764 224204
rect 534540 223304 534592 223310
rect 534540 223246 534592 223252
rect 534356 220516 534408 220522
rect 534356 220458 534408 220464
rect 534368 220114 534396 220458
rect 534356 220108 534408 220114
rect 534356 220050 534408 220056
rect 534552 219450 534580 223246
rect 534736 220522 534764 229570
rect 534920 221338 534948 229706
rect 535288 227050 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 227044 535328 227050
rect 535276 226986 535328 226992
rect 535748 224954 535776 227394
rect 535932 224954 535960 231676
rect 536576 229906 536604 231676
rect 536944 231662 537234 231690
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 535748 224926 535868 224954
rect 535932 224926 536052 224954
rect 535644 224392 535696 224398
rect 535644 224334 535696 224340
rect 535656 224058 535684 224334
rect 535840 224210 535868 224926
rect 536024 224398 536052 224926
rect 536012 224392 536064 224398
rect 536012 224334 536064 224340
rect 535840 224182 535960 224210
rect 535644 224052 535696 224058
rect 535644 223994 535696 224000
rect 534908 221332 534960 221338
rect 534908 221274 534960 221280
rect 534724 220516 534776 220522
rect 534724 220458 534776 220464
rect 535000 220108 535052 220114
rect 535000 220050 535052 220056
rect 534552 219422 534672 219450
rect 533712 219292 533764 219298
rect 533712 219234 533764 219240
rect 534448 219292 534500 219298
rect 534448 219234 534500 219240
rect 533724 219167 533752 219234
rect 533894 219192 533950 219201
rect 533710 219158 533766 219167
rect 533894 219127 533950 219136
rect 534078 219192 534134 219201
rect 534078 219127 534134 219136
rect 534262 219192 534318 219201
rect 534262 219127 534264 219136
rect 533710 219093 533766 219102
rect 533908 218822 533936 219127
rect 534092 219026 534120 219127
rect 534316 219127 534318 219136
rect 534264 219098 534316 219104
rect 534080 219020 534132 219026
rect 534080 218962 534132 218968
rect 534460 218890 534488 219234
rect 534448 218884 534500 218890
rect 534448 218826 534500 218832
rect 533896 218816 533948 218822
rect 533896 218758 533948 218764
rect 534080 218748 534132 218754
rect 534080 218690 534132 218696
rect 534092 218006 534120 218690
rect 534080 218000 534132 218006
rect 534080 217942 534132 217948
rect 534172 217864 534224 217870
rect 534172 217806 534224 217812
rect 534184 217462 534212 217806
rect 534172 217456 534224 217462
rect 534172 217398 534224 217404
rect 534644 217274 534672 219422
rect 533344 217252 533396 217258
rect 533344 217194 533396 217200
rect 534230 217246 534672 217274
rect 533356 217138 533384 217194
rect 532528 217110 532602 217138
rect 533356 217110 533430 217138
rect 532574 216988 532602 217110
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535012 217138 535040 220050
rect 535932 217394 535960 224182
rect 536656 224052 536708 224058
rect 536656 223994 536708 224000
rect 535920 217388 535972 217394
rect 535920 217330 535972 217336
rect 535932 217274 535960 217330
rect 535886 217246 535960 217274
rect 535012 217110 535086 217138
rect 535058 216988 535086 217110
rect 535886 216988 535914 217246
rect 536668 217138 536696 223994
rect 536944 220250 536972 231662
rect 537864 228546 537892 231676
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 537852 228540 537904 228546
rect 537852 228482 537904 228488
rect 537484 221876 537536 221882
rect 537484 221818 537536 221824
rect 536932 220244 536984 220250
rect 536932 220186 536984 220192
rect 537496 219162 537524 221818
rect 538784 221474 538812 231662
rect 543004 230444 543056 230450
rect 543004 230386 543056 230392
rect 541256 230308 541308 230314
rect 541256 230250 541308 230256
rect 540796 228948 540848 228954
rect 540796 228890 540848 228896
rect 538956 226024 539008 226030
rect 538956 225966 539008 225972
rect 538772 221468 538824 221474
rect 538772 221410 538824 221416
rect 537484 219156 537536 219162
rect 537484 219098 537536 219104
rect 537496 217138 537524 219098
rect 538968 218006 538996 225966
rect 540808 224954 540836 228890
rect 540808 224926 540928 224954
rect 539968 223440 540020 223446
rect 539968 223382 540020 223388
rect 539232 220380 539284 220386
rect 539232 220322 539284 220328
rect 538404 218000 538456 218006
rect 538404 217942 538456 217948
rect 538956 218000 539008 218006
rect 538956 217942 539008 217948
rect 538416 217138 538444 217942
rect 539048 217728 539100 217734
rect 539048 217670 539100 217676
rect 538680 217388 538732 217394
rect 538680 217330 538732 217336
rect 538692 217274 538720 217330
rect 539060 217326 539088 217670
rect 539048 217320 539100 217326
rect 538692 217246 538904 217274
rect 539048 217262 539100 217268
rect 536668 217110 536742 217138
rect 537496 217110 537570 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217110
rect 538370 217110 538444 217138
rect 538876 217138 538904 217246
rect 539048 217184 539100 217190
rect 538876 217132 539048 217138
rect 539244 217138 539272 220322
rect 539980 219638 540008 223382
rect 540900 221474 540928 224926
rect 541268 223310 541296 230250
rect 541624 224664 541676 224670
rect 541624 224606 541676 224612
rect 541256 223304 541308 223310
rect 541256 223246 541308 223252
rect 540888 221468 540940 221474
rect 540888 221410 540940 221416
rect 539968 219632 540020 219638
rect 539968 219574 540020 219580
rect 539692 219156 539744 219162
rect 539692 219098 539744 219104
rect 539704 218074 539732 219098
rect 539692 218068 539744 218074
rect 539692 218010 539744 218016
rect 539508 218000 539560 218006
rect 539508 217942 539560 217948
rect 539520 217734 539548 217942
rect 539508 217728 539560 217734
rect 539508 217670 539560 217676
rect 538876 217126 539100 217132
rect 538876 217110 539088 217126
rect 539198 217110 539272 217138
rect 539980 217138 540008 219574
rect 540900 217274 540928 221410
rect 540854 217246 540928 217274
rect 539980 217110 540054 217138
rect 538370 216988 538398 217110
rect 539198 216988 539226 217110
rect 540026 216988 540054 217110
rect 540854 216988 540882 217246
rect 541636 217138 541664 224606
rect 542360 223168 542412 223174
rect 542360 223110 542412 223116
rect 542372 221202 542400 223110
rect 543016 222086 543044 230386
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 545764 228404 545816 228410
rect 545764 228346 545816 228352
rect 544384 227588 544436 227594
rect 544384 227530 544436 227536
rect 543004 222080 543056 222086
rect 543004 222022 543056 222028
rect 542360 221196 542412 221202
rect 542360 221138 542412 221144
rect 543280 221196 543332 221202
rect 543280 221138 543332 221144
rect 542544 219904 542596 219910
rect 542544 219846 542596 219852
rect 542556 217138 542584 219846
rect 541636 217110 541710 217138
rect 541682 216988 541710 217110
rect 542510 217110 542584 217138
rect 543292 217138 543320 221138
rect 544108 220652 544160 220658
rect 544108 220594 544160 220600
rect 544120 217274 544148 220594
rect 544396 219162 544424 227530
rect 545776 221066 545804 228346
rect 547156 221882 547184 230114
rect 552204 230036 552256 230042
rect 552204 229978 552256 229984
rect 550640 228812 550692 228818
rect 550640 228754 550692 228760
rect 549904 226160 549956 226166
rect 549904 226102 549956 226108
rect 547880 225888 547932 225894
rect 547880 225830 547932 225836
rect 547144 221876 547196 221882
rect 547144 221818 547196 221824
rect 546592 221740 546644 221746
rect 546592 221682 546644 221688
rect 545764 221060 545816 221066
rect 545764 221002 545816 221008
rect 544384 219156 544436 219162
rect 544384 219098 544436 219104
rect 545028 219156 545080 219162
rect 545028 219098 545080 219104
rect 544120 217246 544194 217274
rect 543292 217110 543366 217138
rect 542510 216988 542538 217110
rect 543338 216988 543366 217110
rect 544166 216988 544194 217246
rect 545040 217138 545068 219098
rect 545776 217274 545804 221002
rect 546604 217274 546632 221682
rect 546776 221332 546828 221338
rect 546776 221274 546828 221280
rect 546788 219774 546816 221274
rect 546776 219768 546828 219774
rect 546776 219710 546828 219716
rect 547420 219768 547472 219774
rect 547420 219710 547472 219716
rect 547432 217274 547460 219710
rect 547892 219298 547920 225830
rect 548340 224528 548392 224534
rect 548340 224470 548392 224476
rect 548352 221746 548380 224470
rect 548340 221740 548392 221746
rect 548340 221682 548392 221688
rect 548156 219428 548208 219434
rect 548156 219370 548208 219376
rect 547880 219292 547932 219298
rect 547880 219234 547932 219240
rect 548168 219162 548196 219370
rect 548156 219156 548208 219162
rect 548156 219098 548208 219104
rect 548352 217274 548380 221682
rect 549916 219298 549944 226102
rect 549076 219292 549128 219298
rect 549076 219234 549128 219240
rect 549904 219292 549956 219298
rect 549904 219234 549956 219240
rect 548708 219020 548760 219026
rect 548708 218962 548760 218968
rect 548720 218754 548748 218962
rect 548708 218748 548760 218754
rect 548708 218690 548760 218696
rect 545776 217246 545850 217274
rect 546604 217246 546678 217274
rect 547432 217246 547506 217274
rect 544994 217110 545068 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217246
rect 546650 216988 546678 217246
rect 547478 216988 547506 217246
rect 548306 217246 548380 217274
rect 548306 216988 548334 217246
rect 549088 217138 549116 219234
rect 549916 217274 549944 219234
rect 550652 218618 550680 228754
rect 550824 227180 550876 227186
rect 550824 227122 550876 227128
rect 550836 222222 550864 227122
rect 552216 223174 552244 229978
rect 554056 228410 554084 249047
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244594 554544 244695
rect 554504 244588 554556 244594
rect 554504 244530 554556 244536
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 554044 228404 554096 228410
rect 554044 228346 554096 228352
rect 554044 227316 554096 227322
rect 554044 227258 554096 227264
rect 552204 223168 552256 223174
rect 552204 223110 552256 223116
rect 553308 223032 553360 223038
rect 553308 222974 553360 222980
rect 550824 222216 550876 222222
rect 550824 222158 550876 222164
rect 550640 218612 550692 218618
rect 550640 218554 550692 218560
rect 550836 217274 550864 222158
rect 553320 221746 553348 222974
rect 553032 221740 553084 221746
rect 553032 221682 553084 221688
rect 553308 221740 553360 221746
rect 553308 221682 553360 221688
rect 552848 221264 552900 221270
rect 552848 221206 552900 221212
rect 552860 220998 552888 221206
rect 553044 220998 553072 221682
rect 552848 220992 552900 220998
rect 552848 220934 552900 220940
rect 553032 220992 553084 220998
rect 553032 220934 553084 220940
rect 552480 220788 552532 220794
rect 552480 220730 552532 220736
rect 552492 220522 552520 220730
rect 552480 220516 552532 220522
rect 552480 220458 552532 220464
rect 551560 218612 551612 218618
rect 551560 218554 551612 218560
rect 549916 217246 549990 217274
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 216988 549990 217246
rect 550790 217246 550864 217274
rect 550790 216988 550818 217246
rect 551572 217138 551600 218554
rect 552492 217274 552520 220458
rect 553124 220380 553176 220386
rect 553124 220322 553176 220328
rect 553136 219473 553164 220322
rect 553122 219464 553178 219473
rect 552664 219428 552716 219434
rect 553122 219399 553178 219408
rect 552664 219370 552716 219376
rect 552676 218618 552704 219370
rect 552664 218612 552716 218618
rect 552664 218554 552716 218560
rect 553320 217274 553348 221682
rect 553676 220584 553728 220590
rect 553676 220526 553728 220532
rect 553688 218890 553716 220526
rect 553860 219360 553912 219366
rect 553860 219302 553912 219308
rect 553872 218890 553900 219302
rect 553676 218884 553728 218890
rect 553676 218826 553728 218832
rect 553860 218884 553912 218890
rect 553860 218826 553912 218832
rect 552446 217246 552520 217274
rect 553274 217246 553348 217274
rect 554056 217274 554084 227258
rect 555436 225894 555464 251194
rect 556816 230042 556844 255274
rect 558184 246356 558236 246362
rect 558184 246298 558236 246304
rect 558196 236094 558224 246298
rect 559564 244588 559616 244594
rect 559564 244530 559616 244536
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 556804 230036 556856 230042
rect 556804 229978 556856 229984
rect 556988 229900 557040 229906
rect 556988 229842 557040 229848
rect 555424 225888 555476 225894
rect 555424 225830 555476 225836
rect 555884 225616 555936 225622
rect 555884 225558 555936 225564
rect 555896 224954 555924 225558
rect 555804 224926 555924 224954
rect 554872 223304 554924 223310
rect 554872 223246 554924 223252
rect 554228 220380 554280 220386
rect 554228 220322 554280 220328
rect 554240 219201 554268 220322
rect 554226 219192 554282 219201
rect 554884 219162 554912 223246
rect 555424 220380 555476 220386
rect 555424 220322 555476 220328
rect 555436 219774 555464 220322
rect 555804 219842 555832 224926
rect 556068 222352 556120 222358
rect 556068 222294 556120 222300
rect 556080 222018 556108 222294
rect 556068 222012 556120 222018
rect 556068 221954 556120 221960
rect 556252 222012 556304 222018
rect 556252 221954 556304 221960
rect 556264 219978 556292 221954
rect 557000 221610 557028 229842
rect 558276 228676 558328 228682
rect 558276 228618 558328 228624
rect 558288 224954 558316 228618
rect 558288 224926 558684 224954
rect 558656 222766 558684 224926
rect 559576 222902 559604 244530
rect 560956 227594 560984 256702
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 560944 227588 560996 227594
rect 560944 227530 560996 227536
rect 561496 225752 561548 225758
rect 561496 225694 561548 225700
rect 561312 224256 561364 224262
rect 561312 224198 561364 224204
rect 559012 222896 559064 222902
rect 559012 222838 559064 222844
rect 559564 222896 559616 222902
rect 559564 222838 559616 222844
rect 558644 222760 558696 222766
rect 558644 222702 558696 222708
rect 557356 222352 557408 222358
rect 557356 222294 557408 222300
rect 556528 221604 556580 221610
rect 556528 221546 556580 221552
rect 556988 221604 557040 221610
rect 556988 221546 557040 221552
rect 556252 219972 556304 219978
rect 556252 219914 556304 219920
rect 555792 219836 555844 219842
rect 555792 219778 555844 219784
rect 555424 219768 555476 219774
rect 555424 219710 555476 219716
rect 554226 219127 554282 219136
rect 554872 219156 554924 219162
rect 554872 219098 554924 219104
rect 554056 217246 554130 217274
rect 551572 217110 551646 217138
rect 551618 216988 551646 217110
rect 552446 216988 552474 217246
rect 553274 216988 553302 217246
rect 554102 216988 554130 217246
rect 554884 217138 554912 219098
rect 555804 217274 555832 219778
rect 555758 217246 555832 217274
rect 554884 217110 554958 217138
rect 554930 216988 554958 217110
rect 555758 216988 555786 217246
rect 556540 217138 556568 221546
rect 556896 219156 556948 219162
rect 556896 219098 556948 219104
rect 556908 218754 556936 219098
rect 556896 218748 556948 218754
rect 556896 218690 556948 218696
rect 557368 217138 557396 222294
rect 558656 222194 558684 222702
rect 558564 222166 558684 222194
rect 558368 222148 558420 222154
rect 558368 222090 558420 222096
rect 558380 221270 558408 222090
rect 558184 221264 558236 221270
rect 558184 221206 558236 221212
rect 558368 221264 558420 221270
rect 558368 221206 558420 221212
rect 558196 220862 558224 221206
rect 558184 220856 558236 220862
rect 558184 220798 558236 220804
rect 558564 220674 558592 222166
rect 558012 220646 558592 220674
rect 558012 217274 558040 220646
rect 558828 220244 558880 220250
rect 558828 220186 558880 220192
rect 558840 219842 558868 220186
rect 559024 220130 559052 222838
rect 561324 222154 561352 224198
rect 560760 222148 560812 222154
rect 560760 222090 560812 222096
rect 561312 222148 561364 222154
rect 561312 222090 561364 222096
rect 559564 222012 559616 222018
rect 559564 221954 559616 221960
rect 559380 220244 559432 220250
rect 559380 220186 559432 220192
rect 559024 220102 559144 220130
rect 558460 219836 558512 219842
rect 558460 219778 558512 219784
rect 558828 219836 558880 219842
rect 558828 219778 558880 219784
rect 558472 219722 558500 219778
rect 558472 219694 558684 219722
rect 558368 219632 558420 219638
rect 558368 219574 558420 219580
rect 558380 219450 558408 219574
rect 558656 219570 558684 219694
rect 558828 219700 558880 219706
rect 558828 219642 558880 219648
rect 558644 219564 558696 219570
rect 558644 219506 558696 219512
rect 558840 219450 558868 219642
rect 558380 219422 558868 219450
rect 558184 218884 558236 218890
rect 558184 218826 558236 218832
rect 558196 218618 558224 218826
rect 558184 218612 558236 218618
rect 558184 218554 558236 218560
rect 559116 217274 559144 220102
rect 559392 219706 559420 220186
rect 559576 219978 559604 221954
rect 559840 221876 559892 221882
rect 559840 221818 559892 221824
rect 559564 219972 559616 219978
rect 559564 219914 559616 219920
rect 559380 219700 559432 219706
rect 559380 219642 559432 219648
rect 559852 218890 559880 221818
rect 559840 218884 559892 218890
rect 559840 218826 559892 218832
rect 558012 217246 558270 217274
rect 556540 217110 556614 217138
rect 557368 217110 557442 217138
rect 556586 216988 556614 217110
rect 557414 216988 557442 217110
rect 558242 216988 558270 217246
rect 559070 217246 559144 217274
rect 559070 216988 559098 217246
rect 559852 217138 559880 218826
rect 560772 217138 560800 222090
rect 561508 217274 561536 225694
rect 561680 223168 561732 223174
rect 561680 223110 561732 223116
rect 561692 222630 561720 223110
rect 561680 222624 561732 222630
rect 561680 222566 561732 222572
rect 562140 222624 562192 222630
rect 562140 222566 562192 222572
rect 562152 217274 562180 222566
rect 562336 222018 562364 252554
rect 562784 227044 562836 227050
rect 562784 226986 562836 226992
rect 562324 222012 562376 222018
rect 562324 221954 562376 221960
rect 562796 221882 562824 226986
rect 563716 224194 563744 259422
rect 565636 229764 565688 229770
rect 565636 229706 565688 229712
rect 563980 224392 564032 224398
rect 563980 224334 564032 224340
rect 563704 224188 563756 224194
rect 563704 224130 563756 224136
rect 563152 222624 563204 222630
rect 563152 222566 563204 222572
rect 563164 222222 563192 222566
rect 563334 222320 563390 222329
rect 563334 222255 563390 222264
rect 563152 222216 563204 222222
rect 563152 222158 563204 222164
rect 563014 222148 563066 222154
rect 563014 222090 563066 222096
rect 563026 222034 563054 222090
rect 563348 222034 563376 222255
rect 563992 222194 564020 224334
rect 565648 224330 565676 229706
rect 568592 229094 568620 260850
rect 571996 234598 572024 261462
rect 647252 246362 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 606484 245676 606536 245682
rect 606484 245618 606536 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 571984 234592 572036 234598
rect 571984 234534 572036 234540
rect 571340 230036 571392 230042
rect 571340 229978 571392 229984
rect 571352 229094 571380 229978
rect 568592 229066 569448 229094
rect 571352 229066 572300 229094
rect 566096 228540 566148 228546
rect 566096 228482 566148 228488
rect 565636 224324 565688 224330
rect 565636 224266 565688 224272
rect 565452 222624 565504 222630
rect 565452 222566 565504 222572
rect 563992 222166 564664 222194
rect 563026 222006 563376 222034
rect 562784 221876 562836 221882
rect 562784 221818 562836 221824
rect 562796 219434 562824 221818
rect 563060 220720 563112 220726
rect 563112 220680 563652 220708
rect 563060 220662 563112 220668
rect 563428 220516 563480 220522
rect 563428 220458 563480 220464
rect 563440 219774 563468 220458
rect 563624 220368 563652 220680
rect 563624 220340 564204 220368
rect 563428 219768 563480 219774
rect 563428 219710 563480 219716
rect 563796 219700 563848 219706
rect 563796 219642 563848 219648
rect 563520 219632 563572 219638
rect 563026 219558 563192 219586
rect 563808 219586 563836 219642
rect 563572 219580 563836 219586
rect 563520 219574 563836 219580
rect 563532 219558 563836 219574
rect 563026 219502 563054 219558
rect 563014 219496 563066 219502
rect 563014 219438 563066 219444
rect 562796 219406 562916 219434
rect 562888 217274 562916 219406
rect 563164 219280 563192 219558
rect 564176 219502 564204 220340
rect 564348 219768 564400 219774
rect 564348 219710 564400 219716
rect 563704 219496 563756 219502
rect 564164 219496 564216 219502
rect 563756 219456 564020 219484
rect 563704 219438 563756 219444
rect 563992 219416 564020 219456
rect 564164 219438 564216 219444
rect 563992 219388 564112 219416
rect 564084 219314 564112 219388
rect 564360 219314 564388 219710
rect 563428 219292 563480 219298
rect 563164 219252 563428 219280
rect 564084 219286 564388 219314
rect 563428 219234 563480 219240
rect 563026 219014 563468 219042
rect 563026 218890 563054 219014
rect 563014 218884 563066 218890
rect 563014 218826 563066 218832
rect 563152 218884 563204 218890
rect 563152 218826 563204 218832
rect 563164 218090 563192 218826
rect 563026 218074 563192 218090
rect 563014 218068 563192 218074
rect 563066 218062 563192 218068
rect 563014 218010 563066 218016
rect 563152 218000 563204 218006
rect 563072 217948 563152 217954
rect 563072 217942 563204 217948
rect 563072 217926 563192 217942
rect 563072 217569 563100 217926
rect 563440 217870 563468 219014
rect 563244 217864 563296 217870
rect 563244 217806 563296 217812
rect 563428 217864 563480 217870
rect 563428 217806 563480 217812
rect 563256 217569 563284 217806
rect 563058 217560 563114 217569
rect 563058 217495 563114 217504
rect 563242 217560 563298 217569
rect 563242 217495 563298 217504
rect 561508 217246 561582 217274
rect 562152 217246 562410 217274
rect 562888 217246 563238 217274
rect 559852 217110 559926 217138
rect 559898 216988 559926 217110
rect 560726 217110 560800 217138
rect 560726 216988 560754 217110
rect 561554 216988 561582 217246
rect 562382 216988 562410 217246
rect 563210 216988 563238 217246
rect 564636 217138 564664 222166
rect 564900 221604 564952 221610
rect 564900 221546 564952 221552
rect 564912 217138 564940 221546
rect 565464 220522 565492 222566
rect 565648 220522 565676 224266
rect 565452 220516 565504 220522
rect 565452 220458 565504 220464
rect 565636 220516 565688 220522
rect 565636 220458 565688 220464
rect 565464 219434 565492 220458
rect 566108 219434 566136 228482
rect 568120 227588 568172 227594
rect 568120 227530 568172 227536
rect 568132 224954 568160 227530
rect 569420 224954 569448 229066
rect 570788 225888 570840 225894
rect 570788 225830 570840 225836
rect 570800 224954 570828 225830
rect 572272 224954 572300 229066
rect 568132 224926 568436 224954
rect 569420 224926 569816 224954
rect 567844 224052 567896 224058
rect 567844 223994 567896 224000
rect 567856 223786 567884 223994
rect 567844 223780 567896 223786
rect 567844 223722 567896 223728
rect 567108 222624 567160 222630
rect 567108 222566 567160 222572
rect 567660 222624 567712 222630
rect 567660 222566 567712 222572
rect 567120 220674 567148 222566
rect 567672 221610 567700 222566
rect 567660 221604 567712 221610
rect 567660 221546 567712 221552
rect 567844 221604 567896 221610
rect 567844 221546 567896 221552
rect 567856 220862 567884 221546
rect 568408 220946 568436 224926
rect 568580 224324 568632 224330
rect 568580 224266 568632 224272
rect 568592 223786 568620 224266
rect 568948 224188 569000 224194
rect 568948 224130 569000 224136
rect 568580 223780 568632 223786
rect 568580 223722 568632 223728
rect 568764 222760 568816 222766
rect 568764 222702 568816 222708
rect 568408 220918 568528 220946
rect 567844 220856 567896 220862
rect 567844 220798 567896 220804
rect 568028 220788 568080 220794
rect 568028 220730 568080 220736
rect 568040 220674 568068 220730
rect 567120 220646 568068 220674
rect 566372 220516 566424 220522
rect 566372 220458 566424 220464
rect 566832 220516 566884 220522
rect 566832 220458 566884 220464
rect 566384 219586 566412 220458
rect 566556 220380 566608 220386
rect 566844 220368 566872 220458
rect 566608 220340 566872 220368
rect 566556 220322 566608 220328
rect 568304 220040 568356 220046
rect 568304 219982 568356 219988
rect 568316 219858 568344 219982
rect 568500 219858 568528 220918
rect 567672 219830 568344 219858
rect 568408 219830 568528 219858
rect 566384 219558 567332 219586
rect 565464 219406 565860 219434
rect 566108 219406 566228 219434
rect 565832 217274 565860 219406
rect 564038 217110 564664 217138
rect 564866 217110 564940 217138
rect 565694 217246 565860 217274
rect 564038 216988 564066 217110
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566200 217138 566228 219406
rect 566740 219020 566792 219026
rect 566740 218962 566792 218968
rect 566752 218906 566780 218962
rect 566752 218890 567148 218906
rect 566752 218884 567160 218890
rect 566752 218878 567108 218884
rect 567108 218826 567160 218832
rect 567304 217274 567332 219558
rect 567672 218385 567700 219830
rect 568408 219042 568436 219830
rect 568776 219774 568804 222702
rect 568580 219768 568632 219774
rect 568580 219710 568632 219716
rect 568764 219768 568816 219774
rect 568764 219710 568816 219716
rect 568592 219586 568620 219710
rect 568592 219558 568712 219586
rect 568408 219014 568528 219042
rect 567842 218920 567898 218929
rect 567842 218855 567898 218864
rect 568302 218920 568358 218929
rect 568302 218855 568358 218864
rect 567856 218385 567884 218855
rect 567658 218376 567714 218385
rect 567658 218311 567714 218320
rect 567842 218376 567898 218385
rect 567842 218311 567898 218320
rect 568316 218006 568344 218855
rect 568304 218000 568356 218006
rect 568304 217942 568356 217948
rect 567568 217864 567620 217870
rect 567620 217812 568160 217818
rect 567568 217806 568160 217812
rect 567580 217790 568160 217806
rect 568132 217734 568160 217790
rect 568120 217728 568172 217734
rect 568120 217670 568172 217676
rect 568500 217274 568528 219014
rect 568684 218006 568712 219558
rect 568672 218000 568724 218006
rect 568672 217942 568724 217948
rect 567304 217246 567378 217274
rect 566200 217110 566550 217138
rect 566522 216988 566550 217110
rect 567350 216988 567378 217246
rect 568178 217246 568528 217274
rect 568178 216988 568206 217246
rect 568960 217138 568988 224130
rect 569788 217274 569816 224926
rect 570708 224926 570828 224954
rect 571812 224926 572300 224954
rect 570708 217274 570736 224926
rect 571616 222624 571668 222630
rect 571616 222566 571668 222572
rect 571628 222018 571656 222566
rect 571812 222442 571840 224926
rect 571720 222414 571840 222442
rect 571720 222170 571748 222414
rect 571890 222320 571946 222329
rect 571890 222255 571946 222264
rect 571720 222142 571840 222170
rect 571432 222012 571484 222018
rect 571432 221954 571484 221960
rect 571616 222012 571668 222018
rect 571616 221954 571668 221960
rect 569788 217246 569862 217274
rect 568960 217110 569034 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217246
rect 570662 217246 570736 217274
rect 570662 216988 570690 217246
rect 571444 217138 571472 221954
rect 571812 217274 571840 222142
rect 571904 218090 571932 222255
rect 577320 220788 577372 220794
rect 577320 220730 577372 220736
rect 572076 220652 572128 220658
rect 572076 220594 572128 220600
rect 572088 218226 572116 220594
rect 577332 220114 577360 220730
rect 577320 220108 577372 220114
rect 577320 220050 577372 220056
rect 574468 220040 574520 220046
rect 574468 219982 574520 219988
rect 572272 219388 572668 219416
rect 572272 219026 572300 219388
rect 572640 219298 572668 219388
rect 572444 219292 572496 219298
rect 572444 219234 572496 219240
rect 572628 219292 572680 219298
rect 572628 219234 572680 219240
rect 572456 219178 572484 219234
rect 572456 219150 572760 219178
rect 572260 219020 572312 219026
rect 572260 218962 572312 218968
rect 572444 219020 572496 219026
rect 572444 218962 572496 218968
rect 572456 218385 572484 218962
rect 572732 218929 572760 219150
rect 572718 218920 572774 218929
rect 572718 218855 572774 218864
rect 572442 218376 572498 218385
rect 572442 218311 572498 218320
rect 572626 218376 572682 218385
rect 572626 218311 572682 218320
rect 572640 218226 572668 218311
rect 572088 218198 572668 218226
rect 572994 218104 573050 218113
rect 571904 218062 572346 218090
rect 572318 218006 572346 218062
rect 572456 218062 572760 218090
rect 572168 218000 572220 218006
rect 572168 217942 572220 217948
rect 572306 218000 572358 218006
rect 572306 217942 572358 217948
rect 572180 217852 572208 217942
rect 572456 217852 572484 218062
rect 572732 217954 572760 218062
rect 573050 218074 573220 218090
rect 573050 218068 573232 218074
rect 573050 218062 573180 218068
rect 572994 218039 573050 218048
rect 573180 218010 573232 218016
rect 572732 217926 574232 217954
rect 572180 217824 572484 217852
rect 572720 217864 572772 217870
rect 572772 217812 573128 217818
rect 572720 217806 573128 217812
rect 572732 217790 573128 217806
rect 573100 217734 573128 217790
rect 572076 217728 572128 217734
rect 572076 217670 572128 217676
rect 572260 217728 572312 217734
rect 572260 217670 572312 217676
rect 572720 217728 572772 217734
rect 573088 217728 573140 217734
rect 572772 217676 572944 217682
rect 572720 217670 572944 217676
rect 573088 217670 573140 217676
rect 572088 217410 572116 217670
rect 572272 217569 572300 217670
rect 572732 217654 572944 217670
rect 572916 217569 572944 217654
rect 572258 217560 572314 217569
rect 572258 217495 572314 217504
rect 572902 217560 572958 217569
rect 572902 217495 572958 217504
rect 572088 217382 572484 217410
rect 572456 217274 572484 217382
rect 571812 217246 572346 217274
rect 572456 217246 574140 217274
rect 571444 217110 571518 217138
rect 571490 216988 571518 217110
rect 572318 216988 572346 217246
rect 574112 214606 574140 217246
rect 574204 215294 574232 217926
rect 574204 215266 574324 215294
rect 574100 214600 574152 214606
rect 574100 214542 574152 214548
rect 574296 213246 574324 215266
rect 574480 214878 574508 219982
rect 575664 219292 575716 219298
rect 575664 219234 575716 219240
rect 575480 217048 575532 217054
rect 575480 216990 575532 216996
rect 574468 214872 574520 214878
rect 574468 214814 574520 214820
rect 575492 213382 575520 216990
rect 575676 214742 575704 219234
rect 575848 219020 575900 219026
rect 575848 218962 575900 218968
rect 575860 215014 575888 218962
rect 577320 217728 577372 217734
rect 577320 217670 577372 217676
rect 577332 217054 577360 217670
rect 577320 217048 577372 217054
rect 577320 216990 577372 216996
rect 577044 215892 577096 215898
rect 577044 215834 577096 215840
rect 577056 215121 577084 215834
rect 577042 215112 577098 215121
rect 577042 215047 577098 215056
rect 575848 215008 575900 215014
rect 575848 214950 575900 214956
rect 575664 214736 575716 214742
rect 575664 214678 575716 214684
rect 575480 213376 575532 213382
rect 575480 213318 575532 213324
rect 574284 213240 574336 213246
rect 574284 213182 574336 213188
rect 577516 99142 577544 240110
rect 606300 224188 606352 224194
rect 606300 224130 606352 224136
rect 606312 223922 606340 224130
rect 606300 223916 606352 223922
rect 606300 223858 606352 223864
rect 593972 222488 594024 222494
rect 593972 222430 594024 222436
rect 577688 222012 577740 222018
rect 577688 221954 577740 221960
rect 577700 220862 577728 221954
rect 577688 220856 577740 220862
rect 577688 220798 577740 220804
rect 591396 219224 591448 219230
rect 591394 219192 591396 219201
rect 591448 219192 591450 219201
rect 587348 219156 587400 219162
rect 591394 219127 591450 219136
rect 587348 219098 587400 219104
rect 587164 218884 587216 218890
rect 587164 218826 587216 218832
rect 587176 218618 587204 218826
rect 587360 218618 587388 219098
rect 587164 218612 587216 218618
rect 587164 218554 587216 218560
rect 587348 218612 587400 218618
rect 587348 218554 587400 218560
rect 582102 218104 582158 218113
rect 582102 218039 582158 218048
rect 582286 218104 582342 218113
rect 582286 218039 582288 218048
rect 582116 217818 582144 218039
rect 582340 218039 582342 218048
rect 582288 218010 582340 218016
rect 591854 217832 591910 217841
rect 582116 217790 582328 217818
rect 582104 217728 582156 217734
rect 582104 217670 582156 217676
rect 582116 217569 582144 217670
rect 582300 217569 582328 217790
rect 591910 217790 592080 217818
rect 591854 217767 591910 217776
rect 592052 217734 592080 217790
rect 586888 217728 586940 217734
rect 586888 217670 586940 217676
rect 592040 217728 592092 217734
rect 592040 217670 592092 217676
rect 582102 217560 582158 217569
rect 582102 217495 582158 217504
rect 582286 217560 582342 217569
rect 582286 217495 582342 217504
rect 582378 217288 582434 217297
rect 582378 217223 582434 217232
rect 582392 216918 582420 217223
rect 586900 217025 586928 217670
rect 582930 217016 582986 217025
rect 582930 216951 582986 216960
rect 586886 217016 586942 217025
rect 592222 217016 592278 217025
rect 586886 216951 586942 216960
rect 592052 216974 592222 217002
rect 582380 216912 582432 216918
rect 582380 216854 582432 216860
rect 582944 216050 582972 216951
rect 592052 216918 592080 216974
rect 592222 216951 592278 216960
rect 592040 216912 592092 216918
rect 592040 216854 592092 216860
rect 582392 216022 582972 216050
rect 582392 215937 582420 216022
rect 582378 215928 582434 215937
rect 582378 215863 582434 215872
rect 582562 215928 582618 215937
rect 582562 215863 582564 215872
rect 582616 215863 582618 215872
rect 582564 215834 582616 215840
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578238 211712 578294 211721
rect 578238 211647 578294 211656
rect 578252 211342 578280 211647
rect 578240 211336 578292 211342
rect 578240 211278 578292 211284
rect 578896 208350 578924 213959
rect 580448 211336 580500 211342
rect 580448 211278 580500 211284
rect 579252 209840 579304 209846
rect 579250 209808 579252 209817
rect 579304 209808 579306 209817
rect 579250 209743 579306 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 580460 207670 580488 211278
rect 593984 210202 594012 222430
rect 599490 222048 599546 222057
rect 596272 222012 596324 222018
rect 596272 221954 596324 221960
rect 597008 222012 597060 222018
rect 599490 221983 599546 221992
rect 597008 221954 597060 221960
rect 596284 221610 596312 221954
rect 596272 221604 596324 221610
rect 596272 221546 596324 221552
rect 596456 221604 596508 221610
rect 596456 221546 596508 221552
rect 596468 221270 596496 221546
rect 596456 221264 596508 221270
rect 596456 221206 596508 221212
rect 596640 221264 596692 221270
rect 596640 221206 596692 221212
rect 596652 220998 596680 221206
rect 597020 221134 597048 221954
rect 597008 221128 597060 221134
rect 597008 221070 597060 221076
rect 596640 220992 596692 220998
rect 596640 220934 596692 220940
rect 594154 219464 594210 219473
rect 594154 219399 594210 219408
rect 594168 219230 594196 219399
rect 594156 219224 594208 219230
rect 594156 219166 594208 219172
rect 595166 219192 595222 219201
rect 595166 219127 595222 219136
rect 594984 217728 595036 217734
rect 594984 217670 595036 217676
rect 594996 216753 595024 217670
rect 594798 216744 594854 216753
rect 594798 216679 594854 216688
rect 594982 216744 595038 216753
rect 594982 216679 595038 216688
rect 594614 215656 594670 215665
rect 594614 215591 594616 215600
rect 594668 215591 594670 215600
rect 594616 215562 594668 215568
rect 594812 210202 594840 216679
rect 595180 210202 595208 219127
rect 597744 219020 597796 219026
rect 597744 218962 597796 218968
rect 596824 218884 596876 218890
rect 596824 218826 596876 218832
rect 596640 217456 596692 217462
rect 596640 217398 596692 217404
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596652 216918 596680 217398
rect 596640 216912 596692 216918
rect 596640 216854 596692 216860
rect 596362 216200 596418 216209
rect 596362 216135 596418 216144
rect 596180 215348 596232 215354
rect 596180 215294 596232 215296
rect 596100 215290 596232 215294
rect 596100 215266 596220 215290
rect 596100 215121 596128 215266
rect 596086 215112 596142 215121
rect 596086 215047 596142 215056
rect 596376 210202 596404 216135
rect 596836 215966 596864 218826
rect 597558 217832 597614 217841
rect 597558 217767 597614 217776
rect 596824 215960 596876 215966
rect 596824 215902 596876 215908
rect 596824 215348 596876 215354
rect 596824 215290 596876 215296
rect 596836 210202 596864 215290
rect 597572 210202 597600 217767
rect 597756 216102 597784 218962
rect 599030 216744 599086 216753
rect 599030 216679 599086 216688
rect 597744 216096 597796 216102
rect 597744 216038 597796 216044
rect 597926 215656 597982 215665
rect 597926 215591 597982 215600
rect 598480 215620 598532 215626
rect 597940 210202 597968 215591
rect 598480 215562 598532 215568
rect 598492 210202 598520 215562
rect 599044 210202 599072 216679
rect 599504 210202 599532 221983
rect 603354 221776 603410 221785
rect 603354 221711 603410 221720
rect 600318 221504 600374 221513
rect 600318 221439 600374 221448
rect 600332 212430 600360 221439
rect 600778 221232 600834 221241
rect 600778 221167 600834 221176
rect 600594 220960 600650 220969
rect 600594 220895 600650 220904
rect 600608 212534 600636 220895
rect 600792 215294 600820 221167
rect 602066 218648 602122 218657
rect 602066 218583 602122 218592
rect 602080 217598 602108 218583
rect 602068 217592 602120 217598
rect 602068 217534 602120 217540
rect 602344 217456 602396 217462
rect 602344 217398 602396 217404
rect 600516 212506 600636 212534
rect 600700 215266 600820 215294
rect 600320 212424 600372 212430
rect 600320 212366 600372 212372
rect 600516 211070 600544 212506
rect 600504 211064 600556 211070
rect 600504 211006 600556 211012
rect 600700 210882 600728 215266
rect 601792 213376 601844 213382
rect 601792 213318 601844 213324
rect 601240 212424 601292 212430
rect 601240 212366 601292 212372
rect 600872 211064 600924 211070
rect 600872 211006 600924 211012
rect 600516 210854 600728 210882
rect 600516 210202 600544 210854
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600544 210202
rect 600884 210202 600912 211006
rect 601252 210202 601280 212366
rect 601804 210202 601832 213318
rect 602356 210202 602384 217398
rect 603080 217320 603132 217326
rect 603080 217262 603132 217268
rect 603092 210202 603120 217262
rect 603368 210202 603396 221711
rect 606496 221474 606524 245618
rect 648632 242214 648660 277366
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 628564 241528 628616 241534
rect 628564 241470 628616 241476
rect 616880 224052 616932 224058
rect 616880 223994 616932 224000
rect 610532 221876 610584 221882
rect 610532 221818 610584 221824
rect 608600 221740 608652 221746
rect 608600 221682 608652 221688
rect 607312 221604 607364 221610
rect 607312 221546 607364 221552
rect 605472 221468 605524 221474
rect 605472 221410 605524 221416
rect 606484 221468 606536 221474
rect 606484 221410 606536 221416
rect 605288 220652 605340 220658
rect 605288 220594 605340 220600
rect 605300 219638 605328 220594
rect 605288 219632 605340 219638
rect 605288 219574 605340 219580
rect 604368 218476 604420 218482
rect 604368 218418 604420 218424
rect 604380 217462 604408 218418
rect 604368 217456 604420 217462
rect 604368 217398 604420 217404
rect 604552 217184 604604 217190
rect 604552 217126 604604 217132
rect 604000 216912 604052 216918
rect 604000 216854 604052 216860
rect 604012 210202 604040 216854
rect 604564 210202 604592 217126
rect 605104 217048 605156 217054
rect 605104 216990 605156 216996
rect 605116 210202 605144 216990
rect 605484 212534 605512 221410
rect 606944 221128 606996 221134
rect 606944 221070 606996 221076
rect 606208 220992 606260 220998
rect 606128 220940 606208 220946
rect 606128 220934 606260 220940
rect 606128 220918 606248 220934
rect 605656 219768 605708 219774
rect 605656 219710 605708 219716
rect 605668 219366 605696 219710
rect 606128 219450 606156 220918
rect 606484 220516 606536 220522
rect 606484 220458 606536 220464
rect 606300 220380 606352 220386
rect 606300 220322 606352 220328
rect 606312 219638 606340 220322
rect 606496 219774 606524 220458
rect 606484 219768 606536 219774
rect 606484 219710 606536 219716
rect 606300 219632 606352 219638
rect 606300 219574 606352 219580
rect 606128 219422 606340 219450
rect 605656 219360 605708 219366
rect 605656 219302 605708 219308
rect 605748 218204 605800 218210
rect 605748 218146 605800 218152
rect 605760 217734 605788 218146
rect 605748 217728 605800 217734
rect 605748 217670 605800 217676
rect 606312 215294 606340 219422
rect 606758 217560 606814 217569
rect 606758 217495 606814 217504
rect 606772 217025 606800 217495
rect 606758 217016 606814 217025
rect 606758 216951 606814 216960
rect 606220 215266 606340 215294
rect 605484 212506 605880 212534
rect 605852 210202 605880 212506
rect 606220 210202 606248 215266
rect 606956 212534 606984 221070
rect 607324 214606 607352 221546
rect 607496 221264 607548 221270
rect 607496 221206 607548 221212
rect 607312 214600 607364 214606
rect 607312 214542 607364 214548
rect 606772 212506 606984 212534
rect 606772 210202 606800 212506
rect 607508 210202 607536 221206
rect 607864 214600 607916 214606
rect 607864 214542 607916 214548
rect 607876 210202 607904 214542
rect 608612 210202 608640 221682
rect 608968 220652 609020 220658
rect 608968 220594 609020 220600
rect 608784 219360 608836 219366
rect 608784 219302 608836 219308
rect 608796 214606 608824 219302
rect 608784 214600 608836 214606
rect 608784 214542 608836 214548
rect 608980 210202 609008 220594
rect 610072 217864 610124 217870
rect 610072 217806 610124 217812
rect 609520 214600 609572 214606
rect 609520 214542 609572 214548
rect 609532 210202 609560 214542
rect 610084 210202 610112 217806
rect 610544 210202 610572 221818
rect 611360 220108 611412 220114
rect 611360 220050 611412 220056
rect 611372 210202 611400 220050
rect 611544 218612 611596 218618
rect 611544 218554 611596 218560
rect 611556 215354 611584 218554
rect 612738 218376 612794 218385
rect 612738 218311 612794 218320
rect 616144 218340 616196 218346
rect 612752 217326 612780 218311
rect 616144 218282 616196 218288
rect 615040 217728 615092 217734
rect 615040 217670 615092 217676
rect 613384 217592 613436 217598
rect 613384 217534 613436 217540
rect 612740 217320 612792 217326
rect 612740 217262 612792 217268
rect 611726 215928 611782 215937
rect 611726 215863 611782 215872
rect 611544 215348 611596 215354
rect 611544 215290 611596 215296
rect 611740 210202 611768 215863
rect 612280 215008 612332 215014
rect 612280 214950 612332 214956
rect 612292 210202 612320 214950
rect 612832 214872 612884 214878
rect 612832 214814 612884 214820
rect 612844 210202 612872 214814
rect 613396 210202 613424 217534
rect 614120 217456 614172 217462
rect 614120 217398 614172 217404
rect 614132 210202 614160 217398
rect 614488 215348 614540 215354
rect 614488 215290 614540 215296
rect 614500 210202 614528 215290
rect 615052 210202 615080 217670
rect 615592 213240 615644 213246
rect 615592 213182 615644 213188
rect 615604 210202 615632 213182
rect 616156 210202 616184 218282
rect 616892 210202 616920 223994
rect 627920 223780 627972 223786
rect 627920 223722 627972 223728
rect 626540 222352 626592 222358
rect 626540 222294 626592 222300
rect 618810 220552 618866 220561
rect 618810 220487 618866 220496
rect 618168 218748 618220 218754
rect 618168 218690 618220 218696
rect 617798 217560 617854 217569
rect 617798 217495 617854 217504
rect 617246 217288 617302 217297
rect 617246 217223 617302 217232
rect 617260 210202 617288 217223
rect 617812 210202 617840 217495
rect 618180 216714 618208 218690
rect 618168 216708 618220 216714
rect 618168 216650 618220 216656
rect 618350 216472 618406 216481
rect 618350 216407 618406 216416
rect 618364 210202 618392 216407
rect 618824 210202 618852 220487
rect 619638 220280 619694 220289
rect 619638 220215 619694 220224
rect 619652 219434 619680 220215
rect 621112 220108 621164 220114
rect 621112 220050 621164 220056
rect 620466 220008 620522 220017
rect 620466 219943 620522 219952
rect 619822 219736 619878 219745
rect 619822 219671 619878 219680
rect 619652 219406 619772 219434
rect 619744 212534 619772 219406
rect 619652 212506 619772 212534
rect 619652 211070 619680 212506
rect 619640 211064 619692 211070
rect 619640 211006 619692 211012
rect 619836 210746 619864 219671
rect 620008 211064 620060 211070
rect 620008 211006 620060 211012
rect 619836 210718 619956 210746
rect 619928 210202 619956 210718
rect 600884 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602356 210174 602692 210202
rect 603092 210174 603244 210202
rect 603368 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605116 210174 605452 210202
rect 605852 210174 606004 210202
rect 606220 210174 606556 210202
rect 606772 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210174 608764 210202
rect 608980 210174 609316 210202
rect 609532 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611372 210174 611524 210202
rect 611740 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615604 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618364 210174 618700 210202
rect 618824 210174 619252 210202
rect 619804 210174 619956 210202
rect 620020 210202 620048 211006
rect 620480 210202 620508 219943
rect 621124 214606 621152 220050
rect 622492 219904 622544 219910
rect 622492 219846 622544 219852
rect 621294 219464 621350 219473
rect 621294 219399 621350 219408
rect 621112 214600 621164 214606
rect 621112 214542 621164 214548
rect 621308 210202 621336 219399
rect 622308 214736 622360 214742
rect 622308 214678 622360 214684
rect 621664 214600 621716 214606
rect 621664 214542 621716 214548
rect 621676 210202 621704 214542
rect 622320 214418 622348 214678
rect 622504 214606 622532 219846
rect 624332 219768 624384 219774
rect 624332 219710 624384 219716
rect 622676 219632 622728 219638
rect 622676 219574 622728 219580
rect 622492 214600 622544 214606
rect 622492 214542 622544 214548
rect 622320 214390 622532 214418
rect 622504 210202 622532 214390
rect 622688 210202 622716 219574
rect 623872 216708 623924 216714
rect 623872 216650 623924 216656
rect 623320 214600 623372 214606
rect 623320 214542 623372 214548
rect 623332 210202 623360 214542
rect 623884 210202 623912 216650
rect 624344 210202 624372 219710
rect 625160 219496 625212 219502
rect 625160 219438 625212 219444
rect 625172 216050 625200 219438
rect 626080 216096 626132 216102
rect 625172 216022 625476 216050
rect 626080 216038 626132 216044
rect 625252 215960 625304 215966
rect 625252 215902 625304 215908
rect 625264 210202 625292 215902
rect 625448 210202 625476 216022
rect 626092 210202 626120 216038
rect 626552 210202 626580 222294
rect 627734 218104 627790 218113
rect 627734 218039 627790 218048
rect 627184 214464 627236 214470
rect 627184 214406 627236 214412
rect 627196 210202 627224 214406
rect 627748 213994 627776 218039
rect 627932 214606 627960 223722
rect 628196 222216 628248 222222
rect 628196 222158 628248 222164
rect 627920 214600 627972 214606
rect 627920 214542 627972 214548
rect 627736 213988 627788 213994
rect 627736 213930 627788 213936
rect 628208 210202 628236 222158
rect 628380 220856 628432 220862
rect 628380 220798 628432 220804
rect 620020 210174 620356 210202
rect 620480 210174 620908 210202
rect 621308 210174 621460 210202
rect 621676 210174 622012 210202
rect 622504 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624344 210174 624772 210202
rect 625264 210174 625324 210202
rect 625448 210174 625876 210202
rect 626092 210174 626428 210202
rect 626552 210174 626980 210202
rect 627196 210174 627532 210202
rect 628084 210174 628236 210202
rect 628392 210202 628420 220798
rect 628576 214742 628604 241470
rect 639602 229800 639658 229809
rect 639602 229735 639658 229744
rect 632704 228404 632756 228410
rect 632704 228346 632756 228352
rect 630956 223916 631008 223922
rect 630956 223858 631008 223864
rect 629852 223644 629904 223650
rect 629852 223586 629904 223592
rect 629392 217320 629444 217326
rect 629392 217262 629444 217268
rect 628564 214736 628616 214742
rect 628564 214678 628616 214684
rect 628840 214600 628892 214606
rect 628840 214542 628892 214548
rect 628852 210202 628880 214542
rect 629404 210202 629432 217262
rect 629864 210202 629892 223586
rect 630678 218648 630734 218657
rect 630678 218583 630734 218592
rect 630692 210202 630720 218583
rect 630968 210202 630996 223858
rect 631600 213988 631652 213994
rect 631600 213930 631652 213936
rect 631612 210202 631640 213930
rect 632716 212770 632744 228346
rect 633716 222896 633768 222902
rect 633716 222838 633768 222844
rect 633440 221468 633492 221474
rect 633440 221410 633492 221416
rect 632888 214736 632940 214742
rect 632888 214678 632940 214684
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 632900 210202 632928 214678
rect 633452 210202 633480 221410
rect 633728 210202 633756 222838
rect 637578 220144 637634 220153
rect 636476 220108 636528 220114
rect 637578 220079 637634 220088
rect 636476 220050 636528 220056
rect 636292 214600 636344 214606
rect 636292 214542 636344 214548
rect 635556 213512 635608 213518
rect 635556 213454 635608 213460
rect 634360 212764 634412 212770
rect 634360 212706 634412 212712
rect 634372 210202 634400 212706
rect 635568 210202 635596 213454
rect 628392 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631612 210174 631948 210202
rect 632900 210174 633052 210202
rect 633452 210174 633604 210202
rect 633728 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636304 210202 636332 214542
rect 636488 210202 636516 220050
rect 637592 213926 637620 220079
rect 639616 214606 639644 229735
rect 650642 225584 650698 225593
rect 650642 225519 650698 225528
rect 646134 220416 646190 220425
rect 646134 220351 646190 220360
rect 641166 218920 641222 218929
rect 641166 218855 641222 218864
rect 639970 217560 640026 217569
rect 639970 217495 640026 217504
rect 639604 214600 639656 214606
rect 639604 214542 639656 214548
rect 637580 213920 637632 213926
rect 637580 213862 637632 213868
rect 638224 213920 638276 213926
rect 638224 213862 638276 213868
rect 638040 213784 638092 213790
rect 638040 213726 638092 213732
rect 638052 210202 638080 213726
rect 636304 210174 636364 210202
rect 636488 210174 636916 210202
rect 638020 210174 638080 210202
rect 638236 210202 638264 213862
rect 639984 210202 640012 217495
rect 641180 213790 641208 218855
rect 643834 218376 643890 218385
rect 643834 218311 643890 218320
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 641168 213784 641220 213790
rect 641168 213726 641220 213732
rect 641628 213648 641680 213654
rect 641628 213590 641680 213596
rect 640248 213376 640300 213382
rect 640248 213318 640300 213324
rect 640260 210202 640288 213318
rect 641640 210202 641668 213590
rect 642180 213240 642232 213246
rect 642180 213182 642232 213188
rect 642192 210202 642220 213182
rect 643020 210202 643048 215863
rect 643848 210202 643876 218311
rect 644938 217832 644994 217841
rect 644938 217767 644994 217776
rect 644952 210202 644980 217767
rect 646148 213926 646176 220351
rect 648618 219872 648674 219881
rect 648618 219807 648674 219816
rect 648252 218204 648304 218210
rect 648252 218146 648304 218152
rect 646594 216200 646650 216209
rect 646594 216135 646650 216144
rect 645492 213920 645544 213926
rect 645492 213862 645544 213868
rect 646136 213920 646188 213926
rect 646136 213862 646188 213868
rect 645504 210202 645532 213862
rect 646608 210202 646636 216135
rect 647146 213208 647202 213217
rect 647146 213143 647202 213152
rect 647160 210202 647188 213143
rect 648264 210202 648292 218146
rect 648436 214600 648488 214606
rect 648436 214542 648488 214548
rect 638236 210174 638572 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647956 210174 648292 210202
rect 648448 210202 648476 214542
rect 648632 213926 648660 219807
rect 650458 214568 650514 214577
rect 650458 214503 650514 214512
rect 648620 213920 648672 213926
rect 648620 213862 648672 213868
rect 649264 213920 649316 213926
rect 649264 213862 649316 213868
rect 649276 210202 649304 213862
rect 650472 210202 650500 214503
rect 650656 213654 650684 225519
rect 651286 219192 651342 219201
rect 651286 219127 651342 219136
rect 650644 213648 650696 213654
rect 650644 213590 650696 213596
rect 651300 210202 651328 219127
rect 651840 213648 651892 213654
rect 651840 213590 651892 213596
rect 651852 210202 651880 213590
rect 648448 210174 648508 210202
rect 649276 210174 649612 210202
rect 650164 210174 650500 210202
rect 651268 210174 651328 210202
rect 651820 210174 651880 210202
rect 581736 209840 581788 209846
rect 581736 209782 581788 209788
rect 581552 208616 581604 208622
rect 581552 208558 581604 208564
rect 580448 207664 580500 207670
rect 580448 207606 580500 207612
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 581564 200114 581592 208558
rect 581748 206310 581776 209782
rect 652036 209574 652064 338263
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652220 209574 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 411913 660344 550598
rect 661696 491609 661724 603094
rect 663076 538801 663104 656882
rect 664456 580145 664484 709310
rect 665836 626113 665864 749362
rect 666296 711657 666324 778359
rect 666466 742520 666522 742529
rect 666466 742455 666522 742464
rect 666282 711648 666338 711657
rect 666282 711583 666338 711592
rect 666480 665417 666508 742455
rect 667216 671129 667244 803150
rect 668214 789440 668270 789449
rect 668214 789375 668270 789384
rect 668584 789404 668636 789410
rect 667846 743200 667902 743209
rect 667846 743135 667902 743144
rect 667662 688936 667718 688945
rect 667662 688871 667718 688880
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 666466 665408 666522 665417
rect 666466 665343 666522 665352
rect 667204 628584 667256 628590
rect 667204 628526 667256 628532
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 665824 590708 665876 590714
rect 665824 590650 665876 590656
rect 664442 580136 664498 580145
rect 664442 580071 664498 580080
rect 664444 576904 664496 576910
rect 664444 576846 664496 576852
rect 663062 538792 663118 538801
rect 663062 538727 663118 538736
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661682 491600 661738 491609
rect 661682 491535 661738 491544
rect 661684 456816 661736 456822
rect 661684 456758 661736 456764
rect 660302 411904 660358 411913
rect 660302 411839 660358 411848
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 661696 313585 661724 456758
rect 661880 406337 661908 522990
rect 663248 494760 663300 494766
rect 664456 494737 664484 576846
rect 663248 494702 663300 494708
rect 664442 494728 664498 494737
rect 663064 416832 663116 416838
rect 663064 416774 663116 416780
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 661868 364404 661920 364410
rect 661868 364346 661920 364352
rect 661682 313576 661738 313585
rect 661682 313511 661738 313520
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 661880 232626 661908 364346
rect 663076 268161 663104 416774
rect 663260 358601 663288 494702
rect 664442 494663 664498 494672
rect 665836 492153 665864 590650
rect 667216 534177 667244 628526
rect 667676 621217 667704 688871
rect 667860 665961 667888 743135
rect 668228 709617 668256 789375
rect 668584 789346 668636 789352
rect 668400 775600 668452 775606
rect 668400 775542 668452 775548
rect 668412 735321 668440 775542
rect 668398 735312 668454 735321
rect 668398 735247 668454 735256
rect 668214 709608 668270 709617
rect 668214 709543 668270 709552
rect 668398 692880 668454 692889
rect 668398 692815 668454 692824
rect 668214 685536 668270 685545
rect 668214 685471 668270 685480
rect 667846 665952 667902 665961
rect 667846 665887 667902 665896
rect 667846 643240 667902 643249
rect 667846 643175 667902 643184
rect 667662 621208 667718 621217
rect 667662 621143 667718 621152
rect 667860 576065 667888 643175
rect 668228 615641 668256 685471
rect 668412 619993 668440 692815
rect 668596 670585 668624 789346
rect 668872 755313 668900 872199
rect 669042 866688 669098 866697
rect 669042 866623 669098 866632
rect 668858 755304 668914 755313
rect 668858 755239 668914 755248
rect 669056 750825 669084 866623
rect 669240 753545 669268 876279
rect 669778 873488 669834 873497
rect 669778 873423 669834 873432
rect 669594 783864 669650 783873
rect 669594 783799 669650 783808
rect 669226 753536 669282 753545
rect 669226 753471 669282 753480
rect 669042 750816 669098 750825
rect 669042 750751 669098 750760
rect 669226 741160 669282 741169
rect 669226 741095 669282 741104
rect 668766 738984 668822 738993
rect 668766 738919 668822 738928
rect 668582 670576 668638 670585
rect 668582 670511 668638 670520
rect 668780 666233 668808 738919
rect 669042 733680 669098 733689
rect 669042 733615 669098 733624
rect 668766 666224 668822 666233
rect 668766 666159 668822 666168
rect 669056 662561 669084 733615
rect 669240 663921 669268 741095
rect 669608 708801 669636 783799
rect 669792 756129 669820 873423
rect 669964 841832 670016 841838
rect 669964 841774 670016 841780
rect 669778 756120 669834 756129
rect 669778 756055 669834 756064
rect 669778 731504 669834 731513
rect 669778 731439 669834 731448
rect 669594 708792 669650 708801
rect 669594 708727 669650 708736
rect 669594 701176 669650 701185
rect 669594 701111 669650 701120
rect 669226 663912 669282 663921
rect 669226 663847 669282 663856
rect 669042 662552 669098 662561
rect 669042 662487 669098 662496
rect 669226 654256 669282 654265
rect 669226 654191 669282 654200
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668398 619984 668454 619993
rect 668398 619919 668454 619928
rect 668214 615632 668270 615641
rect 668214 615567 668270 615576
rect 668398 593600 668454 593609
rect 668398 593535 668454 593544
rect 667846 576056 667902 576065
rect 667846 575991 667902 576000
rect 667846 564496 667902 564505
rect 667846 564431 667902 564440
rect 667662 554704 667718 554713
rect 667662 554639 667718 554648
rect 667202 534168 667258 534177
rect 667202 534103 667258 534112
rect 665822 492144 665878 492153
rect 665822 492079 665878 492088
rect 667204 484424 667256 484430
rect 667204 484366 667256 484372
rect 665824 470620 665876 470626
rect 665824 470562 665876 470568
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663246 358592 663302 358601
rect 663246 358527 663302 358536
rect 664456 271153 664484 404330
rect 665836 315489 665864 470562
rect 667216 360913 667244 484366
rect 667676 482769 667704 554639
rect 667860 485217 667888 564431
rect 668412 528601 668440 593535
rect 668596 535945 668624 643078
rect 668766 604344 668822 604353
rect 668766 604279 668822 604288
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668780 528873 668808 604279
rect 669042 599312 669098 599321
rect 669042 599247 669098 599256
rect 668766 528864 668822 528873
rect 668766 528799 668822 528808
rect 668398 528592 668454 528601
rect 668398 528527 668454 528536
rect 669056 527377 669084 599247
rect 669240 574161 669268 654191
rect 669608 621625 669636 701111
rect 669792 664193 669820 731439
rect 669976 715737 670004 841774
rect 670330 782504 670386 782513
rect 670330 782439 670386 782448
rect 670146 775704 670202 775713
rect 670146 775639 670202 775648
rect 669962 715728 670018 715737
rect 669962 715663 670018 715672
rect 670160 710025 670188 775639
rect 670146 710016 670202 710025
rect 670146 709951 670202 709960
rect 670344 707169 670372 782439
rect 670620 754633 670648 876823
rect 670790 778424 670846 778433
rect 670790 778359 670846 778368
rect 670804 776529 670832 778359
rect 670790 776520 670846 776529
rect 670790 776455 670846 776464
rect 670988 763065 671016 895630
rect 671158 869136 671214 869145
rect 671158 869071 671214 869080
rect 670974 763056 671030 763065
rect 670974 762991 671030 763000
rect 670974 758296 671030 758305
rect 670974 758231 671030 758240
rect 670606 754624 670662 754633
rect 670606 754559 670662 754568
rect 670790 750136 670846 750145
rect 670790 750071 670846 750080
rect 670606 730552 670662 730561
rect 670606 730487 670662 730496
rect 670330 707160 670386 707169
rect 670330 707095 670386 707104
rect 669964 696992 670016 696998
rect 669964 696934 670016 696940
rect 670422 696960 670478 696969
rect 669778 664184 669834 664193
rect 669778 664119 669834 664128
rect 669778 638616 669834 638625
rect 669778 638551 669834 638560
rect 669594 621616 669650 621625
rect 669594 621551 669650 621560
rect 669594 614952 669650 614961
rect 669594 614887 669650 614896
rect 669226 574152 669282 574161
rect 669226 574087 669282 574096
rect 669226 557560 669282 557569
rect 669226 557495 669282 557504
rect 669042 527368 669098 527377
rect 669042 527303 669098 527312
rect 669240 486033 669268 557495
rect 669226 486024 669282 486033
rect 669226 485959 669282 485968
rect 667846 485208 667902 485217
rect 667846 485143 667902 485152
rect 667662 482760 667718 482769
rect 667662 482695 667718 482704
rect 669608 455025 669636 614887
rect 669792 574433 669820 638551
rect 669976 581097 670004 696934
rect 670422 696895 670478 696904
rect 670146 685944 670202 685953
rect 670146 685879 670202 685888
rect 670160 620401 670188 685879
rect 670436 620673 670464 696895
rect 670620 660113 670648 730487
rect 670804 727977 670832 750071
rect 670790 727968 670846 727977
rect 670790 727903 670846 727912
rect 670988 713697 671016 758231
rect 671172 753409 671200 869071
rect 671448 759529 671476 937479
rect 671618 775024 671674 775033
rect 671618 774959 671674 774968
rect 671434 759520 671490 759529
rect 671434 759455 671490 759464
rect 671158 753400 671214 753409
rect 671158 753335 671214 753344
rect 671158 751360 671214 751369
rect 671158 751295 671214 751304
rect 671172 728249 671200 751295
rect 671342 734904 671398 734913
rect 671342 734839 671398 734848
rect 671158 728240 671214 728249
rect 671158 728175 671214 728184
rect 671158 714096 671214 714105
rect 671158 714031 671214 714040
rect 670974 713688 671030 713697
rect 670974 713623 671030 713632
rect 670974 713280 671030 713289
rect 670974 713215 671030 713224
rect 670988 668273 671016 713215
rect 671172 669905 671200 714031
rect 671158 669896 671214 669905
rect 671158 669831 671214 669840
rect 670974 668264 671030 668273
rect 670974 668199 671030 668208
rect 671066 667992 671122 668001
rect 671066 667927 671122 667936
rect 670606 660104 670662 660113
rect 670606 660039 670662 660048
rect 670606 659696 670662 659705
rect 670606 659631 670662 659640
rect 670422 620664 670478 620673
rect 670422 620599 670478 620608
rect 670146 620392 670202 620401
rect 670146 620327 670202 620336
rect 670422 616176 670478 616185
rect 670422 616111 670478 616120
rect 670146 600400 670202 600409
rect 670146 600335 670202 600344
rect 669962 581088 670018 581097
rect 669962 581023 670018 581032
rect 669778 574424 669834 574433
rect 669778 574359 669834 574368
rect 669962 554024 670018 554033
rect 669962 553959 670018 553968
rect 669778 553480 669834 553489
rect 669778 553415 669834 553424
rect 669792 482361 669820 553415
rect 669976 551585 670004 553959
rect 669962 551576 670018 551585
rect 669962 551511 670018 551520
rect 669964 536852 670016 536858
rect 669964 536794 670016 536800
rect 669778 482352 669834 482361
rect 669778 482287 669834 482296
rect 669594 455016 669650 455025
rect 669594 454951 669650 454960
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667202 360904 667258 360913
rect 667202 360839 667258 360848
rect 667388 350600 667440 350606
rect 667388 350542 667440 350548
rect 665822 315480 665878 315489
rect 665822 315415 665878 315424
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 663062 268152 663118 268161
rect 663062 268087 663118 268096
rect 667018 237144 667074 237153
rect 667018 237079 667074 237088
rect 661868 232620 661920 232626
rect 661868 232562 661920 232568
rect 664996 232212 665048 232218
rect 664996 232154 665048 232160
rect 663798 231296 663854 231305
rect 663798 231231 663854 231240
rect 662328 231124 662380 231130
rect 662328 231066 662380 231072
rect 660946 229528 661002 229537
rect 660946 229463 661002 229472
rect 653402 229120 653458 229129
rect 653402 229055 653458 229064
rect 652390 222864 652446 222873
rect 652390 222799 652446 222808
rect 652404 213518 652432 222799
rect 653034 221504 653090 221513
rect 653034 221439 653090 221448
rect 652852 214736 652904 214742
rect 652852 214678 652904 214684
rect 652392 213512 652444 213518
rect 652392 213454 652444 213460
rect 652864 210202 652892 214678
rect 653048 210202 653076 221439
rect 653416 220114 653444 229055
rect 659476 227792 659528 227798
rect 659476 227734 659528 227740
rect 658922 226672 658978 226681
rect 658922 226607 658978 226616
rect 654782 226400 654838 226409
rect 654782 226335 654838 226344
rect 653404 220108 653456 220114
rect 653404 220050 653456 220056
rect 654796 218210 654824 226335
rect 655610 225312 655666 225321
rect 655610 225247 655666 225256
rect 655624 223650 655652 225247
rect 658186 224224 658242 224233
rect 658186 224159 658242 224168
rect 656898 223952 656954 223961
rect 656898 223887 656954 223896
rect 656162 223680 656218 223689
rect 654968 223644 655020 223650
rect 654968 223586 655020 223592
rect 655612 223644 655664 223650
rect 656162 223615 656218 223624
rect 655612 223586 655664 223592
rect 654784 218204 654836 218210
rect 654784 218146 654836 218152
rect 654980 210202 655008 223586
rect 656176 218074 656204 223615
rect 656912 222306 656940 223887
rect 657542 223136 657598 223145
rect 657542 223071 657598 223080
rect 656728 222278 656940 222306
rect 655428 218068 655480 218074
rect 655428 218010 655480 218016
rect 656164 218068 656216 218074
rect 656164 218010 656216 218016
rect 655440 210202 655468 218010
rect 656530 217288 656586 217297
rect 656530 217223 656586 217232
rect 656544 210202 656572 217223
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654580 210174 655008 210202
rect 655132 210174 655468 210202
rect 656236 210174 656572 210202
rect 656728 210202 656756 222278
rect 657556 213654 657584 223071
rect 657544 213648 657596 213654
rect 657544 213590 657596 213596
rect 658200 210202 658228 224159
rect 658936 214606 658964 226607
rect 659290 214840 659346 214849
rect 659290 214775 659346 214784
rect 658924 214600 658976 214606
rect 658924 214542 658976 214548
rect 658740 212764 658792 212770
rect 658740 212706 658792 212712
rect 658752 210202 658780 212706
rect 656728 210174 656788 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659304 210202 659332 214775
rect 659488 212770 659516 227734
rect 660762 222048 660818 222057
rect 660762 221983 660818 221992
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 659476 212764 659528 212770
rect 659476 212706 659528 212712
rect 660408 210202 660436 213862
rect 660776 213382 660804 221983
rect 660960 213926 660988 229463
rect 661682 225040 661738 225049
rect 661682 224975 661738 224984
rect 661696 214742 661724 224975
rect 662050 215112 662106 215121
rect 662050 215047 662106 215056
rect 661684 214736 661736 214742
rect 661684 214678 661736 214684
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660764 213376 660816 213382
rect 660764 213318 660816 213324
rect 660960 210202 660988 213726
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 215047
rect 662340 210202 662368 231066
rect 663062 230752 663118 230761
rect 663062 230687 663118 230696
rect 663076 213790 663104 230687
rect 663812 228154 663840 231231
rect 663628 228126 663840 228154
rect 663064 213784 663116 213790
rect 663064 213726 663116 213732
rect 663156 213512 663208 213518
rect 663156 213454 663208 213460
rect 663168 210202 663196 213454
rect 663628 210202 663656 228126
rect 665008 224954 665036 232154
rect 665822 231024 665878 231033
rect 665822 230959 665878 230968
rect 665178 230344 665234 230353
rect 665178 230279 665234 230288
rect 665192 227798 665220 230279
rect 665180 227792 665232 227798
rect 665180 227734 665232 227740
rect 665008 224926 665128 224954
rect 664166 221776 664222 221785
rect 664166 221711 664222 221720
rect 664180 213178 664208 221711
rect 664810 213752 664866 213761
rect 664810 213687 664866 213696
rect 664168 213172 664220 213178
rect 664168 213114 664220 213120
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 213687
rect 665100 213042 665128 224926
rect 665836 213518 665864 230959
rect 666836 224460 666888 224466
rect 666836 224402 666888 224408
rect 666848 223961 666876 224402
rect 666834 223952 666890 223961
rect 666834 223887 666890 223896
rect 665824 213512 665876 213518
rect 665824 213454 665876 213460
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 659304 210174 659548 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663656 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 652208 209568 652260 209574
rect 652208 209510 652260 209516
rect 666836 209568 666888 209574
rect 666836 209510 666888 209516
rect 632164 209494 632500 209510
rect 666652 209092 666704 209098
rect 666652 209034 666704 209040
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 207664 589516 207670
rect 589464 207606 589516 207612
rect 589476 206417 589504 207606
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 581736 206304 581788 206310
rect 581736 206246 581788 206252
rect 589648 206304 589700 206310
rect 589648 206246 589700 206252
rect 589660 204785 589688 206246
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 581564 200086 581684 200114
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580448 151836 580500 151842
rect 580448 151778 580500 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 579252 145308 579304 145314
rect 579252 145250 579304 145256
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 579068 136876 579120 136882
rect 579068 136818 579120 136824
rect 579080 132297 579108 136818
rect 579264 136649 579292 145250
rect 579528 144696 579580 144702
rect 579526 144664 579528 144673
rect 579580 144664 579582 144673
rect 579526 144599 579582 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580460 140758 580488 151778
rect 580448 140752 580500 140758
rect 580448 140694 580500 140700
rect 580264 139460 580316 139466
rect 580264 139402 580316 139408
rect 579250 136640 579306 136649
rect 579250 136575 579306 136584
rect 579528 135176 579580 135182
rect 579528 135118 579580 135124
rect 579540 134473 579568 135118
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131300 578936 131306
rect 578884 131242 578936 131248
rect 578332 124160 578384 124166
rect 578332 124102 578384 124108
rect 578344 123593 578372 124102
rect 578330 123584 578386 123593
rect 578330 123519 578386 123528
rect 578700 118584 578752 118590
rect 578700 118526 578752 118532
rect 578712 118425 578740 118526
rect 578698 118416 578754 118425
rect 578698 118351 578754 118360
rect 578700 117224 578752 117230
rect 578700 117166 578752 117172
rect 578712 116929 578740 117166
rect 578698 116920 578754 116929
rect 578698 116855 578754 116864
rect 578896 110401 578924 131242
rect 579068 131164 579120 131170
rect 579068 131106 579120 131112
rect 579080 129713 579108 131106
rect 579066 129704 579122 129713
rect 579066 129639 579122 129648
rect 579160 128308 579212 128314
rect 579160 128250 579212 128256
rect 579172 127809 579200 128250
rect 579158 127800 579214 127809
rect 579158 127735 579214 127744
rect 579068 126268 579120 126274
rect 579068 126210 579120 126216
rect 579080 113174 579108 126210
rect 579528 125384 579580 125390
rect 579526 125352 579528 125361
rect 579580 125352 579582 125361
rect 579526 125287 579582 125296
rect 580276 124166 580304 139402
rect 580632 131776 580684 131782
rect 580632 131718 580684 131724
rect 580264 124160 580316 124166
rect 580264 124102 580316 124108
rect 580448 122868 580500 122874
rect 580448 122810 580500 122816
rect 579528 121440 579580 121446
rect 579528 121382 579580 121388
rect 579540 121145 579568 121382
rect 579526 121136 579582 121145
rect 579526 121071 579582 121080
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 578988 113146 579108 113174
rect 578988 110514 579016 113146
rect 579160 113076 579212 113082
rect 579160 113018 579212 113024
rect 579172 112577 579200 113018
rect 579158 112568 579214 112577
rect 579158 112503 579214 112512
rect 578988 110486 579108 110514
rect 578882 110392 578938 110401
rect 578882 110327 578938 110336
rect 578884 108996 578936 109002
rect 578884 108938 578936 108944
rect 578896 108361 578924 108938
rect 578882 108352 578938 108361
rect 578882 108287 578938 108296
rect 579080 105913 579108 110486
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 579344 105188 579396 105194
rect 579344 105130 579396 105136
rect 578332 103352 578384 103358
rect 578330 103320 578332 103329
rect 578384 103320 578386 103329
rect 578330 103255 578386 103264
rect 578516 102128 578568 102134
rect 578516 102070 578568 102076
rect 578528 101697 578556 102070
rect 578514 101688 578570 101697
rect 578514 101623 578570 101632
rect 579160 99272 579212 99278
rect 579158 99240 579160 99249
rect 579212 99240 579214 99249
rect 579158 99175 579214 99184
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 577504 95940 577556 95946
rect 577504 95882 577556 95888
rect 574928 57384 574980 57390
rect 574928 57326 574980 57332
rect 574744 56024 574796 56030
rect 574744 55966 574796 55972
rect 574560 55888 574612 55894
rect 574560 55830 574612 55836
rect 574572 54126 574600 55830
rect 574756 55049 574784 55966
rect 574742 55040 574798 55049
rect 574742 54975 574798 54984
rect 574560 54120 574612 54126
rect 574560 54062 574612 54068
rect 574940 53990 574968 57326
rect 575480 57248 575532 57254
rect 575480 57190 575532 57196
rect 575492 54233 575520 57190
rect 577516 55214 577544 95882
rect 579160 93424 579212 93430
rect 579160 93366 579212 93372
rect 579172 93129 579200 93366
rect 579158 93120 579214 93129
rect 579158 93055 579214 93064
rect 578516 91724 578568 91730
rect 578516 91666 578568 91672
rect 578528 90953 578556 91666
rect 578514 90944 578570 90953
rect 578514 90879 578570 90888
rect 578516 88324 578568 88330
rect 578516 88266 578568 88272
rect 578528 88097 578556 88266
rect 578514 88088 578570 88097
rect 578514 88023 578570 88032
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 579068 85468 579120 85474
rect 579068 85410 579120 85416
rect 578516 82612 578568 82618
rect 578516 82554 578568 82560
rect 578528 82249 578556 82554
rect 578514 82240 578570 82249
rect 578514 82175 578570 82184
rect 578516 78464 578568 78470
rect 578516 78406 578568 78412
rect 578528 77897 578556 78406
rect 578514 77888 578570 77897
rect 578514 77823 578570 77832
rect 579080 75721 579108 85410
rect 579356 80073 579384 105130
rect 580264 104168 580316 104174
rect 580264 104110 580316 104116
rect 579528 95056 579580 95062
rect 579526 95024 579528 95033
rect 579580 95024 579582 95033
rect 579526 94959 579582 94968
rect 579528 84040 579580 84046
rect 579526 84008 579528 84017
rect 579580 84008 579582 84017
rect 579526 83943 579582 83952
rect 579342 80064 579398 80073
rect 579342 79999 579398 80008
rect 580276 78470 580304 104110
rect 580460 102134 580488 122810
rect 580644 117230 580672 131718
rect 580632 117224 580684 117230
rect 580632 117166 580684 117172
rect 581656 114510 581684 200086
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 666664 178537 666692 209034
rect 666650 178528 666706 178537
rect 666650 178463 666706 178472
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 145314 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 145308 585192 145314
rect 585140 145250 585192 145256
rect 585968 144968 586020 144974
rect 585968 144910 586020 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 584588 143608 584640 143614
rect 584588 143550 584640 143556
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 140820 583076 140826
rect 583024 140762 583076 140768
rect 583036 125390 583064 140762
rect 584404 135312 584456 135318
rect 584404 135254 584456 135260
rect 583024 125384 583076 125390
rect 583024 125326 583076 125332
rect 583208 124908 583260 124914
rect 583208 124850 583260 124856
rect 581828 122120 581880 122126
rect 581828 122062 581880 122068
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 111104 581696 111110
rect 581644 111046 581696 111052
rect 581276 107704 581328 107710
rect 581276 107646 581328 107652
rect 581288 105194 581316 107646
rect 581276 105188 581328 105194
rect 581276 105130 581328 105136
rect 580448 102128 580500 102134
rect 580448 102070 580500 102076
rect 580448 100020 580500 100026
rect 580448 99962 580500 99968
rect 580460 86970 580488 99962
rect 581656 99278 581684 111046
rect 581840 109002 581868 122062
rect 583024 109744 583076 109750
rect 583024 109686 583076 109692
rect 581828 108996 581880 109002
rect 581828 108938 581880 108944
rect 581828 104916 581880 104922
rect 581828 104858 581880 104864
rect 581644 99272 581696 99278
rect 581644 99214 581696 99220
rect 581644 89004 581696 89010
rect 581644 88946 581696 88952
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 580264 78464 580316 78470
rect 580264 78406 580316 78412
rect 580446 77888 580502 77897
rect 580446 77823 580502 77832
rect 579344 76560 579396 76566
rect 579344 76502 579396 76508
rect 579066 75712 579122 75721
rect 579066 75647 579122 75656
rect 578516 71596 578568 71602
rect 578516 71538 578568 71544
rect 578528 71233 578556 71538
rect 578514 71224 578570 71233
rect 578514 71159 578570 71168
rect 579068 58812 579120 58818
rect 579068 58754 579120 58760
rect 577688 58676 577740 58682
rect 577688 58618 577740 58624
rect 577504 55208 577556 55214
rect 577504 55150 577556 55156
rect 575478 54224 575534 54233
rect 575478 54159 575534 54168
rect 574928 53984 574980 53990
rect 577700 53961 577728 58618
rect 578516 56568 578568 56574
rect 578516 56510 578568 56516
rect 578528 56137 578556 56510
rect 578514 56128 578570 56137
rect 578514 56063 578570 56072
rect 579080 54262 579108 58754
rect 579356 57905 579384 76502
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 62076 579580 62082
rect 579528 62018 579580 62024
rect 579540 61849 579568 62018
rect 579526 61840 579582 61849
rect 579526 61775 579582 61784
rect 579528 60716 579580 60722
rect 579528 60658 579580 60664
rect 579540 60353 579568 60658
rect 579526 60344 579582 60353
rect 579526 60279 579582 60288
rect 579342 57896 579398 57905
rect 579342 57831 579398 57840
rect 580460 54398 580488 77823
rect 581656 54505 581684 88946
rect 581840 85474 581868 104858
rect 581828 85468 581880 85474
rect 581828 85410 581880 85416
rect 583036 84046 583064 109686
rect 583220 103358 583248 124850
rect 584416 118590 584444 135254
rect 584600 131170 584628 143550
rect 585980 136882 586008 144910
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 136876 586020 136882
rect 585968 136818 586020 136824
rect 585784 136672 585836 136678
rect 585784 136614 585836 136620
rect 584588 131164 584640 131170
rect 584588 131106 584640 131112
rect 585796 121446 585824 136614
rect 587176 128314 587204 142394
rect 588556 135182 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 135318 589504 136167
rect 589464 135312 589516 135318
rect 589464 135254 589516 135260
rect 588544 135176 588596 135182
rect 588544 135118 588596 135124
rect 590290 134600 590346 134609
rect 590290 134535 590346 134544
rect 588726 132968 588782 132977
rect 588726 132903 588782 132912
rect 587164 128308 587216 128314
rect 587164 128250 587216 128256
rect 587624 127220 587676 127226
rect 587624 127162 587676 127168
rect 587636 126274 587664 127162
rect 587624 126268 587676 126274
rect 587624 126210 587676 126216
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585784 121440 585836 121446
rect 585784 121382 585836 121388
rect 584588 118720 584640 118726
rect 584588 118662 584640 118668
rect 584404 118584 584456 118590
rect 584404 118526 584456 118532
rect 584404 113212 584456 113218
rect 584404 113154 584456 113160
rect 583208 103352 583260 103358
rect 583208 103294 583260 103300
rect 583024 84040 583076 84046
rect 583024 83982 583076 83988
rect 584416 82618 584444 113154
rect 584600 95062 584628 118662
rect 585968 117360 586020 117366
rect 585968 117302 586020 117308
rect 585784 116000 585836 116006
rect 585784 115942 585836 115948
rect 584588 95056 584640 95062
rect 584588 94998 584640 95004
rect 585796 91730 585824 115942
rect 585980 93430 586008 117302
rect 587164 100768 587216 100774
rect 587164 100710 587216 100716
rect 585968 93424 586020 93430
rect 585968 93366 586020 93372
rect 585784 91724 585836 91730
rect 585784 91666 585836 91672
rect 584404 82612 584456 82618
rect 584404 82554 584456 82560
rect 584404 79348 584456 79354
rect 584404 79290 584456 79296
rect 584416 71602 584444 79290
rect 587176 73166 587204 100710
rect 587360 97986 587388 121450
rect 588740 113082 588768 132903
rect 590304 131782 590332 134535
rect 666848 133113 666876 209510
rect 667032 160041 667060 237079
rect 667018 160032 667074 160041
rect 667018 159967 667074 159976
rect 667216 141409 667244 310490
rect 667400 181393 667428 350542
rect 667756 324352 667808 324358
rect 667756 324294 667808 324300
rect 667572 284368 667624 284374
rect 667572 284310 667624 284316
rect 667386 181384 667442 181393
rect 667386 181319 667442 181328
rect 667202 141400 667258 141409
rect 667202 141335 667258 141344
rect 667584 135969 667612 284310
rect 667768 178809 667796 324294
rect 668596 311953 668624 444382
rect 669976 403753 670004 536794
rect 670160 529961 670188 600335
rect 670146 529952 670202 529961
rect 670146 529887 670202 529896
rect 670436 455297 670464 616111
rect 670620 455841 670648 659631
rect 670882 647320 670938 647329
rect 670882 647255 670938 647264
rect 670896 574841 670924 647255
rect 671080 623529 671108 667927
rect 671356 663794 671384 734839
rect 671632 705537 671660 774959
rect 671816 760073 671844 938295
rect 672170 938088 672226 938097
rect 672170 938023 672226 938032
rect 672184 937281 672212 938023
rect 672722 937816 672778 937825
rect 672722 937751 672778 937760
rect 672736 937281 672764 937751
rect 672170 937272 672226 937281
rect 672170 937207 672226 937216
rect 672722 937272 672778 937281
rect 672722 937207 672778 937216
rect 672354 936728 672410 936737
rect 672354 936663 672410 936672
rect 671986 929520 672042 929529
rect 671986 929455 672042 929464
rect 671802 760064 671858 760073
rect 671802 759999 671858 760008
rect 671802 757480 671858 757489
rect 671802 757415 671858 757424
rect 671816 712881 671844 757415
rect 672000 732873 672028 929455
rect 672170 759792 672226 759801
rect 672170 759727 672226 759736
rect 671986 732864 672042 732873
rect 671986 732799 672042 732808
rect 671986 730144 672042 730153
rect 671986 730079 672042 730088
rect 671802 712872 671858 712881
rect 671802 712807 671858 712816
rect 671618 705528 671674 705537
rect 671618 705463 671674 705472
rect 671802 687440 671858 687449
rect 671802 687375 671858 687384
rect 671618 670304 671674 670313
rect 671618 670239 671674 670248
rect 671632 668794 671660 670239
rect 671632 668766 671752 668794
rect 671526 668672 671582 668681
rect 671526 668607 671582 668616
rect 671540 663794 671568 668607
rect 671724 663794 671752 668766
rect 671264 663766 671384 663794
rect 671448 663766 671568 663794
rect 671632 663766 671752 663794
rect 671264 661337 671292 663766
rect 671250 661328 671306 661337
rect 671250 661263 671306 661272
rect 671448 624345 671476 663766
rect 671632 625161 671660 663766
rect 671618 625152 671674 625161
rect 671618 625087 671674 625096
rect 671618 624744 671674 624753
rect 671618 624679 671674 624688
rect 671434 624336 671490 624345
rect 671434 624271 671490 624280
rect 671250 623928 671306 623937
rect 671250 623863 671306 623872
rect 671066 623520 671122 623529
rect 671066 623455 671122 623464
rect 671066 622296 671122 622305
rect 671066 622231 671122 622240
rect 671080 616214 671108 622231
rect 671068 616208 671120 616214
rect 671068 616150 671120 616156
rect 671066 594824 671122 594833
rect 671066 594759 671122 594768
rect 670882 574832 670938 574841
rect 670882 574767 670938 574776
rect 670882 552120 670938 552129
rect 670882 552055 670938 552064
rect 670896 483993 670924 552055
rect 671080 524929 671108 594759
rect 671264 578921 671292 623863
rect 671434 623112 671490 623121
rect 671434 623047 671490 623056
rect 671448 582374 671476 623047
rect 671632 621014 671660 624679
rect 671356 582346 671476 582374
rect 671540 620986 671660 621014
rect 671356 580666 671384 582346
rect 671540 580825 671568 620986
rect 671816 618225 671844 687375
rect 672000 665689 672028 730079
rect 672184 715329 672212 759727
rect 672368 758713 672396 936663
rect 672538 935776 672594 935785
rect 672538 935711 672594 935720
rect 672354 758704 672410 758713
rect 672354 758639 672410 758648
rect 672552 758554 672580 935711
rect 673012 933473 673040 952167
rect 672998 933464 673054 933473
rect 672998 933399 673054 933408
rect 673196 930617 673224 958151
rect 673380 932657 673408 962775
rect 674102 957128 674158 957137
rect 674102 957063 674158 957072
rect 673366 932648 673422 932657
rect 673366 932583 673422 932592
rect 673182 930608 673238 930617
rect 673182 930543 673238 930552
rect 674116 930209 674144 957063
rect 674300 933065 674328 966062
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675298 964744 675354 964753
rect 675298 964679 675354 964688
rect 675312 962418 675340 964679
rect 675496 963393 675524 963595
rect 675482 963384 675538 963393
rect 675482 963319 675538 963328
rect 675496 962849 675524 963016
rect 675482 962840 675538 962849
rect 675482 962775 675538 962784
rect 675312 962390 675418 962418
rect 675220 961741 675418 961769
rect 674470 959440 674526 959449
rect 674470 959375 674526 959384
rect 674484 933881 674512 959375
rect 674930 959168 674986 959177
rect 674986 959112 675064 959114
rect 674930 959103 675064 959112
rect 674944 959086 675064 959103
rect 674654 958896 674710 958905
rect 674654 958831 674710 958840
rect 674668 956354 674696 958831
rect 674576 956326 674696 956354
rect 674576 954122 674604 956326
rect 674576 954094 674696 954122
rect 674470 933872 674526 933881
rect 674470 933807 674526 933816
rect 674286 933056 674342 933065
rect 674286 932991 674342 933000
rect 674668 931025 674696 954094
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 931016 674710 931025
rect 674654 930951 674710 930960
rect 674102 930200 674158 930209
rect 674102 930135 674158 930144
rect 674852 928792 674880 953391
rect 675036 949454 675064 959086
rect 675220 958905 675248 961741
rect 675390 959440 675446 959449
rect 675390 959375 675446 959384
rect 675404 959276 675432 959375
rect 675206 958896 675262 958905
rect 675206 958831 675262 958840
rect 675312 958718 675418 958746
rect 675312 958225 675340 958718
rect 675298 958216 675354 958225
rect 675298 958151 675354 958160
rect 675772 957817 675800 958052
rect 675298 957808 675354 957817
rect 675298 957743 675354 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 675312 955482 675340 957743
rect 675496 957137 675524 957440
rect 675482 957128 675538 957137
rect 675482 957063 675538 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675220 954366 675418 954394
rect 675220 951561 675248 954366
rect 675404 953465 675432 953768
rect 675390 953456 675446 953465
rect 675390 953391 675446 953400
rect 675496 952241 675524 952544
rect 675482 952232 675538 952241
rect 675482 952167 675538 952176
rect 675206 951552 675262 951561
rect 675206 951487 675262 951496
rect 675850 951552 675906 951561
rect 675850 951487 675906 951496
rect 675864 949482 675892 951487
rect 683302 950736 683358 950745
rect 683302 950671 683358 950680
rect 675852 949476 675904 949482
rect 675036 949426 675156 949454
rect 675128 934289 675156 949426
rect 675852 949418 675904 949424
rect 682384 949476 682436 949482
rect 682384 949418 682436 949424
rect 675298 949240 675354 949249
rect 675298 949175 675354 949184
rect 675312 946694 675340 949175
rect 679622 948832 679678 948841
rect 679622 948767 679678 948776
rect 675220 946666 675340 946694
rect 675220 943934 675248 946666
rect 675220 943906 675524 943934
rect 675496 934697 675524 943906
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 679636 935649 679664 948767
rect 679622 935640 679678 935649
rect 679622 935575 679678 935584
rect 682396 935241 682424 949418
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 675482 934688 675538 934697
rect 675482 934623 675538 934632
rect 675114 934280 675170 934289
rect 675114 934215 675170 934224
rect 683316 932385 683344 950671
rect 683486 947336 683542 947345
rect 683486 947271 683542 947280
rect 683500 939729 683528 947271
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683486 939720 683542 939729
rect 683486 939655 683542 939664
rect 683302 932376 683358 932385
rect 683302 932311 683358 932320
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 673182 928296 673238 928305
rect 673182 928231 673238 928240
rect 672998 869408 673054 869417
rect 672998 869343 673054 869352
rect 672814 784408 672870 784417
rect 672814 784343 672870 784352
rect 672828 780722 672856 784343
rect 672828 780694 672948 780722
rect 672722 780600 672778 780609
rect 672722 780535 672778 780544
rect 672736 775690 672764 780535
rect 672460 758526 672580 758554
rect 672644 775662 672764 775690
rect 672460 757897 672488 758526
rect 672446 757888 672502 757897
rect 672446 757823 672502 757832
rect 672354 734224 672410 734233
rect 672354 734159 672410 734168
rect 672170 715320 672226 715329
rect 672170 715255 672226 715264
rect 672170 689072 672226 689081
rect 672170 689007 672226 689016
rect 671986 665680 672042 665689
rect 671986 665615 672042 665624
rect 671986 661056 672042 661065
rect 671986 660991 672042 661000
rect 671802 618216 671858 618225
rect 671802 618151 671858 618160
rect 671712 616208 671764 616214
rect 671712 616150 671764 616156
rect 671724 601694 671752 616150
rect 671724 601666 671844 601694
rect 671526 580816 671582 580825
rect 671526 580751 671582 580760
rect 671356 580638 671660 580666
rect 671434 579320 671490 579329
rect 671434 579255 671490 579264
rect 671250 578912 671306 578921
rect 671250 578847 671306 578856
rect 671448 578082 671476 579255
rect 671632 578270 671660 580638
rect 671620 578264 671672 578270
rect 671620 578206 671672 578212
rect 671264 578054 671476 578082
rect 671264 534721 671292 578054
rect 671436 577992 671488 577998
rect 671436 577934 671488 577940
rect 671448 577833 671476 577934
rect 671434 577824 671490 577833
rect 671434 577759 671490 577768
rect 671618 577552 671674 577561
rect 671618 577487 671674 577496
rect 671434 576872 671490 576881
rect 671434 576807 671490 576816
rect 671250 534712 671306 534721
rect 671250 534647 671306 534656
rect 671448 533089 671476 576807
rect 671434 533080 671490 533089
rect 671434 533015 671490 533024
rect 671632 531457 671660 577487
rect 671816 577289 671844 601666
rect 671802 577280 671858 577289
rect 671802 577215 671858 577224
rect 671802 569528 671858 569537
rect 671802 569463 671858 569472
rect 671618 531448 671674 531457
rect 671618 531383 671674 531392
rect 671066 524920 671122 524929
rect 671066 524855 671122 524864
rect 670882 483984 670938 483993
rect 670882 483919 670938 483928
rect 670606 455832 670662 455841
rect 670606 455767 670662 455776
rect 670422 455288 670478 455297
rect 670422 455223 670478 455232
rect 671816 455054 671844 569463
rect 672000 501673 672028 660991
rect 672184 616593 672212 689007
rect 672368 662833 672396 734159
rect 672644 710433 672672 775662
rect 672920 775574 672948 780694
rect 672736 775546 672948 775574
rect 672736 712094 672764 775546
rect 673012 751777 673040 869343
rect 673196 785234 673224 928231
rect 675220 877662 675524 877690
rect 675220 877554 675248 877662
rect 674944 877526 675248 877554
rect 675496 877540 675524 877662
rect 674944 873497 674972 877526
rect 675312 876982 675432 877010
rect 675114 876888 675170 876897
rect 675312 876874 675340 876982
rect 675170 876846 675340 876874
rect 675404 876860 675432 876982
rect 675114 876823 675170 876832
rect 675114 876344 675170 876353
rect 675114 876279 675170 876288
rect 675128 873882 675156 876279
rect 675680 875945 675708 876248
rect 675666 875936 675722 875945
rect 675666 875871 675722 875880
rect 675772 874177 675800 874412
rect 675758 874168 675814 874177
rect 675758 874103 675814 874112
rect 675128 873854 675340 873882
rect 675312 873746 675340 873854
rect 675404 873746 675432 873868
rect 675312 873718 675432 873746
rect 674930 873488 674986 873497
rect 674930 873423 674986 873432
rect 675114 873216 675170 873225
rect 675170 873174 675418 873202
rect 675114 873151 675170 873160
rect 675588 872273 675616 872576
rect 675114 872264 675170 872273
rect 675114 872199 675170 872208
rect 675574 872264 675630 872273
rect 675574 872199 675630 872208
rect 675128 870074 675156 872199
rect 675128 870046 675418 870074
rect 674116 869502 675418 869530
rect 673918 864784 673974 864793
rect 673918 864719 673974 864728
rect 673196 785206 673316 785234
rect 673288 760345 673316 785206
rect 673734 779240 673790 779249
rect 673734 779175 673790 779184
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673274 760336 673330 760345
rect 673274 760271 673330 760280
rect 673366 759112 673422 759121
rect 673366 759047 673422 759056
rect 672998 751768 673054 751777
rect 672998 751703 673054 751712
rect 673380 734174 673408 759047
rect 673288 734146 673408 734174
rect 672908 734052 672960 734058
rect 672908 733994 672960 734000
rect 672920 725529 672948 733994
rect 673288 733938 673316 734146
rect 673564 734058 673592 777407
rect 673748 765914 673776 779175
rect 673932 772041 673960 864719
rect 673918 772032 673974 772041
rect 673918 771967 673974 771976
rect 673748 765886 673868 765914
rect 673840 746594 673868 765886
rect 674116 754361 674144 869502
rect 675114 869408 675170 869417
rect 675114 869343 675170 869352
rect 674930 869136 674986 869145
rect 674930 869071 674986 869080
rect 674654 868728 674710 868737
rect 674710 868686 674880 868714
rect 674654 868663 674710 868672
rect 674654 868456 674710 868465
rect 674654 868391 674710 868400
rect 674470 788080 674526 788089
rect 674470 788015 674526 788024
rect 674286 778696 674342 778705
rect 674286 778631 674342 778640
rect 674102 754352 674158 754361
rect 674102 754287 674158 754296
rect 673656 746566 673868 746594
rect 673656 743834 673684 746566
rect 673656 743806 674052 743834
rect 673826 741704 673882 741713
rect 673826 741639 673882 741648
rect 673840 738154 673868 741639
rect 673656 738126 673868 738154
rect 673656 734174 673684 738126
rect 674024 734174 674052 743806
rect 673656 734146 673776 734174
rect 674024 734146 674144 734174
rect 673552 734052 673604 734058
rect 673552 733994 673604 734000
rect 673288 733910 673408 733938
rect 673182 733000 673238 733009
rect 673182 732935 673238 732944
rect 673196 728668 673224 732935
rect 673196 728640 673316 728668
rect 673090 728512 673146 728521
rect 673090 728447 673092 728456
rect 673144 728447 673146 728456
rect 673092 728418 673144 728424
rect 672906 725520 672962 725529
rect 672906 725455 672962 725464
rect 673288 717614 673316 728640
rect 673104 717586 673316 717614
rect 672906 714912 672962 714921
rect 672906 714847 672962 714856
rect 672736 712066 672856 712094
rect 672630 710424 672686 710433
rect 672630 710359 672686 710368
rect 672828 710274 672856 712066
rect 672644 710246 672856 710274
rect 672644 709209 672672 710246
rect 672630 709200 672686 709209
rect 672630 709135 672686 709144
rect 672540 707260 672592 707266
rect 672540 707202 672592 707208
rect 672552 667457 672580 707202
rect 672920 702434 672948 714847
rect 672828 702406 672948 702434
rect 672828 669497 672856 702406
rect 672814 669488 672870 669497
rect 672814 669423 672870 669432
rect 672538 667448 672594 667457
rect 672538 667383 672594 667392
rect 672722 666632 672778 666641
rect 672722 666567 672778 666576
rect 672354 662824 672410 662833
rect 672354 662759 672410 662768
rect 672538 647864 672594 647873
rect 672538 647799 672594 647808
rect 672552 640334 672580 647799
rect 672460 640306 672580 640334
rect 672170 616584 672226 616593
rect 672170 616519 672226 616528
rect 672262 607336 672318 607345
rect 672262 607271 672318 607280
rect 672276 538214 672304 607271
rect 672460 571985 672488 640306
rect 672736 635497 672764 666567
rect 673104 661609 673132 717586
rect 673380 714513 673408 733910
rect 673748 732578 673776 734146
rect 673472 732550 673776 732578
rect 673472 717614 673500 732550
rect 674116 728770 674144 734146
rect 673748 728742 674144 728770
rect 673748 724514 673776 728742
rect 674104 728680 674156 728686
rect 674102 728648 674104 728657
rect 674156 728648 674158 728657
rect 674102 728583 674158 728592
rect 673918 728240 673974 728249
rect 673918 728175 673920 728184
rect 673972 728175 673974 728184
rect 673920 728146 673972 728152
rect 674150 728136 674202 728142
rect 674150 728078 674202 728084
rect 674162 727977 674190 728078
rect 674148 727968 674204 727977
rect 674148 727903 674204 727912
rect 674300 726889 674328 778631
rect 674484 746594 674512 788015
rect 674668 770681 674696 868391
rect 674852 866946 674880 868686
rect 674944 867049 674972 869071
rect 675128 868238 675156 869343
rect 675312 868861 675418 868889
rect 675312 868465 675340 868861
rect 675298 868456 675354 868465
rect 675298 868391 675354 868400
rect 675128 868210 675418 868238
rect 674944 867021 675418 867049
rect 674852 866918 675156 866946
rect 674930 866688 674986 866697
rect 674930 866623 674986 866632
rect 674944 864566 674972 866623
rect 675128 865858 675156 866918
rect 675128 865830 675418 865858
rect 675128 865181 675418 865209
rect 675128 864793 675156 865181
rect 675114 864784 675170 864793
rect 675114 864719 675170 864728
rect 674944 864538 675418 864566
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675220 863314 675340 863342
rect 675404 863328 675432 863382
rect 675220 794894 675248 863314
rect 674852 794866 675248 794894
rect 674852 780881 674880 794866
rect 675114 789440 675170 789449
rect 675114 789375 675170 789384
rect 675128 787693 675156 789375
rect 675312 788310 675418 788338
rect 675312 788089 675340 788310
rect 675298 788080 675354 788089
rect 675298 788015 675354 788024
rect 675128 787665 675418 787693
rect 674944 787018 675418 787046
rect 674944 785234 674972 787018
rect 674944 785206 675064 785234
rect 674838 780872 674894 780881
rect 674838 780807 674894 780816
rect 675036 779226 675064 785206
rect 674944 779198 675064 779226
rect 675128 785182 675418 785210
rect 674944 776030 674972 779198
rect 675128 779090 675156 785182
rect 675404 784417 675432 784652
rect 675390 784408 675446 784417
rect 675390 784343 675446 784352
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675404 783057 675432 783360
rect 675390 783048 675446 783057
rect 675390 782983 675446 782992
rect 675482 782504 675538 782513
rect 675312 782462 675482 782490
rect 675312 780450 675340 782462
rect 675482 782439 675538 782448
rect 675496 780609 675524 780844
rect 675482 780600 675538 780609
rect 675482 780535 675538 780544
rect 675312 780422 675432 780450
rect 675404 780300 675432 780422
rect 675312 779674 675418 779702
rect 675312 779249 675340 779674
rect 675298 779240 675354 779249
rect 675298 779175 675354 779184
rect 675036 779062 675156 779090
rect 675036 776506 675064 779062
rect 675206 778968 675262 778977
rect 675206 778903 675262 778912
rect 675220 776642 675248 778903
rect 675496 778705 675524 779008
rect 675482 778696 675538 778705
rect 675482 778631 675538 778640
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675220 776614 675418 776642
rect 675482 776520 675538 776529
rect 675036 776478 675248 776506
rect 674944 776002 675064 776030
rect 674838 775704 674894 775713
rect 674838 775639 674894 775648
rect 674852 774625 674880 775639
rect 674838 774616 674894 774625
rect 674838 774551 674894 774560
rect 675036 772814 675064 776002
rect 674944 772786 675064 772814
rect 675220 772814 675248 776478
rect 675482 776455 675538 776464
rect 675496 776016 675524 776455
rect 675404 775033 675432 775336
rect 675390 775024 675446 775033
rect 675390 774959 675446 774968
rect 675482 774616 675538 774625
rect 675482 774551 675538 774560
rect 675496 774180 675524 774551
rect 675220 772786 675340 772814
rect 674654 770672 674710 770681
rect 674654 770607 674710 770616
rect 674944 766601 674972 772786
rect 674930 766592 674986 766601
rect 675312 766578 675340 772786
rect 683210 772032 683266 772041
rect 683210 771967 683266 771976
rect 678242 771488 678298 771497
rect 678242 771423 678298 771432
rect 676126 766592 676182 766601
rect 675312 766550 676126 766578
rect 674930 766527 674986 766536
rect 676126 766527 676182 766536
rect 676034 763056 676090 763065
rect 676034 762991 676090 763000
rect 676048 760753 676076 762991
rect 676954 761832 677010 761841
rect 676586 761788 676642 761797
rect 676954 761767 677010 761776
rect 676586 761723 676642 761732
rect 676034 760744 676090 760753
rect 676034 760679 676090 760688
rect 676034 756392 676090 756401
rect 676034 756327 676090 756336
rect 675850 754352 675906 754361
rect 675850 754287 675852 754296
rect 675904 754287 675906 754296
rect 675852 754258 675904 754264
rect 676048 753817 676076 756327
rect 676034 753808 676090 753817
rect 676034 753743 676090 753752
rect 676600 753642 676628 761723
rect 676968 755041 676996 761767
rect 678256 757081 678284 771423
rect 682382 768768 682438 768777
rect 682382 768703 682438 768712
rect 678242 757072 678298 757081
rect 678242 757007 678298 757016
rect 682396 755857 682424 768703
rect 683224 756673 683252 771967
rect 683394 770672 683450 770681
rect 683394 770607 683450 770616
rect 683210 756664 683266 756673
rect 683210 756599 683266 756608
rect 682382 755848 682438 755857
rect 682382 755783 682438 755792
rect 676954 755032 677010 755041
rect 676954 754967 677010 754976
rect 683120 754316 683172 754322
rect 683120 754258 683172 754264
rect 676036 753636 676088 753642
rect 676036 753578 676088 753584
rect 676588 753636 676640 753642
rect 676588 753578 676640 753584
rect 676048 752593 676076 753578
rect 676034 752584 676090 752593
rect 676034 752519 676090 752528
rect 683132 752185 683160 754258
rect 683408 753001 683436 770607
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683394 752992 683450 753001
rect 683394 752927 683450 752936
rect 683118 752176 683174 752185
rect 683118 752111 683174 752120
rect 674484 746566 674604 746594
rect 674286 726880 674342 726889
rect 674286 726815 674342 726824
rect 674576 726617 674604 746566
rect 675128 743294 675418 743322
rect 675128 743209 675156 743294
rect 675114 743200 675170 743209
rect 675114 743135 675170 743144
rect 675128 742682 675340 742710
rect 675128 742257 675156 742682
rect 675312 742642 675340 742682
rect 675404 742642 675432 742696
rect 675312 742614 675432 742642
rect 675298 742520 675354 742529
rect 675298 742455 675354 742464
rect 675114 742248 675170 742257
rect 675114 742183 675170 742192
rect 675114 741160 675170 741169
rect 675114 741095 675170 741104
rect 675128 739650 675156 741095
rect 675312 740194 675340 742455
rect 675496 741713 675524 742016
rect 675482 741704 675538 741713
rect 675482 741639 675538 741648
rect 675312 740166 675418 740194
rect 675128 739622 675418 739650
rect 674930 738984 674986 738993
rect 674930 738919 674986 738928
rect 674944 736934 674972 738919
rect 675404 738721 675432 739024
rect 675390 738712 675446 738721
rect 675390 738647 675446 738656
rect 675128 738330 675418 738358
rect 675128 738177 675156 738330
rect 675114 738168 675170 738177
rect 675114 738103 675170 738112
rect 674944 736906 675156 736934
rect 675128 735910 675156 736906
rect 675128 735882 675340 735910
rect 675312 735842 675340 735882
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 674930 735312 674986 735321
rect 674930 735247 674986 735256
rect 675128 735305 675418 735333
rect 674944 731626 674972 735247
rect 675128 734913 675156 735305
rect 675114 734904 675170 734913
rect 675114 734839 675170 734848
rect 675128 734658 675418 734686
rect 675128 734233 675156 734658
rect 675114 734224 675170 734233
rect 675114 734159 675170 734168
rect 675312 734017 675418 734045
rect 675114 733680 675170 733689
rect 675114 733615 675170 733624
rect 675128 732850 675156 733615
rect 675312 733009 675340 734017
rect 675298 733000 675354 733009
rect 675298 732935 675354 732944
rect 675128 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674944 731598 675340 731626
rect 675404 731612 675432 731734
rect 674930 731504 674986 731513
rect 674930 731439 674986 731448
rect 674944 729178 674972 731439
rect 675128 730986 675418 731014
rect 675128 730153 675156 730986
rect 675298 730552 675354 730561
rect 675298 730487 675354 730496
rect 675312 730365 675340 730487
rect 675312 730337 675418 730365
rect 675114 730144 675170 730153
rect 675114 730079 675170 730088
rect 674944 729150 675418 729178
rect 683118 726880 683174 726889
rect 683118 726815 683174 726824
rect 674562 726608 674618 726617
rect 674562 726543 674618 726552
rect 681002 725792 681058 725801
rect 681002 725727 681058 725736
rect 673656 724486 673776 724514
rect 673656 724033 673684 724486
rect 677324 724260 677376 724266
rect 677324 724202 677376 724208
rect 677336 724033 677364 724202
rect 673642 724024 673698 724033
rect 673642 723959 673698 723968
rect 677322 724024 677378 724033
rect 677322 723959 677378 723968
rect 673472 717586 673684 717614
rect 673366 714504 673422 714513
rect 673366 714439 673422 714448
rect 673274 712464 673330 712473
rect 673274 712399 673330 712408
rect 673288 707266 673316 712399
rect 673276 707260 673328 707266
rect 673276 707202 673328 707208
rect 673366 705120 673422 705129
rect 673366 705055 673422 705064
rect 673090 661600 673146 661609
rect 673090 661535 673146 661544
rect 672998 648680 673054 648689
rect 672998 648615 673054 648624
rect 672722 635488 672778 635497
rect 672722 635423 672778 635432
rect 672630 608696 672686 608705
rect 672630 608631 672686 608640
rect 672446 571976 672502 571985
rect 672446 571911 672502 571920
rect 672644 538214 672672 608631
rect 672814 578640 672870 578649
rect 672814 578575 672870 578584
rect 672184 538186 672304 538214
rect 672552 538186 672672 538214
rect 672184 529145 672212 538186
rect 672354 535120 672410 535129
rect 672354 535055 672410 535064
rect 672368 529258 672396 535055
rect 672552 531729 672580 538186
rect 672828 534313 672856 578575
rect 673012 573209 673040 648615
rect 673182 644056 673238 644065
rect 673182 643991 673238 644000
rect 672998 573200 673054 573209
rect 672998 573135 673054 573144
rect 673196 571169 673224 643991
rect 673380 605834 673408 705055
rect 673656 682417 673684 717586
rect 681016 710841 681044 725727
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 683132 706761 683160 726815
rect 683394 726472 683450 726481
rect 683394 726407 683450 726416
rect 683408 711249 683436 726407
rect 683578 725520 683634 725529
rect 683578 725455 683634 725464
rect 683394 711240 683450 711249
rect 683394 711175 683450 711184
rect 683592 708393 683620 725455
rect 683856 724260 683908 724266
rect 683856 724202 683908 724208
rect 683578 708384 683634 708393
rect 683578 708319 683634 708328
rect 683868 707985 683896 724202
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683854 707976 683910 707985
rect 683854 707911 683910 707920
rect 683118 706752 683174 706761
rect 683118 706687 683174 706696
rect 675114 701176 675170 701185
rect 675114 701111 675170 701120
rect 675128 698337 675156 701111
rect 675128 698309 675418 698337
rect 674024 697666 675418 697694
rect 673826 690160 673882 690169
rect 673826 690095 673882 690104
rect 673642 682408 673698 682417
rect 673642 682343 673698 682352
rect 673550 644872 673606 644881
rect 673550 644807 673606 644816
rect 673564 630674 673592 644807
rect 673840 636857 673868 690095
rect 673826 636848 673882 636857
rect 673826 636783 673882 636792
rect 673564 630646 673776 630674
rect 673288 605806 673408 605834
rect 673288 592034 673316 605806
rect 673458 599720 673514 599729
rect 673458 599655 673514 599664
rect 673472 597530 673500 599655
rect 673748 597961 673776 630646
rect 674024 619177 674052 697666
rect 675114 696960 675170 696969
rect 675114 696895 675170 696904
rect 675128 695209 675156 696895
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695181 675418 695209
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 674392 693994 675418 694022
rect 674194 666224 674250 666233
rect 674194 666159 674250 666168
rect 674208 665145 674236 666159
rect 674194 665136 674250 665145
rect 674194 665071 674250 665080
rect 674392 647170 674420 693994
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 674852 693314 675340 693342
rect 675404 693328 675432 693382
rect 674654 689616 674710 689625
rect 674654 689551 674710 689560
rect 674668 689330 674696 689551
rect 674852 689466 674880 693314
rect 675114 692880 675170 692889
rect 675114 692815 675170 692824
rect 675128 690894 675156 692815
rect 675128 690866 675418 690894
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675312 689710 675432 689738
rect 675312 689625 675340 689710
rect 675404 689656 675432 689710
rect 675298 689616 675354 689625
rect 675298 689551 675354 689560
rect 674208 647142 674420 647170
rect 674484 689302 674696 689330
rect 674760 689438 674880 689466
rect 674208 642433 674236 647142
rect 674194 642424 674250 642433
rect 674194 642359 674250 642368
rect 674194 641744 674250 641753
rect 674194 641679 674250 641688
rect 674010 619168 674066 619177
rect 674010 619103 674066 619112
rect 673918 603528 673974 603537
rect 673918 603463 673974 603472
rect 673734 597952 673790 597961
rect 673734 597887 673790 597896
rect 673932 597802 673960 603463
rect 673840 597774 673960 597802
rect 673472 597502 673684 597530
rect 673458 597408 673514 597417
rect 673458 597343 673514 597352
rect 673288 592006 673408 592034
rect 673182 571160 673238 571169
rect 673182 571095 673238 571104
rect 672998 570344 673054 570353
rect 672998 570279 673054 570288
rect 672814 534304 672870 534313
rect 672814 534239 672870 534248
rect 672814 532808 672870 532817
rect 672814 532743 672870 532752
rect 672828 532114 672856 532743
rect 672828 532086 672948 532114
rect 672722 531992 672778 532001
rect 672722 531927 672778 531936
rect 672538 531720 672594 531729
rect 672538 531655 672594 531664
rect 672368 529230 672488 529258
rect 672170 529136 672226 529145
rect 672170 529071 672226 529080
rect 671986 501664 672042 501673
rect 671986 501599 672042 501608
rect 672460 490929 672488 529230
rect 672736 495434 672764 531927
rect 672920 528554 672948 532086
rect 672644 495406 672764 495434
rect 672828 528526 672948 528554
rect 672446 490920 672502 490929
rect 672446 490855 672502 490864
rect 672446 489696 672502 489705
rect 672446 489631 672502 489640
rect 672264 455388 672316 455394
rect 672264 455330 672316 455336
rect 671804 455048 671856 455054
rect 672276 455025 672304 455330
rect 671804 454990 671856 454996
rect 672262 455016 672318 455025
rect 672262 454951 672318 454960
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 671344 430636 671396 430642
rect 671344 430578 671396 430584
rect 669962 403744 670018 403753
rect 669962 403679 670018 403688
rect 670606 393544 670662 393553
rect 670606 393479 670662 393488
rect 670422 347304 670478 347313
rect 670422 347239 670478 347248
rect 668582 311944 668638 311953
rect 668582 311879 668638 311888
rect 669226 302288 669282 302297
rect 669226 302223 669282 302232
rect 668952 236904 669004 236910
rect 668952 236846 669004 236852
rect 668676 235952 668728 235958
rect 668676 235894 668728 235900
rect 668308 234592 668360 234598
rect 668308 234534 668360 234540
rect 668124 231464 668176 231470
rect 668124 231406 668176 231412
rect 667940 225684 667992 225690
rect 667940 225626 667992 225632
rect 667952 223145 667980 225626
rect 667938 223136 667994 223145
rect 667938 223071 667994 223080
rect 667938 222048 667994 222057
rect 667938 221983 667994 221992
rect 667952 220969 667980 221983
rect 667938 220960 667994 220969
rect 667938 220895 667994 220904
rect 668136 219434 668164 231406
rect 668044 219406 668164 219434
rect 668044 202473 668072 219406
rect 668030 202464 668086 202473
rect 668030 202399 668086 202408
rect 667940 199232 667992 199238
rect 667938 199200 667940 199209
rect 667992 199200 667994 199209
rect 667938 199135 667994 199144
rect 668122 198792 668178 198801
rect 668122 198727 668178 198736
rect 667940 194336 667992 194342
rect 667938 194304 667940 194313
rect 667992 194304 667994 194313
rect 667938 194239 667994 194248
rect 667940 189440 667992 189446
rect 667938 189408 667940 189417
rect 667992 189408 667994 189417
rect 667938 189343 667994 189352
rect 668136 187649 668164 198727
rect 668122 187640 668178 187649
rect 668122 187575 668178 187584
rect 668122 184920 668178 184929
rect 668122 184855 668178 184864
rect 667754 178800 667810 178809
rect 667754 178735 667810 178744
rect 667940 174752 667992 174758
rect 667938 174720 667940 174729
rect 667992 174720 667994 174729
rect 667938 174655 667994 174664
rect 667940 169720 667992 169726
rect 667938 169688 667940 169697
rect 667992 169688 667994 169697
rect 667938 169623 667994 169632
rect 668136 168201 668164 184855
rect 668320 182889 668348 234534
rect 668490 234288 668546 234297
rect 668490 234223 668546 234232
rect 668306 182880 668362 182889
rect 668306 182815 668362 182824
rect 668122 168192 668178 168201
rect 668122 168127 668178 168136
rect 668308 150272 668360 150278
rect 668306 150240 668308 150249
rect 668360 150240 668362 150249
rect 668306 150175 668362 150184
rect 668504 148617 668532 234223
rect 668688 224954 668716 235894
rect 668964 230602 668992 236846
rect 669240 234614 669268 302223
rect 670146 264072 670202 264081
rect 670146 264007 670202 264016
rect 669962 259584 670018 259593
rect 669962 259519 670018 259528
rect 669976 245857 670004 259519
rect 669962 245848 670018 245857
rect 669962 245783 670018 245792
rect 670160 235929 670188 264007
rect 670146 235920 670202 235929
rect 670146 235855 670202 235864
rect 669148 234586 669268 234614
rect 668964 230574 669084 230602
rect 668860 230444 668912 230450
rect 668860 230386 668912 230392
rect 668688 224926 668808 224954
rect 668780 153513 668808 224926
rect 668872 205634 668900 230386
rect 669056 219434 669084 230574
rect 669148 224954 669176 234586
rect 669780 234388 669832 234394
rect 669780 234330 669832 234336
rect 669594 232792 669650 232801
rect 669594 232727 669650 232736
rect 669412 228268 669464 228274
rect 669412 228210 669464 228216
rect 669424 225729 669452 228210
rect 669410 225720 669466 225729
rect 669410 225655 669466 225664
rect 669318 225312 669374 225321
rect 669318 225247 669374 225256
rect 669332 225162 669360 225247
rect 669332 225134 669452 225162
rect 669424 225078 669452 225134
rect 669412 225072 669464 225078
rect 669412 225014 669464 225020
rect 669148 224926 669268 224954
rect 668964 219406 669084 219434
rect 668964 209774 668992 219406
rect 669240 215665 669268 224926
rect 669412 224868 669464 224874
rect 669412 224810 669464 224816
rect 669424 223689 669452 224810
rect 669410 223680 669466 223689
rect 669410 223615 669466 223624
rect 669410 216608 669466 216617
rect 669410 216543 669466 216552
rect 669226 215656 669282 215665
rect 669226 215591 669282 215600
rect 669226 214568 669282 214577
rect 669226 214503 669282 214512
rect 669240 214146 669268 214503
rect 669148 214118 669268 214146
rect 669148 209774 669176 214118
rect 668964 209746 669084 209774
rect 669148 209746 669268 209774
rect 668872 205606 668992 205634
rect 668964 192681 668992 205606
rect 669056 192794 669084 209746
rect 669240 207278 669268 209746
rect 669148 207250 669268 207278
rect 669148 202450 669176 207250
rect 669424 205634 669452 216543
rect 669608 215294 669636 232727
rect 669792 224954 669820 234330
rect 670054 233200 670110 233209
rect 670054 233135 670110 233144
rect 669792 224926 669912 224954
rect 669332 205606 669452 205634
rect 669516 215266 669636 215294
rect 669332 202609 669360 205606
rect 669318 202600 669374 202609
rect 669318 202535 669374 202544
rect 669148 202422 669268 202450
rect 669240 201657 669268 202422
rect 669226 201648 669282 201657
rect 669226 201583 669282 201592
rect 669056 192766 669176 192794
rect 668950 192672 669006 192681
rect 668950 192607 669006 192616
rect 669148 186314 669176 192766
rect 669056 186286 669176 186314
rect 669056 180794 669084 186286
rect 669228 184544 669280 184550
rect 669226 184512 669228 184521
rect 669280 184512 669282 184521
rect 669226 184447 669282 184456
rect 668964 180766 669084 180794
rect 668964 163305 668992 180766
rect 669134 167104 669190 167113
rect 669134 167039 669190 167048
rect 668950 163296 669006 163305
rect 668950 163231 669006 163240
rect 668766 153504 668822 153513
rect 668766 153439 668822 153448
rect 668766 153096 668822 153105
rect 668766 153031 668822 153040
rect 668490 148608 668546 148617
rect 668490 148543 668546 148552
rect 667938 137456 667994 137465
rect 667938 137391 667994 137400
rect 667570 135960 667626 135969
rect 667570 135895 667626 135904
rect 667952 135561 667980 137391
rect 667938 135552 667994 135561
rect 667938 135487 667994 135496
rect 666834 133104 666890 133113
rect 666834 133039 666890 133048
rect 590292 131776 590344 131782
rect 590292 131718 590344 131724
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 589646 129704 589702 129713
rect 589646 129639 589702 129648
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127226 589504 128007
rect 589464 127220 589516 127226
rect 589464 127162 589516 127168
rect 589660 124914 589688 129639
rect 590106 126440 590162 126449
rect 590106 126375 590162 126384
rect 589648 124908 589700 124914
rect 589648 124850 589700 124856
rect 589922 124808 589978 124817
rect 589922 124743 589978 124752
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 589462 119912 589518 119921
rect 589462 119847 589518 119856
rect 589476 118726 589504 119847
rect 589464 118720 589516 118726
rect 589464 118662 589516 118668
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 588728 113076 588780 113082
rect 588728 113018 588780 113024
rect 588544 111852 588596 111858
rect 588544 111794 588596 111800
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 588556 88330 588584 111794
rect 589370 111752 589426 111761
rect 589370 111687 589426 111696
rect 589384 109750 589412 111687
rect 589936 111110 589964 124743
rect 590120 122126 590148 126375
rect 668780 125769 668808 153031
rect 669148 143721 669176 167039
rect 669516 164937 669544 215266
rect 669686 214568 669742 214577
rect 669686 214503 669742 214512
rect 669700 200569 669728 214503
rect 669686 200560 669742 200569
rect 669686 200495 669742 200504
rect 669884 195974 669912 224926
rect 669792 195946 669912 195974
rect 669792 184550 669820 195946
rect 669780 184544 669832 184550
rect 669780 184486 669832 184492
rect 670068 169726 670096 233135
rect 670240 232892 670292 232898
rect 670240 232834 670292 232840
rect 670252 174758 670280 232834
rect 670436 211177 670464 347239
rect 670620 214033 670648 393479
rect 671356 275369 671384 430578
rect 672460 401713 672488 489631
rect 672644 488481 672672 495406
rect 672828 489297 672856 528526
rect 673012 500993 673040 570279
rect 673182 559056 673238 559065
rect 673182 558991 673238 559000
rect 672998 500984 673054 500993
rect 672998 500919 673054 500928
rect 672814 489288 672870 489297
rect 672814 489223 672870 489232
rect 672630 488472 672686 488481
rect 672630 488407 672686 488416
rect 672630 488064 672686 488073
rect 672630 487999 672686 488008
rect 672446 401704 672502 401713
rect 672446 401639 672502 401648
rect 672644 400081 672672 487999
rect 673196 484809 673224 558991
rect 673182 484800 673238 484809
rect 673182 484735 673238 484744
rect 673090 457056 673146 457065
rect 673090 456991 673146 457000
rect 673104 455002 673132 456991
rect 673380 456634 673408 592006
rect 673472 580530 673500 597343
rect 673656 596034 673684 597502
rect 673564 596006 673684 596034
rect 673564 589274 673592 596006
rect 673840 594130 673868 597774
rect 674010 596592 674066 596601
rect 674010 596527 674066 596536
rect 673840 594102 673960 594130
rect 673564 589246 673684 589274
rect 673656 587894 673684 589246
rect 673656 587866 673776 587894
rect 673748 582593 673776 587866
rect 673734 582584 673790 582593
rect 673734 582519 673790 582528
rect 673932 582374 673960 594102
rect 673840 582346 673960 582374
rect 673472 580502 673776 580530
rect 673550 580408 673606 580417
rect 673550 580343 673606 580352
rect 673564 553394 673592 580343
rect 673748 575474 673776 580502
rect 673472 553366 673592 553394
rect 673656 575446 673776 575474
rect 673472 538214 673500 553366
rect 673656 547097 673684 575446
rect 673642 547088 673698 547097
rect 673642 547023 673698 547032
rect 673840 545850 673868 582346
rect 674024 553394 674052 596527
rect 674208 591297 674236 641679
rect 674484 639826 674512 689302
rect 674760 685874 674788 689438
rect 674930 689344 674986 689353
rect 674930 689279 674986 689288
rect 674944 688922 674972 689279
rect 675114 689072 675170 689081
rect 675170 689030 675418 689058
rect 675114 689007 675170 689016
rect 674944 688894 675248 688922
rect 674930 688800 674986 688809
rect 674930 688735 674986 688744
rect 674944 687290 674972 688735
rect 675220 688634 675248 688894
rect 675220 688606 675340 688634
rect 674944 687262 675156 687290
rect 674930 687168 674986 687177
rect 674930 687103 674986 687112
rect 674576 685846 674788 685874
rect 674576 683114 674604 685846
rect 674944 683114 674972 687103
rect 675128 686474 675156 687262
rect 675312 686610 675340 688606
rect 675496 687449 675524 687820
rect 675482 687440 675538 687449
rect 675482 687375 675538 687384
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675128 686446 675432 686474
rect 675404 685984 675432 686446
rect 675206 685944 675262 685953
rect 675036 685902 675206 685930
rect 675036 684162 675064 685902
rect 675206 685879 675262 685888
rect 675482 685536 675538 685545
rect 675482 685471 675538 685480
rect 675496 685372 675524 685471
rect 675036 684134 675418 684162
rect 674576 683086 674696 683114
rect 674944 683086 675248 683114
rect 674300 639798 674512 639826
rect 674300 637574 674328 639798
rect 674668 637922 674696 683086
rect 675022 670168 675078 670177
rect 675022 670103 675078 670112
rect 675036 669225 675064 670103
rect 675022 669216 675078 669225
rect 675022 669151 675078 669160
rect 674838 666224 674894 666233
rect 674838 666159 674894 666168
rect 674852 665689 674880 666159
rect 674838 665680 674894 665689
rect 674838 665615 674894 665624
rect 674838 664728 674894 664737
rect 674838 664663 674894 664672
rect 674852 664193 674880 664663
rect 674838 664184 674894 664193
rect 674838 664119 674894 664128
rect 674838 663096 674894 663105
rect 674838 663031 674894 663040
rect 674852 662561 674880 663031
rect 674838 662552 674894 662561
rect 674838 662487 674894 662496
rect 674838 661872 674894 661881
rect 674838 661807 674894 661816
rect 674852 661337 674880 661807
rect 674838 661328 674894 661337
rect 674838 661263 674894 661272
rect 675220 650162 675248 683086
rect 683210 682408 683266 682417
rect 683210 682343 683266 682352
rect 676494 673160 676550 673169
rect 676494 673095 676550 673104
rect 676508 671129 676536 673095
rect 676494 671120 676550 671129
rect 676494 671055 676550 671064
rect 683224 667049 683252 682343
rect 683394 681048 683450 681057
rect 683394 680983 683450 680992
rect 683210 667040 683266 667049
rect 683210 666975 683266 666984
rect 683408 663785 683436 680983
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683394 663776 683450 663785
rect 683394 663711 683450 663720
rect 675390 654256 675446 654265
rect 675390 654191 675446 654200
rect 675404 654134 675432 654191
rect 675312 654106 675432 654134
rect 675312 653018 675340 654106
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675588 651545 675616 651848
rect 675574 651536 675630 651545
rect 675574 651471 675630 651480
rect 675220 650134 675340 650162
rect 675312 649994 675340 650134
rect 674852 649966 675340 649994
rect 674852 645854 674880 649966
rect 675404 649618 675432 650012
rect 674806 645833 674880 645854
rect 674792 645826 674880 645833
rect 674944 649590 675432 649618
rect 674944 645854 674972 649590
rect 675496 648961 675524 649468
rect 675482 648952 675538 648961
rect 675482 648887 675538 648896
rect 675496 648689 675524 648788
rect 675482 648680 675538 648689
rect 675482 648615 675538 648624
rect 675496 647873 675524 648176
rect 675482 647864 675538 647873
rect 675482 647799 675538 647808
rect 675298 647320 675354 647329
rect 675298 647255 675354 647264
rect 675312 646218 675340 647255
rect 675312 646190 675432 646218
rect 674944 645826 675064 645854
rect 674792 645824 674848 645826
rect 674792 645759 674848 645768
rect 675036 644858 675064 645826
rect 675404 645660 675432 646190
rect 675496 644881 675524 645116
rect 674852 644830 675064 644858
rect 675482 644872 675538 644881
rect 674852 643498 674880 644830
rect 675482 644807 675538 644816
rect 675772 644337 675800 644475
rect 675758 644328 675814 644337
rect 675758 644263 675814 644272
rect 675482 644056 675538 644065
rect 675482 643991 675538 644000
rect 675496 643824 675524 643991
rect 674806 643470 674880 643498
rect 675298 643512 675354 643521
rect 674806 643226 674834 643470
rect 675298 643447 675354 643456
rect 674760 643198 674834 643226
rect 674760 642546 674788 643198
rect 675312 643090 675340 643447
rect 675128 643062 675340 643090
rect 674760 642518 674972 642546
rect 674576 637894 674696 637922
rect 674576 637574 674604 637894
rect 674746 637800 674802 637809
rect 674746 637735 674802 637744
rect 674300 637546 674512 637574
rect 674576 637546 674696 637574
rect 674484 617817 674512 637546
rect 674668 619585 674696 637546
rect 674760 635882 674788 637735
rect 674944 636041 674972 642518
rect 675128 641458 675156 643062
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675206 641336 675262 641345
rect 675206 641271 675262 641280
rect 675220 640809 675248 641271
rect 675220 640781 675418 640809
rect 675128 640138 675418 640166
rect 675128 638330 675156 640138
rect 675298 639432 675354 639441
rect 675298 639367 675354 639376
rect 675128 638302 675248 638330
rect 675220 638058 675248 638302
rect 675036 638030 675248 638058
rect 675036 637574 675064 638030
rect 675312 637922 675340 639367
rect 675496 638625 675524 638928
rect 675482 638616 675538 638625
rect 675482 638551 675538 638560
rect 675574 637936 675630 637945
rect 675312 637894 675432 637922
rect 675404 637650 675432 637894
rect 675574 637871 675630 637880
rect 675312 637622 675432 637650
rect 675036 637546 675248 637574
rect 674930 636032 674986 636041
rect 674930 635967 674986 635976
rect 674760 635854 674972 635882
rect 674944 635769 674972 635854
rect 674930 635760 674986 635769
rect 674930 635695 674986 635704
rect 675220 631417 675248 637546
rect 675312 631666 675340 637622
rect 675312 631638 675432 631666
rect 674838 631408 674894 631417
rect 674838 631343 674894 631352
rect 675206 631408 675262 631417
rect 675206 631343 675262 631352
rect 674852 626534 674880 631343
rect 675404 629785 675432 631638
rect 675588 631417 675616 637871
rect 682382 637664 682438 637673
rect 682382 637599 682438 637608
rect 675574 631408 675630 631417
rect 675574 631343 675630 631352
rect 675390 629776 675446 629785
rect 675390 629711 675446 629720
rect 675206 629504 675262 629513
rect 675206 629439 675262 629448
rect 675220 626534 675248 629439
rect 676494 628552 676550 628561
rect 676494 628487 676550 628496
rect 674852 626506 675064 626534
rect 674654 619576 674710 619585
rect 674654 619511 674710 619520
rect 674470 617808 674526 617817
rect 674470 617743 674526 617752
rect 674838 608696 674894 608705
rect 674838 608631 674894 608640
rect 674852 607073 674880 608631
rect 674838 607064 674894 607073
rect 674838 606999 674894 607008
rect 674470 604616 674526 604625
rect 674470 604551 674526 604560
rect 674194 591288 674250 591297
rect 674194 591223 674250 591232
rect 674194 558376 674250 558385
rect 674194 558311 674250 558320
rect 673748 545822 673868 545850
rect 673932 553366 674052 553394
rect 673748 543734 673776 545822
rect 673932 545737 673960 553366
rect 673918 545728 673974 545737
rect 673918 545663 673974 545672
rect 673748 543706 673868 543734
rect 673472 538186 673592 538214
rect 673564 526969 673592 538186
rect 673840 528329 673868 543706
rect 674010 535392 674066 535401
rect 674010 535327 674066 535336
rect 674024 534041 674052 535327
rect 674010 534032 674066 534041
rect 674010 533967 674066 533976
rect 674010 533488 674066 533497
rect 674010 533423 674066 533432
rect 673826 528320 673882 528329
rect 673826 528255 673882 528264
rect 673550 526960 673606 526969
rect 673550 526895 673606 526904
rect 674024 490113 674052 533423
rect 674010 490104 674066 490113
rect 674010 490039 674066 490048
rect 674208 484401 674236 558311
rect 674484 538214 674512 604551
rect 675036 600114 675064 626506
rect 674668 600086 675064 600114
rect 675128 626506 675248 626534
rect 674668 598934 674696 600086
rect 675128 599434 675156 626506
rect 676508 625705 676536 628487
rect 676494 625696 676550 625705
rect 676494 625631 676550 625640
rect 682396 622033 682424 637599
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 683210 635488 683266 635497
rect 683210 635423 683266 635432
rect 683224 622849 683252 635423
rect 683210 622840 683266 622849
rect 683210 622775 683266 622784
rect 682382 622024 682438 622033
rect 682382 621959 682438 621968
rect 676494 621616 676550 621625
rect 676494 621551 676550 621560
rect 676508 621217 676536 621551
rect 676494 621208 676550 621217
rect 676494 621143 676550 621152
rect 676494 620392 676550 620401
rect 676494 620327 676550 620336
rect 676508 619993 676536 620327
rect 676494 619984 676550 619993
rect 676494 619919 676550 619928
rect 677230 619576 677286 619585
rect 677230 619511 677286 619520
rect 677244 619177 677272 619511
rect 677230 619168 677286 619177
rect 677230 619103 677286 619112
rect 683118 619168 683174 619177
rect 683118 619103 683174 619112
rect 683132 617545 683160 619103
rect 683118 617536 683174 617545
rect 683118 617471 683174 617480
rect 683408 617137 683436 636783
rect 683762 635760 683818 635769
rect 683762 635695 683818 635704
rect 683776 618769 683804 635695
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683762 618760 683818 618769
rect 683762 618695 683818 618704
rect 683394 617128 683450 617137
rect 683394 617063 683450 617072
rect 675496 607889 675524 608124
rect 675482 607880 675538 607889
rect 675482 607815 675538 607824
rect 675312 607465 675418 607493
rect 675312 607345 675340 607465
rect 675298 607336 675354 607345
rect 675298 607271 675354 607280
rect 675298 607064 675354 607073
rect 675298 606999 675354 607008
rect 675312 606846 675340 606999
rect 675312 606818 675418 606846
rect 675312 604982 675418 605010
rect 675312 604625 675340 604982
rect 675298 604616 675354 604625
rect 675298 604551 675354 604560
rect 675312 604438 675418 604466
rect 675312 604353 675340 604438
rect 675298 604344 675354 604353
rect 675298 604279 675354 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675312 603146 675418 603174
rect 675312 602993 675340 603146
rect 675298 602984 675354 602993
rect 675298 602919 675354 602928
rect 675496 600409 675524 600644
rect 675482 600400 675538 600409
rect 675482 600335 675538 600344
rect 675312 600222 675432 600250
rect 675312 599729 675340 600222
rect 675404 600100 675432 600222
rect 675298 599720 675354 599729
rect 675298 599655 675354 599664
rect 674576 598906 674696 598934
rect 675036 599406 675156 599434
rect 675220 599474 675418 599502
rect 674576 596306 674604 598906
rect 675036 597554 675064 599406
rect 675220 599321 675248 599474
rect 675206 599312 675262 599321
rect 675206 599247 675262 599256
rect 675312 598862 675432 598890
rect 675312 598822 675340 598862
rect 674944 597526 675064 597554
rect 675220 598794 675340 598822
rect 675404 598808 675432 598862
rect 674576 596278 674788 596306
rect 674760 592385 674788 596278
rect 674746 592376 674802 592385
rect 674746 592311 674802 592320
rect 674944 589274 674972 597526
rect 675220 596601 675248 598794
rect 675404 597417 675432 597652
rect 675390 597408 675446 597417
rect 675390 597343 675446 597352
rect 675390 596864 675446 596873
rect 675390 596799 675446 596808
rect 675206 596592 675262 596601
rect 675206 596527 675262 596536
rect 675404 596428 675432 596799
rect 675404 595354 675432 595816
rect 675312 595326 675432 595354
rect 675312 589274 675340 595326
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675496 593609 675524 593980
rect 675482 593600 675538 593609
rect 675482 593535 675538 593544
rect 675574 593192 675630 593201
rect 675574 593127 675630 593136
rect 674944 589246 675156 589274
rect 675312 589246 675432 589274
rect 675128 581641 675156 589246
rect 675114 581632 675170 581641
rect 675114 581567 675170 581576
rect 675404 581482 675432 589246
rect 675588 586265 675616 593127
rect 676034 592920 676090 592929
rect 676034 592855 676090 592864
rect 675850 592376 675906 592385
rect 675850 592311 675906 592320
rect 675864 591394 675892 592311
rect 675852 591388 675904 591394
rect 675852 591330 675904 591336
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 675850 581632 675906 581641
rect 675850 581567 675906 581576
rect 675220 581454 675432 581482
rect 675022 580816 675078 580825
rect 675022 580751 675078 580760
rect 675036 579873 675064 580751
rect 675022 579864 675078 579873
rect 675022 579799 675078 579808
rect 675022 577688 675078 577697
rect 675022 577623 675078 577632
rect 675036 576881 675064 577623
rect 675022 576872 675078 576881
rect 675022 576807 675078 576816
rect 674838 559464 674894 559473
rect 674838 559399 674894 559408
rect 674654 548312 674710 548321
rect 674654 548247 674710 548256
rect 674668 543734 674696 548247
rect 674852 546281 674880 559399
rect 675220 550633 675248 581454
rect 675482 578368 675538 578377
rect 675482 578303 675538 578312
rect 675496 577017 675524 578303
rect 675482 577008 675538 577017
rect 675482 576943 675538 576952
rect 675864 575385 675892 581567
rect 676048 576609 676076 592855
rect 683118 592648 683174 592657
rect 683118 592583 683174 592592
rect 682384 591388 682436 591394
rect 682384 591330 682436 591336
rect 676034 576600 676090 576609
rect 676034 576535 676090 576544
rect 675850 575376 675906 575385
rect 675850 575311 675906 575320
rect 682396 570761 682424 591330
rect 683132 571985 683160 592583
rect 683394 591288 683450 591297
rect 683394 591223 683450 591232
rect 683408 573209 683436 591223
rect 683670 589928 683726 589937
rect 683670 589863 683726 589872
rect 683684 574025 683712 589863
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683670 574016 683726 574025
rect 683670 573951 683726 573960
rect 683394 573200 683450 573209
rect 683394 573135 683450 573144
rect 683118 571976 683174 571985
rect 683118 571911 683174 571920
rect 682382 570752 682438 570761
rect 682382 570687 682438 570696
rect 675390 564496 675446 564505
rect 675390 564431 675446 564440
rect 675404 564346 675432 564431
rect 675312 564318 675432 564346
rect 675312 562306 675340 564318
rect 675588 562737 675616 562904
rect 675574 562728 675630 562737
rect 675574 562663 675630 562672
rect 675312 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675496 559473 675524 559776
rect 675482 559464 675538 559473
rect 675482 559399 675538 559408
rect 675404 559065 675432 559232
rect 675390 559056 675446 559065
rect 675390 558991 675446 559000
rect 675404 558385 675432 558620
rect 675390 558376 675446 558385
rect 675390 558311 675446 558320
rect 675772 557569 675800 557940
rect 675482 557560 675538 557569
rect 675312 557518 675482 557546
rect 675312 555370 675340 557518
rect 675482 557495 675538 557504
rect 675758 557560 675814 557569
rect 675758 557495 675814 557504
rect 675404 555370 675432 555492
rect 675312 555342 675432 555370
rect 675404 554713 675432 554919
rect 675390 554704 675446 554713
rect 675390 554639 675446 554648
rect 675772 553897 675800 554268
rect 675758 553888 675814 553897
rect 675758 553823 675814 553832
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 675390 551576 675446 551585
rect 675390 551511 675446 551520
rect 675404 551239 675432 551511
rect 675206 550624 675262 550633
rect 675206 550559 675262 550568
rect 675772 550361 675800 550596
rect 675758 550352 675814 550361
rect 675758 550287 675814 550296
rect 675128 549937 675418 549965
rect 675128 547754 675156 549937
rect 675404 548321 675432 548760
rect 675390 548312 675446 548321
rect 675390 548247 675446 548256
rect 675036 547726 675156 547754
rect 674838 546272 674894 546281
rect 674838 546207 674894 546216
rect 674838 546000 674894 546009
rect 674838 545935 674894 545944
rect 674668 543706 674788 543734
rect 674392 538186 674512 538214
rect 674392 530641 674420 538186
rect 674562 532264 674618 532273
rect 674562 532199 674618 532208
rect 674576 531457 674604 532199
rect 674562 531448 674618 531457
rect 674562 531383 674618 531392
rect 674378 530632 674434 530641
rect 674378 530567 674434 530576
rect 674562 529408 674618 529417
rect 674562 529343 674618 529352
rect 674576 528601 674604 529343
rect 674562 528592 674618 528601
rect 674562 528527 674618 528536
rect 674760 485625 674788 543706
rect 674852 540974 674880 545935
rect 674852 540946 674972 540974
rect 674944 511994 674972 540946
rect 674852 511966 674972 511994
rect 674852 503282 674880 511966
rect 675036 510241 675064 547726
rect 675944 547664 675996 547670
rect 675942 547632 675944 547641
rect 678244 547664 678296 547670
rect 675996 547632 675998 547641
rect 675942 547567 675998 547576
rect 677414 547632 677470 547641
rect 678244 547606 678296 547612
rect 677414 547567 677470 547576
rect 675390 546272 675446 546281
rect 675390 546207 675446 546216
rect 675206 545456 675262 545465
rect 675206 545391 675262 545400
rect 675220 540974 675248 545391
rect 675404 540974 675432 546207
rect 675128 540946 675248 540974
rect 675312 540946 675432 540974
rect 675128 510354 675156 540946
rect 675312 511994 675340 540946
rect 676494 538792 676550 538801
rect 676494 538727 676550 538736
rect 676508 535945 676536 538727
rect 676494 535936 676550 535945
rect 676494 535871 676550 535880
rect 675758 535120 675814 535129
rect 675758 535055 675814 535064
rect 675772 534517 675800 535055
rect 675758 534508 675814 534517
rect 675758 534443 675814 534452
rect 676864 520328 676916 520334
rect 676864 520270 676916 520276
rect 676036 518832 676088 518838
rect 676036 518774 676088 518780
rect 675312 511966 675616 511994
rect 675128 510326 675432 510354
rect 675022 510232 675078 510241
rect 675022 510167 675078 510176
rect 675206 503704 675262 503713
rect 675206 503639 675262 503648
rect 675220 503282 675248 503639
rect 674852 503254 675248 503282
rect 675404 503169 675432 510326
rect 675022 503160 675078 503169
rect 675022 503095 675078 503104
rect 675390 503160 675446 503169
rect 675390 503095 675446 503104
rect 675036 502334 675064 503095
rect 675588 502334 675616 511966
rect 675850 510232 675906 510241
rect 675036 502306 675156 502334
rect 675128 487665 675156 502306
rect 675312 502306 675616 502334
rect 675680 510190 675850 510218
rect 675680 502334 675708 510190
rect 675850 510167 675906 510176
rect 675850 503704 675906 503713
rect 675850 503639 675852 503648
rect 675904 503639 675906 503648
rect 675852 503610 675904 503616
rect 675680 502306 675892 502334
rect 675312 499574 675340 502306
rect 675666 500984 675722 500993
rect 675864 500954 675892 502306
rect 675666 500919 675722 500928
rect 675852 500948 675904 500954
rect 675220 499546 675340 499574
rect 675680 499574 675708 500919
rect 675852 500890 675904 500896
rect 675680 499546 675984 499574
rect 675220 495434 675248 499546
rect 675220 495406 675340 495434
rect 675114 487656 675170 487665
rect 675114 487591 675170 487600
rect 675312 486441 675340 495406
rect 675574 490512 675630 490521
rect 675574 490447 675630 490456
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 674746 485616 674802 485625
rect 674746 485551 674802 485560
rect 674194 484392 674250 484401
rect 674194 484327 674250 484336
rect 675588 480254 675616 490447
rect 675758 481944 675814 481953
rect 675758 481879 675814 481888
rect 674944 480226 675616 480254
rect 673380 456618 673500 456634
rect 673380 456612 673512 456618
rect 673380 456606 673460 456612
rect 673460 456554 673512 456560
rect 673826 456104 673882 456113
rect 673826 456039 673828 456048
rect 673880 456039 673882 456048
rect 673828 456010 673880 456016
rect 673734 455832 673790 455841
rect 673734 455767 673736 455776
rect 673788 455767 673790 455776
rect 673736 455738 673788 455744
rect 673598 455592 673650 455598
rect 673596 455560 673598 455569
rect 673650 455560 673652 455569
rect 673596 455495 673652 455504
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673388 455194 673440 455200
rect 673058 454974 673132 455002
rect 673058 454918 673086 454974
rect 673046 454912 673098 454918
rect 672906 454880 672962 454889
rect 673046 454854 673098 454860
rect 672906 454815 672962 454824
rect 672920 454714 672948 454815
rect 672908 454708 672960 454714
rect 672908 454650 672960 454656
rect 673164 454640 673216 454646
rect 673162 454608 673164 454617
rect 673216 454608 673218 454617
rect 673162 454543 673218 454552
rect 672816 454232 672868 454238
rect 672814 454200 672816 454209
rect 672868 454200 672870 454209
rect 672814 454135 672870 454144
rect 674944 453937 674972 480226
rect 675482 480040 675538 480049
rect 675482 479975 675538 479984
rect 675496 466454 675524 479975
rect 675772 466454 675800 481879
rect 675496 466426 675616 466454
rect 675588 454209 675616 466426
rect 675680 466426 675800 466454
rect 675680 454322 675708 466426
rect 675956 455682 675984 499546
rect 676048 480254 676076 518774
rect 676048 480226 676168 480254
rect 676140 457065 676168 480226
rect 676402 474872 676458 474881
rect 676402 474807 676458 474816
rect 676126 457056 676182 457065
rect 676126 456991 676182 457000
rect 676416 456113 676444 474807
rect 676402 456104 676458 456113
rect 676402 456039 676458 456048
rect 675956 455654 676076 455682
rect 675852 455592 675904 455598
rect 675850 455560 675852 455569
rect 675904 455560 675906 455569
rect 675850 455495 675906 455504
rect 676048 454617 676076 455654
rect 676876 454889 676904 520270
rect 677046 501664 677102 501673
rect 677046 501599 677102 501608
rect 677060 455598 677088 501599
rect 677428 489938 677456 547567
rect 678256 531457 678284 547606
rect 683210 547088 683266 547097
rect 683210 547023 683266 547032
rect 682382 546816 682438 546825
rect 682382 546751 682438 546760
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 682396 531049 682424 546751
rect 682382 531040 682438 531049
rect 682382 530975 682438 530984
rect 683224 528193 683252 547023
rect 683394 545728 683450 545737
rect 683394 545663 683450 545672
rect 683210 528184 683266 528193
rect 683210 528119 683266 528128
rect 683408 526561 683436 545663
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683578 533896 683634 533905
rect 683578 533831 683634 533840
rect 683592 527377 683620 533831
rect 683578 527368 683634 527377
rect 683578 527303 683634 527312
rect 683394 526552 683450 526561
rect 683394 526487 683450 526496
rect 683118 525736 683174 525745
rect 683118 525671 683174 525680
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 677888 518838 677916 524447
rect 683132 520334 683160 525671
rect 683120 520328 683172 520334
rect 683120 520270 683172 520276
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683578 503704 683634 503713
rect 679624 503668 679676 503674
rect 683578 503639 683634 503648
rect 679624 503610 679676 503616
rect 677416 489932 677468 489938
rect 677416 489874 677468 489880
rect 679636 486849 679664 503610
rect 683394 503432 683450 503441
rect 683394 503367 683450 503376
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 679622 486840 679678 486849
rect 679622 486775 679678 486784
rect 681016 481545 681044 500890
rect 683118 494728 683174 494737
rect 683118 494663 683174 494672
rect 683132 491337 683160 494663
rect 683118 491328 683174 491337
rect 683118 491263 683174 491272
rect 683120 489932 683172 489938
rect 683120 489874 683172 489880
rect 683132 483177 683160 489874
rect 683408 483585 683436 503367
rect 683592 487257 683620 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 487248 683634 487257
rect 683578 487183 683634 487192
rect 683394 483576 683450 483585
rect 683394 483511 683450 483520
rect 683118 483168 683174 483177
rect 683118 483103 683174 483112
rect 681002 481536 681058 481545
rect 681002 481471 681058 481480
rect 677048 455592 677100 455598
rect 677048 455534 677100 455540
rect 676862 454880 676918 454889
rect 676862 454815 676918 454824
rect 676034 454608 676090 454617
rect 676034 454543 676090 454552
rect 675680 454294 675800 454322
rect 675574 454200 675630 454209
rect 675574 454135 675630 454144
rect 674746 453928 674802 453937
rect 674746 453863 674802 453872
rect 674930 453928 674986 453937
rect 674930 453863 674986 453872
rect 674760 453778 674788 453863
rect 675772 453778 675800 454294
rect 674760 453750 675800 453778
rect 683302 411904 683358 411913
rect 683302 411839 683358 411848
rect 676034 410544 676090 410553
rect 676034 410479 676090 410488
rect 676048 402665 676076 410479
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 683132 403345 683160 406263
rect 683316 403753 683344 411839
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683302 403744 683358 403753
rect 683302 403679 683358 403688
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 676034 402656 676090 402665
rect 676034 402591 676090 402600
rect 674654 402248 674710 402257
rect 674654 402183 674710 402192
rect 674194 401432 674250 401441
rect 674194 401367 674250 401376
rect 673274 400480 673330 400489
rect 673274 400415 673330 400424
rect 672630 400072 672686 400081
rect 672630 400007 672686 400016
rect 672538 398848 672594 398857
rect 672538 398783 672594 398792
rect 672170 392320 672226 392329
rect 672170 392255 672226 392264
rect 671986 348936 672042 348945
rect 671986 348871 672042 348880
rect 672000 329769 672028 348871
rect 671986 329760 672042 329769
rect 671986 329695 672042 329704
rect 671342 275360 671398 275369
rect 671342 275295 671398 275304
rect 671710 262032 671766 262041
rect 671710 261967 671766 261976
rect 671526 259176 671582 259185
rect 671526 259111 671582 259120
rect 671342 257952 671398 257961
rect 671342 257887 671398 257896
rect 671356 241505 671384 257887
rect 671540 242865 671568 259111
rect 671724 245041 671752 261967
rect 671986 256728 672042 256737
rect 671986 256663 672042 256672
rect 671710 245032 671766 245041
rect 671710 244967 671766 244976
rect 671526 242856 671582 242865
rect 671526 242791 671582 242800
rect 671342 241496 671398 241505
rect 671342 241431 671398 241440
rect 672000 238105 672028 256663
rect 672184 253934 672212 392255
rect 672552 355065 672580 398783
rect 672722 397216 672778 397225
rect 672722 397151 672778 397160
rect 672736 377913 672764 397151
rect 673090 394224 673146 394233
rect 673090 394159 673146 394168
rect 672906 393952 672962 393961
rect 672906 393887 672962 393896
rect 672722 377904 672778 377913
rect 672722 377839 672778 377848
rect 672920 376961 672948 393887
rect 672906 376952 672962 376961
rect 672906 376887 672962 376896
rect 673104 376281 673132 394159
rect 673090 376272 673146 376281
rect 673090 376207 673146 376216
rect 672722 357096 672778 357105
rect 672722 357031 672778 357040
rect 672538 355056 672594 355065
rect 672538 354991 672594 355000
rect 672538 352200 672594 352209
rect 672538 352135 672594 352144
rect 672354 349752 672410 349761
rect 672354 349687 672410 349696
rect 672368 335617 672396 349687
rect 672552 335889 672580 352135
rect 672538 335880 672594 335889
rect 672538 335815 672594 335824
rect 672354 335608 672410 335617
rect 672354 335543 672410 335552
rect 672736 312497 672764 357031
rect 673288 355881 673316 400415
rect 674010 396128 674066 396137
rect 674010 396063 674066 396072
rect 673826 395720 673882 395729
rect 673826 395655 673882 395664
rect 673458 378176 673514 378185
rect 673458 378111 673514 378120
rect 673274 355872 673330 355881
rect 673274 355807 673330 355816
rect 673274 355464 673330 355473
rect 673274 355399 673330 355408
rect 673090 354648 673146 354657
rect 673090 354583 673146 354592
rect 672906 352608 672962 352617
rect 672906 352543 672962 352552
rect 672920 333985 672948 352543
rect 672906 333976 672962 333985
rect 672906 333911 672962 333920
rect 672906 312760 672962 312769
rect 672906 312695 672962 312704
rect 672722 312488 672778 312497
rect 672722 312423 672778 312432
rect 672446 304736 672502 304745
rect 672446 304671 672502 304680
rect 672460 290193 672488 304671
rect 672630 304328 672686 304337
rect 672630 304263 672686 304272
rect 672446 290184 672502 290193
rect 672446 290119 672502 290128
rect 672644 287881 672672 304263
rect 672920 292574 672948 312695
rect 673104 310049 673132 354583
rect 673288 310865 673316 355399
rect 673274 310856 673330 310865
rect 673274 310791 673330 310800
rect 673090 310040 673146 310049
rect 673090 309975 673146 309984
rect 673090 309632 673146 309641
rect 673090 309567 673146 309576
rect 672828 292546 672948 292574
rect 672630 287872 672686 287881
rect 672630 287807 672686 287816
rect 672828 267345 672856 292546
rect 672814 267336 672870 267345
rect 672814 267271 672870 267280
rect 672538 265704 672594 265713
rect 672538 265639 672594 265648
rect 672184 253906 672304 253934
rect 671986 238096 672042 238105
rect 671986 238031 672042 238040
rect 671712 237856 671764 237862
rect 671712 237798 671764 237804
rect 671528 237312 671580 237318
rect 671528 237254 671580 237260
rect 671344 236088 671396 236094
rect 671344 236030 671396 236036
rect 671160 235816 671212 235822
rect 671160 235758 671212 235764
rect 670790 233608 670846 233617
rect 670790 233543 670846 233552
rect 670804 231854 670832 233543
rect 670976 233368 671028 233374
rect 670976 233310 671028 233316
rect 670712 231826 670832 231854
rect 670712 224346 670740 231826
rect 670988 225457 671016 233310
rect 671172 233209 671200 235758
rect 671158 233200 671214 233209
rect 671158 233135 671214 233144
rect 671160 233028 671212 233034
rect 671160 232970 671212 232976
rect 670974 225448 671030 225457
rect 670974 225383 671030 225392
rect 670974 224768 671030 224777
rect 670974 224703 670976 224712
rect 671028 224703 671030 224712
rect 670976 224674 671028 224680
rect 670712 224318 671108 224346
rect 670928 224224 670984 224233
rect 670928 224159 670930 224168
rect 670982 224159 670984 224168
rect 670930 224130 670982 224136
rect 670790 223952 670846 223961
rect 670790 223887 670846 223896
rect 670606 214024 670662 214033
rect 670606 213959 670662 213968
rect 670606 211440 670662 211449
rect 670606 211375 670662 211384
rect 670422 211168 670478 211177
rect 670422 211103 670478 211112
rect 670620 190369 670648 211375
rect 670804 199238 670832 223887
rect 671080 215294 671108 224318
rect 670988 215266 671108 215294
rect 670792 199232 670844 199238
rect 670792 199174 670844 199180
rect 670988 194426 671016 215266
rect 670804 194398 671016 194426
rect 670804 194342 670832 194398
rect 670792 194336 670844 194342
rect 670792 194278 670844 194284
rect 671172 190454 671200 232970
rect 671356 227066 671384 236030
rect 671540 230081 671568 237254
rect 671724 234297 671752 237798
rect 671896 237652 671948 237658
rect 671896 237594 671948 237600
rect 671908 234954 671936 237594
rect 672080 237448 672132 237454
rect 672080 237390 672132 237396
rect 672092 235958 672120 237390
rect 672080 235952 672132 235958
rect 672080 235894 672132 235900
rect 671908 234926 672120 234954
rect 671894 234832 671950 234841
rect 671894 234767 671950 234776
rect 671908 234410 671936 234767
rect 672092 234569 672120 234926
rect 672078 234560 672134 234569
rect 672078 234495 672134 234504
rect 671908 234382 672120 234410
rect 671710 234288 671766 234297
rect 671710 234223 671766 234232
rect 671712 233232 671764 233238
rect 671712 233174 671764 233180
rect 671526 230072 671582 230081
rect 671526 230007 671582 230016
rect 671356 227038 671568 227066
rect 671344 226976 671396 226982
rect 671344 226918 671396 226924
rect 671356 222194 671384 226918
rect 671540 225434 671568 227038
rect 671724 226982 671752 233174
rect 671896 227248 671948 227254
rect 671896 227190 671948 227196
rect 671712 226976 671764 226982
rect 671908 226953 671936 227190
rect 671712 226918 671764 226924
rect 671894 226944 671950 226953
rect 672092 226930 672120 234382
rect 672276 231577 672304 253906
rect 672552 244274 672580 265639
rect 673104 265033 673132 309567
rect 673274 303512 673330 303521
rect 673274 303447 673330 303456
rect 673090 265024 673146 265033
rect 673090 264959 673146 264968
rect 672906 263800 672962 263809
rect 672906 263735 672962 263744
rect 672920 258074 672948 263735
rect 673090 260400 673146 260409
rect 673090 260335 673146 260344
rect 673104 258074 673132 260335
rect 672920 258046 673040 258074
rect 673104 258046 673224 258074
rect 672722 257136 672778 257145
rect 672722 257071 672778 257080
rect 672736 244274 672764 257071
rect 673012 244274 673040 258046
rect 673196 245313 673224 258046
rect 673288 245426 673316 303447
rect 673472 246265 673500 378111
rect 673840 375465 673868 395655
rect 674024 381449 674052 396063
rect 674010 381440 674066 381449
rect 674010 381375 674066 381384
rect 673826 375456 673882 375465
rect 673826 375391 673882 375400
rect 674208 356697 674236 401367
rect 674378 396536 674434 396545
rect 674378 396471 674434 396480
rect 674392 382265 674420 396471
rect 674378 382256 674434 382265
rect 674378 382191 674434 382200
rect 674668 357513 674696 402183
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 674838 394496 674894 394505
rect 674838 394431 674894 394440
rect 674852 393961 674880 394431
rect 674838 393952 674894 393961
rect 674838 393887 674894 393896
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 683026 392728 683082 392737
rect 683026 392663 683082 392672
rect 683040 389065 683068 392663
rect 683026 389056 683082 389065
rect 683026 388991 683082 389000
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675114 378040 675170 378049
rect 675114 377975 675170 377984
rect 675128 373994 675156 377975
rect 675404 377210 675432 377740
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675312 377182 675432 377210
rect 675312 376961 675340 377182
rect 675772 377060 675800 377295
rect 675298 376952 675354 376961
rect 675298 376887 675354 376896
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675298 375456 675354 375465
rect 675298 375391 675354 375400
rect 675312 375238 675340 375391
rect 675312 375210 675418 375238
rect 675128 373966 675340 373994
rect 675312 373402 675340 373966
rect 675312 373374 675418 373402
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372776 675708 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 357504 674710 357513
rect 674654 357439 674710 357448
rect 674194 356688 674250 356697
rect 674194 356623 674250 356632
rect 674194 356280 674250 356289
rect 674194 356215 674250 356224
rect 673642 353424 673698 353433
rect 673642 353359 673698 353368
rect 673656 340785 673684 353359
rect 673826 350568 673882 350577
rect 673826 350503 673882 350512
rect 673642 340776 673698 340785
rect 673642 340711 673698 340720
rect 673840 331129 673868 350503
rect 674010 349480 674066 349489
rect 674010 349415 674066 349424
rect 674024 332761 674052 349415
rect 674010 332752 674066 332761
rect 674010 332687 674066 332696
rect 673826 331120 673882 331129
rect 673826 331055 673882 331064
rect 674208 311681 674236 356215
rect 675850 351792 675906 351801
rect 675850 351727 675906 351736
rect 674746 351384 674802 351393
rect 674746 351319 674802 351328
rect 674562 347712 674618 347721
rect 674562 347647 674618 347656
rect 674576 327570 674604 347647
rect 674760 336857 674788 351319
rect 675864 350305 675892 351727
rect 675850 350296 675906 350305
rect 675850 350231 675906 350240
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 346633 676076 350095
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675666 339416 675722 339425
rect 675666 339351 675722 339360
rect 675680 339252 675708 339351
rect 675404 337249 675432 337416
rect 675390 337240 675446 337249
rect 675390 337175 675446 337184
rect 674760 336829 675418 336857
rect 675758 336560 675814 336569
rect 675758 336495 675814 336504
rect 675772 336192 675800 336495
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675758 332344 675814 332353
rect 675758 332279 675814 332288
rect 675772 331875 675800 332279
rect 675128 331214 675418 331242
rect 675128 329769 675156 331214
rect 675298 331120 675354 331129
rect 675298 331055 675354 331064
rect 675312 330049 675340 331055
rect 675312 330021 675418 330049
rect 675114 329760 675170 329769
rect 675114 329695 675170 329704
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 674576 327542 675418 327570
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 313032 674710 313041
rect 674654 312967 674710 312976
rect 674668 311953 674696 312967
rect 674838 312760 674894 312769
rect 674838 312695 674894 312704
rect 674852 312089 674880 312695
rect 674838 312080 674894 312089
rect 674838 312015 674894 312024
rect 674654 311944 674710 311953
rect 674654 311879 674710 311888
rect 674194 311672 674250 311681
rect 674194 311607 674250 311616
rect 674654 311264 674710 311273
rect 674654 311199 674710 311208
rect 674286 310448 674342 310457
rect 674286 310383 674342 310392
rect 674102 305552 674158 305561
rect 674102 305487 674158 305496
rect 674116 285569 674144 305487
rect 674102 285560 674158 285569
rect 674102 285495 674158 285504
rect 674010 267064 674066 267073
rect 674010 266999 674066 267008
rect 673826 260944 673882 260953
rect 673826 260879 673882 260888
rect 673642 258496 673698 258505
rect 673642 258431 673698 258440
rect 673458 246256 673514 246265
rect 673458 246191 673514 246200
rect 673288 245398 673408 245426
rect 673182 245304 673238 245313
rect 673182 245239 673238 245248
rect 672368 244246 672580 244274
rect 672644 244246 672764 244274
rect 672920 244246 673040 244274
rect 672368 234054 672396 244246
rect 672644 239442 672672 244246
rect 672460 239414 672672 239442
rect 672460 234138 672488 239414
rect 672722 237416 672778 237425
rect 672722 237351 672778 237360
rect 672736 237182 672764 237351
rect 672724 237176 672776 237182
rect 672724 237118 672776 237124
rect 672630 236464 672686 236473
rect 672630 236399 672686 236408
rect 672460 234110 672580 234138
rect 672368 234048 672432 234054
rect 672368 233996 672380 234048
rect 672368 233990 672432 233996
rect 672368 233974 672420 233990
rect 672262 231568 672318 231577
rect 672262 231503 672318 231512
rect 672356 228064 672408 228070
rect 672356 228006 672408 228012
rect 672368 227089 672396 228006
rect 672354 227080 672410 227089
rect 672354 227015 672410 227024
rect 672092 226902 672304 226930
rect 671894 226879 671950 226888
rect 671712 226840 671764 226846
rect 671712 226782 671764 226788
rect 672080 226840 672132 226846
rect 672080 226782 672132 226788
rect 671724 225865 671752 226782
rect 671818 226672 671874 226681
rect 671816 226616 671818 226658
rect 671816 226607 671874 226616
rect 671942 226636 671994 226642
rect 671816 226522 671844 226607
rect 671942 226578 671994 226584
rect 671816 226506 671860 226522
rect 671816 226500 671872 226506
rect 671816 226494 671820 226500
rect 671820 226442 671872 226448
rect 671954 226409 671982 226578
rect 671940 226400 671996 226409
rect 671940 226335 671996 226344
rect 672092 226250 672120 226782
rect 672092 226222 672212 226250
rect 672034 226160 672086 226166
rect 672032 226128 672034 226137
rect 672086 226128 672088 226137
rect 672032 226063 672088 226072
rect 671942 225956 671994 225962
rect 671942 225898 671994 225904
rect 671710 225856 671766 225865
rect 671710 225791 671766 225800
rect 671820 225752 671872 225758
rect 671818 225720 671820 225729
rect 671872 225720 671874 225729
rect 671818 225655 671874 225664
rect 671954 225570 671982 225898
rect 671954 225542 672028 225570
rect 672000 225457 672028 225542
rect 671986 225448 672042 225457
rect 671540 225406 671844 225434
rect 671596 225344 671648 225350
rect 671596 225286 671648 225292
rect 671608 225185 671636 225286
rect 671594 225176 671650 225185
rect 671482 225140 671534 225146
rect 671594 225111 671650 225120
rect 671482 225082 671534 225088
rect 671494 224954 671522 225082
rect 671264 222166 671384 222194
rect 671448 224926 671522 224954
rect 671264 215294 671292 222166
rect 671448 221513 671476 224926
rect 671618 224088 671674 224097
rect 671618 224023 671674 224032
rect 671434 221504 671490 221513
rect 671434 221439 671490 221448
rect 671632 215294 671660 224023
rect 671816 221354 671844 225406
rect 671986 225383 672042 225392
rect 671986 225176 672042 225185
rect 672184 225162 672212 226222
rect 672042 225134 672212 225162
rect 671986 225111 672042 225120
rect 672078 224768 672134 224777
rect 672078 224703 672134 224712
rect 671264 215266 671384 215294
rect 670804 190426 671200 190454
rect 670606 190360 670662 190369
rect 670606 190295 670662 190304
rect 670804 189446 670832 190426
rect 670792 189440 670844 189446
rect 670792 189382 670844 189388
rect 670240 174752 670292 174758
rect 670240 174694 670292 174700
rect 670606 172000 670662 172009
rect 670606 171935 670662 171944
rect 670056 169720 670108 169726
rect 670056 169662 670108 169668
rect 669778 169552 669834 169561
rect 669778 169487 669834 169496
rect 669502 164928 669558 164937
rect 669502 164863 669558 164872
rect 669792 154873 669820 169487
rect 670146 168328 670202 168337
rect 670146 168263 670202 168272
rect 669778 154864 669834 154873
rect 669778 154799 669834 154808
rect 669134 143712 669190 143721
rect 669134 143647 669190 143656
rect 669042 142216 669098 142225
rect 669042 142151 669098 142160
rect 669056 138825 669084 142151
rect 669042 138816 669098 138825
rect 669042 138751 669098 138760
rect 668950 128208 669006 128217
rect 668950 128143 669006 128152
rect 668766 125760 668822 125769
rect 668766 125695 668822 125704
rect 590108 122120 590160 122126
rect 590108 122062 590160 122068
rect 668964 120873 668992 128143
rect 669226 122224 669282 122233
rect 669226 122159 669282 122168
rect 668950 120864 669006 120873
rect 668950 120799 669006 120808
rect 668582 120592 668638 120601
rect 668582 120527 668638 120536
rect 667940 120148 667992 120154
rect 667940 120090 667992 120096
rect 667952 119241 667980 120090
rect 667938 119232 667994 119241
rect 667938 119167 667994 119176
rect 668032 118584 668084 118590
rect 668032 118526 668084 118532
rect 668044 117609 668072 118526
rect 668030 117600 668086 117609
rect 668030 117535 668086 117544
rect 590382 115016 590438 115025
rect 590382 114951 590438 114960
rect 590396 111858 590424 114951
rect 590384 111852 590436 111858
rect 590384 111794 590436 111800
rect 589924 111104 589976 111110
rect 668596 111081 668624 120527
rect 669240 114345 669268 122159
rect 670160 120154 670188 168263
rect 670330 165608 670386 165617
rect 670330 165543 670386 165552
rect 670148 120148 670200 120154
rect 670148 120090 670200 120096
rect 670344 118590 670372 165543
rect 670620 149025 670648 171935
rect 671356 151814 671384 215266
rect 671540 215266 671660 215294
rect 671724 221326 671844 221354
rect 671540 158409 671568 215266
rect 671724 173097 671752 221326
rect 671894 221232 671950 221241
rect 671894 221167 671950 221176
rect 671908 176497 671936 221167
rect 672092 217297 672120 224703
rect 672276 222194 672304 226902
rect 672380 226704 672432 226710
rect 672380 226646 672432 226652
rect 672392 226545 672420 226646
rect 672378 226536 672434 226545
rect 672378 226471 672434 226480
rect 672552 226114 672580 234110
rect 672184 222166 672304 222194
rect 672368 226086 672580 226114
rect 672368 222194 672396 226086
rect 672644 225672 672672 236399
rect 672744 235272 672796 235278
rect 672736 235220 672744 235226
rect 672736 235214 672796 235220
rect 672736 235198 672784 235214
rect 672736 231854 672764 235198
rect 672920 233510 672948 244246
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 672908 233504 672960 233510
rect 672908 233446 672960 233452
rect 673104 233322 673132 237458
rect 673380 234614 673408 245398
rect 673526 237144 673582 237153
rect 673526 237079 673582 237088
rect 673540 236910 673568 237079
rect 673528 236904 673580 236910
rect 673528 236846 673580 236852
rect 673656 236722 673684 258431
rect 673840 246537 673868 260879
rect 673826 246528 673882 246537
rect 673826 246463 673882 246472
rect 674024 244274 674052 266999
rect 674300 266121 674328 310383
rect 674470 303920 674526 303929
rect 674470 303855 674526 303864
rect 674484 286657 674512 303855
rect 674470 286648 674526 286657
rect 674470 286583 674526 286592
rect 674668 266665 674696 311199
rect 675022 309224 675078 309233
rect 675022 309159 675078 309168
rect 674838 308000 674894 308009
rect 674838 307935 674894 307944
rect 674852 292913 674880 307935
rect 675036 294250 675064 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 676232 305266 676260 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 675864 305238 676260 305266
rect 675864 302234 675892 305238
rect 675680 302206 675892 302234
rect 675680 299474 675708 302206
rect 675312 299446 675708 299474
rect 675312 295542 675340 299446
rect 675852 298104 675904 298110
rect 675852 298046 675904 298052
rect 675864 296585 675892 298046
rect 676036 297968 676088 297974
rect 676036 297910 676088 297916
rect 676048 296857 676076 297910
rect 678256 297401 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 681016 297974 681044 307527
rect 683026 302696 683082 302705
rect 683026 302631 683082 302640
rect 683040 299441 683068 302631
rect 683026 299432 683082 299441
rect 683026 299367 683082 299376
rect 681004 297968 681056 297974
rect 681004 297910 681056 297916
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 676034 296848 676090 296857
rect 676034 296783 676090 296792
rect 675850 296576 675906 296585
rect 675850 296511 675906 296520
rect 675312 295514 675418 295542
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675036 294222 675418 294250
rect 674838 292904 674894 292913
rect 674838 292839 674894 292848
rect 675390 292904 675446 292913
rect 675390 292839 675446 292848
rect 675404 292400 675432 292839
rect 675574 292088 675630 292097
rect 675574 292023 675630 292032
rect 675588 291856 675616 292023
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675404 290193 675432 290564
rect 675390 290184 675446 290193
rect 675390 290119 675446 290128
rect 675298 289912 675354 289921
rect 675298 289847 675354 289856
rect 675312 288538 675340 289847
rect 675312 288510 675432 288538
rect 675404 288048 675432 288510
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286648 675446 286657
rect 675390 286583 675446 286592
rect 675404 286212 675432 286583
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675680 281217 675708 281355
rect 675666 281208 675722 281217
rect 675666 281143 675722 281152
rect 683302 275360 683358 275369
rect 683302 275295 683358 275304
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 683132 268161 683160 271079
rect 683316 268569 683344 275295
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683302 268560 683358 268569
rect 683302 268495 683358 268504
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 674654 266656 674710 266665
rect 674654 266591 674710 266600
rect 674286 266112 674342 266121
rect 674286 266047 674342 266056
rect 676494 266112 676550 266121
rect 676494 266047 676550 266056
rect 676508 265305 676536 266047
rect 674562 265296 674618 265305
rect 674562 265231 674618 265240
rect 676494 265296 676550 265305
rect 676494 265231 676550 265240
rect 674576 253934 674604 265231
rect 674838 264480 674894 264489
rect 674838 264415 674894 264424
rect 674852 263809 674880 264415
rect 676494 264072 676550 264081
rect 676494 264007 676550 264016
rect 674838 263800 674894 263809
rect 674838 263735 674894 263744
rect 676508 263673 676536 264007
rect 676494 263664 676550 263673
rect 676494 263599 676550 263608
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 260522 676260 262783
rect 676140 260494 676260 260522
rect 675942 258768 675998 258777
rect 675942 258703 675998 258712
rect 675956 258233 675984 258703
rect 675942 258224 675998 258233
rect 675942 258159 675998 258168
rect 675298 257544 675354 257553
rect 675298 257479 675354 257488
rect 675312 256737 675340 257479
rect 675298 256728 675354 256737
rect 675298 256663 675354 256672
rect 676140 255921 676168 260494
rect 675206 255912 675262 255921
rect 675206 255847 675262 255856
rect 676126 255912 676182 255921
rect 676126 255847 676182 255856
rect 674576 253906 674788 253934
rect 674286 249656 674342 249665
rect 674286 249591 674342 249600
rect 673472 236694 673684 236722
rect 673932 244246 674052 244274
rect 674300 244274 674328 249591
rect 674300 244246 674696 244274
rect 673472 236314 673500 236694
rect 673644 236496 673696 236502
rect 673642 236464 673644 236473
rect 673696 236464 673698 236473
rect 673642 236399 673698 236408
rect 673752 236360 673804 236366
rect 673472 236286 673592 236314
rect 673752 236302 673804 236308
rect 673564 236076 673592 236286
rect 673012 233294 673132 233322
rect 673196 234586 673408 234614
rect 673472 236048 673592 236076
rect 673012 233238 673040 233294
rect 673000 233232 673052 233238
rect 673000 233174 673052 233180
rect 672736 231826 673040 231854
rect 672816 229016 672868 229022
rect 672816 228958 672868 228964
rect 672828 228857 672856 228958
rect 672814 228848 672870 228857
rect 672814 228783 672870 228792
rect 672814 228576 672870 228585
rect 672814 228511 672816 228520
rect 672868 228511 672870 228520
rect 672816 228482 672868 228488
rect 672816 228404 672868 228410
rect 672816 228346 672868 228352
rect 672828 227866 672856 228346
rect 672816 227860 672868 227866
rect 672816 227802 672868 227808
rect 672816 227520 672868 227526
rect 672552 225644 672672 225672
rect 672736 227468 672816 227474
rect 672736 227462 672868 227468
rect 672736 227446 672856 227462
rect 672552 225570 672580 225644
rect 672460 225542 672580 225570
rect 672460 223802 672488 225542
rect 672736 224641 672764 227446
rect 673012 226250 673040 231826
rect 673196 226817 673224 234586
rect 673472 230081 673500 236048
rect 673764 236042 673792 236302
rect 673748 236014 673792 236042
rect 673748 232801 673776 236014
rect 673932 234614 673960 244246
rect 674196 235476 674248 235482
rect 674196 235418 674248 235424
rect 674208 234954 674236 235418
rect 674426 235136 674478 235142
rect 674424 235104 674426 235113
rect 674478 235104 674480 235113
rect 674424 235039 674480 235048
rect 673840 234586 673960 234614
rect 674116 234926 674236 234954
rect 673840 232914 673868 234586
rect 674116 232914 674144 234926
rect 674286 234832 674342 234841
rect 674286 234767 674342 234776
rect 674300 234666 674328 234767
rect 674288 234660 674340 234666
rect 674288 234602 674340 234608
rect 674380 234252 674432 234258
rect 674380 234194 674432 234200
rect 673840 232886 673960 232914
rect 674116 232898 674236 232914
rect 674116 232892 674248 232898
rect 674116 232886 674196 232892
rect 673734 232792 673790 232801
rect 673734 232727 673790 232736
rect 673932 232642 673960 232886
rect 674196 232834 674248 232840
rect 673932 232614 674236 232642
rect 673642 232520 673698 232529
rect 673642 232455 673698 232464
rect 673656 230976 673684 232455
rect 673828 232008 673880 232014
rect 673828 231950 673880 231956
rect 673840 231130 673868 231950
rect 673828 231124 673880 231130
rect 673828 231066 673880 231072
rect 673656 230948 674144 230976
rect 673644 230852 673696 230858
rect 673644 230794 673696 230800
rect 673458 230072 673514 230081
rect 673458 230007 673514 230016
rect 673656 229537 673684 230794
rect 673918 230480 673974 230489
rect 673918 230415 673974 230424
rect 673932 229974 673960 230415
rect 674116 230058 674144 230948
rect 674070 230030 674144 230058
rect 674208 230058 674236 232614
rect 674392 230994 674420 234194
rect 674534 234152 674590 234161
rect 674534 234087 674536 234096
rect 674588 234087 674590 234096
rect 674536 234058 674588 234064
rect 674536 233640 674588 233646
rect 674588 233588 674604 233594
rect 674536 233582 674604 233588
rect 674548 233566 674604 233582
rect 674576 231962 674604 233566
rect 674484 231934 674604 231962
rect 674484 231554 674512 231934
rect 674668 231849 674696 244246
rect 674760 234546 674788 253906
rect 675022 251832 675078 251841
rect 675022 251767 675078 251776
rect 675036 249506 675064 251767
rect 675036 249478 675156 249506
rect 674930 249384 674986 249393
rect 674930 249319 674986 249328
rect 674944 246650 674972 249319
rect 675128 246854 675156 249478
rect 675220 247398 675248 255847
rect 676036 252408 676088 252414
rect 676036 252350 676088 252356
rect 675852 252272 675904 252278
rect 675312 252220 675852 252226
rect 675312 252214 675904 252220
rect 675312 252198 675892 252214
rect 675312 250526 675340 252198
rect 676048 251841 676076 252350
rect 678256 252278 678284 263191
rect 679622 261216 679678 261225
rect 679622 261151 679678 261160
rect 679636 252414 679664 261151
rect 679624 252408 679676 252414
rect 679624 252350 679676 252356
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 676034 251832 676090 251841
rect 676034 251767 676090 251776
rect 675312 250498 675418 250526
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249656 675446 249665
rect 675390 249591 675446 249600
rect 675404 249220 675432 249591
rect 675220 247370 675418 247398
rect 675128 246826 675418 246854
rect 674944 246622 675248 246650
rect 674930 245576 674986 245585
rect 674930 245511 674986 245520
rect 674944 241890 674972 245511
rect 675220 243085 675248 246622
rect 675390 246528 675446 246537
rect 675390 246463 675446 246472
rect 675404 246199 675432 246463
rect 675390 245848 675446 245857
rect 675390 245783 675446 245792
rect 675404 245548 675432 245783
rect 675220 243057 675418 243085
rect 675114 242856 675170 242865
rect 675114 242791 675170 242800
rect 675128 242533 675156 242791
rect 675128 242505 675418 242533
rect 674944 241862 675418 241890
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675036 238190 675418 238218
rect 675036 235929 675064 238190
rect 675390 238096 675446 238105
rect 675390 238031 675446 238040
rect 675404 237524 675432 238031
rect 675206 237280 675262 237289
rect 675206 237215 675262 237224
rect 675220 236382 675248 237215
rect 675220 236354 675418 236382
rect 675022 235920 675078 235929
rect 675022 235855 675078 235864
rect 674760 234530 675892 234546
rect 674760 234524 675904 234530
rect 674760 234518 675852 234524
rect 675852 234466 675904 234472
rect 679808 234524 679860 234530
rect 679808 234466 679860 234472
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674898 234002 674926 234262
rect 675850 234152 675906 234161
rect 675850 234087 675852 234096
rect 675904 234087 675906 234096
rect 679624 234116 679676 234122
rect 675852 234058 675904 234064
rect 679624 234058 679676 234064
rect 674852 233974 674926 234002
rect 674852 233034 674880 233974
rect 674978 233912 675030 233918
rect 675030 233860 675892 233866
rect 674978 233854 675892 233860
rect 674990 233850 675892 233854
rect 674990 233844 675904 233850
rect 674990 233838 675852 233844
rect 675852 233786 675904 233792
rect 677876 233844 677928 233850
rect 677876 233786 677928 233792
rect 675116 233776 675168 233782
rect 675116 233718 675168 233724
rect 675128 233617 675156 233718
rect 675114 233608 675170 233617
rect 675114 233543 675170 233552
rect 675208 233436 675260 233442
rect 675208 233378 675260 233384
rect 675220 233322 675248 233378
rect 675220 233306 675892 233322
rect 675220 233300 675904 233306
rect 675220 233294 675852 233300
rect 675852 233242 675904 233248
rect 674840 233028 674892 233034
rect 674840 232970 674892 232976
rect 675496 232626 675892 232642
rect 675484 232620 675892 232626
rect 675536 232614 675892 232620
rect 675484 232562 675536 232568
rect 675864 232558 675892 232614
rect 675852 232552 675904 232558
rect 675852 232494 675904 232500
rect 674654 231840 674710 231849
rect 674654 231775 674710 231784
rect 674840 231804 674892 231810
rect 674840 231746 674892 231752
rect 674654 231568 674710 231577
rect 674484 231526 674558 231554
rect 674530 231470 674558 231526
rect 674654 231503 674710 231512
rect 674518 231464 674570 231470
rect 674518 231406 674570 231412
rect 674668 231198 674696 231503
rect 674656 231192 674708 231198
rect 674656 231134 674708 231140
rect 674732 231056 674784 231062
rect 674730 231024 674732 231033
rect 674784 231024 674786 231033
rect 674380 230988 674432 230994
rect 674730 230959 674786 230968
rect 674380 230930 674432 230936
rect 674852 230761 674880 231746
rect 675850 231568 675906 231577
rect 675070 231532 675122 231538
rect 675850 231503 675852 231512
rect 675070 231474 675122 231480
rect 675904 231503 675906 231512
rect 677600 231532 677652 231538
rect 675852 231474 675904 231480
rect 677600 231474 677652 231480
rect 674956 231328 675008 231334
rect 675082 231305 675110 231474
rect 674956 231270 675008 231276
rect 675068 231296 675124 231305
rect 674968 231146 674996 231270
rect 675068 231231 675124 231240
rect 674968 231130 675892 231146
rect 674968 231124 675904 231130
rect 674968 231118 675852 231124
rect 675852 231066 675904 231072
rect 674838 230752 674894 230761
rect 674838 230687 674894 230696
rect 675022 230752 675078 230761
rect 675022 230687 675078 230696
rect 675850 230752 675906 230761
rect 675850 230687 675906 230696
rect 674380 230648 674432 230654
rect 675036 230602 675064 230687
rect 674432 230596 675064 230602
rect 674380 230590 675064 230596
rect 674392 230574 675064 230590
rect 674518 230512 674570 230518
rect 674518 230454 674570 230460
rect 674396 230308 674448 230314
rect 674396 230250 674448 230256
rect 674408 230183 674436 230250
rect 674530 230194 674558 230454
rect 674654 230208 674710 230217
rect 674394 230174 674450 230183
rect 674530 230166 674654 230194
rect 674654 230143 674710 230152
rect 674394 230109 674450 230118
rect 674208 230030 674328 230058
rect 675864 230042 675892 230687
rect 676218 230480 676274 230489
rect 676218 230415 676274 230424
rect 673920 229968 673972 229974
rect 673920 229910 673972 229916
rect 673826 229800 673882 229809
rect 674070 229786 674098 230030
rect 674172 229968 674224 229974
rect 674170 229936 674172 229945
rect 674224 229936 674226 229945
rect 674170 229871 674226 229880
rect 674070 229758 674236 229786
rect 673826 229735 673882 229744
rect 673642 229528 673698 229537
rect 673840 229498 673868 229735
rect 673948 229560 674000 229566
rect 673946 229528 673948 229537
rect 674000 229528 674002 229537
rect 673642 229463 673698 229472
rect 673828 229492 673880 229498
rect 673946 229463 674002 229472
rect 673828 229434 673880 229440
rect 673918 229256 673974 229265
rect 673472 229214 673918 229242
rect 673472 229158 673500 229214
rect 673918 229191 673974 229200
rect 673460 229152 673512 229158
rect 673736 229152 673788 229158
rect 673460 229094 673512 229100
rect 673734 229120 673736 229129
rect 673788 229120 673790 229129
rect 673734 229055 673790 229064
rect 673598 228948 673650 228954
rect 673598 228890 673650 228896
rect 673610 228834 673638 228890
rect 673610 228806 673960 228834
rect 673506 228744 673558 228750
rect 673558 228704 673776 228732
rect 673506 228686 673558 228692
rect 673182 226808 673238 226817
rect 673182 226743 673238 226752
rect 673012 226222 673132 226250
rect 672722 224632 672778 224641
rect 672722 224567 672778 224576
rect 672906 224088 672962 224097
rect 672906 224023 672962 224032
rect 672722 223952 672778 223961
rect 672722 223887 672778 223896
rect 672460 223774 672672 223802
rect 672368 222166 672580 222194
rect 672184 217546 672212 222166
rect 672552 222034 672580 222166
rect 672276 222006 672580 222034
rect 672276 220814 672304 222006
rect 672446 221912 672502 221921
rect 672446 221847 672502 221856
rect 672460 221762 672488 221847
rect 672644 221762 672672 223774
rect 672460 221734 672672 221762
rect 672276 220786 672580 220814
rect 672552 219042 672580 220786
rect 672736 220674 672764 223887
rect 672920 220969 672948 224023
rect 672906 220960 672962 220969
rect 672906 220895 672962 220904
rect 672736 220646 672856 220674
rect 672828 220402 672856 220646
rect 672644 220374 672856 220402
rect 672644 220130 672672 220374
rect 672644 220102 672764 220130
rect 672736 219201 672764 220102
rect 672722 219192 672778 219201
rect 672722 219127 672778 219136
rect 672552 219014 672764 219042
rect 672184 217518 672396 217546
rect 672078 217288 672134 217297
rect 672078 217223 672134 217232
rect 672078 213752 672134 213761
rect 672078 213687 672134 213696
rect 672092 200841 672120 213687
rect 672368 205634 672396 217518
rect 672538 214024 672594 214033
rect 672538 213959 672594 213968
rect 672552 211154 672580 213959
rect 672736 211154 672764 219014
rect 673104 218498 673132 226222
rect 673458 226128 673514 226137
rect 673458 226063 673514 226072
rect 673472 224954 673500 226063
rect 673748 225570 673776 228704
rect 673932 226273 673960 228806
rect 673918 226264 673974 226273
rect 673918 226199 673974 226208
rect 673918 225584 673974 225593
rect 673748 225542 673918 225570
rect 673918 225519 673974 225528
rect 673734 225448 673790 225457
rect 674208 225434 674236 229758
rect 673734 225383 673790 225392
rect 674116 225406 674236 225434
rect 673472 224926 673592 224954
rect 673274 224632 673330 224641
rect 673274 224567 673330 224576
rect 673288 222194 673316 224567
rect 672276 205606 672396 205634
rect 672460 211126 672580 211154
rect 672644 211126 672764 211154
rect 673012 218470 673132 218498
rect 673196 222166 673316 222194
rect 672078 200832 672134 200841
rect 672078 200767 672134 200776
rect 672276 198801 672304 205606
rect 672262 198792 672318 198801
rect 672262 198727 672318 198736
rect 672460 184929 672488 211126
rect 672446 184920 672502 184929
rect 672446 184855 672502 184864
rect 672078 183560 672134 183569
rect 672078 183495 672134 183504
rect 671894 176488 671950 176497
rect 671894 176423 671950 176432
rect 671710 173088 671766 173097
rect 671710 173023 671766 173032
rect 671894 169960 671950 169969
rect 671894 169895 671950 169904
rect 671710 166968 671766 166977
rect 671710 166903 671766 166912
rect 671526 158400 671582 158409
rect 671526 158335 671582 158344
rect 670804 151786 671384 151814
rect 670804 150278 670832 151786
rect 670792 150272 670844 150278
rect 670792 150214 670844 150220
rect 670606 149016 670662 149025
rect 670606 148951 670662 148960
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670332 118584 670384 118590
rect 670332 118526 670384 118532
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 671356 113174 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670712 113146 671384 113174
rect 589924 111046 589976 111052
rect 668582 111072 668638 111081
rect 668582 111007 668638 111016
rect 668122 110800 668178 110809
rect 668122 110735 668178 110744
rect 590106 110120 590162 110129
rect 590106 110055 590162 110064
rect 589372 109744 589424 109750
rect 589372 109686 589424 109692
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589646 106856 589702 106865
rect 589646 106791 589702 106800
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589660 104174 589688 106791
rect 589648 104168 589700 104174
rect 589648 104110 589700 104116
rect 589922 101960 589978 101969
rect 589922 101895 589978 101904
rect 588544 88324 588596 88330
rect 588544 88266 588596 88272
rect 589936 79354 589964 101895
rect 590120 100026 590148 110055
rect 666560 106140 666612 106146
rect 666836 106140 666888 106146
rect 666560 106082 666612 106088
rect 666834 106108 666836 106117
rect 666888 106108 666890 106117
rect 590290 103592 590346 103601
rect 590290 103527 590346 103536
rect 590304 100774 590332 103527
rect 590292 100768 590344 100774
rect 590292 100710 590344 100716
rect 624792 100156 624844 100162
rect 624792 100098 624844 100104
rect 590108 100020 590160 100026
rect 590108 99962 590160 99968
rect 594064 100020 594116 100026
rect 594064 99962 594116 99968
rect 595272 100014 595608 100042
rect 591304 97708 591356 97714
rect 591304 97650 591356 97656
rect 589924 79348 589976 79354
rect 589924 79290 589976 79296
rect 587164 73160 587216 73166
rect 587164 73102 587216 73108
rect 584404 71596 584456 71602
rect 584404 71538 584456 71544
rect 584404 68332 584456 68338
rect 584404 68274 584456 68280
rect 584416 54777 584444 68274
rect 591316 55078 591344 97650
rect 594076 64870 594104 99962
rect 595272 99142 595300 100014
rect 596330 99770 596358 100028
rect 596284 99742 596358 99770
rect 596468 100014 597080 100042
rect 597572 100014 597816 100042
rect 598216 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601712 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 594064 64864 594116 64870
rect 594064 64806 594116 64812
rect 591304 55072 591356 55078
rect 591304 55014 591356 55020
rect 596284 54806 596312 99742
rect 596468 54942 596496 100014
rect 597572 58818 597600 100014
rect 598216 97714 598244 100014
rect 598204 97708 598256 97714
rect 598204 97650 598256 97656
rect 597560 58812 597612 58818
rect 597560 58754 597612 58760
rect 598952 56030 598980 100014
rect 599504 84194 599532 100014
rect 600424 95946 600452 100014
rect 600412 95940 600464 95946
rect 600412 95882 600464 95888
rect 600884 84194 600912 100014
rect 601712 89010 601740 100014
rect 601700 89004 601752 89010
rect 601700 88946 601752 88952
rect 602356 84194 602384 100014
rect 599136 84166 599532 84194
rect 600516 84166 600912 84194
rect 601896 84166 602384 84194
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 599136 55894 599164 84166
rect 600516 57390 600544 84166
rect 600504 57384 600556 57390
rect 600504 57326 600556 57332
rect 601896 57254 601924 84166
rect 603092 58682 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 604426 99742 604500 99770
rect 604472 68338 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 94518 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 94512 606996 94518
rect 606944 94454 606996 94460
rect 607140 75342 607168 96902
rect 607692 94654 607720 100014
rect 607680 94648 607732 94654
rect 607680 94590 607732 94596
rect 608520 84182 608548 100014
rect 609164 95946 609192 100014
rect 609152 95940 609204 95946
rect 609152 95882 609204 95888
rect 609900 85542 609928 100014
rect 610636 96966 610664 100014
rect 610624 96960 610676 96966
rect 610624 96902 610676 96908
rect 611084 96960 611136 96966
rect 611084 96902 611136 96908
rect 611096 93158 611124 96902
rect 611084 93152 611136 93158
rect 611084 93094 611136 93100
rect 611280 91050 611308 100014
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 613384 97300 613436 97306
rect 613384 97242 613436 97248
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 612002 95840 612058 95849
rect 612002 95775 612058 95784
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 607128 75336 607180 75342
rect 607128 75278 607180 75284
rect 604460 68332 604512 68338
rect 604460 68274 604512 68280
rect 612016 62082 612044 95775
rect 612660 79490 612688 96834
rect 612648 79484 612700 79490
rect 612648 79426 612700 79432
rect 613396 75206 613424 97242
rect 613580 96830 613608 100014
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 615480 100014 615816 100042
rect 616216 100014 616644 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 614040 96966 614068 99742
rect 614028 96960 614080 96966
rect 614028 96902 614080 96908
rect 614764 96960 614816 96966
rect 614764 96902 614816 96908
rect 613568 96824 613620 96830
rect 613568 96766 613620 96772
rect 614028 96824 614080 96830
rect 614028 96766 614080 96772
rect 614040 77994 614068 96766
rect 614776 79354 614804 96902
rect 615052 93854 615080 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 615052 93826 615448 93854
rect 615420 80850 615448 93826
rect 616616 91798 616644 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616604 91792 616656 91798
rect 616604 91734 616656 91740
rect 615408 80844 615460 80850
rect 615408 80786 615460 80792
rect 614764 79348 614816 79354
rect 614764 79290 614816 79296
rect 614028 77988 614080 77994
rect 614028 77930 614080 77936
rect 616800 76702 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91186 618208 96834
rect 619560 93838 619588 100014
rect 620204 97714 620232 100014
rect 620192 97708 620244 97714
rect 620192 97650 620244 97656
rect 620284 97436 620336 97442
rect 620284 97378 620336 97384
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618536 93152 618588 93158
rect 618536 93094 618588 93100
rect 618168 91180 618220 91186
rect 618168 91122 618220 91128
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618180 88330 618208 90986
rect 618168 88324 618220 88330
rect 618168 88266 618220 88272
rect 618548 86358 618576 93094
rect 618536 86352 618588 86358
rect 618536 86294 618588 86300
rect 616788 76696 616840 76702
rect 616788 76638 616840 76644
rect 620296 75478 620324 97378
rect 620940 95198 620968 100014
rect 621676 97306 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 623148 97442 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97436 623188 97442
rect 623136 97378 623188 97384
rect 621664 97300 621716 97306
rect 621664 97242 621716 97248
rect 624620 97034 624648 100014
rect 624608 97028 624660 97034
rect 624608 96970 624660 96976
rect 621664 95940 621716 95946
rect 621664 95882 621716 95888
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620928 94648 620980 94654
rect 620928 94590 620980 94596
rect 620940 89690 620968 94590
rect 620928 89684 620980 89690
rect 620928 89626 620980 89632
rect 621676 85406 621704 95882
rect 623044 94512 623096 94518
rect 623044 94454 623096 94460
rect 623056 88194 623084 94454
rect 623044 88188 623096 88194
rect 623044 88130 623096 88136
rect 621664 85400 621716 85406
rect 621664 85342 621716 85348
rect 624804 84194 624832 100098
rect 625034 99770 625062 100028
rect 625784 100014 626212 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 625816 92041 625844 97922
rect 625988 97708 626040 97714
rect 625988 97650 626040 97656
rect 626000 93673 626028 97650
rect 626184 97578 626212 100014
rect 626828 97714 626856 100014
rect 627564 98938 627592 100014
rect 627552 98932 627604 98938
rect 627552 98874 627604 98880
rect 628300 97850 628328 100014
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 628288 97844 628340 97850
rect 628288 97786 628340 97792
rect 626816 97708 626868 97714
rect 626816 97650 626868 97656
rect 626172 97572 626224 97578
rect 626172 97514 626224 97520
rect 629300 97300 629352 97306
rect 629300 97242 629352 97248
rect 629312 95826 629340 97242
rect 630784 95826 630812 99282
rect 631244 96354 631272 100014
rect 631416 98252 631468 98258
rect 631416 98194 631468 98200
rect 631428 97850 631456 98194
rect 631416 97844 631468 97850
rect 631416 97786 631468 97792
rect 631600 97844 631652 97850
rect 631600 97786 631652 97792
rect 631612 97578 631640 97786
rect 631980 97578 632008 100014
rect 631600 97572 631652 97578
rect 631600 97514 631652 97520
rect 631968 97572 632020 97578
rect 631968 97514 632020 97520
rect 632716 97442 632744 100014
rect 632060 97436 632112 97442
rect 632060 97378 632112 97384
rect 632704 97436 632756 97442
rect 632704 97378 632756 97384
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97378
rect 633268 97306 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 633256 97300 633308 97306
rect 633256 97242 633308 97248
rect 633452 95826 633480 99146
rect 634188 96898 634216 100014
rect 634740 97170 634768 100014
rect 634728 97164 634780 97170
rect 634728 97106 634780 97112
rect 635004 97028 635056 97034
rect 635004 96970 635056 96976
rect 634176 96892 634228 96898
rect 634176 96834 634228 96840
rect 635016 95826 635044 96970
rect 635568 96393 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635554 96384 635610 96393
rect 635554 96319 635610 96328
rect 635752 96121 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 635738 96112 635794 96121
rect 635738 96047 635794 96056
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97844 637816 97850
rect 637764 97786 637816 97792
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97786
rect 638604 97034 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 638592 97028 638644 97034
rect 638592 96970 638644 96976
rect 639064 96626 639092 99742
rect 639236 97708 639288 97714
rect 639236 97650 639288 97656
rect 639052 96620 639104 96626
rect 639052 96562 639104 96568
rect 639248 95826 639276 97650
rect 640076 96490 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640536 96626 640564 99742
rect 640708 98932 640760 98938
rect 640708 98874 640760 98880
rect 640340 96620 640392 96626
rect 640340 96562 640392 96568
rect 640524 96620 640576 96626
rect 640524 96562 640576 96568
rect 640064 96484 640116 96490
rect 640064 96426 640116 96432
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639248 95798 639584 95826
rect 640352 95470 640380 96562
rect 640720 95826 640748 98874
rect 641548 96082 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96121 642036 99742
rect 642180 98184 642232 98190
rect 642180 98126 642232 98132
rect 641994 96112 642050 96121
rect 641536 96076 641588 96082
rect 641994 96047 642050 96056
rect 641536 96018 641588 96024
rect 642192 95826 642220 98126
rect 643020 97714 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97708 643060 97714
rect 643008 97650 643060 97656
rect 640720 95798 641056 95826
rect 642192 95798 642528 95826
rect 643480 95470 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643664 95826 643692 98738
rect 644308 97850 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644860 99742 644934 99770
rect 644296 97844 644348 97850
rect 644296 97786 644348 97792
rect 644860 95946 644888 99742
rect 645124 98048 645176 98054
rect 645124 97990 645176 97996
rect 644848 95940 644900 95946
rect 644848 95882 644900 95888
rect 645136 95826 645164 97990
rect 643664 95798 644000 95826
rect 645136 95798 645472 95826
rect 645780 95810 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648292 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 95804 645820 95810
rect 645768 95746 645820 95752
rect 646424 95674 646452 99742
rect 647160 98802 647188 99742
rect 647148 98796 647200 98802
rect 647148 98738 647200 98744
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646608 95826 646636 98602
rect 647792 97028 647844 97034
rect 647792 96970 647844 96976
rect 647804 96778 647832 96970
rect 647976 96892 648028 96898
rect 647976 96834 648028 96840
rect 647988 96778 648016 96834
rect 647712 96750 647832 96778
rect 647896 96750 648016 96778
rect 647422 96384 647478 96393
rect 647148 96348 647200 96354
rect 647422 96319 647478 96328
rect 647148 96290 647200 96296
rect 646608 95798 646944 95826
rect 646412 95668 646464 95674
rect 646412 95610 646464 95616
rect 640340 95464 640392 95470
rect 640340 95406 640392 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 626460 94489 626488 95134
rect 647160 95033 647188 96290
rect 647146 95024 647202 95033
rect 647146 94959 647202 94968
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 625986 93664 626042 93673
rect 625986 93599 626042 93608
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626264 91792 626316 91798
rect 626264 91734 626316 91740
rect 626276 89593 626304 91734
rect 626460 91225 626488 92414
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626262 89584 626318 89593
rect 626262 89519 626318 89528
rect 626460 88777 626488 89626
rect 626446 88768 626502 88777
rect 626446 88703 626502 88712
rect 625620 88324 625672 88330
rect 625620 88266 625672 88272
rect 625632 87145 625660 88266
rect 626448 88188 626500 88194
rect 626448 88130 626500 88136
rect 626460 87961 626488 88130
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 625618 87136 625674 87145
rect 625618 87071 625674 87080
rect 626448 86352 626500 86358
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 624436 84166 624832 84194
rect 626448 84176 626500 84182
rect 621664 75948 621716 75954
rect 621664 75890 621716 75896
rect 620284 75472 620336 75478
rect 620284 75414 620336 75420
rect 613384 75200 613436 75206
rect 613384 75142 613436 75148
rect 612004 62076 612056 62082
rect 612004 62018 612056 62024
rect 603080 58676 603132 58682
rect 603080 58618 603132 58624
rect 601884 57248 601936 57254
rect 601884 57190 601936 57196
rect 621676 56574 621704 75890
rect 623044 66292 623096 66298
rect 623044 66234 623096 66240
rect 621664 56568 621716 56574
rect 621664 56510 621716 56516
rect 599124 55888 599176 55894
rect 599124 55830 599176 55836
rect 596456 54936 596508 54942
rect 596456 54878 596508 54884
rect 596272 54800 596324 54806
rect 584402 54768 584458 54777
rect 596272 54742 596324 54748
rect 584402 54703 584458 54712
rect 581642 54496 581698 54505
rect 581642 54431 581698 54440
rect 580448 54392 580500 54398
rect 580448 54334 580500 54340
rect 579068 54256 579120 54262
rect 579068 54198 579120 54204
rect 574928 53926 574980 53932
rect 577686 53952 577742 53961
rect 577686 53887 577742 53896
rect 459466 53680 459522 53689
rect 459466 53615 459522 53624
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 462594 53680 462650 53689
rect 461674 53615 461730 53624
rect 462136 53644 462188 53650
rect 129188 53372 129240 53378
rect 129188 53314 129240 53320
rect 129004 53100 129056 53106
rect 129004 53042 129056 53048
rect 129016 51074 129044 53042
rect 129016 51046 129136 51074
rect 128728 50516 128780 50522
rect 128728 50458 128780 50464
rect 128544 50380 128596 50386
rect 128544 50322 128596 50328
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 47768 49020 47820 49026
rect 47768 48962 47820 48968
rect 128556 44198 128584 50322
rect 128740 47734 128768 50458
rect 128912 49156 128964 49162
rect 128912 49098 128964 49104
rect 128924 47870 128952 49098
rect 128912 47864 128964 47870
rect 128912 47806 128964 47812
rect 128728 47728 128780 47734
rect 128728 47670 128780 47676
rect 129108 44826 129136 51046
rect 129016 44798 129136 44826
rect 129016 44538 129044 44798
rect 129200 44674 129228 53314
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 129556 52012 129608 52018
rect 129556 51954 129608 51960
rect 129372 51876 129424 51882
rect 129372 51818 129424 51824
rect 129384 44810 129412 51818
rect 129568 45082 129596 51954
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129372 44804 129424 44810
rect 129372 44746 129424 44752
rect 129188 44668 129240 44674
rect 129188 44610 129240 44616
rect 129004 44532 129056 44538
rect 129004 44474 129056 44480
rect 128544 44192 128596 44198
rect 128544 44134 128596 44140
rect 130396 44062 130424 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 306024 51746 306052 53108
rect 130568 51740 130620 51746
rect 130568 51682 130620 51688
rect 145380 51740 145432 51746
rect 145380 51682 145432 51688
rect 306012 51740 306064 51746
rect 306012 51682 306064 51688
rect 130580 44334 130608 51682
rect 145392 50810 145420 51682
rect 145084 50782 145420 50810
rect 131028 49020 131080 49026
rect 131028 48962 131080 48968
rect 130568 44328 130620 44334
rect 130568 44270 130620 44276
rect 130384 44056 130436 44062
rect 130384 43998 130436 44004
rect 131040 43926 131068 48962
rect 308048 48929 308076 53108
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53615
rect 459848 52578 459876 53615
rect 460066 52828 460118 52834
rect 460066 52770 460118 52776
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460078 52564 460106 52770
rect 460768 52578 460796 53615
rect 461308 53508 461360 53514
rect 461308 53450 461360 53456
rect 461320 52578 461348 53450
rect 461688 52578 461716 53615
rect 462594 53615 462650 53624
rect 463332 53644 463384 53650
rect 462136 53586 462188 53592
rect 462148 52578 462176 53586
rect 462608 52578 462636 53615
rect 463332 53586 463384 53592
rect 464068 53644 464120 53650
rect 464068 53586 464120 53592
rect 464988 53644 465040 53650
rect 464988 53586 465040 53592
rect 465908 53644 465960 53650
rect 465908 53586 465960 53592
rect 467932 53644 467984 53650
rect 467932 53586 467984 53592
rect 468576 53644 468628 53650
rect 468576 53586 468628 53592
rect 468760 53644 468812 53650
rect 468760 53586 468812 53592
rect 463148 53372 463200 53378
rect 463148 53314 463200 53320
rect 463160 52578 463188 53314
rect 463344 52578 463372 53586
rect 464080 52578 464108 53586
rect 464206 52828 464258 52834
rect 464206 52770 464258 52776
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462176 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463372 52578
rect 463772 52550 464108 52578
rect 464218 52564 464246 52770
rect 465000 52578 465028 53586
rect 465448 53168 465500 53174
rect 465448 53110 465500 53116
rect 465460 52578 465488 53110
rect 465920 52578 465948 53586
rect 467944 52970 467972 53586
rect 468588 53174 468616 53586
rect 468576 53168 468628 53174
rect 468576 53110 468628 53116
rect 467932 52964 467984 52970
rect 467932 52906 467984 52912
rect 468772 52834 468800 53586
rect 468760 52828 468812 52834
rect 468760 52770 468812 52776
rect 464692 52550 465028 52578
rect 465152 52550 465488 52578
rect 465612 52550 465948 52578
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 308034 48920 308090 48929
rect 308034 48855 308090 48864
rect 131580 47864 131632 47870
rect 131580 47806 131632 47812
rect 131592 44810 131620 47806
rect 132040 47728 132092 47734
rect 132040 47670 132092 47676
rect 131580 44804 131632 44810
rect 131580 44746 131632 44752
rect 132052 44538 132080 47670
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460796 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132040 44532 132092 44538
rect 132040 44474 132092 44480
rect 132408 44464 132460 44470
rect 132236 44412 132408 44418
rect 132236 44406 132460 44412
rect 132236 44390 132448 44406
rect 132236 44198 132264 44390
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 132224 44192 132276 44198
rect 132224 44134 132276 44140
rect 307298 44160 307354 44169
rect 307298 44095 307354 44104
rect 131028 43920 131080 43926
rect 131028 43862 131080 43868
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 43444 42832 43496 42838
rect 43444 42774 43496 42780
rect 187344 42092 187372 43522
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 44095
rect 419722 43888 419778 43897
rect 419722 43823 419778 43832
rect 415398 43616 415454 43625
rect 415398 43551 415454 43560
rect 310428 42764 310480 42770
rect 310428 42706 310480 42712
rect 310440 42106 310468 42706
rect 415412 42364 415440 43551
rect 419736 42500 419764 43823
rect 431236 43654 431264 44775
rect 456062 43888 456118 43897
rect 456062 43823 456118 43832
rect 431224 43648 431276 43654
rect 439596 43648 439648 43654
rect 431224 43590 431276 43596
rect 439594 43616 439596 43625
rect 441620 43648 441672 43654
rect 439648 43616 439650 43625
rect 439594 43551 439650 43560
rect 441618 43616 441620 43625
rect 441672 43616 441674 43625
rect 441618 43551 441674 43560
rect 456076 43353 456104 43823
rect 456062 43344 456118 43353
rect 456062 43279 456118 43288
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405556 42356 405608 42362
rect 405556 42298 405608 42304
rect 420736 42356 420788 42362
rect 420736 42298 420788 42304
rect 427084 42356 427136 42362
rect 427084 42298 427136 42304
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 194322 42055 194378 42064
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 365166 41848 365222 41857
rect 364918 41806 365166 41834
rect 361946 41783 362002 41792
rect 365166 41783 365222 41792
rect 404464 41478 404492 42298
rect 405568 42092 405596 42298
rect 416686 42256 416742 42265
rect 416686 42191 416742 42200
rect 416700 42106 416728 42191
rect 416622 42078 416728 42106
rect 420748 41478 420776 42298
rect 427096 41478 427124 42298
rect 431236 42090 431264 42706
rect 446402 42256 446458 42265
rect 446402 42191 446458 42200
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 446416 41585 446444 42191
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 446402 41576 446458 41585
rect 446402 41511 446458 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460768 43081 460796 47654
rect 460998 47410 461026 47668
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 460952 47382 461026 47410
rect 460754 43072 460810 43081
rect 460754 43007 460810 43016
rect 460952 42401 460980 47382
rect 461780 43625 461808 47654
rect 461964 43897 461992 47654
rect 462700 43897 462728 47654
rect 461950 43888 462006 43897
rect 461950 43823 462006 43832
rect 462686 43888 462742 43897
rect 462686 43823 462742 43832
rect 461766 43616 461822 43625
rect 461766 43551 461822 43560
rect 462884 43353 462912 47654
rect 463068 47654 463312 47682
rect 462870 43344 462926 43353
rect 462870 43279 462926 43288
rect 463068 42770 463096 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464356 47654 464692 47682
rect 463712 44441 463740 47382
rect 463698 44432 463754 44441
rect 463698 44367 463754 44376
rect 463896 44169 463924 47654
rect 464356 44305 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 623056 46510 623084 66234
rect 624436 60722 624464 84166
rect 626448 84118 626500 84124
rect 626460 83881 626488 84118
rect 626446 83872 626502 83881
rect 626446 83807 626502 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 80986 628788 83263
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 80980 628800 80986
rect 628748 80922 628800 80928
rect 629220 80034 629248 81631
rect 632808 80974 633144 81002
rect 642456 80980 642508 80986
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 628472 77444 628524 77450
rect 628472 77386 628524 77392
rect 625804 77308 625856 77314
rect 625804 77250 625856 77256
rect 624424 60716 624476 60722
rect 624424 60658 624476 60664
rect 625816 54534 625844 77250
rect 625986 75984 626042 75993
rect 628484 75954 628512 77386
rect 631060 77314 631088 78066
rect 632808 77450 632836 80974
rect 643080 80974 643140 81002
rect 642456 80922 642508 80928
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78266 633480 79970
rect 633440 78260 633492 78266
rect 633440 78202 633492 78208
rect 633898 77616 633954 77625
rect 633898 77551 633954 77560
rect 632796 77444 632848 77450
rect 632796 77386 632848 77392
rect 631048 77308 631100 77314
rect 631048 77250 631100 77256
rect 625986 75919 626042 75928
rect 628472 75948 628524 75954
rect 626000 54670 626028 75919
rect 628472 75890 628524 75896
rect 628484 75290 628512 75890
rect 631060 75290 631088 77250
rect 633912 75993 633940 77551
rect 633898 75984 633954 75993
rect 633898 75919 633954 75928
rect 633912 75290 633940 75919
rect 636764 75290 636792 80650
rect 639602 77888 639658 77897
rect 639602 77823 639658 77832
rect 639616 75290 639644 77823
rect 642468 75290 642496 80922
rect 643112 78130 643140 80974
rect 646136 80844 646188 80850
rect 646136 80786 646188 80792
rect 645952 79484 646004 79490
rect 645952 79426 646004 79432
rect 645308 78260 645360 78266
rect 645308 78202 645360 78208
rect 643100 78124 643152 78130
rect 643100 78066 643152 78072
rect 645320 75290 645348 78202
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 645964 64874 645992 79426
rect 646148 69193 646176 80786
rect 647240 77988 647292 77994
rect 647240 77930 647292 77936
rect 646504 76696 646556 76702
rect 646504 76638 646556 76644
rect 646320 75336 646372 75342
rect 646320 75278 646372 75284
rect 646332 74225 646360 75278
rect 646318 74216 646374 74225
rect 646318 74151 646374 74160
rect 646516 71777 646544 76638
rect 646502 71768 646558 71777
rect 646502 71703 646558 71712
rect 646134 69184 646190 69193
rect 646134 69119 646190 69128
rect 645964 64846 646176 64874
rect 646148 59401 646176 64846
rect 647252 64433 647280 77930
rect 647238 64424 647294 64433
rect 647238 64359 647294 64368
rect 646134 59392 646190 59401
rect 646134 59327 646190 59336
rect 647436 57361 647464 96319
rect 647712 91730 647740 96750
rect 647896 95826 647924 96750
rect 648068 95940 648120 95946
rect 648068 95882 648120 95888
rect 647896 95798 648016 95826
rect 647988 95282 648016 95798
rect 648080 95554 648108 95882
rect 648264 95826 648292 100014
rect 648620 97572 648672 97578
rect 648620 97514 648672 97520
rect 648436 96620 648488 96626
rect 648436 96562 648488 96568
rect 648448 95946 648476 96562
rect 648436 95940 648488 95946
rect 648436 95882 648488 95888
rect 648264 95798 648476 95826
rect 648080 95526 648200 95554
rect 648172 95402 648200 95526
rect 648160 95396 648212 95402
rect 648160 95338 648212 95344
rect 647988 95254 648108 95282
rect 648080 95198 648108 95254
rect 647884 95192 647936 95198
rect 647884 95134 647936 95140
rect 648068 95192 648120 95198
rect 648068 95134 648120 95140
rect 647700 91724 647752 91730
rect 647700 91666 647752 91672
rect 647896 86766 647924 95134
rect 648448 93906 648476 95798
rect 648436 93900 648488 93906
rect 648436 93842 648488 93848
rect 648632 92041 648660 97514
rect 648908 96354 648936 100014
rect 649080 97164 649132 97170
rect 649080 97106 649132 97112
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 648804 95056 648856 95062
rect 648804 94998 648856 95004
rect 648618 92032 648674 92041
rect 648618 91967 648674 91976
rect 648816 90710 648844 94998
rect 648804 90704 648856 90710
rect 648804 90646 648856 90652
rect 649092 89714 649120 97106
rect 648908 89686 649120 89714
rect 647884 86760 647936 86766
rect 647884 86702 647936 86708
rect 648908 82249 648936 89686
rect 649736 88806 649764 100014
rect 650380 97578 650408 100014
rect 650368 97572 650420 97578
rect 650368 97514 650420 97520
rect 650276 97436 650328 97442
rect 650276 97378 650328 97384
rect 650000 95192 650052 95198
rect 650000 95134 650052 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650012 84697 650040 95134
rect 650288 89593 650316 97378
rect 650552 97300 650604 97306
rect 650552 97242 650604 97248
rect 650274 89584 650330 89593
rect 650274 89519 650330 89528
rect 650564 87145 650592 97242
rect 651300 93566 651328 100014
rect 651852 97442 651880 100014
rect 651840 97436 651892 97442
rect 651840 97378 651892 97384
rect 652588 96490 652616 100014
rect 653324 96626 653352 100014
rect 653968 97986 653996 100014
rect 653956 97980 654008 97986
rect 653956 97922 654008 97928
rect 654796 96966 654824 100014
rect 655210 99770 655238 100028
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655210 99742 655284 99770
rect 655060 97980 655112 97986
rect 655060 97922 655112 97928
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 653312 96620 653364 96626
rect 653312 96562 653364 96568
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652576 96484 652628 96490
rect 652576 96426 652628 96432
rect 651288 93560 651340 93566
rect 651288 93502 651340 93508
rect 650550 87136 650606 87145
rect 650550 87071 650606 87080
rect 652036 86630 652064 96426
rect 652208 95804 652260 95810
rect 652208 95746 652260 95752
rect 652220 86902 652248 95746
rect 653404 95668 653456 95674
rect 653404 95610 653456 95616
rect 652208 86896 652260 86902
rect 652208 86838 652260 86844
rect 652024 86624 652076 86630
rect 652024 86566 652076 86572
rect 653416 86222 653444 95610
rect 655072 94217 655100 97922
rect 655256 96830 655284 99742
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655244 96824 655296 96830
rect 655244 96766 655296 96772
rect 655058 94208 655114 94217
rect 655058 94143 655114 94152
rect 654784 93900 654836 93906
rect 655440 93854 655468 96902
rect 654836 93848 654916 93854
rect 654784 93842 654916 93848
rect 654796 93826 654916 93842
rect 654692 91724 654744 91730
rect 654692 91666 654744 91672
rect 654704 91497 654732 91666
rect 654690 91488 654746 91497
rect 654690 91423 654746 91432
rect 654888 86358 654916 93826
rect 655256 93826 655468 93854
rect 655256 88330 655284 93826
rect 655428 93560 655480 93566
rect 655428 93502 655480 93508
rect 655440 93401 655468 93502
rect 655426 93392 655482 93401
rect 655426 93327 655482 93336
rect 655428 90704 655480 90710
rect 655426 90672 655428 90681
rect 655480 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97238 656848 100014
rect 656808 97232 656860 97238
rect 656808 97174 656860 97180
rect 656164 95804 656216 95810
rect 656164 95746 656216 95752
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86494 656204 95746
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97714 658228 99742
rect 658832 97844 658884 97850
rect 658832 97786 658884 97792
rect 658004 97708 658056 97714
rect 658004 97650 658056 97656
rect 658188 97708 658240 97714
rect 658188 97650 658240 97656
rect 658016 97102 658044 97650
rect 658280 97572 658332 97578
rect 658280 97514 658332 97520
rect 658004 97096 658056 97102
rect 658004 97038 658056 97044
rect 658292 95132 658320 97514
rect 658844 95132 658872 97786
rect 659212 97578 659240 100014
rect 659200 97572 659252 97578
rect 659200 97514 659252 97520
rect 659948 97442 659976 100014
rect 659568 97436 659620 97442
rect 659568 97378 659620 97384
rect 659936 97436 659988 97442
rect 659936 97378 659988 97384
rect 659580 95132 659608 97378
rect 660120 97096 660172 97102
rect 660120 97038 660172 97044
rect 660132 95132 660160 97038
rect 660684 96966 660712 100014
rect 661960 98796 662012 98802
rect 661960 98738 662012 98744
rect 661408 97232 661460 97238
rect 661408 97174 661460 97180
rect 660672 96960 660724 96966
rect 660672 96902 660724 96908
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 660684 95132 660712 96154
rect 661420 95132 661448 97174
rect 661972 95132 662000 98738
rect 663064 97708 663116 97714
rect 663064 97650 663116 97656
rect 662512 96824 662564 96830
rect 662512 96766 662564 96772
rect 662524 95132 662552 96766
rect 663076 95132 663104 97650
rect 663892 97572 663944 97578
rect 663892 97514 663944 97520
rect 663248 96960 663300 96966
rect 663248 96902 663300 96908
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656164 86488 656216 86494
rect 656164 86430 656216 86436
rect 654876 86352 654928 86358
rect 654876 86294 654928 86300
rect 657188 86222 657216 88196
rect 657740 86902 657768 88196
rect 659580 86970 659608 88196
rect 659568 86964 659620 86970
rect 659568 86906 659620 86912
rect 657728 86896 657780 86902
rect 657728 86838 657780 86844
rect 660132 86630 660160 88196
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 660684 86494 660712 88196
rect 661420 86766 661448 88196
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660672 86488 660724 86494
rect 660672 86430 660724 86436
rect 662524 86358 662552 88196
rect 663260 86970 663288 96902
rect 663708 96076 663760 96082
rect 663708 96018 663760 96024
rect 663720 95962 663748 96018
rect 663720 95934 663840 95962
rect 663812 92970 663840 95934
rect 663720 92942 663840 92970
rect 663720 92857 663748 92942
rect 663706 92848 663762 92857
rect 663706 92783 663762 92792
rect 663904 88806 663932 97514
rect 665364 97436 665416 97442
rect 665364 97378 665416 97384
rect 665180 96620 665232 96626
rect 665180 96562 665232 96568
rect 664168 96484 664220 96490
rect 664168 96426 664220 96432
rect 664180 90681 664208 96426
rect 664352 96348 664404 96354
rect 664352 96290 664404 96296
rect 664166 90672 664222 90681
rect 664166 90607 664222 90616
rect 664364 89865 664392 96290
rect 664536 95940 664588 95946
rect 664536 95882 664588 95888
rect 664548 91769 664576 95882
rect 664534 91760 664590 91769
rect 664534 91695 664590 91704
rect 664350 89856 664406 89865
rect 664350 89791 664406 89800
rect 665192 89049 665220 96562
rect 665376 93401 665404 97378
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663248 86964 663300 86970
rect 663248 86906 663300 86912
rect 662512 86352 662564 86358
rect 662512 86294 662564 86300
rect 653404 86216 653456 86222
rect 653404 86158 653456 86164
rect 657176 86216 657228 86222
rect 657176 86158 657228 86164
rect 649998 84688 650054 84697
rect 649998 84623 650054 84632
rect 648894 82240 648950 82249
rect 648894 82175 648950 82184
rect 648712 79348 648764 79354
rect 648712 79290 648764 79296
rect 648724 67153 648752 79290
rect 666572 76566 666600 106082
rect 666834 106043 666890 106052
rect 668136 104417 668164 110735
rect 668398 109304 668454 109313
rect 668398 109239 668454 109248
rect 668122 104408 668178 104417
rect 668122 104343 668178 104352
rect 667938 102776 667994 102785
rect 667938 102711 667994 102720
rect 667952 100026 667980 102711
rect 667940 100020 667992 100026
rect 667940 99962 667992 99968
rect 668136 95849 668164 104343
rect 668412 100162 668440 109239
rect 670712 106146 670740 113146
rect 671540 107817 671568 130863
rect 671724 115841 671752 166903
rect 671908 151881 671936 169895
rect 671894 151872 671950 151881
rect 671894 151807 671950 151816
rect 672092 140457 672120 183495
rect 672644 153105 672672 211126
rect 672814 210352 672870 210361
rect 672814 210287 672870 210296
rect 672630 153096 672686 153105
rect 672630 153031 672686 153040
rect 672078 140448 672134 140457
rect 672078 140383 672134 140392
rect 672354 125624 672410 125633
rect 672354 125559 672410 125568
rect 671710 115832 671766 115841
rect 671710 115767 671766 115776
rect 672368 111353 672396 125559
rect 672828 124137 672856 210287
rect 673012 177993 673040 218470
rect 673196 218385 673224 222166
rect 673366 221912 673422 221921
rect 673366 221847 673422 221856
rect 673182 218376 673238 218385
rect 673182 218311 673238 218320
rect 672998 177984 673054 177993
rect 672998 177919 673054 177928
rect 673380 177313 673408 221847
rect 673564 219881 673592 224926
rect 673550 219872 673606 219881
rect 673550 219807 673606 219816
rect 673550 219464 673606 219473
rect 673550 219399 673606 219408
rect 673366 177304 673422 177313
rect 673366 177239 673422 177248
rect 673366 176896 673422 176905
rect 673366 176831 673422 176840
rect 673182 176080 673238 176089
rect 673182 176015 673238 176024
rect 672998 169144 673054 169153
rect 672998 169079 673054 169088
rect 673012 152561 673040 169079
rect 672998 152552 673054 152561
rect 672998 152487 673054 152496
rect 673196 131345 673224 176015
rect 673380 132161 673408 176831
rect 673564 174865 673592 219399
rect 673748 214305 673776 225383
rect 673918 223680 673974 223689
rect 673918 223615 673974 223624
rect 673734 214296 673790 214305
rect 673734 214231 673790 214240
rect 673932 212945 673960 223615
rect 673918 212936 673974 212945
rect 673918 212871 673974 212880
rect 673734 211168 673790 211177
rect 673734 211103 673790 211112
rect 673748 203969 673776 211103
rect 673918 209672 673974 209681
rect 673918 209607 673974 209616
rect 673734 203960 673790 203969
rect 673734 203895 673790 203904
rect 673932 197441 673960 209607
rect 673918 197432 673974 197441
rect 673918 197367 673974 197376
rect 673550 174856 673606 174865
rect 673550 174791 673606 174800
rect 673918 168736 673974 168745
rect 673918 168671 673974 168680
rect 673932 151065 673960 168671
rect 674116 154601 674144 225406
rect 674300 222329 674328 230030
rect 675852 230036 675904 230042
rect 675852 229978 675904 229984
rect 675114 229936 675170 229945
rect 675170 229906 675892 229922
rect 675170 229900 675904 229906
rect 675170 229894 675852 229900
rect 675114 229871 675170 229880
rect 675852 229842 675904 229848
rect 675114 229256 675170 229265
rect 675114 229191 675170 229200
rect 674838 227080 674894 227089
rect 674838 227015 674894 227024
rect 674470 226536 674526 226545
rect 674470 226471 674526 226480
rect 674484 223689 674512 226471
rect 674470 223680 674526 223689
rect 674470 223615 674526 223624
rect 674470 222728 674526 222737
rect 674470 222663 674526 222672
rect 674286 222320 674342 222329
rect 674286 222255 674342 222264
rect 674484 220130 674512 222663
rect 674852 221649 674880 227015
rect 675128 226386 675156 229191
rect 675128 226358 675340 226386
rect 675022 225856 675078 225865
rect 675022 225791 675078 225800
rect 674838 221640 674894 221649
rect 674838 221575 674894 221584
rect 675036 220561 675064 225791
rect 675022 220552 675078 220561
rect 675022 220487 675078 220496
rect 674654 220280 674710 220289
rect 674654 220215 674710 220224
rect 674300 220102 674512 220130
rect 674300 179489 674328 220102
rect 674470 217424 674526 217433
rect 674470 217359 674526 217368
rect 674484 198257 674512 217359
rect 674470 198248 674526 198257
rect 674470 198183 674526 198192
rect 674286 179480 674342 179489
rect 674286 179415 674342 179424
rect 674668 175681 674696 220215
rect 675114 219872 675170 219881
rect 675114 219807 675170 219816
rect 675128 218929 675156 219807
rect 675114 218920 675170 218929
rect 675114 218855 675170 218864
rect 675312 218226 675340 226358
rect 675666 225176 675722 225185
rect 675666 225111 675722 225120
rect 675482 224360 675538 224369
rect 675482 224295 675538 224304
rect 675496 222194 675524 224295
rect 675036 218198 675340 218226
rect 675404 222166 675524 222194
rect 674838 217832 674894 217841
rect 674838 217767 674894 217776
rect 674852 202065 674880 217767
rect 675036 215393 675064 218198
rect 675206 218104 675262 218113
rect 675404 218090 675432 222166
rect 675262 218062 675432 218090
rect 675206 218039 675262 218048
rect 675206 216200 675262 216209
rect 675206 216135 675262 216144
rect 675022 215384 675078 215393
rect 675022 215319 675078 215328
rect 675220 202874 675248 216135
rect 675680 215937 675708 225111
rect 676232 219994 676260 230415
rect 677046 230208 677102 230217
rect 677046 230143 677102 230152
rect 676772 229900 676824 229906
rect 676772 229842 676824 229848
rect 676402 226264 676458 226273
rect 676402 226199 676458 226208
rect 676416 224954 676444 226199
rect 675864 219966 676260 219994
rect 676324 224926 676444 224954
rect 675666 215928 675722 215937
rect 675666 215863 675722 215872
rect 675864 215294 675892 219966
rect 676034 219872 676090 219881
rect 676324 219858 676352 224926
rect 676496 220108 676548 220114
rect 676496 220050 676548 220056
rect 676090 219830 676352 219858
rect 676034 219807 676090 219816
rect 676220 219700 676272 219706
rect 676220 219642 676272 219648
rect 675496 215266 675892 215294
rect 675496 207369 675524 215266
rect 676036 215144 676088 215150
rect 676034 215112 676036 215121
rect 676088 215112 676090 215121
rect 676034 215047 676090 215056
rect 675852 214872 675904 214878
rect 675666 214840 675722 214849
rect 675722 214820 675852 214826
rect 675722 214814 675904 214820
rect 675722 214798 675892 214814
rect 675666 214775 675722 214784
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 676048 213654 676076 214503
rect 676036 213648 676088 213654
rect 676036 213590 676088 213596
rect 676034 213480 676090 213489
rect 676232 213466 676260 219642
rect 676090 213438 676260 213466
rect 676034 213415 676090 213424
rect 676034 213208 676090 213217
rect 676508 213194 676536 220050
rect 676090 213166 676536 213194
rect 676034 213143 676090 213152
rect 676784 211177 676812 229842
rect 677060 220114 677088 230143
rect 677416 230036 677468 230042
rect 677416 229978 677468 229984
rect 677048 220108 677100 220114
rect 677048 220050 677100 220056
rect 677428 215294 677456 229978
rect 677336 215266 677456 215294
rect 677336 214878 677364 215266
rect 677612 215150 677640 231474
rect 677600 215144 677652 215150
rect 677600 215086 677652 215092
rect 677324 214872 677376 214878
rect 677324 214814 677376 214820
rect 676956 213648 677008 213654
rect 676956 213590 677008 213596
rect 676968 211177 676996 213590
rect 676770 211168 676826 211177
rect 676770 211103 676826 211112
rect 676954 211168 677010 211177
rect 676954 211103 677010 211112
rect 677888 209681 677916 233786
rect 678428 231124 678480 231130
rect 678428 231066 678480 231072
rect 678440 219706 678468 231066
rect 679636 220697 679664 234058
rect 679820 221513 679848 234466
rect 683210 233880 683266 233889
rect 683210 233815 683266 233824
rect 683224 223145 683252 233815
rect 683396 233300 683448 233306
rect 683396 233242 683448 233248
rect 683210 223136 683266 223145
rect 683210 223071 683266 223080
rect 679806 221504 679862 221513
rect 679806 221439 679862 221448
rect 679622 220688 679678 220697
rect 679622 220623 679678 220632
rect 683408 219881 683436 233242
rect 683672 232552 683724 232558
rect 683672 232494 683724 232500
rect 683684 222737 683712 232494
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683670 222728 683726 222737
rect 683670 222663 683726 222672
rect 683394 219872 683450 219881
rect 683394 219807 683450 219816
rect 678428 219700 678480 219706
rect 678428 219642 678480 219648
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 677874 209672 677930 209681
rect 677874 209607 677930 209616
rect 675482 207360 675538 207369
rect 675482 207295 675538 207304
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675036 202846 675248 202874
rect 675312 204666 675418 204694
rect 674838 202056 674894 202065
rect 674838 201991 674894 202000
rect 675036 201906 675064 202846
rect 675312 202722 675340 204666
rect 675482 204232 675538 204241
rect 675482 204167 675538 204176
rect 675496 204035 675524 204167
rect 675312 202694 675524 202722
rect 675496 202609 675524 202694
rect 675482 202600 675538 202609
rect 675482 202535 675538 202544
rect 675496 202065 675524 202195
rect 675482 202056 675538 202065
rect 675482 201991 675538 202000
rect 675036 201878 675432 201906
rect 675114 201648 675170 201657
rect 675404 201620 675432 201878
rect 675114 201583 675170 201592
rect 675128 201022 675156 201583
rect 675128 200994 675418 201022
rect 674930 200832 674986 200841
rect 674930 200767 674986 200776
rect 674944 196058 674972 200767
rect 675758 200696 675814 200705
rect 675758 200631 675814 200640
rect 675298 200560 675354 200569
rect 675298 200495 675354 200504
rect 675312 197282 675340 200495
rect 675772 200328 675800 200631
rect 675482 198248 675538 198257
rect 675482 198183 675538 198192
rect 675496 197880 675524 198183
rect 675404 197282 675432 197336
rect 675312 197254 675432 197282
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 674944 196030 675418 196058
rect 675666 195256 675722 195265
rect 675666 195191 675722 195200
rect 675680 194820 675708 195191
rect 675128 192970 675418 192998
rect 675128 189825 675156 192970
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190369 675340 191950
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675298 190360 675354 190369
rect 675298 190295 675354 190304
rect 675114 189816 675170 189825
rect 675114 189751 675170 189760
rect 675850 181384 675906 181393
rect 675850 181319 675906 181328
rect 675864 178129 675892 181319
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676034 178800 676090 178809
rect 676034 178735 676090 178744
rect 675850 178120 675906 178129
rect 675850 178055 675906 178064
rect 676048 177721 676076 178735
rect 676034 177712 676090 177721
rect 676034 177647 676090 177656
rect 674654 175672 674710 175681
rect 674654 175607 674710 175616
rect 674654 175264 674710 175273
rect 674654 175199 674710 175208
rect 674378 174448 674434 174457
rect 674378 174383 674434 174392
rect 674102 154592 674158 154601
rect 674102 154527 674158 154536
rect 673918 151056 673974 151065
rect 673918 150991 673974 151000
rect 673366 132152 673422 132161
rect 673366 132087 673422 132096
rect 673182 131336 673238 131345
rect 673182 131271 673238 131280
rect 674392 129713 674420 174383
rect 674668 130529 674696 175199
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674852 157593 674880 172751
rect 675022 171184 675078 171193
rect 675022 171119 675078 171128
rect 675036 166994 675064 171119
rect 676232 169674 676260 173182
rect 681002 171592 681058 171601
rect 681002 171527 681058 171536
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 675864 169646 676260 169674
rect 675864 166994 675892 169646
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 674944 166966 675064 166994
rect 675496 166966 675892 166994
rect 674944 164234 674972 166966
rect 674944 164206 675064 164234
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675036 156657 675064 164206
rect 675206 161392 675262 161401
rect 675206 161327 675262 161336
rect 675220 159678 675248 161327
rect 675496 161106 675524 166966
rect 676048 165617 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 681016 162586 681044 171527
rect 675852 162580 675904 162586
rect 675852 162522 675904 162528
rect 681004 162580 681056 162586
rect 681004 162522 681056 162528
rect 675864 161401 675892 162522
rect 675850 161392 675906 161401
rect 675850 161327 675906 161336
rect 675312 161078 675524 161106
rect 675312 160290 675340 161078
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 675758 159352 675814 159361
rect 675758 159287 675814 159296
rect 675772 159052 675800 159287
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675036 156629 675418 156657
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675128 155366 675340 155394
rect 675128 154873 675156 155366
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675312 155230 675432 155258
rect 675114 154864 675170 154873
rect 675114 154799 675170 154808
rect 675312 152850 675418 152878
rect 675312 151609 675340 152850
rect 675482 152552 675538 152561
rect 675482 152487 675538 152496
rect 675496 152320 675524 152487
rect 675482 151872 675538 151881
rect 675482 151807 675538 151816
rect 675496 151675 675524 151807
rect 675298 151600 675354 151609
rect 675298 151535 675354 151544
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675666 150376 675722 150385
rect 675666 150311 675722 150320
rect 675680 149835 675708 150311
rect 675298 149016 675354 149025
rect 675298 148951 675354 148960
rect 675312 146690 675340 148951
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 683302 141400 683358 141409
rect 683302 141335 683358 141344
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 683132 132705 683160 135895
rect 683316 133113 683344 141335
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683302 133104 683358 133113
rect 683302 133039 683358 133048
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674654 130520 674710 130529
rect 674654 130455 674710 130464
rect 676034 130112 676090 130121
rect 676034 130047 676090 130056
rect 674378 129704 674434 129713
rect 674378 129639 674434 129648
rect 674102 129296 674158 129305
rect 674102 129231 674158 129240
rect 673918 125216 673974 125225
rect 673918 125151 673974 125160
rect 673182 124400 673238 124409
rect 673182 124335 673238 124344
rect 672814 124128 672870 124137
rect 672814 124063 672870 124072
rect 672722 122496 672778 122505
rect 672722 122431 672778 122440
rect 672736 112713 672764 122431
rect 672722 112704 672778 112713
rect 672722 112639 672778 112648
rect 672354 111344 672410 111353
rect 672354 111279 672410 111288
rect 673196 110401 673224 124335
rect 673366 123720 673422 123729
rect 673366 123655 673422 123664
rect 673182 110392 673238 110401
rect 673182 110327 673238 110336
rect 671526 107808 671582 107817
rect 671526 107743 671582 107752
rect 673380 106865 673408 123655
rect 673366 106856 673422 106865
rect 673366 106791 673422 106800
rect 670700 106140 670752 106146
rect 670700 106082 670752 106088
rect 673932 104689 673960 125151
rect 674116 111081 674144 129231
rect 676048 128353 676076 130047
rect 674286 128344 674342 128353
rect 674286 128279 674342 128288
rect 676034 128344 676090 128353
rect 676034 128279 676090 128288
rect 674102 111072 674158 111081
rect 674102 111007 674158 111016
rect 673918 104680 673974 104689
rect 673918 104615 673974 104624
rect 674300 102377 674328 128279
rect 679622 128208 679678 128217
rect 679622 128143 679678 128152
rect 678242 127800 678298 127809
rect 678242 127735 678298 127744
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 126032 674710 126041
rect 674654 125967 674710 125976
rect 674470 120048 674526 120057
rect 674470 119983 674526 119992
rect 674484 105822 674512 119983
rect 674668 111466 674696 125967
rect 674852 112010 674880 127599
rect 676218 126984 676274 126993
rect 676218 126919 676274 126928
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 676232 124953 676260 126919
rect 676218 124944 676274 124953
rect 676218 124879 676274 124888
rect 676678 123312 676734 123321
rect 676678 123247 676734 123256
rect 676692 120057 676720 123247
rect 676678 120048 676734 120057
rect 676678 119983 676734 119992
rect 678256 117298 678284 127735
rect 679636 117337 679664 128143
rect 679622 117328 679678 117337
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 678244 117292 678296 117298
rect 679622 117263 679678 117272
rect 678244 117234 678296 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 674668 111438 675418 111466
rect 675390 111344 675446 111353
rect 675390 111279 675446 111288
rect 675404 110772 675432 111279
rect 675114 110392 675170 110401
rect 675114 110327 675170 110336
rect 675128 110174 675156 110327
rect 675128 110146 675418 110174
rect 675206 109032 675262 109041
rect 675206 108967 675262 108976
rect 675220 106502 675248 108967
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675496 106865 675524 107100
rect 675482 106856 675538 106865
rect 675482 106791 675538 106800
rect 675220 106474 675418 106502
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674484 105794 675340 105822
rect 675404 105808 675432 105862
rect 675114 104680 675170 104689
rect 675170 104638 675340 104666
rect 675114 104615 675170 104624
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675666 103184 675722 103193
rect 675666 103119 675722 103128
rect 675680 102816 675708 103119
rect 675758 102504 675814 102513
rect 675758 102439 675814 102448
rect 674286 102368 674342 102377
rect 674286 102303 674342 102312
rect 675772 102136 675800 102439
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668400 100156 668452 100162
rect 668400 100098 668452 100104
rect 668122 95840 668178 95849
rect 668122 95775 668178 95784
rect 666560 76560 666612 76566
rect 666560 76502 666612 76508
rect 648896 75472 648948 75478
rect 648896 75414 648948 75420
rect 648710 67144 648766 67153
rect 648710 67079 648766 67088
rect 648908 62121 648936 75414
rect 662604 75200 662656 75206
rect 662604 75142 662656 75148
rect 648894 62112 648950 62121
rect 648894 62047 648950 62056
rect 647422 57352 647478 57361
rect 647422 57287 647478 57296
rect 625988 54664 626040 54670
rect 625988 54606 626040 54612
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 662418 48512 662474 48521
rect 662418 48447 662474 48456
rect 661590 47789 661646 47798
rect 661590 47724 661646 47733
rect 661604 46510 661632 47724
rect 623044 46504 623096 46510
rect 623044 46446 623096 46452
rect 661592 46504 661644 46510
rect 661592 46446 661644 46452
rect 464342 44296 464398 44305
rect 464342 44231 464398 44240
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 465814 43888 465870 43897
rect 465814 43823 465870 43832
rect 463698 43616 463754 43625
rect 463698 43551 463754 43560
rect 463056 42764 463108 42770
rect 463056 42706 463108 42712
rect 460938 42392 460994 42401
rect 463712 42378 463740 43551
rect 465828 42500 465856 43823
rect 471150 42800 471206 42809
rect 471150 42735 471206 42744
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 463712 42350 464036 42378
rect 460938 42327 460994 42336
rect 471164 42106 471192 42735
rect 518820 42364 518848 42735
rect 662432 42231 662460 48447
rect 662616 47433 662644 75142
rect 662602 47424 662658 47433
rect 662602 47359 662658 47368
rect 662420 42225 662472 42231
rect 662420 42167 662472 42173
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471164 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 427084 41472 427136 41478
rect 427084 41414 427136 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40488 141754 40497
rect 141698 40423 141754 40432
rect 141712 39984 141740 40423
<< via2 >>
rect 428002 1006868 428058 1006904
rect 428002 1006848 428004 1006868
rect 428004 1006848 428056 1006868
rect 428056 1006848 428058 1006868
rect 504546 1006868 504602 1006904
rect 504546 1006848 504548 1006868
rect 504548 1006848 504600 1006868
rect 504600 1006848 504602 1006868
rect 559654 1006868 559710 1006904
rect 559654 1006848 559656 1006868
rect 559656 1006848 559708 1006868
rect 559708 1006848 559710 1006868
rect 428370 1006732 428426 1006768
rect 428370 1006712 428372 1006732
rect 428372 1006712 428424 1006732
rect 428424 1006712 428426 1006732
rect 505374 1006732 505430 1006768
rect 505374 1006712 505376 1006732
rect 505376 1006712 505428 1006732
rect 505428 1006712 505430 1006732
rect 152922 1006596 152978 1006632
rect 152922 1006576 152924 1006596
rect 152924 1006576 152976 1006596
rect 152976 1006576 152978 1006596
rect 308126 1006596 308182 1006632
rect 308126 1006576 308128 1006596
rect 308128 1006576 308180 1006596
rect 308180 1006576 308182 1006596
rect 357714 1006612 357716 1006632
rect 357716 1006612 357768 1006632
rect 357768 1006612 357770 1006632
rect 357714 1006576 357770 1006612
rect 103978 1006460 104034 1006496
rect 103978 1006440 103980 1006460
rect 103980 1006440 104032 1006460
rect 104032 1006440 104034 1006460
rect 74446 996920 74502 996976
rect 74630 996920 74686 996976
rect 80426 995696 80482 995752
rect 84658 995696 84714 995752
rect 87878 995696 87934 995752
rect 88982 995696 89038 995752
rect 89626 995696 89682 995752
rect 77942 995424 77998 995480
rect 77022 995152 77078 995208
rect 42154 968768 42210 968824
rect 41970 967136 42026 967192
rect 42338 966728 42394 966784
rect 43810 968768 43866 968824
rect 43442 966728 43498 966784
rect 42430 964688 42486 964744
rect 42430 963872 42486 963928
rect 42430 963328 42486 963384
rect 42338 963056 42394 963112
rect 41786 962104 41842 962160
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42430 958704 42486 958760
rect 42062 957888 42118 957944
rect 41786 955440 41842 955496
rect 28538 952856 28594 952912
rect 35806 943064 35862 943120
rect 28538 942656 28594 942712
rect 35806 941840 35862 941896
rect 35806 940208 35862 940264
rect 43166 963328 43222 963384
rect 42798 963056 42854 963112
rect 39302 952176 39358 952232
rect 37922 938984 37978 939040
rect 36542 938406 36598 938462
rect 41602 951904 41658 951960
rect 40038 951768 40094 951824
rect 39302 937352 39358 937408
rect 41418 951632 41474 951688
rect 40406 943744 40462 943800
rect 41602 944288 41658 944344
rect 42246 943744 42302 943800
rect 41418 938576 41474 938632
rect 40038 934326 40094 934382
rect 41326 932864 41382 932920
rect 42246 935720 42302 935776
rect 43626 958704 43682 958760
rect 43442 952856 43498 952912
rect 44638 964688 44694 964744
rect 44270 963872 44326 963928
rect 43810 936944 43866 937000
rect 43626 936128 43682 936184
rect 43166 934904 43222 934960
rect 42890 934088 42946 934144
rect 44454 941024 44510 941080
rect 44270 933680 44326 933736
rect 43626 933272 43682 933328
rect 42246 911920 42302 911976
rect 41786 911784 41842 911840
rect 42936 892254 42992 892256
rect 42936 892202 42938 892254
rect 42938 892202 42990 892254
rect 42990 892202 42992 892254
rect 42936 892200 42992 892202
rect 43074 891948 43130 891984
rect 43074 891928 43076 891948
rect 43076 891928 43128 891948
rect 43128 891928 43130 891948
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 35806 817264 35862 817320
rect 35806 816448 35862 816504
rect 35806 814816 35862 814872
rect 42062 884584 42118 884640
rect 43074 815224 43130 815280
rect 41142 813184 41198 813240
rect 40958 812368 41014 812424
rect 39302 811552 39358 811608
rect 33046 811144 33102 811200
rect 41326 812776 41382 812832
rect 42522 808968 42578 809024
rect 41786 808288 41842 808344
rect 41142 805568 41198 805624
rect 40958 805296 41014 805352
rect 42246 806656 42302 806712
rect 41786 805024 41842 805080
rect 41602 801660 41604 801680
rect 41604 801660 41656 801680
rect 41656 801660 41658 801680
rect 41602 801624 41658 801660
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42522 804344 42578 804400
rect 42706 801624 42762 801680
rect 42522 799584 42578 799640
rect 42522 796728 42578 796784
rect 41970 796048 42026 796104
rect 42246 796048 42302 796104
rect 42430 794280 42486 794336
rect 42246 792512 42302 792568
rect 42614 792240 42670 792296
rect 42430 791696 42486 791752
rect 42154 790064 42210 790120
rect 42614 790064 42670 790120
rect 41786 788568 41842 788624
rect 42706 788568 42762 788624
rect 42246 787888 42302 787944
rect 42062 786392 42118 786448
rect 41786 785576 41842 785632
rect 35806 773472 35862 773528
rect 43258 810328 43314 810384
rect 43442 807608 43498 807664
rect 43258 791696 43314 791752
rect 43074 772384 43130 772440
rect 35346 769392 35402 769448
rect 35530 769004 35586 769040
rect 35530 768984 35532 769004
rect 35532 768984 35584 769004
rect 35584 768984 35586 769004
rect 35806 768984 35862 769040
rect 35622 768168 35678 768224
rect 31022 767760 31078 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 35806 763292 35862 763328
rect 35806 763272 35808 763292
rect 35808 763272 35860 763292
rect 35860 763272 35862 763292
rect 36542 759056 36598 759112
rect 42798 766672 42854 766728
rect 41326 765312 41382 765368
rect 42614 765312 42670 765368
rect 40590 764088 40646 764144
rect 42522 764088 42578 764144
rect 40406 763680 40462 763736
rect 42338 763680 42394 763736
rect 40590 758396 40646 758432
rect 40590 758376 40592 758396
rect 40592 758376 40644 758396
rect 40644 758376 40646 758396
rect 42338 758784 42394 758840
rect 42338 758376 42394 758432
rect 39302 757696 39358 757752
rect 41786 757016 41842 757072
rect 41878 755384 41934 755440
rect 42154 754568 42210 754624
rect 42062 754160 42118 754216
rect 42338 753888 42394 753944
rect 42154 753344 42210 753400
rect 41970 752936 42026 752992
rect 42430 752392 42486 752448
rect 43350 764632 43406 764688
rect 43166 763000 43222 763056
rect 42890 752120 42946 752176
rect 42154 751712 42210 751768
rect 41786 751032 41842 751088
rect 41786 750352 41842 750408
rect 42154 749672 42210 749728
rect 42062 749128 42118 749184
rect 42154 746816 42210 746872
rect 42890 749672 42946 749728
rect 42154 745456 42210 745512
rect 42338 744912 42394 744968
rect 42706 745184 42762 745240
rect 42798 744368 42854 744424
rect 42890 742736 42946 742792
rect 43350 753888 43406 753944
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 33782 725192 33838 725248
rect 31666 724376 31722 724432
rect 36542 724784 36598 724840
rect 34518 723968 34574 724024
rect 40682 723152 40738 723208
rect 38750 720296 38806 720352
rect 31666 715400 31722 715456
rect 40314 715672 40370 715728
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41694 715128 41750 715184
rect 42062 715672 42118 715728
rect 41878 714584 41934 714640
rect 42706 715128 42762 715184
rect 42430 714584 42486 714640
rect 42062 714312 42118 714368
rect 38750 714176 38806 714232
rect 40682 714176 40738 714232
rect 41418 714176 41474 714232
rect 41786 713496 41842 713552
rect 42246 713224 42302 713280
rect 41786 712136 41842 712192
rect 42246 711048 42302 711104
rect 42706 714040 42762 714096
rect 42614 713224 42670 713280
rect 41786 709824 41842 709880
rect 42062 709008 42118 709064
rect 41786 708464 41842 708520
rect 42062 707784 42118 707840
rect 42246 706696 42302 706752
rect 41970 706424 42026 706480
rect 42246 705200 42302 705256
rect 42246 704520 42302 704576
rect 42154 703432 42210 703488
rect 42706 709960 42762 710016
rect 42062 702752 42118 702808
rect 42706 702752 42762 702808
rect 42614 702344 42670 702400
rect 41786 700440 41842 700496
rect 41786 699760 41842 699816
rect 35622 691328 35678 691384
rect 41418 689288 41474 689344
rect 35806 687656 35862 687712
rect 35622 687248 35678 687304
rect 35806 683576 35862 683632
rect 35806 683188 35862 683224
rect 35806 683168 35808 683188
rect 35808 683168 35860 683188
rect 35860 683168 35862 683188
rect 35438 682760 35494 682816
rect 35622 682352 35678 682408
rect 35806 681980 35808 682000
rect 35808 681980 35860 682000
rect 35860 681980 35862 682000
rect 35806 681944 35862 681980
rect 32402 681536 32458 681592
rect 31022 681128 31078 681184
rect 35622 680720 35678 680776
rect 37186 677048 37242 677104
rect 31022 671336 31078 671392
rect 41694 681844 41696 681864
rect 41696 681844 41748 681864
rect 41748 681844 41750 681864
rect 41694 681808 41750 681844
rect 42614 681808 42670 681864
rect 41786 677592 41842 677648
rect 40958 675960 41014 676016
rect 42890 679904 42946 679960
rect 42522 673512 42578 673568
rect 40590 673140 40592 673160
rect 40592 673140 40644 673160
rect 40644 673140 40646 673160
rect 40590 673104 40646 673140
rect 42338 673104 42394 673160
rect 39670 671880 39726 671936
rect 40130 670964 40132 670984
rect 40132 670964 40184 670984
rect 40184 670964 40186 670984
rect 40130 670928 40186 670964
rect 42338 671880 42394 671936
rect 42154 670928 42210 670984
rect 42062 668208 42118 668264
rect 42246 667800 42302 667856
rect 42246 666984 42302 667040
rect 42062 666576 42118 666632
rect 41786 665352 41842 665408
rect 41786 664128 41842 664184
rect 42338 663312 42394 663368
rect 42430 662904 42486 662960
rect 42062 662768 42118 662824
rect 42154 659776 42210 659832
rect 42890 666576 42946 666632
rect 42154 658960 42210 659016
rect 42706 658960 42762 659016
rect 42614 658552 42670 658608
rect 42430 658280 42486 658336
rect 41970 657328 42026 657384
rect 42614 655424 42670 655480
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35346 639784 35402 639840
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 35806 638560 35862 638616
rect 33782 638152 33838 638208
rect 40038 638560 40094 638616
rect 41786 638152 41842 638208
rect 41786 637540 41842 637596
rect 36542 630672 36598 630728
rect 41418 629992 41474 630048
rect 42890 636248 42946 636304
rect 42522 633800 42578 633856
rect 42062 625776 42118 625832
rect 42706 629992 42762 630048
rect 42522 625776 42578 625832
rect 42430 624144 42486 624200
rect 42246 623736 42302 623792
rect 42430 623736 42486 623792
rect 42062 623328 42118 623384
rect 42062 620880 42118 620936
rect 42798 623736 42854 623792
rect 42246 620064 42302 620120
rect 42706 619792 42762 619848
rect 42522 619520 42578 619576
rect 42522 618704 42578 618760
rect 42430 615984 42486 616040
rect 41786 615712 41842 615768
rect 42154 613536 42210 613592
rect 41786 612720 41842 612776
rect 43350 633392 43406 633448
rect 43074 612312 43130 612368
rect 43810 932048 43866 932104
rect 44086 892764 44142 892800
rect 44086 892744 44088 892764
rect 44088 892744 44140 892764
rect 44140 892744 44142 892764
rect 44086 892472 44142 892528
rect 46294 943472 46350 943528
rect 44822 941432 44878 941488
rect 44638 935312 44694 935368
rect 48962 942248 49018 942304
rect 50342 940616 50398 940672
rect 51722 939800 51778 939856
rect 47582 891928 47638 891984
rect 44914 816040 44970 816096
rect 44454 815632 44510 815688
rect 44638 814408 44694 814464
rect 44178 807880 44234 807936
rect 43994 806248 44050 806304
rect 44178 796320 44234 796376
rect 44178 772792 44234 772848
rect 44454 771976 44510 772032
rect 44178 730088 44234 730144
rect 44270 729680 44326 729736
rect 45466 813592 45522 813648
rect 45098 810736 45154 810792
rect 44822 809512 44878 809568
rect 44822 797680 44878 797736
rect 44638 771568 44694 771624
rect 44638 771160 44694 771216
rect 44454 729272 44510 729328
rect 44178 722744 44234 722800
rect 44178 707784 44234 707840
rect 45282 809920 45338 809976
rect 45282 792240 45338 792296
rect 45190 786392 45246 786448
rect 45006 773200 45062 773256
rect 45466 770752 45522 770808
rect 45006 770344 45062 770400
rect 44822 731312 44878 731368
rect 44638 728456 44694 728512
rect 44822 728048 44878 728104
rect 44638 727232 44694 727288
rect 44362 686840 44418 686896
rect 44362 686432 44418 686488
rect 44178 684800 44234 684856
rect 45190 766264 45246 766320
rect 45190 754840 45246 754896
rect 46938 764360 46994 764416
rect 46202 754160 46258 754216
rect 45190 728864 45246 728920
rect 45006 727640 45062 727696
rect 45006 723560 45062 723616
rect 45006 705200 45062 705256
rect 45558 721112 45614 721168
rect 45190 686024 45246 686080
rect 45190 685616 45246 685672
rect 44822 685208 44878 685264
rect 44638 684392 44694 684448
rect 45006 683984 45062 684040
rect 44546 680312 44602 680368
rect 44730 679496 44786 679552
rect 44730 666984 44786 667040
rect 44546 662904 44602 662960
rect 44362 643592 44418 643648
rect 44822 643320 44878 643376
rect 44638 642504 44694 642560
rect 44178 642232 44234 642288
rect 44270 636520 44326 636576
rect 44454 635704 44510 635760
rect 44270 623328 44326 623384
rect 44454 620064 44510 620120
rect 43718 612332 43774 612368
rect 43718 612312 43720 612332
rect 43720 612312 43772 612332
rect 43772 612312 43774 612332
rect 43350 610952 43406 611008
rect 44086 610952 44142 611008
rect 44270 610972 44326 611008
rect 44270 610952 44272 610972
rect 44272 610952 44324 610972
rect 44324 610952 44326 610972
rect 45190 643048 45246 643104
rect 45006 641416 45062 641472
rect 45374 641144 45430 641200
rect 45190 640872 45246 640928
rect 45006 635296 45062 635352
rect 45006 620880 45062 620936
rect 44822 600480 44878 600536
rect 44822 600072 44878 600128
rect 44638 599664 44694 599720
rect 44638 598440 44694 598496
rect 42982 596944 43038 597000
rect 41326 596808 41382 596864
rect 41142 595992 41198 596048
rect 33046 595584 33102 595640
rect 31022 594360 31078 594416
rect 35162 595176 35218 595232
rect 40682 594768 40738 594824
rect 39946 590688 40002 590744
rect 40498 589600 40554 589656
rect 39946 585928 40002 585984
rect 40130 584840 40186 584896
rect 41694 594496 41750 594552
rect 41786 593544 41842 593600
rect 39394 584568 39450 584624
rect 40682 584568 40738 584624
rect 41786 593136 41842 593192
rect 41786 592728 41842 592784
rect 41878 592320 41934 592376
rect 41418 589464 41474 589520
rect 42522 594496 42578 594552
rect 42798 593952 42854 594008
rect 41878 589328 41934 589384
rect 42338 585928 42394 585984
rect 41786 584296 41842 584352
rect 42430 581984 42486 582040
rect 41970 580760 42026 580816
rect 42246 580760 42302 580816
rect 41970 580216 42026 580272
rect 41786 578176 41842 578232
rect 41786 577496 41842 577552
rect 42338 576680 42394 576736
rect 42062 576544 42118 576600
rect 42154 573824 42210 573880
rect 42706 581304 42762 581360
rect 42706 576680 42762 576736
rect 42706 573824 42762 573880
rect 42614 573280 42670 573336
rect 42522 572056 42578 572112
rect 41786 570152 41842 570208
rect 42338 569200 42394 569256
rect 41326 558048 41382 558104
rect 41326 554804 41382 554840
rect 41326 554784 41328 554804
rect 41328 554784 41380 554804
rect 41380 554784 41382 554804
rect 44178 591912 44234 591968
rect 43442 590280 43498 590336
rect 32402 551928 32458 551984
rect 31758 548086 31814 548142
rect 41234 553352 41290 553408
rect 41142 552744 41198 552800
rect 42890 552336 42946 552392
rect 41786 551928 41842 551984
rect 41786 551112 41842 551168
rect 40774 550296 40830 550352
rect 41234 549480 41290 549536
rect 41234 548140 41290 548142
rect 41234 548088 41236 548140
rect 41236 548088 41288 548140
rect 41288 548088 41290 548140
rect 41234 548086 41290 548088
rect 40774 545672 40830 545728
rect 40590 545400 40646 545456
rect 41878 550160 41934 550216
rect 41786 549888 41842 549944
rect 41694 548140 41750 548176
rect 41694 548120 41696 548140
rect 41696 548120 41748 548140
rect 41748 548120 41750 548140
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42614 540232 42670 540288
rect 42522 537376 42578 537432
rect 41786 536968 41842 537024
rect 42062 536968 42118 537024
rect 41786 535200 41842 535256
rect 42154 533840 42210 533896
rect 43074 550160 43130 550216
rect 42890 534112 42946 534168
rect 42522 532616 42578 532672
rect 42430 529760 42486 529816
rect 42246 529488 42302 529544
rect 41878 529352 41934 529408
rect 42706 529080 42762 529136
rect 41326 425992 41382 426048
rect 40958 425584 41014 425640
rect 33690 424360 33746 424416
rect 41326 423952 41382 424008
rect 41786 423816 41842 423872
rect 41326 422340 41382 422376
rect 41326 422320 41328 422340
rect 41328 422320 41380 422340
rect 41380 422320 41382 422340
rect 41786 422320 41842 422376
rect 41786 421232 41842 421288
rect 41326 421096 41382 421152
rect 41786 420960 41842 421016
rect 42798 423816 42854 423872
rect 42154 422728 42210 422784
rect 42338 421912 42394 421968
rect 42154 418784 42210 418840
rect 42522 419872 42578 419928
rect 42338 418512 42394 418568
rect 42062 411848 42118 411904
rect 42614 411848 42670 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42430 407088 42486 407144
rect 42430 406816 42486 406872
rect 41786 406272 41842 406328
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 42430 399744 42486 399800
rect 43166 422320 43222 422376
rect 42982 420960 43038 421016
rect 42982 407768 43038 407824
rect 43166 407088 43222 407144
rect 41786 398792 41842 398848
rect 41142 387116 41198 387152
rect 41142 387096 41144 387116
rect 41144 387096 41196 387116
rect 41196 387096 41198 387116
rect 41878 386960 41934 387016
rect 41326 386688 41382 386744
rect 41510 386688 41566 386744
rect 41326 383016 41382 383072
rect 41142 382608 41198 382664
rect 40222 382200 40278 382256
rect 40038 381792 40094 381848
rect 35806 379344 35862 379400
rect 41326 380976 41382 381032
rect 41694 379344 41750 379400
rect 41326 378528 41382 378584
rect 42338 378528 42394 378584
rect 40222 376896 40278 376952
rect 35806 376488 35862 376544
rect 40038 376488 40094 376544
rect 28906 376080 28962 376136
rect 39578 375672 39634 375728
rect 41694 371884 41750 371920
rect 41694 371864 41696 371884
rect 41696 371864 41748 371884
rect 41748 371864 41750 371884
rect 41786 368600 41842 368656
rect 42430 366968 42486 367024
rect 42430 365744 42486 365800
rect 41786 364248 41842 364304
rect 41786 363568 41842 363624
rect 41878 362888 41934 362944
rect 42430 361528 42486 361584
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 42062 358672 42118 358728
rect 42430 357312 42486 357368
rect 44178 581032 44234 581088
rect 45006 599256 45062 599312
rect 44822 557232 44878 557288
rect 46110 719888 46166 719944
rect 45742 676640 45798 676696
rect 45926 637744 45982 637800
rect 45926 613536 45982 613592
rect 46294 636928 46350 636984
rect 46478 626592 46534 626648
rect 46478 624144 46534 624200
rect 46294 619520 46350 619576
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47582 712136 47638 712192
rect 47214 677864 47270 677920
rect 53286 892472 53342 892528
rect 85026 994880 85082 994936
rect 90270 995424 90326 995480
rect 92662 995696 92718 995752
rect 92478 995424 92534 995480
rect 86314 995152 86370 995208
rect 92662 994880 92718 994936
rect 93490 997192 93546 997248
rect 101126 1006324 101182 1006360
rect 101126 1006304 101128 1006324
rect 101128 1006304 101180 1006324
rect 101180 1006304 101182 1006324
rect 94502 996920 94558 996976
rect 98274 1006188 98330 1006224
rect 98274 1006168 98276 1006188
rect 98276 1006168 98328 1006188
rect 98328 1006168 98330 1006188
rect 107658 1006188 107714 1006224
rect 107658 1006168 107660 1006188
rect 107660 1006168 107712 1006188
rect 107712 1006168 107714 1006188
rect 99470 1006052 99526 1006088
rect 99470 1006032 99472 1006052
rect 99472 1006032 99524 1006052
rect 99524 1006032 99526 1006052
rect 104806 1006052 104862 1006088
rect 104806 1006032 104808 1006052
rect 104808 1006032 104860 1006052
rect 104860 1006032 104862 1006052
rect 108486 1006052 108542 1006088
rect 108486 1006032 108488 1006052
rect 108488 1006032 108540 1006052
rect 108540 1006032 108542 1006052
rect 101494 1002516 101550 1002552
rect 101494 1002496 101496 1002516
rect 101496 1002496 101548 1002516
rect 101548 1002496 101550 1002516
rect 94686 996648 94742 996704
rect 93306 996376 93362 996432
rect 93306 995968 93362 996024
rect 93122 995152 93178 995208
rect 86038 994336 86094 994392
rect 92846 994336 92902 994392
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 99102 1002244 99158 1002280
rect 99102 1002224 99104 1002244
rect 99104 1002224 99156 1002244
rect 99156 1002224 99158 1002244
rect 100298 1002108 100354 1002144
rect 100298 1002088 100300 1002108
rect 100300 1002088 100352 1002108
rect 100352 1002088 100354 1002108
rect 101954 1002244 102010 1002280
rect 101954 1002224 101956 1002244
rect 101956 1002224 102008 1002244
rect 102008 1002224 102010 1002244
rect 101126 1001972 101182 1002008
rect 101126 1001952 101128 1001972
rect 101128 1001952 101180 1001972
rect 101180 1001952 101182 1001972
rect 102322 1001972 102378 1002008
rect 102322 1001952 102324 1001972
rect 102324 1001952 102376 1001972
rect 102376 1001952 102378 1001972
rect 101402 995152 101458 995208
rect 104806 1003892 104808 1003912
rect 104808 1003892 104860 1003912
rect 104860 1003892 104862 1003912
rect 104806 1003856 104862 1003892
rect 106830 1002652 106886 1002688
rect 106830 1002632 106832 1002652
rect 106832 1002632 106884 1002652
rect 106884 1002632 106886 1002652
rect 108026 1002516 108082 1002552
rect 108026 1002496 108028 1002516
rect 108028 1002496 108080 1002516
rect 108080 1002496 108082 1002516
rect 103150 1002380 103206 1002416
rect 103150 1002360 103152 1002380
rect 103152 1002360 103204 1002380
rect 103204 1002360 103206 1002380
rect 106830 1002380 106886 1002416
rect 106830 1002360 106832 1002380
rect 106832 1002360 106884 1002380
rect 106884 1002360 106886 1002380
rect 106002 1002244 106058 1002280
rect 106002 1002224 106004 1002244
rect 106004 1002224 106056 1002244
rect 106056 1002224 106058 1002244
rect 108854 1002244 108910 1002280
rect 108854 1002224 108856 1002244
rect 108856 1002224 108908 1002244
rect 108908 1002224 108910 1002244
rect 103150 1002108 103206 1002144
rect 103150 1002088 103152 1002108
rect 103152 1002088 103204 1002108
rect 103204 1002088 103206 1002108
rect 105634 1002108 105690 1002144
rect 105634 1002088 105636 1002108
rect 105636 1002088 105688 1002108
rect 105688 1002088 105690 1002108
rect 103978 1001952 104034 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 108854 1001972 108910 1002008
rect 108854 1001952 108856 1001972
rect 108856 1001952 108908 1001972
rect 108908 1001952 108910 1001972
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 117226 997192 117282 997248
rect 116306 996920 116362 996976
rect 126242 996240 126298 996296
rect 143998 996920 144054 996976
rect 131854 995696 131910 995752
rect 132958 995696 133014 995752
rect 140410 995696 140466 995752
rect 141054 995696 141110 995752
rect 144182 995832 144238 995888
rect 141790 995560 141846 995616
rect 124862 995016 124918 995072
rect 132406 995288 132462 995344
rect 132130 994744 132186 994800
rect 137374 995424 137430 995480
rect 135902 994336 135958 994392
rect 137558 994084 137614 994120
rect 137558 994064 137560 994084
rect 137560 994064 137612 994084
rect 137612 994064 137614 994084
rect 137742 993928 137798 993984
rect 144826 997192 144882 997248
rect 144826 996532 144882 996568
rect 144826 996512 144828 996532
rect 144828 996512 144880 996532
rect 144880 996512 144882 996532
rect 144366 994744 144422 994800
rect 144550 994744 144606 994800
rect 142158 994472 142214 994528
rect 141974 994336 142030 994392
rect 133142 993656 133198 993712
rect 139214 993656 139270 993712
rect 139398 993656 139454 993712
rect 152094 1006460 152150 1006496
rect 152094 1006440 152096 1006460
rect 152096 1006440 152148 1006460
rect 152148 1006440 152150 1006460
rect 157430 1006460 157486 1006496
rect 157430 1006440 157432 1006460
rect 157432 1006440 157484 1006460
rect 157484 1006440 157486 1006460
rect 158258 1006324 158314 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 151266 1006188 151322 1006224
rect 151266 1006168 151268 1006188
rect 151268 1006168 151320 1006188
rect 151320 1006168 151322 1006188
rect 153750 1006188 153806 1006224
rect 153750 1006168 153752 1006188
rect 153752 1006168 153804 1006188
rect 153804 1006168 153806 1006188
rect 160282 1006188 160338 1006224
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 147126 1006032 147182 1006088
rect 148874 1006052 148930 1006088
rect 148874 1006032 148876 1006052
rect 148876 1006032 148928 1006052
rect 148928 1006032 148930 1006052
rect 145746 996104 145802 996160
rect 142342 993928 142398 993984
rect 145562 993928 145618 993984
rect 142158 993656 142214 993712
rect 142342 993384 142398 993440
rect 150070 1006052 150126 1006088
rect 150070 1006032 150072 1006052
rect 150072 1006032 150124 1006052
rect 150124 1006032 150126 1006052
rect 159454 1006052 159510 1006088
rect 159454 1006032 159456 1006052
rect 159456 1006032 159508 1006052
rect 159508 1006032 159510 1006052
rect 152922 1005100 152978 1005136
rect 152922 1005080 152924 1005100
rect 152924 1005080 152976 1005100
rect 152976 1005080 152978 1005100
rect 158626 1005100 158682 1005136
rect 158626 1005080 158628 1005100
rect 158628 1005080 158680 1005100
rect 158680 1005080 158682 1005100
rect 147126 995560 147182 995616
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 153750 1004964 153806 1005000
rect 153750 1004944 153752 1004964
rect 153752 1004944 153804 1004964
rect 153804 1004944 153806 1004964
rect 150898 1002380 150954 1002416
rect 150898 1002360 150900 1002380
rect 150900 1002360 150952 1002380
rect 150952 1002360 150954 1002380
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 149886 994744 149942 994800
rect 151726 1004828 151782 1004864
rect 151726 1004808 151728 1004828
rect 151728 1004808 151780 1004828
rect 151780 1004808 151782 1004828
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 154118 1004692 154174 1004728
rect 154118 1004672 154120 1004692
rect 154120 1004672 154172 1004692
rect 154172 1004672 154174 1004692
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 156602 1002244 156658 1002280
rect 156602 1002224 156604 1002244
rect 156604 1002224 156656 1002244
rect 156656 1002224 156658 1002244
rect 148506 994200 148562 994256
rect 154578 1001972 154634 1002008
rect 154578 1001952 154580 1001972
rect 154580 1001952 154632 1001972
rect 154632 1001952 154634 1001972
rect 154946 1001972 155002 1002008
rect 154946 1001952 154948 1001972
rect 154948 1001952 155000 1001972
rect 155000 1001952 155002 1001972
rect 155774 1001952 155830 1002008
rect 155130 995560 155186 995616
rect 155130 995016 155186 995072
rect 156602 1001952 156658 1002008
rect 157798 1001972 157854 1002008
rect 157798 1001952 157800 1001972
rect 157800 1001952 157852 1001972
rect 157852 1001952 157854 1001972
rect 157338 994472 157394 994528
rect 152462 993928 152518 993984
rect 170310 997192 170366 997248
rect 210054 1006324 210110 1006360
rect 210054 1006304 210056 1006324
rect 210056 1006304 210108 1006324
rect 210108 1006304 210110 1006324
rect 254122 1006324 254178 1006360
rect 254122 1006304 254124 1006324
rect 254124 1006304 254176 1006324
rect 254176 1006304 254178 1006324
rect 172334 996240 172390 996296
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 195058 996920 195114 996976
rect 183834 995696 183890 995752
rect 188802 995560 188858 995616
rect 190458 995560 190514 995616
rect 175922 995016 175978 995072
rect 180154 994744 180210 994800
rect 183282 994200 183338 994256
rect 188158 995288 188214 995344
rect 187606 994472 187662 994528
rect 192482 995288 192538 995344
rect 192942 995324 192944 995344
rect 192944 995324 192996 995344
rect 192996 995324 192998 995344
rect 192942 995288 192998 995324
rect 195702 996376 195758 996432
rect 195886 995288 195942 995344
rect 202694 1001972 202750 1002008
rect 202694 1001952 202696 1001972
rect 202696 1001952 202748 1001972
rect 202748 1001952 202750 1001972
rect 200670 997908 200672 997928
rect 200672 997908 200724 997928
rect 200724 997908 200726 997928
rect 200670 997872 200726 997908
rect 202694 998300 202750 998336
rect 202694 998280 202696 998300
rect 202696 998280 202748 998300
rect 202748 998280 202750 998300
rect 201866 998044 201868 998064
rect 201868 998044 201920 998064
rect 201920 998044 201922 998064
rect 201866 998008 201922 998044
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 200762 995560 200818 995616
rect 202326 995832 202382 995888
rect 203522 1002108 203578 1002144
rect 203522 1002088 203524 1002108
rect 203524 1002088 203576 1002108
rect 203576 1002088 203578 1002108
rect 203890 998572 203946 998608
rect 203890 998552 203892 998572
rect 203892 998552 203944 998572
rect 203944 998552 203946 998572
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 204718 998028 204774 998064
rect 204718 998008 204720 998028
rect 204720 998008 204772 998028
rect 204772 998008 204774 998028
rect 203522 997892 203578 997928
rect 203522 997872 203524 997892
rect 203524 997872 203576 997892
rect 203576 997872 203578 997892
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 208398 1006052 208454 1006088
rect 208398 1006032 208400 1006052
rect 208400 1006032 208452 1006052
rect 208452 1006032 208454 1006052
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 207570 1004828 207626 1004864
rect 207570 1004808 207572 1004828
rect 207572 1004808 207624 1004828
rect 207624 1004808 207626 1004828
rect 211250 1004828 211306 1004864
rect 211250 1004808 211252 1004828
rect 211252 1004808 211304 1004828
rect 211304 1004808 211306 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002244 206430 1002280
rect 206374 1002224 206376 1002244
rect 206376 1002224 206428 1002244
rect 206428 1002224 206430 1002244
rect 206742 1002108 206798 1002144
rect 206742 1002088 206744 1002108
rect 206744 1002088 206796 1002108
rect 206796 1002088 206798 1002108
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 205546 998164 205602 998200
rect 205546 998144 205548 998164
rect 205548 998144 205600 998164
rect 205600 998144 205602 998164
rect 207202 1001952 207258 1002008
rect 207570 1001972 207626 1002008
rect 207570 1001952 207572 1001972
rect 207572 1001952 207624 1001972
rect 207624 1001952 207626 1001972
rect 207018 994744 207074 994800
rect 203338 994472 203394 994528
rect 196806 993928 196862 993984
rect 210882 1002380 210938 1002416
rect 210882 1002360 210884 1002380
rect 210884 1002360 210936 1002380
rect 210936 1002360 210938 1002380
rect 210882 1002108 210938 1002144
rect 210882 1002088 210884 1002108
rect 210884 1002088 210936 1002108
rect 210936 1002088 210938 1002108
rect 212538 1004692 212594 1004728
rect 212538 1004672 212540 1004692
rect 212540 1004672 212592 1004692
rect 212592 1004672 212594 1004692
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 208398 994200 208454 994256
rect 229006 997736 229062 997792
rect 229374 997736 229430 997792
rect 228822 997192 228878 997248
rect 229190 997192 229246 997248
rect 239586 995696 239642 995752
rect 242070 995696 242126 995752
rect 235262 994472 235318 994528
rect 236550 994744 236606 994800
rect 240046 995424 240102 995480
rect 243266 995424 243322 995480
rect 243910 995152 243966 995208
rect 247038 995696 247094 995752
rect 240874 994200 240930 994256
rect 247406 995152 247462 995208
rect 246762 994472 246818 994528
rect 255318 1006188 255374 1006224
rect 255318 1006168 255320 1006188
rect 255320 1006168 255372 1006188
rect 255372 1006168 255374 1006188
rect 261850 1006188 261906 1006224
rect 261850 1006168 261852 1006188
rect 261852 1006168 261904 1006188
rect 261904 1006168 261906 1006188
rect 252466 1006052 252522 1006088
rect 252466 1006032 252468 1006052
rect 252468 1006032 252520 1006052
rect 252520 1006032 252522 1006052
rect 260194 1006052 260250 1006088
rect 260194 1006032 260196 1006052
rect 260196 1006032 260248 1006052
rect 260248 1006032 260250 1006052
rect 263046 1005100 263102 1005136
rect 263046 1005080 263048 1005100
rect 263048 1005080 263100 1005100
rect 263100 1005080 263102 1005100
rect 256146 1002652 256202 1002688
rect 256146 1002632 256148 1002652
rect 256148 1002632 256200 1002652
rect 256200 1002632 256202 1002652
rect 261022 1002652 261078 1002688
rect 261022 1002632 261024 1002652
rect 261024 1002632 261076 1002652
rect 261076 1002632 261078 1002652
rect 250442 997192 250498 997248
rect 249246 995968 249302 996024
rect 252466 997892 252522 997928
rect 252466 997872 252468 997892
rect 252468 997872 252520 997892
rect 252520 997872 252522 997892
rect 251638 996240 251694 996296
rect 251454 994744 251510 994800
rect 249062 994200 249118 994256
rect 253294 998028 253350 998064
rect 253294 998008 253296 998028
rect 253296 998008 253348 998028
rect 253348 998008 253350 998028
rect 255318 1002516 255374 1002552
rect 255318 1002496 255320 1002516
rect 255320 1002496 255372 1002516
rect 255372 1002496 255374 1002516
rect 256146 1002380 256202 1002416
rect 256146 1002360 256148 1002380
rect 256148 1002360 256200 1002380
rect 256200 1002360 256202 1002380
rect 261022 1002396 261024 1002416
rect 261024 1002396 261076 1002416
rect 261076 1002396 261078 1002416
rect 261022 1002360 261078 1002396
rect 254490 1002244 254546 1002280
rect 254490 1002224 254492 1002244
rect 254492 1002224 254544 1002244
rect 254544 1002224 254546 1002244
rect 262678 1002260 262680 1002280
rect 262680 1002260 262732 1002280
rect 262732 1002260 262734 1002280
rect 262678 1002224 262734 1002260
rect 263506 1001988 263508 1002008
rect 263508 1001988 263560 1002008
rect 263560 1001988 263562 1002008
rect 263506 1001952 263562 1001988
rect 258170 999132 258172 999152
rect 258172 999132 258224 999152
rect 258224 999132 258226 999152
rect 253662 998164 253718 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 256514 997908 256516 997928
rect 256516 997908 256568 997928
rect 256568 997908 256570 997928
rect 256514 997872 256570 997908
rect 258170 999096 258226 999132
rect 258998 998436 259054 998472
rect 258998 998416 259000 998436
rect 259000 998416 259052 998436
rect 259052 998416 259054 998436
rect 257342 998164 257398 998200
rect 257342 998144 257344 998164
rect 257344 998144 257396 998164
rect 257396 998144 257398 998164
rect 258998 997908 259000 997928
rect 259000 997908 259052 997928
rect 259052 997908 259054 997928
rect 256974 997772 256976 997792
rect 256976 997772 257028 997792
rect 257028 997772 257030 997792
rect 256974 997736 257030 997772
rect 258998 997872 259054 997908
rect 259826 997908 259828 997928
rect 259828 997908 259880 997928
rect 259880 997908 259882 997928
rect 259826 997872 259882 997908
rect 258170 997772 258172 997792
rect 258172 997772 258224 997792
rect 258224 997772 258226 997792
rect 258170 997736 258226 997772
rect 260194 997772 260196 997792
rect 260196 997772 260248 997792
rect 260248 997772 260250 997792
rect 260194 997736 260250 997772
rect 261850 997736 261906 997792
rect 263874 1002124 263876 1002144
rect 263876 1002124 263928 1002144
rect 263928 1002124 263930 1002144
rect 263874 1002088 263930 1002124
rect 298466 999096 298522 999152
rect 298282 998416 298338 998472
rect 298098 998008 298154 998064
rect 282734 995696 282790 995752
rect 290646 995696 290702 995752
rect 294786 995696 294842 995752
rect 295062 995696 295118 995752
rect 290462 995560 290518 995616
rect 280802 995288 280858 995344
rect 279422 995016 279478 995072
rect 292302 995324 292304 995344
rect 292304 995324 292356 995344
rect 292356 995324 292358 995344
rect 292302 995288 292358 995324
rect 292486 995288 292542 995344
rect 291842 994744 291898 994800
rect 288070 994472 288126 994528
rect 295706 995288 295762 995344
rect 296718 995288 296774 995344
rect 298650 996648 298706 996704
rect 293314 994472 293370 994528
rect 298650 994472 298706 994528
rect 299662 1002632 299718 1002688
rect 299294 997736 299350 997792
rect 299110 997192 299166 997248
rect 299662 996920 299718 996976
rect 299386 996396 299442 996432
rect 299386 996376 299388 996396
rect 299388 996376 299440 996396
rect 299440 996376 299442 996396
rect 359738 1006476 359740 1006496
rect 359740 1006476 359792 1006496
rect 359792 1006476 359794 1006496
rect 359738 1006440 359794 1006476
rect 358542 1006324 358598 1006360
rect 358542 1006304 358544 1006324
rect 358544 1006304 358596 1006324
rect 358596 1006304 358598 1006324
rect 306102 1006188 306158 1006224
rect 306102 1006168 306104 1006188
rect 306104 1006168 306156 1006188
rect 306156 1006168 306158 1006188
rect 361394 1006188 361450 1006224
rect 361394 1006168 361396 1006188
rect 361396 1006168 361448 1006188
rect 361448 1006168 361450 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006032 311862 1006088
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 354862 1006032 354918 1006088
rect 304078 1005796 304080 1005816
rect 304080 1005796 304132 1005816
rect 304132 1005796 304134 1005816
rect 304078 1005760 304134 1005796
rect 313830 1004964 313886 1005000
rect 313830 1004944 313832 1004964
rect 313832 1004944 313884 1004964
rect 313884 1004944 313886 1004964
rect 314658 1004828 314714 1004864
rect 314658 1004808 314660 1004828
rect 314660 1004808 314712 1004828
rect 314712 1004808 314714 1004828
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 303250 1002652 303306 1002688
rect 303250 1002632 303252 1002652
rect 303252 1002632 303304 1002652
rect 303304 1002632 303306 1002652
rect 306930 1002652 306986 1002688
rect 306930 1002632 306932 1002652
rect 306932 1002632 306984 1002652
rect 306984 1002632 306986 1002652
rect 304906 1002108 304962 1002144
rect 304906 1002088 304908 1002108
rect 304908 1002088 304960 1002108
rect 304960 1002088 304962 1002108
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 301686 999096 301742 999152
rect 308954 998588 308956 998608
rect 308956 998588 309008 998608
rect 309008 998588 309010 998608
rect 308954 998552 309010 998588
rect 303250 998452 303252 998472
rect 303252 998452 303304 998472
rect 303304 998452 303306 998472
rect 303250 998416 303306 998452
rect 305274 998452 305276 998472
rect 305276 998452 305328 998472
rect 305328 998452 305330 998472
rect 305274 998416 305330 998452
rect 307298 998300 307354 998336
rect 307298 998280 307300 998300
rect 307300 998280 307352 998300
rect 307352 998280 307354 998300
rect 303066 998008 303122 998064
rect 301502 996104 301558 996160
rect 301502 995560 301558 995616
rect 303250 996684 303252 996704
rect 303252 996684 303304 996704
rect 303304 996684 303306 996704
rect 303250 996648 303306 996684
rect 302882 994744 302938 994800
rect 306930 998164 306986 998200
rect 306930 998144 306932 998164
rect 306932 998144 306984 998164
rect 306984 998144 306986 998164
rect 306102 998028 306158 998064
rect 306102 998008 306104 998028
rect 306104 998008 306156 998028
rect 306156 998008 306158 998028
rect 308954 998028 309010 998064
rect 308954 998008 308956 998028
rect 308956 998008 309008 998028
rect 309008 998008 309010 998028
rect 307758 997892 307814 997928
rect 307758 997872 307760 997892
rect 307760 997872 307812 997892
rect 307812 997872 307814 997892
rect 310610 997892 310666 997928
rect 310610 997872 310612 997892
rect 310612 997872 310664 997892
rect 310664 997872 310666 997892
rect 307022 995560 307078 995616
rect 309782 997736 309838 997792
rect 316406 994200 316462 994256
rect 363418 1005932 363420 1005952
rect 363420 1005932 363472 1005952
rect 363472 1005932 363474 1005952
rect 363418 1005896 363474 1005932
rect 360566 1005524 360568 1005544
rect 360568 1005524 360620 1005544
rect 360620 1005524 360622 1005544
rect 360566 1005488 360622 1005524
rect 358542 1005388 358544 1005408
rect 358544 1005388 358596 1005408
rect 358596 1005388 358598 1005408
rect 358542 1005352 358598 1005388
rect 356518 1005100 356574 1005136
rect 356518 1005080 356520 1005100
rect 356520 1005080 356572 1005100
rect 356572 1005080 356574 1005100
rect 361394 1005100 361450 1005136
rect 361394 1005080 361396 1005100
rect 361396 1005080 361448 1005100
rect 361448 1005080 361450 1005100
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 355690 1004964 355746 1005000
rect 355690 1004944 355692 1004964
rect 355692 1004944 355744 1004964
rect 355744 1004944 355746 1004964
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 356886 1003892 356888 1003912
rect 356888 1003892 356940 1003912
rect 356940 1003892 356942 1003912
rect 356886 1003856 356942 1003892
rect 359370 1002516 359426 1002552
rect 359370 1002496 359372 1002516
rect 359372 1002496 359424 1002516
rect 359424 1002496 359426 1002516
rect 357346 1002380 357402 1002416
rect 357346 1002360 357348 1002380
rect 357348 1002360 357400 1002380
rect 357400 1002360 357402 1002380
rect 357714 1002244 357770 1002280
rect 357714 1002224 357716 1002244
rect 357716 1002224 357768 1002244
rect 357768 1002224 357770 1002244
rect 355690 1001972 355746 1002008
rect 355690 1001952 355692 1001972
rect 355692 1001952 355744 1001972
rect 355744 1001952 355746 1001972
rect 360566 1002108 360622 1002144
rect 360566 1002088 360568 1002108
rect 360568 1002088 360620 1002108
rect 360620 1002088 360622 1002108
rect 360198 1001972 360254 1002008
rect 360198 1001952 360200 1001972
rect 360200 1001952 360252 1001972
rect 360252 1001952 360254 1001972
rect 365074 1002260 365076 1002280
rect 365076 1002260 365128 1002280
rect 365128 1002260 365130 1002280
rect 365074 1002224 365130 1002260
rect 365074 1001988 365076 1002008
rect 365076 1001988 365128 1002008
rect 365128 1001988 365130 1002008
rect 365074 1001952 365130 1001988
rect 365902 1002124 365904 1002144
rect 365904 1002124 365956 1002144
rect 365956 1002124 365958 1002144
rect 365902 1002088 365958 1002124
rect 372526 996920 372582 996976
rect 372342 996376 372398 996432
rect 373262 996104 373318 996160
rect 375378 995288 375434 995344
rect 372986 995016 373042 995072
rect 380162 996648 380218 996704
rect 382278 995968 382334 996024
rect 383566 997192 383622 997248
rect 383474 996648 383530 996704
rect 399942 996920 399998 996976
rect 388166 995696 388222 995752
rect 389362 995288 389418 995344
rect 388994 995016 389050 995072
rect 392398 995424 392454 995480
rect 378046 994472 378102 994528
rect 392122 994472 392178 994528
rect 394974 995424 395030 995480
rect 422666 1006032 422722 1006088
rect 425518 1006052 425574 1006088
rect 425518 1006032 425520 1006052
rect 425520 1006032 425572 1006052
rect 425572 1006032 425574 1006052
rect 426346 1005780 426402 1005816
rect 426346 1005760 426348 1005780
rect 426348 1005760 426400 1005780
rect 426400 1005760 426402 1005780
rect 426346 1005524 426348 1005544
rect 426348 1005524 426400 1005544
rect 426400 1005524 426402 1005544
rect 426346 1005488 426402 1005524
rect 423494 1005252 423496 1005272
rect 423496 1005252 423548 1005272
rect 423548 1005252 423550 1005272
rect 423494 1005216 423550 1005252
rect 423494 1004964 423550 1005000
rect 423494 1004944 423496 1004964
rect 423496 1004944 423548 1004964
rect 423548 1004944 423550 1004964
rect 415950 995696 416006 995752
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 424322 1002804 424324 1002824
rect 424324 1002804 424376 1002824
rect 424376 1002804 424378 1002824
rect 424322 1002768 424378 1002804
rect 431682 1006460 431738 1006496
rect 431682 1006440 431684 1006460
rect 431684 1006440 431736 1006460
rect 431736 1006440 431738 1006460
rect 429198 1006188 429254 1006224
rect 429198 1006168 429200 1006188
rect 429200 1006168 429252 1006188
rect 429252 1006168 429254 1006188
rect 431682 1006204 431684 1006224
rect 431684 1006204 431736 1006224
rect 431736 1006204 431738 1006224
rect 431682 1006168 431738 1006204
rect 430854 1005932 430856 1005952
rect 430856 1005932 430908 1005952
rect 430908 1005932 430910 1005952
rect 430854 1005896 430910 1005932
rect 506202 1006460 506258 1006496
rect 506202 1006440 506204 1006460
rect 506204 1006440 506256 1006460
rect 506256 1006440 506258 1006460
rect 430026 1005388 430028 1005408
rect 430028 1005388 430080 1005408
rect 430080 1005388 430082 1005408
rect 430026 1005352 430082 1005388
rect 430026 1005100 430082 1005136
rect 430026 1005080 430028 1005100
rect 430028 1005080 430080 1005100
rect 430080 1005080 430082 1005100
rect 431222 1004964 431278 1005000
rect 431222 1004944 431224 1004964
rect 431224 1004944 431276 1004964
rect 431276 1004944 431278 1004964
rect 427174 1003892 427176 1003912
rect 427176 1003892 427228 1003912
rect 427228 1003892 427230 1003912
rect 427174 1003856 427230 1003892
rect 421470 1002108 421526 1002144
rect 421470 1002088 421472 1002108
rect 421472 1002088 421524 1002108
rect 421524 1002088 421526 1002108
rect 427542 1002108 427598 1002144
rect 427542 1002088 427544 1002108
rect 427544 1002088 427596 1002108
rect 427596 1002088 427598 1002108
rect 424322 1001972 424378 1002008
rect 424322 1001952 424324 1001972
rect 424324 1001952 424376 1001972
rect 424376 1001952 424378 1001972
rect 425150 1001952 425206 1002008
rect 425518 1001972 425574 1002008
rect 425518 1001952 425520 1001972
rect 425520 1001952 425572 1001972
rect 425572 1001952 425574 1001972
rect 428370 1002244 428426 1002280
rect 428370 1002224 428372 1002244
rect 428372 1002224 428424 1002244
rect 428424 1002224 428426 1002244
rect 429198 1001972 429254 1002008
rect 429198 1001952 429200 1001972
rect 429200 1001952 429252 1001972
rect 429252 1001952 429254 1001972
rect 432050 1002244 432106 1002280
rect 432050 1002224 432052 1002244
rect 432052 1002224 432104 1002244
rect 432104 1002224 432106 1002244
rect 433338 1002108 433394 1002144
rect 433338 1002088 433340 1002108
rect 433340 1002088 433392 1002108
rect 433392 1002088 433394 1002108
rect 432878 1001972 432934 1002008
rect 432878 1001952 432880 1001972
rect 432880 1001952 432932 1001972
rect 432932 1001952 432934 1001972
rect 439870 997192 439926 997248
rect 439686 996920 439742 996976
rect 453210 996240 453266 996296
rect 449162 995560 449218 995616
rect 458822 998144 458878 998200
rect 446402 994744 446458 994800
rect 508226 1006188 508282 1006224
rect 508226 1006168 508228 1006188
rect 508228 1006168 508280 1006188
rect 508280 1006168 508282 1006188
rect 461122 994472 461178 994528
rect 469862 995560 469918 995616
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 509054 1006052 509110 1006088
rect 509054 1006032 509056 1006052
rect 509056 1006032 509108 1006052
rect 509108 1006032 509110 1006052
rect 471242 995016 471298 995072
rect 472438 998144 472494 998200
rect 472438 996512 472494 996568
rect 472254 995968 472310 996024
rect 472438 995560 472494 995616
rect 488906 997192 488962 997248
rect 489090 996920 489146 996976
rect 489550 996648 489606 996704
rect 490102 996648 490158 996704
rect 472898 995696 472954 995752
rect 474002 995696 474058 995752
rect 476946 995696 477002 995752
rect 480810 995696 480866 995752
rect 485594 995696 485650 995752
rect 474738 995560 474794 995616
rect 478326 995560 478382 995616
rect 480258 995560 480314 995616
rect 476072 995016 476128 995072
rect 472070 994200 472126 994256
rect 478234 995288 478290 995344
rect 480258 994744 480314 994800
rect 476762 994200 476818 994256
rect 482650 994472 482706 994528
rect 494702 996376 494758 996432
rect 502154 1005388 502156 1005408
rect 502156 1005388 502208 1005408
rect 502208 1005388 502210 1005408
rect 502154 1005352 502210 1005388
rect 499670 1005252 499672 1005272
rect 499672 1005252 499724 1005272
rect 499724 1005252 499726 1005272
rect 499670 1005216 499726 1005252
rect 507030 1004964 507086 1005000
rect 507030 1004944 507032 1004964
rect 507032 1004944 507084 1004964
rect 507084 1004944 507086 1004964
rect 507858 1004828 507914 1004864
rect 507858 1004808 507860 1004828
rect 507860 1004808 507912 1004828
rect 507912 1004808 507914 1004828
rect 501326 1004692 501382 1004728
rect 501326 1004672 501328 1004692
rect 501328 1004672 501380 1004692
rect 501380 1004672 501382 1004692
rect 498474 1001972 498530 1002008
rect 498474 1001952 498476 1001972
rect 498476 1001952 498528 1001972
rect 498528 1001952 498530 1001972
rect 505374 1004572 505376 1004592
rect 505376 1004572 505428 1004592
rect 505428 1004572 505430 1004592
rect 505374 1004536 505430 1004572
rect 505006 1003892 505008 1003912
rect 505008 1003892 505060 1003912
rect 505060 1003892 505062 1003912
rect 505006 1003856 505062 1003892
rect 504178 1002668 504180 1002688
rect 504180 1002668 504232 1002688
rect 504232 1002668 504234 1002688
rect 504178 1002632 504234 1002668
rect 501694 1002532 501696 1002552
rect 501696 1002532 501748 1002552
rect 501748 1002532 501750 1002552
rect 501694 1002496 501750 1002532
rect 503350 1002380 503406 1002416
rect 503350 1002360 503352 1002380
rect 503352 1002360 503404 1002380
rect 503404 1002360 503406 1002380
rect 500498 1002244 500554 1002280
rect 500498 1002224 500500 1002244
rect 500500 1002224 500552 1002244
rect 500552 1002224 500554 1002244
rect 500498 1001972 500554 1002008
rect 500498 1001952 500500 1001972
rect 500500 1001952 500552 1001972
rect 500552 1001952 500554 1001972
rect 502154 1001972 502210 1002008
rect 502154 1001952 502156 1001972
rect 502156 1001952 502208 1001972
rect 502208 1001952 502210 1001972
rect 502522 1001972 502578 1002008
rect 502522 1001952 502524 1001972
rect 502524 1001952 502576 1001972
rect 502576 1001952 502578 1001972
rect 503350 1002108 503406 1002144
rect 503350 1002088 503352 1002108
rect 503352 1002088 503404 1002108
rect 503404 1002088 503406 1002108
rect 506202 1001952 506258 1002008
rect 507398 1001952 507454 1002008
rect 509882 1002244 509938 1002280
rect 509882 1002224 509884 1002244
rect 509884 1002224 509936 1002244
rect 509936 1002224 509938 1002244
rect 510342 1002108 510398 1002144
rect 510342 1002088 510344 1002108
rect 510344 1002088 510396 1002108
rect 510396 1002088 510398 1002108
rect 503810 995560 503866 995616
rect 503810 995016 503866 995072
rect 554318 1006732 554374 1006768
rect 554318 1006712 554320 1006732
rect 554320 1006712 554372 1006732
rect 554372 1006712 554374 1006732
rect 555974 1006460 556030 1006496
rect 555974 1006440 555976 1006460
rect 555976 1006440 556028 1006460
rect 556028 1006440 556030 1006460
rect 516690 998552 516746 998608
rect 516690 997192 516746 997248
rect 517058 996920 517114 996976
rect 516874 995560 516930 995616
rect 519818 996240 519874 996296
rect 550270 1006052 550326 1006088
rect 550270 1006032 550272 1006052
rect 550272 1006032 550324 1006052
rect 550324 1006032 550326 1006052
rect 553950 1006052 554006 1006088
rect 553950 1006032 553952 1006052
rect 553952 1006032 554004 1006052
rect 554004 1006032 554006 1006052
rect 522302 996240 522358 996296
rect 520922 995832 520978 995888
rect 520186 995016 520242 995072
rect 517518 994472 517574 994528
rect 522946 995288 523002 995344
rect 523406 998552 523462 998608
rect 524050 997736 524106 997792
rect 540334 997192 540390 997248
rect 540518 996920 540574 996976
rect 523866 995968 523922 996024
rect 523406 995016 523462 995072
rect 532238 995696 532294 995752
rect 525338 995288 525394 995344
rect 529846 995560 529902 995616
rect 536930 995560 536986 995616
rect 528558 995288 528614 995344
rect 528926 995288 528982 995344
rect 526074 995016 526130 995072
rect 527914 995016 527970 995072
rect 526534 994744 526590 994800
rect 523222 994200 523278 994256
rect 533710 994744 533766 994800
rect 533066 994472 533122 994528
rect 526534 994200 526590 994256
rect 551466 1005388 551468 1005408
rect 551468 1005388 551520 1005408
rect 551520 1005388 551522 1005408
rect 551466 1005352 551522 1005388
rect 551466 1005116 551468 1005136
rect 551468 1005116 551520 1005136
rect 551520 1005116 551522 1005136
rect 551466 1005080 551522 1005116
rect 556802 1004964 556858 1005000
rect 556802 1004944 556804 1004964
rect 556804 1004944 556856 1004964
rect 556856 1004944 556858 1004964
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 552294 1003892 552296 1003912
rect 552296 1003892 552348 1003912
rect 552348 1003892 552350 1003912
rect 552294 1003856 552350 1003892
rect 552294 1002108 552350 1002144
rect 552294 1002088 552296 1002108
rect 552296 1002088 552348 1002108
rect 552348 1002088 552350 1002108
rect 554318 1001952 554374 1002008
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 553122 998028 553178 998064
rect 553122 998008 553124 998028
rect 553124 998008 553176 998028
rect 553176 998008 553178 998028
rect 553122 997772 553124 997792
rect 553124 997772 553176 997792
rect 553176 997772 553178 997792
rect 553122 997736 553178 997772
rect 554778 1002224 554834 1002280
rect 555146 1001972 555202 1002008
rect 555146 1001952 555148 1001972
rect 555148 1001952 555200 1001972
rect 555200 1001952 555202 1001972
rect 557170 1006188 557226 1006224
rect 557170 1006168 557172 1006188
rect 557172 1006168 557224 1006188
rect 557224 1006168 557226 1006188
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002108 558054 1002144
rect 557998 1002088 558000 1002108
rect 558000 1002088 558052 1002108
rect 558052 1002088 558054 1002108
rect 558826 1002516 558882 1002552
rect 558826 1002496 558828 1002516
rect 558828 1002496 558880 1002516
rect 558880 1002496 558882 1002516
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 557170 998044 557172 998064
rect 557172 998044 557224 998064
rect 557224 998044 557226 998064
rect 557170 998008 557226 998044
rect 552662 995560 552718 995616
rect 552662 995016 552718 995072
rect 560850 1002380 560906 1002416
rect 560850 1002360 560852 1002380
rect 560852 1002360 560904 1002380
rect 560904 1002360 560906 1002380
rect 560022 1002244 560078 1002280
rect 560022 1002224 560024 1002244
rect 560024 1002224 560076 1002244
rect 560076 1002224 560078 1002244
rect 560850 1002108 560906 1002144
rect 560850 1002088 560852 1002108
rect 560852 1002088 560904 1002108
rect 560904 1002088 560906 1002108
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 599950 996920 600006 996976
rect 590566 996648 590622 996704
rect 591302 996376 591358 996432
rect 599950 996376 600006 996432
rect 618166 996376 618222 996432
rect 590566 995016 590622 995072
rect 620098 995968 620154 996024
rect 623686 995968 623742 996024
rect 635186 995696 635242 995752
rect 625526 995424 625582 995480
rect 627182 995424 627238 995480
rect 627918 995424 627974 995480
rect 631506 995424 631562 995480
rect 633990 995424 634046 995480
rect 634726 995424 634782 995480
rect 631690 995288 631746 995344
rect 568210 993656 568266 993712
rect 576306 990936 576362 990992
rect 660578 995035 660634 995072
rect 660578 995016 660580 995035
rect 660580 995016 660632 995035
rect 660632 995016 660634 995035
rect 641718 993656 641774 993712
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 937216 660358 937272
rect 663062 941704 663118 941760
rect 667202 947280 667258 947336
rect 665822 939800 665878 939856
rect 675666 966456 675722 966512
rect 673366 962784 673422 962840
rect 673182 958160 673238 958216
rect 672998 952176 673054 952232
rect 669962 938712 670018 938768
rect 671802 938304 671858 938360
rect 668582 937760 668638 937816
rect 671434 937488 671490 937544
rect 658922 935992 658978 936048
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 55862 892744 55918 892800
rect 54482 892200 54538 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62762 858608 62818 858664
rect 62118 845552 62174 845608
rect 53102 799584 53158 799640
rect 62118 832496 62174 832552
rect 54482 774288 54538 774344
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793620 62174 793656
rect 62118 793600 62120 793620
rect 62120 793600 62172 793620
rect 62172 793600 62174 793620
rect 651470 856296 651526 856352
rect 651838 842968 651894 843024
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 651470 789928 651526 789984
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 55862 772792 55918 772848
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 50342 730496 50398 730552
rect 48962 669296 49018 669352
rect 47398 638152 47454 638208
rect 47398 618704 47454 618760
rect 47214 610952 47270 611008
rect 45374 598848 45430 598904
rect 45190 598032 45246 598088
rect 652390 776600 652446 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62762 743008 62818 743064
rect 62118 741240 62174 741296
rect 51722 691328 51778 691384
rect 652022 736752 652078 736808
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 50342 626592 50398 626648
rect 51722 601704 51778 601760
rect 48962 601296 49018 601352
rect 651470 723424 651526 723480
rect 651470 710232 651526 710288
rect 651470 696940 651472 696960
rect 651472 696940 651524 696960
rect 651524 696940 651526 696960
rect 651470 696904 651526 696940
rect 62762 689424 62818 689480
rect 62118 689152 62174 689208
rect 651654 683576 651710 683632
rect 62762 676096 62818 676152
rect 62118 663040 62174 663096
rect 651470 670384 651526 670440
rect 651470 657056 651526 657112
rect 62762 656104 62818 656160
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 651562 630536 651618 630592
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652022 628496 652078 628552
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 54482 600888 54538 600944
rect 47582 580488 47638 580544
rect 50342 558456 50398 558512
rect 48962 557640 49018 557696
rect 45558 556824 45614 556880
rect 45006 556416 45062 556472
rect 44914 556008 44970 556064
rect 44638 555600 44694 555656
rect 44730 555192 44786 555248
rect 44362 554376 44418 554432
rect 44178 549072 44234 549128
rect 43626 548120 43682 548176
rect 43810 547032 43866 547088
rect 42982 379344 43038 379400
rect 43350 371864 43406 371920
rect 42982 365744 43038 365800
rect 42430 356088 42486 356144
rect 43350 355816 43406 355872
rect 41786 355680 41842 355736
rect 44178 537376 44234 537432
rect 44546 550704 44602 550760
rect 44546 532752 44602 532808
rect 44546 429256 44602 429312
rect 44362 427624 44418 427680
rect 44178 427216 44234 427272
rect 44178 421504 44234 421560
rect 43994 419464 44050 419520
rect 44178 406816 44234 406872
rect 45098 551520 45154 551576
rect 45282 548664 45338 548720
rect 45282 536968 45338 537024
rect 45098 529760 45154 529816
rect 45558 429664 45614 429720
rect 44914 428848 44970 428904
rect 45006 428440 45062 428496
rect 44730 428032 44786 428088
rect 44822 420688 44878 420744
rect 44546 386688 44602 386744
rect 44638 386008 44694 386064
rect 44638 385192 44694 385248
rect 44362 384784 44418 384840
rect 44454 379888 44510 379944
rect 44270 377440 44326 377496
rect 45190 426808 45246 426864
rect 45374 423136 45430 423192
rect 45374 402872 45430 402928
rect 45098 385600 45154 385656
rect 44454 359896 44510 359952
rect 44270 356632 44326 356688
rect 45190 384376 45246 384432
rect 45374 383968 45430 384024
rect 45190 383560 45246 383616
rect 43902 354184 43958 354240
rect 44730 353776 44786 353832
rect 28538 351192 28594 351248
rect 40222 345480 40278 345536
rect 28538 343848 28594 343904
rect 35806 343848 35862 343904
rect 45006 343304 45062 343360
rect 45558 380296 45614 380352
rect 47582 430072 47638 430128
rect 46938 426400 46994 426456
rect 47122 423544 47178 423600
rect 47122 400152 47178 400208
rect 46938 399744 46994 399800
rect 46938 380704 46994 380760
rect 46202 366968 46258 367024
rect 45558 357312 45614 357368
rect 45650 356632 45706 356688
rect 45926 355816 45982 355872
rect 45374 341672 45430 341728
rect 45466 341264 45522 341320
rect 45190 340856 45246 340912
rect 35806 339768 35862 339824
rect 36634 336504 36690 336560
rect 42798 334600 42854 334656
rect 43074 334600 43130 334656
rect 41602 334464 41658 334520
rect 41602 333648 41658 333704
rect 41786 326712 41842 326768
rect 41786 325352 41842 325408
rect 41878 324808 41934 324864
rect 42062 322768 42118 322824
rect 42522 321408 42578 321464
rect 42246 321136 42302 321192
rect 42430 320864 42486 320920
rect 44178 334328 44234 334384
rect 43258 333648 43314 333704
rect 43074 322768 43130 322824
rect 43258 321136 43314 321192
rect 44178 320864 44234 320920
rect 41786 319912 41842 319968
rect 42246 317464 42302 317520
rect 41786 316648 41842 316704
rect 42154 315968 42210 316024
rect 42154 315424 42210 315480
rect 42154 313656 42210 313712
rect 42430 312704 42486 312760
rect 42154 312296 42210 312352
rect 44546 311480 44602 311536
rect 44362 311208 44418 311264
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 44546 300056 44602 300112
rect 44638 299648 44694 299704
rect 44362 299240 44418 299296
rect 42890 298016 42946 298072
rect 41786 296792 41842 296848
rect 37922 294752 37978 294808
rect 42062 295976 42118 296032
rect 41786 292712 41842 292768
rect 42062 292304 42118 292360
rect 42246 291080 42302 291136
rect 42062 290400 42118 290456
rect 41326 290264 41382 290320
rect 42062 289856 42118 289912
rect 42246 289856 42302 289912
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42430 278704 42486 278760
rect 42430 278160 42486 278216
rect 41786 277888 41842 277944
rect 42338 277616 42394 277672
rect 42154 277344 42210 277400
rect 42062 276528 42118 276584
rect 41786 274216 41842 274272
rect 42062 273400 42118 273456
rect 42062 272856 42118 272912
rect 41786 270408 41842 270464
rect 42430 270408 42486 270464
rect 41786 269048 41842 269104
rect 40682 267008 40738 267064
rect 35806 259936 35862 259992
rect 35806 258304 35862 258360
rect 35806 257080 35862 257136
rect 43258 297200 43314 297256
rect 43074 293528 43130 293584
rect 43074 273400 43130 273456
rect 42890 255176 42946 255232
rect 42890 254768 42946 254824
rect 35806 253408 35862 253464
rect 35622 253000 35678 253056
rect 35806 252612 35862 252648
rect 35806 252592 35808 252612
rect 35808 252592 35860 252612
rect 35860 252592 35862 252612
rect 35806 252184 35862 252240
rect 41326 252184 41382 252240
rect 42522 252184 42578 252240
rect 41694 242836 41696 242856
rect 41696 242836 41748 242856
rect 41748 242836 41750 242856
rect 41694 242800 41750 242836
rect 40682 242528 40738 242584
rect 41786 240080 41842 240136
rect 42062 238448 42118 238504
rect 42706 242800 42762 242856
rect 42522 237360 42578 237416
rect 41786 235864 41842 235920
rect 42430 235864 42486 235920
rect 42246 234096 42302 234152
rect 42154 233280 42210 233336
rect 42430 232464 42486 232520
rect 42430 231784 42486 231840
rect 42154 230424 42210 230480
rect 42430 229336 42486 229392
rect 43442 294344 43498 294400
rect 44362 293936 44418 293992
rect 43626 293120 43682 293176
rect 43810 291896 43866 291952
rect 43626 279792 43682 279848
rect 44178 291488 44234 291544
rect 44178 278160 44234 278216
rect 43810 277344 43866 277400
rect 44362 272856 44418 272912
rect 43442 270408 43498 270464
rect 45190 298832 45246 298888
rect 45006 295160 45062 295216
rect 44822 291896 44878 291952
rect 44638 256808 44694 256864
rect 43626 256400 43682 256456
rect 43442 255584 43498 255640
rect 43258 254360 43314 254416
rect 43074 250280 43130 250336
rect 43258 242528 43314 242584
rect 43074 230424 43130 230480
rect 41970 227296 42026 227352
rect 42154 226616 42210 226672
rect 42430 225664 42486 225720
rect 41694 224440 41750 224496
rect 28538 222808 28594 222864
rect 28538 214240 28594 214296
rect 35806 214240 35862 214296
rect 43258 225664 43314 225720
rect 35622 212200 35678 212256
rect 44178 253952 44234 254008
rect 43810 249056 43866 249112
rect 43810 231784 43866 231840
rect 43626 213696 43682 213752
rect 43442 212880 43498 212936
rect 42890 212064 42946 212120
rect 35806 211384 35862 211440
rect 44362 251912 44418 251968
rect 44546 248648 44602 248704
rect 44546 234096 44602 234152
rect 44362 233280 44418 233336
rect 45006 276528 45062 276584
rect 45834 340040 45890 340096
rect 45650 339224 45706 339280
rect 46018 338816 46074 338872
rect 46018 315424 46074 315480
rect 45834 313656 45890 313712
rect 45650 312296 45706 312352
rect 45466 298424 45522 298480
rect 45466 291896 45522 291952
rect 47122 379072 47178 379128
rect 47122 361528 47178 361584
rect 46938 356088 46994 356144
rect 47582 333104 47638 333160
rect 46386 303048 46442 303104
rect 46202 259936 46258 259992
rect 45098 255992 45154 256048
rect 45558 251096 45614 251152
rect 45006 248240 45062 248296
rect 45006 235864 45062 235920
rect 45834 250688 45890 250744
rect 46018 249464 46074 249520
rect 46202 247832 46258 247888
rect 46018 232464 46074 232520
rect 45834 229336 45890 229392
rect 45558 226616 45614 226672
rect 44822 214920 44878 214976
rect 35806 209788 35808 209808
rect 35808 209788 35860 209808
rect 35860 209788 35862 209808
rect 35806 209752 35862 209788
rect 41694 208936 41750 208992
rect 41326 205672 41382 205728
rect 41142 204040 41198 204096
rect 41326 203632 41382 203688
rect 41326 202136 41382 202192
rect 44178 211248 44234 211304
rect 44178 210432 44234 210488
rect 42798 209616 42854 209672
rect 41878 201456 41934 201512
rect 41142 200640 41198 200696
rect 41786 197104 41842 197160
rect 41786 195744 41842 195800
rect 42246 195336 42302 195392
rect 41970 195064 42026 195120
rect 42246 193160 42302 193216
rect 42430 193160 42486 193216
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41786 187176 41842 187232
rect 42062 186360 42118 186416
rect 42154 185816 42210 185872
rect 42430 184864 42486 184920
rect 42430 183096 42486 183152
rect 43258 207984 43314 208040
rect 42982 206352 43038 206408
rect 42982 191120 43038 191176
rect 43626 206760 43682 206816
rect 43442 200640 43498 200696
rect 43258 183096 43314 183152
rect 43810 205264 43866 205320
rect 43626 193160 43682 193216
rect 43994 204856 44050 204912
rect 43994 191664 44050 191720
rect 43810 190440 43866 190496
rect 44546 208528 44602 208584
rect 44362 205944 44418 206000
rect 44822 204448 44878 204504
rect 44546 189896 44602 189952
rect 44362 187584 44418 187640
rect 44178 184864 44234 184920
rect 46938 247016 46994 247072
rect 46938 238448 46994 238504
rect 46386 203496 46442 203552
rect 50342 430888 50398 430944
rect 48962 386824 49018 386880
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 213288 48006 213344
rect 48134 210840 48190 210896
rect 48134 194384 48190 194440
rect 47950 190440 48006 190496
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 62118 597896 62174 597952
rect 652390 590708 652446 590744
rect 652390 590688 652392 590708
rect 652392 590688 652444 590708
rect 652444 590688 652446 590708
rect 62118 584840 62174 584896
rect 664442 868672 664498 868728
rect 663062 760416 663118 760472
rect 670606 876832 670662 876888
rect 669226 876288 669282 876344
rect 668858 872208 668914 872264
rect 666282 778368 666338 778424
rect 665822 761504 665878 761560
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661682 673104 661738 673160
rect 661682 643728 661738 643784
rect 660302 625232 660358 625288
rect 660302 599528 660358 599584
rect 658922 579672 658978 579728
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 658922 553968 658978 554024
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 652574 497664 652630 497720
rect 62118 493584 62174 493640
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62946 415384 63002 415440
rect 55862 408448 55918 408504
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51722 301280 51778 301336
rect 49146 290400 49202 290456
rect 50342 290128 50398 290184
rect 49606 208936 49662 208992
rect 49422 201456 49478 201512
rect 49606 196424 49662 196480
rect 49422 192344 49478 192400
rect 51722 289856 51778 289912
rect 50526 246472 50582 246528
rect 53286 257488 53342 257544
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 62118 376216 62174 376272
rect 62118 363296 62174 363352
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 55862 278704 55918 278760
rect 651470 404640 651526 404696
rect 652574 391448 652630 391504
rect 651838 364792 651894 364848
rect 652390 351600 652446 351656
rect 62946 345616 63002 345672
rect 652022 338272 652078 338328
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 651470 285232 651526 285288
rect 62946 285096 63002 285152
rect 62762 267008 62818 267064
rect 54482 222808 54538 222864
rect 58990 224168 59046 224224
rect 102046 269728 102102 269784
rect 75918 267008 75974 267064
rect 138110 267008 138166 267064
rect 161294 269728 161350 269784
rect 468482 269728 468538 269784
rect 470966 269184 471022 269240
rect 477590 266328 477646 266384
rect 479706 271360 479762 271416
rect 479706 266328 479762 266384
rect 484122 267008 484178 267064
rect 497462 269456 497518 269512
rect 506110 268368 506166 268424
rect 507766 271088 507822 271144
rect 507950 267008 508006 267064
rect 513194 274080 513250 274136
rect 517150 267008 517206 267064
rect 519818 267280 519874 267336
rect 521474 272992 521530 273048
rect 530950 270272 531006 270328
rect 533434 273808 533490 273864
rect 533894 272720 533950 272776
rect 535734 275168 535790 275224
rect 539322 272448 539378 272504
rect 538034 270000 538090 270056
rect 537666 269728 537722 269784
rect 540518 269728 540574 269784
rect 539506 269184 539562 269240
rect 551742 271360 551798 271416
rect 563702 267280 563758 267336
rect 568578 269456 568634 269512
rect 591118 268368 591174 268424
rect 585782 267008 585838 267064
rect 593142 271088 593198 271144
rect 602526 274080 602582 274136
rect 614394 272992 614450 273048
rect 626630 270272 626686 270328
rect 630954 273808 631010 273864
rect 633346 275168 633402 275224
rect 632150 272720 632206 272776
rect 639234 272448 639290 272504
rect 637578 270000 637634 270056
rect 640706 269728 640762 269784
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553766 255584 553822 255640
rect 554410 253408 554466 253464
rect 553490 251252 553546 251288
rect 553490 251232 553492 251252
rect 553492 251232 553544 251252
rect 553544 251232 553546 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553674 242528 553730 242584
rect 71042 230016 71098 230072
rect 65522 229744 65578 229800
rect 62946 224440 63002 224496
rect 64786 222808 64842 222864
rect 66902 224440 66958 224496
rect 73710 228248 73766 228304
rect 72422 224712 72478 224768
rect 71410 223080 71466 223136
rect 79966 226888 80022 226944
rect 77206 218592 77262 218648
rect 82726 225528 82782 225584
rect 89626 227160 89682 227216
rect 89442 225800 89498 225856
rect 92110 223352 92166 223408
rect 95422 221448 95478 221504
rect 97722 221720 97778 221776
rect 108670 221992 108726 222048
rect 112994 228520 113050 228576
rect 117778 220088 117834 220144
rect 125230 226072 125286 226128
rect 124402 220360 124458 220416
rect 136546 227432 136602 227488
rect 145010 224168 145066 224224
rect 148230 229744 148286 229800
rect 146942 224168 146998 224224
rect 146666 222808 146722 222864
rect 150806 230016 150862 230072
rect 149794 224440 149850 224496
rect 147586 220632 147642 220688
rect 150898 222808 150954 222864
rect 152738 224712 152794 224768
rect 152094 223080 152150 223136
rect 155314 228248 155370 228304
rect 157706 218592 157762 218648
rect 160466 226888 160522 226944
rect 159822 218592 159878 218648
rect 163042 225528 163098 225584
rect 166906 227160 166962 227216
rect 168930 228248 168986 228304
rect 168194 225800 168250 225856
rect 170770 223352 170826 223408
rect 171046 221176 171102 221232
rect 172702 221720 172758 221776
rect 172978 221448 173034 221504
rect 175922 224168 175978 224224
rect 176566 224440 176622 224496
rect 183650 221992 183706 222048
rect 184938 228520 184994 228576
rect 185214 224612 185216 224632
rect 185216 224612 185268 224632
rect 185268 224612 185270 224632
rect 185214 224576 185270 224612
rect 186226 224612 186228 224632
rect 186228 224612 186280 224632
rect 186280 224612 186282 224632
rect 186226 224576 186282 224612
rect 187882 220088 187938 220144
rect 193310 220360 193366 220416
rect 196530 226072 196586 226128
rect 200762 218592 200818 218648
rect 202970 227432 203026 227488
rect 204902 224168 204958 224224
rect 211342 220632 211398 220688
rect 213918 222808 213974 222864
rect 223578 228248 223634 228304
rect 229558 221176 229614 221232
rect 484582 218048 484638 218104
rect 485042 218048 485098 218104
rect 487802 218320 487858 218376
rect 489090 217096 489146 217152
rect 490286 218592 490342 218648
rect 491942 219408 491998 219464
rect 493690 218864 493746 218920
rect 494702 219136 494758 219192
rect 495254 217232 495310 217288
rect 497002 218592 497058 218648
rect 497554 218592 497610 218648
rect 499210 218864 499266 218920
rect 499210 217776 499266 217832
rect 499578 218320 499634 218376
rect 499762 218320 499818 218376
rect 499762 217776 499818 217832
rect 501050 217504 501106 217560
rect 502982 217504 503038 217560
rect 503350 217504 503406 217560
rect 503626 217504 503682 217560
rect 505098 219136 505154 219192
rect 505282 219136 505338 219192
rect 505466 217504 505522 217560
rect 506110 217504 506166 217560
rect 507766 217776 507822 217832
rect 508686 217504 508742 217560
rect 510986 217776 511042 217832
rect 513562 221992 513618 222048
rect 515770 221176 515826 221232
rect 514942 217796 514998 217832
rect 514942 217776 514944 217796
rect 514944 217776 514996 217796
rect 514996 217776 514998 217796
rect 515126 217776 515182 217832
rect 517518 220904 517574 220960
rect 518530 220904 518586 220960
rect 518346 217776 518402 217832
rect 518898 219680 518954 219736
rect 518898 218048 518954 218104
rect 519082 218048 519138 218104
rect 518714 217796 518770 217832
rect 518714 217776 518716 217796
rect 518716 217776 518768 217796
rect 518768 217776 518770 217796
rect 518898 217504 518954 217560
rect 519082 217524 519138 217560
rect 519082 217504 519084 217524
rect 519084 217504 519136 217524
rect 519136 217504 519138 217524
rect 521014 221448 521070 221504
rect 522578 220496 522634 220552
rect 524970 219952 525026 220008
rect 524418 218048 524474 218104
rect 524602 218048 524658 218104
rect 527546 220224 527602 220280
rect 528466 219680 528522 219736
rect 530858 221720 530914 221776
rect 530030 219952 530086 220008
rect 533710 219102 533766 219158
rect 533894 219136 533950 219192
rect 534078 219136 534134 219192
rect 534262 219156 534318 219192
rect 534262 219136 534264 219156
rect 534264 219136 534316 219156
rect 534316 219136 534318 219156
rect 554502 244704 554558 244760
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 553122 219408 553178 219464
rect 554226 219136 554282 219192
rect 563334 222264 563390 222320
rect 563058 217504 563114 217560
rect 563242 217504 563298 217560
rect 567842 218864 567898 218920
rect 568302 218864 568358 218920
rect 567658 218320 567714 218376
rect 567842 218320 567898 218376
rect 571890 222264 571946 222320
rect 572718 218864 572774 218920
rect 572442 218320 572498 218376
rect 572626 218320 572682 218376
rect 572994 218048 573050 218104
rect 572258 217504 572314 217560
rect 572902 217504 572958 217560
rect 577042 215056 577098 215112
rect 591394 219172 591396 219192
rect 591396 219172 591448 219192
rect 591448 219172 591450 219192
rect 591394 219136 591450 219172
rect 582102 218048 582158 218104
rect 582286 218068 582342 218104
rect 582286 218048 582288 218068
rect 582288 218048 582340 218068
rect 582340 218048 582342 218068
rect 591854 217776 591910 217832
rect 582102 217504 582158 217560
rect 582286 217504 582342 217560
rect 582378 217232 582434 217288
rect 582930 216960 582986 217016
rect 586886 216960 586942 217016
rect 592222 216960 592278 217016
rect 582378 215872 582434 215928
rect 582562 215892 582618 215928
rect 582562 215872 582564 215892
rect 582564 215872 582616 215892
rect 582616 215872 582618 215892
rect 578882 213968 578938 214024
rect 578238 211656 578294 211712
rect 579250 209788 579252 209808
rect 579252 209788 579304 209808
rect 579304 209788 579306 209808
rect 579250 209752 579306 209788
rect 599490 221992 599546 222048
rect 594154 219408 594210 219464
rect 595166 219136 595222 219192
rect 594798 216688 594854 216744
rect 594982 216688 595038 216744
rect 594614 215620 594670 215656
rect 594614 215600 594616 215620
rect 594616 215600 594668 215620
rect 594668 215600 594670 215620
rect 595718 216960 595774 217016
rect 596362 216144 596418 216200
rect 596086 215056 596142 215112
rect 597558 217776 597614 217832
rect 599030 216688 599086 216744
rect 597926 215600 597982 215656
rect 603354 221720 603410 221776
rect 600318 221448 600374 221504
rect 600778 221176 600834 221232
rect 600594 220904 600650 220960
rect 602066 218592 602122 218648
rect 606758 217504 606814 217560
rect 606758 216960 606814 217016
rect 612738 218320 612794 218376
rect 611726 215872 611782 215928
rect 618810 220496 618866 220552
rect 617798 217504 617854 217560
rect 617246 217232 617302 217288
rect 618350 216416 618406 216472
rect 619638 220224 619694 220280
rect 620466 219952 620522 220008
rect 619822 219680 619878 219736
rect 621294 219408 621350 219464
rect 627734 218048 627790 218104
rect 639602 229744 639658 229800
rect 630678 218592 630734 218648
rect 637578 220088 637634 220144
rect 650642 225528 650698 225584
rect 646134 220360 646190 220416
rect 641166 218864 641222 218920
rect 639970 217504 640026 217560
rect 643834 218320 643890 218376
rect 643006 215872 643062 215928
rect 644938 217776 644994 217832
rect 648618 219816 648674 219872
rect 646594 216144 646650 216200
rect 647146 213152 647202 213208
rect 650458 214512 650514 214568
rect 651286 219136 651342 219192
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 652206 298424 652262 298480
rect 666466 742464 666522 742520
rect 666282 711592 666338 711648
rect 668214 789384 668270 789440
rect 667846 743144 667902 743200
rect 667662 688880 667718 688936
rect 667202 671064 667258 671120
rect 666466 665352 666522 665408
rect 665822 626048 665878 626104
rect 664442 580080 664498 580136
rect 663062 538736 663118 538792
rect 661682 491544 661738 491600
rect 660302 411848 660358 411904
rect 659106 360032 659162 360088
rect 661866 406272 661922 406328
rect 661682 313520 661738 313576
rect 658922 233824 658978 233880
rect 664442 494672 664498 494728
rect 668398 735256 668454 735312
rect 668214 709552 668270 709608
rect 668398 692824 668454 692880
rect 668214 685480 668270 685536
rect 667846 665896 667902 665952
rect 667846 643184 667902 643240
rect 667662 621152 667718 621208
rect 669042 866632 669098 866688
rect 668858 755248 668914 755304
rect 669778 873432 669834 873488
rect 669594 783808 669650 783864
rect 669226 753480 669282 753536
rect 669042 750760 669098 750816
rect 669226 741104 669282 741160
rect 668766 738928 668822 738984
rect 668582 670520 668638 670576
rect 669042 733624 669098 733680
rect 668766 666168 668822 666224
rect 669778 756064 669834 756120
rect 669778 731448 669834 731504
rect 669594 708736 669650 708792
rect 669594 701120 669650 701176
rect 669226 663856 669282 663912
rect 669042 662496 669098 662552
rect 669226 654200 669282 654256
rect 668398 619928 668454 619984
rect 668214 615576 668270 615632
rect 668398 593544 668454 593600
rect 667846 576000 667902 576056
rect 667846 564440 667902 564496
rect 667662 554648 667718 554704
rect 667202 534112 667258 534168
rect 665822 492088 665878 492144
rect 663246 358536 663302 358592
rect 668766 604288 668822 604344
rect 668582 535880 668638 535936
rect 669042 599256 669098 599312
rect 668766 528808 668822 528864
rect 668398 528536 668454 528592
rect 670330 782448 670386 782504
rect 670146 775648 670202 775704
rect 669962 715672 670018 715728
rect 670146 709960 670202 710016
rect 670790 778368 670846 778424
rect 670790 776464 670846 776520
rect 671158 869080 671214 869136
rect 670974 763000 671030 763056
rect 670974 758240 671030 758296
rect 670606 754568 670662 754624
rect 670790 750080 670846 750136
rect 670606 730496 670662 730552
rect 670330 707104 670386 707160
rect 669778 664128 669834 664184
rect 669778 638560 669834 638616
rect 669594 621560 669650 621616
rect 669594 614896 669650 614952
rect 669226 574096 669282 574152
rect 669226 557504 669282 557560
rect 669042 527312 669098 527368
rect 669226 485968 669282 486024
rect 667846 485152 667902 485208
rect 667662 482704 667718 482760
rect 670422 696904 670478 696960
rect 670146 685888 670202 685944
rect 670790 727912 670846 727968
rect 671618 774968 671674 775024
rect 671434 759464 671490 759520
rect 671158 753344 671214 753400
rect 671158 751304 671214 751360
rect 671342 734848 671398 734904
rect 671158 728184 671214 728240
rect 671158 714040 671214 714096
rect 670974 713632 671030 713688
rect 670974 713224 671030 713280
rect 671158 669840 671214 669896
rect 670974 668208 671030 668264
rect 671066 667936 671122 667992
rect 670606 660048 670662 660104
rect 670606 659640 670662 659696
rect 670422 620608 670478 620664
rect 670146 620336 670202 620392
rect 670422 616120 670478 616176
rect 670146 600344 670202 600400
rect 669962 581032 670018 581088
rect 669778 574368 669834 574424
rect 669962 553968 670018 554024
rect 669778 553424 669834 553480
rect 669962 551520 670018 551576
rect 669778 482296 669834 482352
rect 669594 454960 669650 455016
rect 667202 360848 667258 360904
rect 665822 315424 665878 315480
rect 664442 271088 664498 271144
rect 663062 268096 663118 268152
rect 667018 237088 667074 237144
rect 663798 231240 663854 231296
rect 660946 229472 661002 229528
rect 653402 229064 653458 229120
rect 652390 222808 652446 222864
rect 653034 221448 653090 221504
rect 658922 226616 658978 226672
rect 654782 226344 654838 226400
rect 655610 225256 655666 225312
rect 658186 224168 658242 224224
rect 656898 223896 656954 223952
rect 656162 223624 656218 223680
rect 657542 223080 657598 223136
rect 656530 217232 656586 217288
rect 659290 214784 659346 214840
rect 660762 221992 660818 222048
rect 661682 224984 661738 225040
rect 662050 215056 662106 215112
rect 661498 213424 661554 213480
rect 663062 230696 663118 230752
rect 665822 230968 665878 231024
rect 665178 230288 665234 230344
rect 664166 221720 664222 221776
rect 664810 213696 664866 213752
rect 666834 223896 666890 223952
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579526 144644 579528 144664
rect 579528 144644 579580 144664
rect 579580 144644 579582 144664
rect 579526 144608 579582 144644
rect 579526 142976 579582 143032
rect 579250 136584 579306 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578330 123528 578386 123584
rect 578698 118360 578754 118416
rect 578698 116864 578754 116920
rect 579066 129648 579122 129704
rect 579158 127744 579214 127800
rect 579526 125332 579528 125352
rect 579528 125332 579580 125352
rect 579580 125332 579582 125352
rect 579526 125296 579582 125332
rect 579526 121080 579582 121136
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579158 112512 579214 112568
rect 578882 110336 578938 110392
rect 578882 108296 578938 108352
rect 579066 105848 579122 105904
rect 578330 103300 578332 103320
rect 578332 103300 578384 103320
rect 578384 103300 578386 103320
rect 578330 103264 578386 103300
rect 578514 101632 578570 101688
rect 579158 99220 579160 99240
rect 579160 99220 579212 99240
rect 579212 99220 579214 99240
rect 579158 99184 579214 99220
rect 578330 97416 578386 97472
rect 574742 54984 574798 55040
rect 579158 93064 579214 93120
rect 578514 90888 578570 90944
rect 578514 88032 578570 88088
rect 578330 86400 578386 86456
rect 578514 82184 578570 82240
rect 578514 77832 578570 77888
rect 579526 95004 579528 95024
rect 579528 95004 579580 95024
rect 579580 95004 579582 95024
rect 579526 94968 579582 95004
rect 579526 83988 579528 84008
rect 579528 83988 579580 84008
rect 579580 83988 579582 84008
rect 579526 83952 579582 83988
rect 579342 80008 579398 80064
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 666650 178472 666706 178528
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 580446 77832 580502 77888
rect 579066 75656 579122 75712
rect 578514 71168 578570 71224
rect 575478 54168 575534 54224
rect 578514 56072 578570 56128
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579526 64504 579582 64560
rect 579526 61784 579582 61840
rect 579526 60288 579582 60344
rect 579342 57840 579398 57896
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590290 134544 590346 134600
rect 588726 132912 588782 132968
rect 667018 159976 667074 160032
rect 667386 181328 667442 181384
rect 667202 141344 667258 141400
rect 670146 529896 670202 529952
rect 670882 647264 670938 647320
rect 672170 938032 672226 938088
rect 672722 937760 672778 937816
rect 672170 937216 672226 937272
rect 672722 937216 672778 937272
rect 672354 936672 672410 936728
rect 671986 929464 672042 929520
rect 671802 760008 671858 760064
rect 671802 757424 671858 757480
rect 672170 759736 672226 759792
rect 671986 732808 672042 732864
rect 671986 730088 672042 730144
rect 671802 712816 671858 712872
rect 671618 705472 671674 705528
rect 671802 687384 671858 687440
rect 671618 670248 671674 670304
rect 671526 668616 671582 668672
rect 671250 661272 671306 661328
rect 671618 625096 671674 625152
rect 671618 624688 671674 624744
rect 671434 624280 671490 624336
rect 671250 623872 671306 623928
rect 671066 623464 671122 623520
rect 671066 622240 671122 622296
rect 671066 594768 671122 594824
rect 670882 574776 670938 574832
rect 670882 552064 670938 552120
rect 671434 623056 671490 623112
rect 672538 935720 672594 935776
rect 672354 758648 672410 758704
rect 672998 933408 673054 933464
rect 674102 957072 674158 957128
rect 673366 932592 673422 932648
rect 673182 930552 673238 930608
rect 675758 965096 675814 965152
rect 675298 964688 675354 964744
rect 675482 963328 675538 963384
rect 675482 962784 675538 962840
rect 674470 959384 674526 959440
rect 674930 959112 674986 959168
rect 674654 958840 674710 958896
rect 674470 933816 674526 933872
rect 674286 933000 674342 933056
rect 674838 953400 674894 953456
rect 674654 930960 674710 931016
rect 674102 930144 674158 930200
rect 675390 959384 675446 959440
rect 675206 958840 675262 958896
rect 675298 958160 675354 958216
rect 675298 957752 675354 957808
rect 675758 957752 675814 957808
rect 675482 957072 675538 957128
rect 675758 956392 675814 956448
rect 675390 953400 675446 953456
rect 675482 952176 675538 952232
rect 675206 951496 675262 951552
rect 675850 951496 675906 951552
rect 683302 950680 683358 950736
rect 675298 949184 675354 949240
rect 679622 948776 679678 948832
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 679622 935584 679678 935640
rect 682382 935176 682438 935232
rect 675482 934632 675538 934688
rect 675114 934224 675170 934280
rect 683486 947280 683542 947336
rect 683486 939664 683542 939720
rect 683302 932320 683358 932376
rect 683118 929056 683174 929112
rect 673182 928240 673238 928296
rect 672998 869352 673054 869408
rect 672814 784352 672870 784408
rect 672722 780544 672778 780600
rect 672446 757832 672502 757888
rect 672354 734168 672410 734224
rect 672170 715264 672226 715320
rect 672170 689016 672226 689072
rect 671986 665624 672042 665680
rect 671986 661000 672042 661056
rect 671802 618160 671858 618216
rect 671526 580760 671582 580816
rect 671434 579264 671490 579320
rect 671250 578856 671306 578912
rect 671434 577768 671490 577824
rect 671618 577496 671674 577552
rect 671434 576816 671490 576872
rect 671250 534656 671306 534712
rect 671434 533024 671490 533080
rect 671802 577224 671858 577280
rect 671802 569472 671858 569528
rect 671618 531392 671674 531448
rect 671066 524864 671122 524920
rect 670882 483928 670938 483984
rect 670606 455776 670662 455832
rect 670422 455232 670478 455288
rect 675114 876832 675170 876888
rect 675114 876288 675170 876344
rect 675666 875880 675722 875936
rect 675758 874112 675814 874168
rect 674930 873432 674986 873488
rect 675114 873160 675170 873216
rect 675114 872208 675170 872264
rect 675574 872208 675630 872264
rect 673918 864728 673974 864784
rect 673734 779184 673790 779240
rect 673550 777416 673606 777472
rect 673274 760280 673330 760336
rect 673366 759056 673422 759112
rect 672998 751712 673054 751768
rect 673918 771976 673974 772032
rect 675114 869352 675170 869408
rect 674930 869080 674986 869136
rect 674654 868672 674710 868728
rect 674654 868400 674710 868456
rect 674470 788024 674526 788080
rect 674286 778640 674342 778696
rect 674102 754296 674158 754352
rect 673826 741648 673882 741704
rect 673182 732944 673238 733000
rect 673090 728476 673146 728512
rect 673090 728456 673092 728476
rect 673092 728456 673144 728476
rect 673144 728456 673146 728476
rect 672906 725464 672962 725520
rect 672906 714856 672962 714912
rect 672630 710368 672686 710424
rect 672630 709144 672686 709200
rect 672814 669432 672870 669488
rect 672538 667392 672594 667448
rect 672722 666576 672778 666632
rect 672354 662768 672410 662824
rect 672538 647808 672594 647864
rect 672170 616528 672226 616584
rect 672262 607280 672318 607336
rect 674102 728628 674104 728648
rect 674104 728628 674156 728648
rect 674156 728628 674158 728648
rect 674102 728592 674158 728628
rect 673918 728204 673974 728240
rect 673918 728184 673920 728204
rect 673920 728184 673972 728204
rect 673972 728184 673974 728204
rect 674148 727912 674204 727968
rect 675298 868400 675354 868456
rect 674930 866632 674986 866688
rect 675114 864728 675170 864784
rect 675114 789384 675170 789440
rect 675298 788024 675354 788080
rect 674838 780816 674894 780872
rect 675390 784352 675446 784408
rect 675482 783808 675538 783864
rect 675390 782992 675446 783048
rect 675482 782448 675538 782504
rect 675482 780544 675538 780600
rect 675298 779184 675354 779240
rect 675206 778912 675262 778968
rect 675482 778640 675538 778696
rect 675482 777416 675538 777472
rect 674838 775648 674894 775704
rect 674838 774560 674894 774616
rect 675482 776464 675538 776520
rect 675390 774968 675446 775024
rect 675482 774560 675538 774616
rect 674654 770616 674710 770672
rect 674930 766536 674986 766592
rect 683210 771976 683266 772032
rect 678242 771432 678298 771488
rect 676126 766536 676182 766592
rect 676034 763000 676090 763056
rect 676586 761732 676642 761788
rect 676954 761776 677010 761832
rect 676034 760688 676090 760744
rect 676034 756336 676090 756392
rect 675850 754316 675906 754352
rect 675850 754296 675852 754316
rect 675852 754296 675904 754316
rect 675904 754296 675906 754316
rect 676034 753752 676090 753808
rect 682382 768712 682438 768768
rect 678242 757016 678298 757072
rect 683394 770616 683450 770672
rect 683210 756608 683266 756664
rect 682382 755792 682438 755848
rect 676954 754976 677010 755032
rect 676034 752528 676090 752584
rect 683394 752936 683450 752992
rect 683118 752120 683174 752176
rect 674286 726824 674342 726880
rect 675114 743144 675170 743200
rect 675298 742464 675354 742520
rect 675114 742192 675170 742248
rect 675114 741104 675170 741160
rect 675482 741648 675538 741704
rect 674930 738928 674986 738984
rect 675390 738656 675446 738712
rect 675114 738112 675170 738168
rect 674930 735256 674986 735312
rect 675114 734848 675170 734904
rect 675114 734168 675170 734224
rect 675114 733624 675170 733680
rect 675298 732944 675354 733000
rect 674930 731448 674986 731504
rect 675298 730496 675354 730552
rect 675114 730088 675170 730144
rect 683118 726824 683174 726880
rect 674562 726552 674618 726608
rect 681002 725736 681058 725792
rect 673642 723968 673698 724024
rect 677322 723968 677378 724024
rect 673366 714448 673422 714504
rect 673274 712408 673330 712464
rect 673366 705064 673422 705120
rect 673090 661544 673146 661600
rect 672998 648624 673054 648680
rect 672722 635432 672778 635488
rect 672630 608640 672686 608696
rect 672446 571920 672502 571976
rect 672814 578584 672870 578640
rect 672354 535064 672410 535120
rect 673182 644000 673238 644056
rect 672998 573144 673054 573200
rect 681002 710776 681058 710832
rect 683394 726416 683450 726472
rect 683578 725464 683634 725520
rect 683394 711184 683450 711240
rect 683578 708328 683634 708384
rect 683854 707920 683910 707976
rect 683118 706696 683174 706752
rect 675114 701120 675170 701176
rect 673826 690104 673882 690160
rect 673642 682352 673698 682408
rect 673550 644816 673606 644872
rect 673826 636792 673882 636848
rect 673458 599664 673514 599720
rect 675114 696904 675170 696960
rect 675390 696768 675446 696824
rect 675666 694320 675722 694376
rect 674194 666168 674250 666224
rect 674194 665080 674250 665136
rect 674654 689560 674710 689616
rect 675114 692824 675170 692880
rect 675390 690104 675446 690160
rect 675298 689560 675354 689616
rect 674194 642368 674250 642424
rect 674194 641688 674250 641744
rect 674010 619112 674066 619168
rect 673918 603472 673974 603528
rect 673734 597896 673790 597952
rect 673458 597352 673514 597408
rect 673182 571104 673238 571160
rect 672998 570288 673054 570344
rect 672814 534248 672870 534304
rect 672814 532752 672870 532808
rect 672722 531936 672778 531992
rect 672538 531664 672594 531720
rect 672170 529080 672226 529136
rect 671986 501608 672042 501664
rect 672446 490864 672502 490920
rect 672446 489640 672502 489696
rect 672262 454960 672318 455016
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 669962 403688 670018 403744
rect 670606 393488 670662 393544
rect 670422 347248 670478 347304
rect 668582 311888 668638 311944
rect 669226 302232 669282 302288
rect 667938 223080 667994 223136
rect 667938 221992 667994 222048
rect 667938 220904 667994 220960
rect 668030 202408 668086 202464
rect 667938 199180 667940 199200
rect 667940 199180 667992 199200
rect 667992 199180 667994 199200
rect 667938 199144 667994 199180
rect 668122 198736 668178 198792
rect 667938 194284 667940 194304
rect 667940 194284 667992 194304
rect 667992 194284 667994 194304
rect 667938 194248 667994 194284
rect 667938 189388 667940 189408
rect 667940 189388 667992 189408
rect 667992 189388 667994 189408
rect 667938 189352 667994 189388
rect 668122 187584 668178 187640
rect 668122 184864 668178 184920
rect 667754 178744 667810 178800
rect 667938 174700 667940 174720
rect 667940 174700 667992 174720
rect 667992 174700 667994 174720
rect 667938 174664 667994 174700
rect 667938 169668 667940 169688
rect 667940 169668 667992 169688
rect 667992 169668 667994 169688
rect 667938 169632 667994 169668
rect 668490 234232 668546 234288
rect 668306 182824 668362 182880
rect 668122 168136 668178 168192
rect 668306 150220 668308 150240
rect 668308 150220 668360 150240
rect 668360 150220 668362 150240
rect 668306 150184 668362 150220
rect 670146 264016 670202 264072
rect 669962 259528 670018 259584
rect 669962 245792 670018 245848
rect 670146 235864 670202 235920
rect 669594 232736 669650 232792
rect 669410 225664 669466 225720
rect 669318 225256 669374 225312
rect 669410 223624 669466 223680
rect 669410 216552 669466 216608
rect 669226 215600 669282 215656
rect 669226 214512 669282 214568
rect 670054 233144 670110 233200
rect 669318 202544 669374 202600
rect 669226 201592 669282 201648
rect 668950 192616 669006 192672
rect 669226 184492 669228 184512
rect 669228 184492 669280 184512
rect 669280 184492 669282 184512
rect 669226 184456 669282 184492
rect 669134 167048 669190 167104
rect 668950 163240 669006 163296
rect 668766 153448 668822 153504
rect 668766 153040 668822 153096
rect 668490 148552 668546 148608
rect 667938 137400 667994 137456
rect 667570 135904 667626 135960
rect 667938 135496 667994 135552
rect 666834 133048 666890 133104
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 589646 129648 589702 129704
rect 589462 128016 589518 128072
rect 590106 126384 590162 126440
rect 589922 124752 589978 124808
rect 589462 123120 589518 123176
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 589462 119856 589518 119912
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 589462 113328 589518 113384
rect 589370 111696 589426 111752
rect 669686 214512 669742 214568
rect 669686 200504 669742 200560
rect 673182 559000 673238 559056
rect 672998 500928 673054 500984
rect 672814 489232 672870 489288
rect 672630 488416 672686 488472
rect 672630 488008 672686 488064
rect 672446 401648 672502 401704
rect 673182 484744 673238 484800
rect 673090 457000 673146 457056
rect 674010 596536 674066 596592
rect 673734 582528 673790 582584
rect 673550 580352 673606 580408
rect 673642 547032 673698 547088
rect 674930 689288 674986 689344
rect 675114 689016 675170 689072
rect 674930 688744 674986 688800
rect 674930 687112 674986 687168
rect 675482 687384 675538 687440
rect 675206 685888 675262 685944
rect 675482 685480 675538 685536
rect 675022 670112 675078 670168
rect 675022 669160 675078 669216
rect 674838 666168 674894 666224
rect 674838 665624 674894 665680
rect 674838 664672 674894 664728
rect 674838 664128 674894 664184
rect 674838 663040 674894 663096
rect 674838 662496 674894 662552
rect 674838 661816 674894 661872
rect 674838 661272 674894 661328
rect 683210 682352 683266 682408
rect 676494 673104 676550 673160
rect 676494 671064 676550 671120
rect 683394 680992 683450 681048
rect 683210 666984 683266 667040
rect 683394 663720 683450 663776
rect 675390 654200 675446 654256
rect 675574 652840 675630 652896
rect 675574 651480 675630 651536
rect 675482 648896 675538 648952
rect 675482 648624 675538 648680
rect 675482 647808 675538 647864
rect 675298 647264 675354 647320
rect 674792 645768 674848 645824
rect 675482 644816 675538 644872
rect 675758 644272 675814 644328
rect 675482 644000 675538 644056
rect 675298 643456 675354 643512
rect 674746 637744 674802 637800
rect 675298 641688 675354 641744
rect 675206 641280 675262 641336
rect 675298 639376 675354 639432
rect 675482 638560 675538 638616
rect 675574 637880 675630 637936
rect 674930 635976 674986 636032
rect 674930 635704 674986 635760
rect 674838 631352 674894 631408
rect 675206 631352 675262 631408
rect 682382 637608 682438 637664
rect 675574 631352 675630 631408
rect 675390 629720 675446 629776
rect 675206 629448 675262 629504
rect 676494 628496 676550 628552
rect 674654 619520 674710 619576
rect 674470 617752 674526 617808
rect 674838 608640 674894 608696
rect 674838 607008 674894 607064
rect 674470 604560 674526 604616
rect 674194 591232 674250 591288
rect 674194 558320 674250 558376
rect 673918 545672 673974 545728
rect 674010 535336 674066 535392
rect 674010 533976 674066 534032
rect 674010 533432 674066 533488
rect 673826 528264 673882 528320
rect 673550 526904 673606 526960
rect 674010 490048 674066 490104
rect 676494 625640 676550 625696
rect 683394 636792 683450 636848
rect 683210 635432 683266 635488
rect 683210 622784 683266 622840
rect 682382 621968 682438 622024
rect 676494 621560 676550 621616
rect 676494 621152 676550 621208
rect 676494 620336 676550 620392
rect 676494 619928 676550 619984
rect 677230 619520 677286 619576
rect 677230 619112 677286 619168
rect 683118 619112 683174 619168
rect 683118 617480 683174 617536
rect 683762 635704 683818 635760
rect 683762 618704 683818 618760
rect 683394 617072 683450 617128
rect 675482 607824 675538 607880
rect 675298 607280 675354 607336
rect 675298 607008 675354 607064
rect 675298 604560 675354 604616
rect 675298 604288 675354 604344
rect 675482 603472 675538 603528
rect 675298 602928 675354 602984
rect 675482 600344 675538 600400
rect 675298 599664 675354 599720
rect 675206 599256 675262 599312
rect 674746 592320 674802 592376
rect 675390 597352 675446 597408
rect 675390 596808 675446 596864
rect 675206 596536 675262 596592
rect 675482 594768 675538 594824
rect 675482 593544 675538 593600
rect 675574 593136 675630 593192
rect 675114 581576 675170 581632
rect 676034 592864 676090 592920
rect 675850 592320 675906 592376
rect 675574 586200 675630 586256
rect 675850 581576 675906 581632
rect 675022 580760 675078 580816
rect 675022 579808 675078 579864
rect 675022 577632 675078 577688
rect 675022 576816 675078 576872
rect 674838 559408 674894 559464
rect 674654 548256 674710 548312
rect 675482 578312 675538 578368
rect 675482 576952 675538 577008
rect 683118 592592 683174 592648
rect 676034 576544 676090 576600
rect 675850 575320 675906 575376
rect 683394 591232 683450 591288
rect 683670 589872 683726 589928
rect 683670 573960 683726 574016
rect 683394 573144 683450 573200
rect 683118 571920 683174 571976
rect 682382 570696 682438 570752
rect 675390 564440 675446 564496
rect 675574 562672 675630 562728
rect 675482 561176 675538 561232
rect 675482 559408 675538 559464
rect 675390 559000 675446 559056
rect 675390 558320 675446 558376
rect 675482 557504 675538 557560
rect 675758 557504 675814 557560
rect 675390 554648 675446 554704
rect 675758 553832 675814 553888
rect 675390 553424 675446 553480
rect 675390 552064 675446 552120
rect 675390 551520 675446 551576
rect 675206 550568 675262 550624
rect 675758 550296 675814 550352
rect 675390 548256 675446 548312
rect 674838 546216 674894 546272
rect 674838 545944 674894 546000
rect 674562 532208 674618 532264
rect 674562 531392 674618 531448
rect 674378 530576 674434 530632
rect 674562 529352 674618 529408
rect 674562 528536 674618 528592
rect 675942 547612 675944 547632
rect 675944 547612 675996 547632
rect 675996 547612 675998 547632
rect 675942 547576 675998 547612
rect 677414 547576 677470 547632
rect 675390 546216 675446 546272
rect 675206 545400 675262 545456
rect 676494 538736 676550 538792
rect 676494 535880 676550 535936
rect 675758 535064 675814 535120
rect 675758 534452 675814 534508
rect 675022 510176 675078 510232
rect 675206 503648 675262 503704
rect 675022 503104 675078 503160
rect 675390 503104 675446 503160
rect 675850 510176 675906 510232
rect 675850 503668 675906 503704
rect 675850 503648 675852 503668
rect 675852 503648 675904 503668
rect 675904 503648 675906 503668
rect 675666 500928 675722 500984
rect 675114 487600 675170 487656
rect 675574 490456 675630 490512
rect 675298 486376 675354 486432
rect 674746 485560 674802 485616
rect 674194 484336 674250 484392
rect 675758 481888 675814 481944
rect 673826 456068 673882 456104
rect 673826 456048 673828 456068
rect 673828 456048 673880 456068
rect 673880 456048 673882 456068
rect 673734 455796 673790 455832
rect 673734 455776 673736 455796
rect 673736 455776 673788 455796
rect 673788 455776 673790 455796
rect 673596 455540 673598 455560
rect 673598 455540 673650 455560
rect 673650 455540 673652 455560
rect 673596 455504 673652 455540
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 672906 454824 672962 454880
rect 673162 454588 673164 454608
rect 673164 454588 673216 454608
rect 673216 454588 673218 454608
rect 673162 454552 673218 454588
rect 672814 454180 672816 454200
rect 672816 454180 672868 454200
rect 672868 454180 672870 454200
rect 672814 454144 672870 454180
rect 675482 479984 675538 480040
rect 676402 474816 676458 474872
rect 676126 457000 676182 457056
rect 676402 456048 676458 456104
rect 675850 455540 675852 455560
rect 675852 455540 675904 455560
rect 675904 455540 675906 455560
rect 675850 455504 675906 455540
rect 677046 501608 677102 501664
rect 683210 547032 683266 547088
rect 682382 546760 682438 546816
rect 678242 531392 678298 531448
rect 682382 530984 682438 531040
rect 683394 545672 683450 545728
rect 683210 528128 683266 528184
rect 683578 533840 683634 533896
rect 683578 527312 683634 527368
rect 683394 526496 683450 526552
rect 683118 525680 683174 525736
rect 677874 524456 677930 524512
rect 683578 503648 683634 503704
rect 683394 503376 683450 503432
rect 679622 486784 679678 486840
rect 683118 494672 683174 494728
rect 683118 491272 683174 491328
rect 683578 487192 683634 487248
rect 683394 483520 683450 483576
rect 683118 483112 683174 483168
rect 681002 481480 681058 481536
rect 676862 454824 676918 454880
rect 676034 454552 676090 454608
rect 675574 454144 675630 454200
rect 674746 453872 674802 453928
rect 674930 453872 674986 453928
rect 683302 411848 683358 411904
rect 676034 410488 676090 410544
rect 683118 406272 683174 406328
rect 683302 403688 683358 403744
rect 683118 403280 683174 403336
rect 676034 402600 676090 402656
rect 674654 402192 674710 402248
rect 674194 401376 674250 401432
rect 673274 400424 673330 400480
rect 672630 400016 672686 400072
rect 672538 398792 672594 398848
rect 672170 392264 672226 392320
rect 671986 348880 672042 348936
rect 671986 329704 672042 329760
rect 671342 275304 671398 275360
rect 671710 261976 671766 262032
rect 671526 259120 671582 259176
rect 671342 257896 671398 257952
rect 671986 256672 672042 256728
rect 671710 244976 671766 245032
rect 671526 242800 671582 242856
rect 671342 241440 671398 241496
rect 672722 397160 672778 397216
rect 673090 394168 673146 394224
rect 672906 393896 672962 393952
rect 672722 377848 672778 377904
rect 672906 376896 672962 376952
rect 673090 376216 673146 376272
rect 672722 357040 672778 357096
rect 672538 355000 672594 355056
rect 672538 352144 672594 352200
rect 672354 349696 672410 349752
rect 672538 335824 672594 335880
rect 672354 335552 672410 335608
rect 674010 396072 674066 396128
rect 673826 395664 673882 395720
rect 673458 378120 673514 378176
rect 673274 355816 673330 355872
rect 673274 355408 673330 355464
rect 673090 354592 673146 354648
rect 672906 352552 672962 352608
rect 672906 333920 672962 333976
rect 672906 312704 672962 312760
rect 672722 312432 672778 312488
rect 672446 304680 672502 304736
rect 672630 304272 672686 304328
rect 672446 290128 672502 290184
rect 673274 310800 673330 310856
rect 673090 309984 673146 310040
rect 673090 309576 673146 309632
rect 672630 287816 672686 287872
rect 672814 267280 672870 267336
rect 672538 265648 672594 265704
rect 671986 238040 672042 238096
rect 670790 233552 670846 233608
rect 671158 233144 671214 233200
rect 670974 225392 671030 225448
rect 670974 224732 671030 224768
rect 670974 224712 670976 224732
rect 670976 224712 671028 224732
rect 671028 224712 671030 224732
rect 670928 224188 670984 224224
rect 670928 224168 670930 224188
rect 670930 224168 670982 224188
rect 670982 224168 670984 224188
rect 670790 223896 670846 223952
rect 670606 213968 670662 214024
rect 670606 211384 670662 211440
rect 670422 211112 670478 211168
rect 671894 234776 671950 234832
rect 672078 234504 672134 234560
rect 671710 234232 671766 234288
rect 671526 230016 671582 230072
rect 671894 226888 671950 226944
rect 673274 303456 673330 303512
rect 673090 264968 673146 265024
rect 672906 263744 672962 263800
rect 673090 260344 673146 260400
rect 672722 257080 672778 257136
rect 674010 381384 674066 381440
rect 673826 375400 673882 375456
rect 674378 396480 674434 396536
rect 674378 382200 674434 382256
rect 676034 399336 676090 399392
rect 674838 394440 674894 394496
rect 674838 393896 674894 393952
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 683026 392672 683082 392728
rect 683026 389000 683082 389056
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675114 377984 675170 378040
rect 675758 377304 675814 377360
rect 675298 376896 675354 376952
rect 675390 376216 675446 376272
rect 675298 375400 675354 375456
rect 675666 372952 675722 373008
rect 675114 372544 675170 372600
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 357448 674710 357504
rect 674194 356632 674250 356688
rect 674194 356224 674250 356280
rect 673642 353368 673698 353424
rect 673826 350512 673882 350568
rect 673642 340720 673698 340776
rect 674010 349424 674066 349480
rect 674010 332696 674066 332752
rect 673826 331064 673882 331120
rect 675850 351736 675906 351792
rect 674746 351328 674802 351384
rect 674562 347656 674618 347712
rect 675850 350240 675906 350296
rect 676034 350104 676090 350160
rect 676034 346568 676090 346624
rect 675114 340720 675170 340776
rect 675758 340312 675814 340368
rect 675666 339360 675722 339416
rect 675390 337184 675446 337240
rect 675758 336504 675814 336560
rect 675114 335552 675170 335608
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675758 332288 675814 332344
rect 675298 331064 675354 331120
rect 675114 329704 675170 329760
rect 675758 328344 675814 328400
rect 675390 326848 675446 326904
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 312976 674710 313032
rect 674838 312704 674894 312760
rect 674838 312024 674894 312080
rect 674654 311888 674710 311944
rect 674194 311616 674250 311672
rect 674654 311208 674710 311264
rect 674286 310392 674342 310448
rect 674102 305496 674158 305552
rect 674102 285504 674158 285560
rect 674010 267008 674066 267064
rect 673826 260888 673882 260944
rect 673642 258440 673698 258496
rect 673458 246200 673514 246256
rect 673182 245248 673238 245304
rect 672722 237360 672778 237416
rect 672630 236408 672686 236464
rect 672262 231512 672318 231568
rect 672354 227024 672410 227080
rect 671818 226616 671874 226672
rect 671940 226344 671996 226400
rect 672032 226108 672034 226128
rect 672034 226108 672086 226128
rect 672086 226108 672088 226128
rect 672032 226072 672088 226108
rect 671710 225800 671766 225856
rect 671818 225700 671820 225720
rect 671820 225700 671872 225720
rect 671872 225700 671874 225720
rect 671818 225664 671874 225700
rect 671594 225120 671650 225176
rect 671618 224032 671674 224088
rect 671434 221448 671490 221504
rect 671986 225392 672042 225448
rect 671986 225120 672042 225176
rect 672078 224712 672134 224768
rect 670606 190304 670662 190360
rect 670606 171944 670662 172000
rect 669778 169496 669834 169552
rect 669502 164872 669558 164928
rect 670146 168272 670202 168328
rect 669778 154808 669834 154864
rect 669134 143656 669190 143712
rect 669042 142160 669098 142216
rect 669042 138760 669098 138816
rect 668950 128152 669006 128208
rect 668766 125704 668822 125760
rect 669226 122168 669282 122224
rect 668950 120808 669006 120864
rect 668582 120536 668638 120592
rect 667938 119176 667994 119232
rect 668030 117544 668086 117600
rect 590382 114960 590438 115016
rect 670330 165552 670386 165608
rect 671894 221176 671950 221232
rect 672378 226480 672434 226536
rect 673526 237088 673582 237144
rect 673826 246472 673882 246528
rect 674470 303864 674526 303920
rect 674470 286592 674526 286648
rect 675022 309168 675078 309224
rect 674838 307944 674894 308000
rect 676034 308352 676090 308408
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 678978 306312 679034 306368
rect 683026 302640 683082 302696
rect 683026 299376 683082 299432
rect 678242 297336 678298 297392
rect 676034 296792 676090 296848
rect 675850 296520 675906 296576
rect 675758 295160 675814 295216
rect 674838 292848 674894 292904
rect 675390 292848 675446 292904
rect 675574 292032 675630 292088
rect 675758 291488 675814 291544
rect 675390 290128 675446 290184
rect 675298 289856 675354 289912
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286592 675446 286648
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281152 675722 281208
rect 683302 275304 683358 275360
rect 683118 271088 683174 271144
rect 683302 268504 683358 268560
rect 683118 268096 683174 268152
rect 674654 266600 674710 266656
rect 674286 266056 674342 266112
rect 676494 266056 676550 266112
rect 674562 265240 674618 265296
rect 676494 265240 676550 265296
rect 674838 264424 674894 264480
rect 676494 264016 676550 264072
rect 674838 263744 674894 263800
rect 676494 263608 676550 263664
rect 678242 263200 678298 263256
rect 676218 262792 676274 262848
rect 675942 258712 675998 258768
rect 675942 258168 675998 258224
rect 675298 257488 675354 257544
rect 675298 256672 675354 256728
rect 675206 255856 675262 255912
rect 676126 255856 676182 255912
rect 674286 249600 674342 249656
rect 673642 236444 673644 236464
rect 673644 236444 673696 236464
rect 673696 236444 673698 236464
rect 673642 236408 673698 236444
rect 672814 228792 672870 228848
rect 672814 228540 672870 228576
rect 672814 228520 672816 228540
rect 672816 228520 672868 228540
rect 672868 228520 672870 228540
rect 674424 235084 674426 235104
rect 674426 235084 674478 235104
rect 674478 235084 674480 235104
rect 674424 235048 674480 235084
rect 674286 234776 674342 234832
rect 673734 232736 673790 232792
rect 673642 232464 673698 232520
rect 673458 230016 673514 230072
rect 673918 230424 673974 230480
rect 674534 234116 674590 234152
rect 674534 234096 674536 234116
rect 674536 234096 674588 234116
rect 674588 234096 674590 234116
rect 675022 251776 675078 251832
rect 674930 249328 674986 249384
rect 679622 261160 679678 261216
rect 676034 251776 676090 251832
rect 675758 250280 675814 250336
rect 675390 249600 675446 249656
rect 674930 245520 674986 245576
rect 675390 246472 675446 246528
rect 675390 245792 675446 245848
rect 675114 242800 675170 242856
rect 675114 241440 675170 241496
rect 675390 240216 675446 240272
rect 675390 238040 675446 238096
rect 675206 237224 675262 237280
rect 675022 235864 675078 235920
rect 675850 234116 675906 234152
rect 675850 234096 675852 234116
rect 675852 234096 675904 234116
rect 675904 234096 675906 234116
rect 675114 233552 675170 233608
rect 674654 231784 674710 231840
rect 674654 231512 674710 231568
rect 674730 231004 674732 231024
rect 674732 231004 674784 231024
rect 674784 231004 674786 231024
rect 674730 230968 674786 231004
rect 675850 231532 675906 231568
rect 675850 231512 675852 231532
rect 675852 231512 675904 231532
rect 675904 231512 675906 231532
rect 675068 231240 675124 231296
rect 674838 230696 674894 230752
rect 675022 230696 675078 230752
rect 675850 230696 675906 230752
rect 674394 230118 674450 230174
rect 674654 230152 674710 230208
rect 676218 230424 676274 230480
rect 673826 229744 673882 229800
rect 674170 229916 674172 229936
rect 674172 229916 674224 229936
rect 674224 229916 674226 229936
rect 674170 229880 674226 229916
rect 673642 229472 673698 229528
rect 673946 229508 673948 229528
rect 673948 229508 674000 229528
rect 674000 229508 674002 229528
rect 673946 229472 674002 229508
rect 673918 229200 673974 229256
rect 673734 229100 673736 229120
rect 673736 229100 673788 229120
rect 673788 229100 673790 229120
rect 673734 229064 673790 229100
rect 673182 226752 673238 226808
rect 672722 224576 672778 224632
rect 672906 224032 672962 224088
rect 672722 223896 672778 223952
rect 672446 221856 672502 221912
rect 672906 220904 672962 220960
rect 672722 219136 672778 219192
rect 672078 217232 672134 217288
rect 672078 213696 672134 213752
rect 672538 213968 672594 214024
rect 673458 226072 673514 226128
rect 673918 226208 673974 226264
rect 673918 225528 673974 225584
rect 673734 225392 673790 225448
rect 673274 224576 673330 224632
rect 672078 200776 672134 200832
rect 672262 198736 672318 198792
rect 672446 184864 672502 184920
rect 672078 183504 672134 183560
rect 671894 176432 671950 176488
rect 671710 173032 671766 173088
rect 671894 169904 671950 169960
rect 671710 166912 671766 166968
rect 671526 158344 671582 158400
rect 670606 148960 670662 149016
rect 671342 131688 671398 131744
rect 669226 114280 669282 114336
rect 671526 130872 671582 130928
rect 668582 111016 668638 111072
rect 668122 110744 668178 110800
rect 590106 110064 590162 110120
rect 589462 108432 589518 108488
rect 589646 106800 589702 106856
rect 589462 105168 589518 105224
rect 589922 101904 589978 101960
rect 666834 106088 666836 106108
rect 666836 106088 666888 106108
rect 666888 106088 666890 106108
rect 590290 103536 590346 103592
rect 612002 95784 612058 95840
rect 635554 96328 635610 96384
rect 635738 96056 635794 96112
rect 637026 96872 637082 96928
rect 641994 96056 642050 96112
rect 647422 96328 647478 96384
rect 647146 94968 647202 95024
rect 626446 94424 626502 94480
rect 625986 93608 626042 93664
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 626262 89528 626318 89584
rect 626446 88712 626502 88768
rect 626446 87896 626502 87952
rect 625618 87080 625674 87136
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 584402 54712 584458 54768
rect 581642 54440 581698 54496
rect 577686 53896 577742 53952
rect 459466 53624 459522 53680
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 308034 48864 308090 48920
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 458362 46688 458418 46744
rect 431222 44784 431278 44840
rect 142618 44240 142674 44296
rect 307298 44104 307354 44160
rect 194322 42064 194378 42120
rect 419722 43832 419778 43888
rect 415398 43560 415454 43616
rect 456062 43832 456118 43888
rect 439594 43596 439596 43616
rect 439596 43596 439648 43616
rect 439648 43596 439650 43616
rect 439594 43560 439650 43596
rect 441618 43596 441620 43616
rect 441620 43596 441672 43616
rect 441672 43596 441674 43616
rect 441618 43560 441674 43596
rect 456062 43288 456118 43344
rect 361946 41792 362002 41848
rect 365166 41792 365222 41848
rect 416686 42200 416742 42256
rect 446402 42200 446458 42256
rect 446402 41520 446458 41576
rect 460110 44784 460166 44840
rect 460754 43016 460810 43072
rect 461950 43832 462006 43888
rect 462686 43832 462742 43888
rect 461766 43560 461822 43616
rect 462870 43288 462926 43344
rect 463698 44376 463754 44432
rect 549994 48864 550050 48920
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 626446 83816 626502 83872
rect 628746 83272 628802 83328
rect 629206 81640 629262 81696
rect 625986 75928 626042 75984
rect 633898 77560 633954 77616
rect 633898 75928 633954 75984
rect 639602 77832 639658 77888
rect 646318 74160 646374 74216
rect 646502 71712 646558 71768
rect 646134 69128 646190 69184
rect 647238 64368 647294 64424
rect 646134 59336 646190 59392
rect 648618 91976 648674 92032
rect 650274 89528 650330 89584
rect 650550 87080 650606 87136
rect 655058 94152 655114 94208
rect 654690 91432 654746 91488
rect 655426 93336 655482 93392
rect 655426 90652 655428 90672
rect 655428 90652 655480 90672
rect 655480 90652 655482 90672
rect 655426 90616 655482 90652
rect 655794 89800 655850 89856
rect 663706 92792 663762 92848
rect 664166 90616 664222 90672
rect 664534 91704 664590 91760
rect 664350 89800 664406 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 649998 84632 650054 84688
rect 648894 82184 648950 82240
rect 666834 106052 666890 106088
rect 668398 109248 668454 109304
rect 668122 104352 668178 104408
rect 667938 102720 667994 102776
rect 671894 151816 671950 151872
rect 672814 210296 672870 210352
rect 672630 153040 672686 153096
rect 672078 140392 672134 140448
rect 672354 125568 672410 125624
rect 671710 115776 671766 115832
rect 673366 221856 673422 221912
rect 673182 218320 673238 218376
rect 672998 177928 673054 177984
rect 673550 219816 673606 219872
rect 673550 219408 673606 219464
rect 673366 177248 673422 177304
rect 673366 176840 673422 176896
rect 673182 176024 673238 176080
rect 672998 169088 673054 169144
rect 672998 152496 673054 152552
rect 673918 223624 673974 223680
rect 673734 214240 673790 214296
rect 673918 212880 673974 212936
rect 673734 211112 673790 211168
rect 673918 209616 673974 209672
rect 673734 203904 673790 203960
rect 673918 197376 673974 197432
rect 673550 174800 673606 174856
rect 673918 168680 673974 168736
rect 675114 229880 675170 229936
rect 675114 229200 675170 229256
rect 674838 227024 674894 227080
rect 674470 226480 674526 226536
rect 674470 223624 674526 223680
rect 674470 222672 674526 222728
rect 674286 222264 674342 222320
rect 675022 225800 675078 225856
rect 674838 221584 674894 221640
rect 675022 220496 675078 220552
rect 674654 220224 674710 220280
rect 674470 217368 674526 217424
rect 674470 198192 674526 198248
rect 674286 179424 674342 179480
rect 675114 219816 675170 219872
rect 675114 218864 675170 218920
rect 675666 225120 675722 225176
rect 675482 224304 675538 224360
rect 674838 217776 674894 217832
rect 675206 218048 675262 218104
rect 675206 216144 675262 216200
rect 675022 215328 675078 215384
rect 677046 230152 677102 230208
rect 676402 226208 676458 226264
rect 675666 215872 675722 215928
rect 676034 219816 676090 219872
rect 676034 215092 676036 215112
rect 676036 215092 676088 215112
rect 676088 215092 676090 215112
rect 676034 215056 676090 215092
rect 675666 214784 675722 214840
rect 676034 214512 676090 214568
rect 676034 213424 676090 213480
rect 676034 213152 676090 213208
rect 676770 211112 676826 211168
rect 676954 211112 677010 211168
rect 683210 233824 683266 233880
rect 683210 223080 683266 223136
rect 679806 221448 679862 221504
rect 679622 220632 679678 220688
rect 683670 222672 683726 222728
rect 683394 219816 683450 219872
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 677874 209616 677930 209672
rect 675482 207304 675538 207360
rect 675758 205536 675814 205592
rect 674838 202000 674894 202056
rect 675482 204176 675538 204232
rect 675482 202544 675538 202600
rect 675482 202000 675538 202056
rect 675114 201592 675170 201648
rect 674930 200776 674986 200832
rect 675758 200640 675814 200696
rect 675298 200504 675354 200560
rect 675482 198192 675538 198248
rect 675758 197104 675814 197160
rect 675666 195200 675722 195256
rect 675758 191528 675814 191584
rect 675298 190304 675354 190360
rect 675114 189760 675170 189816
rect 675850 181328 675906 181384
rect 676034 178744 676090 178800
rect 675850 178064 675906 178120
rect 676034 177656 676090 177712
rect 674654 175616 674710 175672
rect 674654 175208 674710 175264
rect 674378 174392 674434 174448
rect 674102 154536 674158 154592
rect 673918 151000 673974 151056
rect 673366 132096 673422 132152
rect 673182 131280 673238 131336
rect 676034 173168 676090 173224
rect 674838 172760 674894 172816
rect 675022 171128 675078 171184
rect 681002 171536 681058 171592
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 674838 157528 674894 157584
rect 675206 161336 675262 161392
rect 676586 166368 676642 166424
rect 676034 165552 676090 165608
rect 675850 161336 675906 161392
rect 675758 159296 675814 159352
rect 675482 157528 675538 157584
rect 675758 156304 675814 156360
rect 675114 154808 675170 154864
rect 675482 152496 675538 152552
rect 675482 151816 675538 151872
rect 675298 151544 675354 151600
rect 675114 151000 675170 151056
rect 675666 150320 675722 150376
rect 675298 148960 675354 149016
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 683302 141344 683358 141400
rect 683118 135904 683174 135960
rect 683302 133048 683358 133104
rect 683118 132640 683174 132696
rect 674654 130464 674710 130520
rect 676034 130056 676090 130112
rect 674378 129648 674434 129704
rect 674102 129240 674158 129296
rect 673918 125160 673974 125216
rect 673182 124344 673238 124400
rect 672814 124072 672870 124128
rect 672722 122440 672778 122496
rect 672722 112648 672778 112704
rect 672354 111288 672410 111344
rect 673366 123664 673422 123720
rect 673182 110336 673238 110392
rect 671526 107752 671582 107808
rect 673366 106800 673422 106856
rect 674286 128288 674342 128344
rect 676034 128288 676090 128344
rect 674102 111016 674158 111072
rect 673918 104624 673974 104680
rect 679622 128152 679678 128208
rect 678242 127744 678298 127800
rect 674838 127608 674894 127664
rect 674654 125976 674710 126032
rect 674470 119992 674526 120048
rect 676218 126928 676274 126984
rect 675022 126384 675078 126440
rect 676218 124888 676274 124944
rect 676678 123256 676734 123312
rect 676678 119992 676734 120048
rect 679622 117272 679678 117328
rect 675298 113056 675354 113112
rect 675390 111288 675446 111344
rect 675114 110336 675170 110392
rect 675206 108976 675262 109032
rect 675666 108024 675722 108080
rect 675482 106800 675538 106856
rect 675114 104624 675170 104680
rect 675666 103128 675722 103184
rect 675758 102448 675814 102504
rect 674286 102312 674342 102368
rect 675758 101360 675814 101416
rect 668122 95784 668178 95840
rect 648710 67088 648766 67144
rect 648894 62056 648950 62112
rect 647422 57296 647478 57352
rect 662418 48456 662474 48512
rect 661590 47733 661646 47789
rect 464342 44240 464398 44296
rect 463882 44104 463938 44160
rect 465814 43832 465870 43888
rect 463698 43560 463754 43616
rect 460938 42336 460994 42392
rect 471150 42744 471206 42800
rect 518806 42744 518862 42800
rect 662602 47368 662658 47424
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40432 141754 40488
<< metal3 >>
rect 427997 1006906 428063 1006909
rect 504541 1006906 504607 1006909
rect 559649 1006906 559715 1006909
rect 427800 1006904 428063 1006906
rect 427800 1006848 428002 1006904
rect 428058 1006848 428063 1006904
rect 427800 1006846 428063 1006848
rect 504436 1006904 504607 1006906
rect 504436 1006848 504546 1006904
rect 504602 1006848 504607 1006904
rect 504436 1006846 504607 1006848
rect 559452 1006904 559715 1006906
rect 559452 1006848 559654 1006904
rect 559710 1006848 559715 1006904
rect 559452 1006846 559715 1006848
rect 427997 1006843 428063 1006846
rect 504541 1006843 504607 1006846
rect 559649 1006843 559715 1006846
rect 428365 1006770 428431 1006773
rect 505369 1006770 505435 1006773
rect 554313 1006770 554379 1006773
rect 428365 1006768 428628 1006770
rect 428365 1006712 428370 1006768
rect 428426 1006712 428628 1006768
rect 428365 1006710 428628 1006712
rect 505172 1006768 505435 1006770
rect 505172 1006712 505374 1006768
rect 505430 1006712 505435 1006768
rect 505172 1006710 505435 1006712
rect 554116 1006768 554379 1006770
rect 554116 1006712 554318 1006768
rect 554374 1006712 554379 1006768
rect 554116 1006710 554379 1006712
rect 428365 1006707 428431 1006710
rect 505369 1006707 505435 1006710
rect 554313 1006707 554379 1006710
rect 152917 1006634 152983 1006637
rect 152720 1006632 152983 1006634
rect 152720 1006576 152922 1006632
rect 152978 1006576 152983 1006632
rect 152720 1006574 152983 1006576
rect 152917 1006571 152983 1006574
rect 308121 1006634 308187 1006637
rect 357709 1006634 357775 1006637
rect 308121 1006632 308384 1006634
rect 308121 1006576 308126 1006632
rect 308182 1006576 308384 1006632
rect 308121 1006574 308384 1006576
rect 357709 1006632 357972 1006634
rect 357709 1006576 357714 1006632
rect 357770 1006576 357972 1006632
rect 357709 1006574 357972 1006576
rect 308121 1006571 308187 1006574
rect 357709 1006571 357775 1006574
rect 103973 1006498 104039 1006501
rect 152089 1006498 152155 1006501
rect 157425 1006498 157491 1006501
rect 359733 1006498 359799 1006501
rect 431677 1006498 431743 1006501
rect 506197 1006498 506263 1006501
rect 103973 1006496 104236 1006498
rect 103973 1006440 103978 1006496
rect 104034 1006440 104236 1006496
rect 103973 1006438 104236 1006440
rect 152089 1006496 152352 1006498
rect 152089 1006440 152094 1006496
rect 152150 1006440 152352 1006496
rect 152089 1006438 152352 1006440
rect 157228 1006496 157491 1006498
rect 157228 1006440 157430 1006496
rect 157486 1006440 157491 1006496
rect 157228 1006438 157491 1006440
rect 359628 1006496 359799 1006498
rect 359628 1006440 359738 1006496
rect 359794 1006440 359799 1006496
rect 359628 1006438 359799 1006440
rect 431480 1006496 431743 1006498
rect 431480 1006440 431682 1006496
rect 431738 1006440 431743 1006496
rect 431480 1006438 431743 1006440
rect 506000 1006496 506263 1006498
rect 506000 1006440 506202 1006496
rect 506258 1006440 506263 1006496
rect 506000 1006438 506263 1006440
rect 103973 1006435 104039 1006438
rect 152089 1006435 152155 1006438
rect 157425 1006435 157491 1006438
rect 359733 1006435 359799 1006438
rect 431677 1006435 431743 1006438
rect 506197 1006435 506263 1006438
rect 555969 1006498 556035 1006501
rect 555969 1006496 556232 1006498
rect 555969 1006440 555974 1006496
rect 556030 1006440 556232 1006496
rect 555969 1006438 556232 1006440
rect 555969 1006435 556035 1006438
rect 101121 1006362 101187 1006365
rect 158253 1006362 158319 1006365
rect 210049 1006362 210115 1006365
rect 101121 1006360 101292 1006362
rect 101121 1006304 101126 1006360
rect 101182 1006304 101292 1006360
rect 101121 1006302 101292 1006304
rect 158056 1006360 158319 1006362
rect 158056 1006304 158258 1006360
rect 158314 1006304 158319 1006360
rect 158056 1006302 158319 1006304
rect 209852 1006360 210115 1006362
rect 209852 1006304 210054 1006360
rect 210110 1006304 210115 1006360
rect 209852 1006302 210115 1006304
rect 101121 1006299 101187 1006302
rect 158253 1006299 158319 1006302
rect 210049 1006299 210115 1006302
rect 254117 1006362 254183 1006365
rect 358537 1006362 358603 1006365
rect 254117 1006360 254380 1006362
rect 254117 1006304 254122 1006360
rect 254178 1006304 254380 1006360
rect 254117 1006302 254380 1006304
rect 358537 1006360 358800 1006362
rect 358537 1006304 358542 1006360
rect 358598 1006304 358800 1006360
rect 358537 1006302 358800 1006304
rect 254117 1006299 254183 1006302
rect 358537 1006299 358603 1006302
rect 98269 1006226 98335 1006229
rect 107653 1006226 107719 1006229
rect 98269 1006224 98532 1006226
rect 98269 1006168 98274 1006224
rect 98330 1006196 98532 1006224
rect 107456 1006224 107719 1006226
rect 98330 1006168 98562 1006196
rect 98269 1006166 98562 1006168
rect 107456 1006168 107658 1006224
rect 107714 1006168 107719 1006224
rect 107456 1006166 107719 1006168
rect 98269 1006163 98335 1006166
rect 98502 1006090 98562 1006166
rect 107653 1006163 107719 1006166
rect 151261 1006226 151327 1006229
rect 153745 1006226 153811 1006229
rect 160277 1006226 160343 1006229
rect 210417 1006226 210483 1006229
rect 151261 1006224 151524 1006226
rect 151261 1006168 151266 1006224
rect 151322 1006168 151524 1006224
rect 151261 1006166 151524 1006168
rect 153548 1006224 153811 1006226
rect 153548 1006168 153750 1006224
rect 153806 1006168 153811 1006224
rect 153548 1006166 153811 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 210220 1006224 210483 1006226
rect 210220 1006168 210422 1006224
rect 210478 1006168 210483 1006224
rect 210220 1006166 210483 1006168
rect 151261 1006163 151327 1006166
rect 153745 1006163 153811 1006166
rect 160277 1006163 160343 1006166
rect 210417 1006163 210483 1006166
rect 255313 1006226 255379 1006229
rect 261845 1006226 261911 1006229
rect 306097 1006226 306163 1006229
rect 361389 1006226 361455 1006229
rect 255313 1006224 255576 1006226
rect 255313 1006168 255318 1006224
rect 255374 1006168 255576 1006224
rect 255313 1006166 255576 1006168
rect 261648 1006224 261911 1006226
rect 261648 1006168 261850 1006224
rect 261906 1006168 261911 1006224
rect 261648 1006166 261911 1006168
rect 305900 1006224 306163 1006226
rect 305900 1006168 306102 1006224
rect 306158 1006168 306163 1006224
rect 305900 1006166 306163 1006168
rect 361192 1006224 361455 1006226
rect 361192 1006168 361394 1006224
rect 361450 1006168 361455 1006224
rect 361192 1006166 361455 1006168
rect 255313 1006163 255379 1006166
rect 261845 1006163 261911 1006166
rect 306097 1006163 306163 1006166
rect 361389 1006163 361455 1006166
rect 429193 1006226 429259 1006229
rect 431677 1006226 431743 1006229
rect 508221 1006226 508287 1006229
rect 557165 1006226 557231 1006229
rect 429193 1006224 429456 1006226
rect 429193 1006168 429198 1006224
rect 429254 1006168 429456 1006224
rect 429193 1006166 429456 1006168
rect 431677 1006224 431940 1006226
rect 431677 1006168 431682 1006224
rect 431738 1006168 431940 1006224
rect 431677 1006166 431940 1006168
rect 508221 1006224 508484 1006226
rect 508221 1006168 508226 1006224
rect 508282 1006168 508484 1006224
rect 508221 1006166 508484 1006168
rect 557060 1006224 557231 1006226
rect 557060 1006168 557170 1006224
rect 557226 1006168 557231 1006224
rect 557060 1006166 557231 1006168
rect 429193 1006163 429259 1006166
rect 431677 1006163 431743 1006166
rect 508221 1006163 508287 1006166
rect 557165 1006163 557231 1006166
rect 99465 1006090 99531 1006093
rect 104801 1006090 104867 1006093
rect 108481 1006090 108547 1006093
rect 98502 1006060 98900 1006090
rect 98532 1006030 98900 1006060
rect 99465 1006088 99728 1006090
rect 99465 1006032 99470 1006088
rect 99526 1006032 99728 1006088
rect 99465 1006030 99728 1006032
rect 104801 1006088 104972 1006090
rect 104801 1006032 104806 1006088
rect 104862 1006032 104972 1006088
rect 104801 1006030 104972 1006032
rect 108284 1006088 108547 1006090
rect 108284 1006032 108486 1006088
rect 108542 1006032 108547 1006088
rect 108284 1006030 108547 1006032
rect 99465 1006027 99531 1006030
rect 104801 1006027 104867 1006030
rect 108481 1006027 108547 1006030
rect 147121 1006090 147187 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 159449 1006090 159515 1006093
rect 201033 1006090 201099 1006093
rect 208393 1006090 208459 1006093
rect 252461 1006090 252527 1006093
rect 260189 1006090 260255 1006093
rect 147121 1006088 148935 1006090
rect 147121 1006032 147126 1006088
rect 147182 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 147121 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 159449 1006088 159712 1006090
rect 159449 1006032 159454 1006088
rect 159510 1006032 159712 1006088
rect 159449 1006030 159712 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 208393 1006088 208656 1006090
rect 208393 1006032 208398 1006088
rect 208454 1006032 208656 1006088
rect 208393 1006030 208656 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 260084 1006088 260255 1006090
rect 260084 1006032 260194 1006088
rect 260250 1006032 260255 1006088
rect 260084 1006030 260255 1006032
rect 147121 1006027 147187 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 159449 1006027 159515 1006030
rect 201033 1006027 201099 1006030
rect 208393 1006027 208459 1006030
rect 252461 1006027 252527 1006030
rect 260189 1006027 260255 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 354857 1006090 354923 1006093
rect 422661 1006090 422727 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314653 1006088 314916 1006090
rect 314653 1006032 314658 1006088
rect 314714 1006032 314916 1006088
rect 314653 1006030 314916 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 422096 1006088 422727 1006090
rect 422096 1006032 422666 1006088
rect 422722 1006032 422727 1006088
rect 422096 1006030 422727 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 354857 1006027 354923 1006030
rect 422661 1006027 422727 1006030
rect 425513 1006090 425579 1006093
rect 498837 1006090 498903 1006093
rect 509049 1006090 509115 1006093
rect 550265 1006090 550331 1006093
rect 553945 1006090 554011 1006093
rect 425513 1006088 425776 1006090
rect 425513 1006032 425518 1006088
rect 425574 1006032 425776 1006088
rect 425513 1006030 425776 1006032
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 509049 1006088 509312 1006090
rect 509049 1006032 509054 1006088
rect 509110 1006032 509312 1006088
rect 509049 1006030 509312 1006032
rect 550265 1006088 550896 1006090
rect 550265 1006032 550270 1006088
rect 550326 1006032 550896 1006088
rect 550265 1006030 550896 1006032
rect 553748 1006088 554011 1006090
rect 553748 1006032 553950 1006088
rect 554006 1006032 554011 1006088
rect 553748 1006030 554011 1006032
rect 425513 1006027 425579 1006030
rect 498837 1006027 498903 1006030
rect 509049 1006027 509115 1006030
rect 550265 1006027 550331 1006030
rect 553945 1006027 554011 1006030
rect 363413 1005954 363479 1005957
rect 430849 1005954 430915 1005957
rect 363308 1005952 363479 1005954
rect 363308 1005896 363418 1005952
rect 363474 1005896 363479 1005952
rect 363308 1005894 363479 1005896
rect 430652 1005952 430915 1005954
rect 430652 1005896 430854 1005952
rect 430910 1005896 430915 1005952
rect 430652 1005894 430915 1005896
rect 363413 1005891 363479 1005894
rect 430849 1005891 430915 1005894
rect 304073 1005818 304139 1005821
rect 303876 1005816 304139 1005818
rect 303876 1005760 304078 1005816
rect 304134 1005760 304139 1005816
rect 303876 1005758 304139 1005760
rect 304073 1005755 304139 1005758
rect 426341 1005818 426407 1005821
rect 426341 1005816 426604 1005818
rect 426341 1005760 426346 1005816
rect 426402 1005760 426604 1005816
rect 426341 1005758 426604 1005760
rect 426341 1005755 426407 1005758
rect 360561 1005546 360627 1005549
rect 426341 1005546 426407 1005549
rect 360364 1005544 360627 1005546
rect 360364 1005488 360566 1005544
rect 360622 1005488 360627 1005544
rect 360364 1005486 360627 1005488
rect 426144 1005544 426407 1005546
rect 426144 1005488 426346 1005544
rect 426402 1005488 426407 1005544
rect 426144 1005486 426407 1005488
rect 360561 1005483 360627 1005486
rect 426341 1005483 426407 1005486
rect 358537 1005410 358603 1005413
rect 358340 1005408 358603 1005410
rect 358340 1005352 358542 1005408
rect 358598 1005352 358603 1005408
rect 358340 1005350 358603 1005352
rect 358537 1005347 358603 1005350
rect 430021 1005410 430087 1005413
rect 502149 1005410 502215 1005413
rect 430021 1005408 430284 1005410
rect 430021 1005352 430026 1005408
rect 430082 1005352 430284 1005408
rect 430021 1005350 430284 1005352
rect 501952 1005408 502215 1005410
rect 501952 1005352 502154 1005408
rect 502210 1005352 502215 1005408
rect 501952 1005350 502215 1005352
rect 430021 1005347 430087 1005350
rect 502149 1005347 502215 1005350
rect 551461 1005410 551527 1005413
rect 551461 1005408 551724 1005410
rect 551461 1005352 551466 1005408
rect 551522 1005352 551724 1005408
rect 551461 1005350 551724 1005352
rect 551461 1005347 551527 1005350
rect 423489 1005274 423555 1005277
rect 499665 1005274 499731 1005277
rect 423489 1005272 423752 1005274
rect 423489 1005216 423494 1005272
rect 423550 1005216 423752 1005272
rect 423489 1005214 423752 1005216
rect 499665 1005272 499928 1005274
rect 499665 1005216 499670 1005272
rect 499726 1005216 499928 1005272
rect 499665 1005214 499928 1005216
rect 423489 1005211 423555 1005214
rect 499665 1005211 499731 1005214
rect 152917 1005138 152983 1005141
rect 158621 1005138 158687 1005141
rect 263041 1005138 263107 1005141
rect 356513 1005138 356579 1005141
rect 152917 1005136 153180 1005138
rect 152917 1005080 152922 1005136
rect 152978 1005080 153180 1005136
rect 152917 1005078 153180 1005080
rect 158621 1005136 158884 1005138
rect 158621 1005080 158626 1005136
rect 158682 1005080 158884 1005136
rect 158621 1005078 158884 1005080
rect 262844 1005136 263107 1005138
rect 262844 1005080 263046 1005136
rect 263102 1005080 263107 1005136
rect 262844 1005078 263107 1005080
rect 356316 1005136 356579 1005138
rect 356316 1005080 356518 1005136
rect 356574 1005080 356579 1005136
rect 356316 1005078 356579 1005080
rect 152917 1005075 152983 1005078
rect 158621 1005075 158687 1005078
rect 263041 1005075 263107 1005078
rect 356513 1005075 356579 1005078
rect 361389 1005138 361455 1005141
rect 430021 1005138 430087 1005141
rect 551461 1005138 551527 1005141
rect 361389 1005136 361652 1005138
rect 361389 1005080 361394 1005136
rect 361450 1005080 361652 1005136
rect 361389 1005078 361652 1005080
rect 429824 1005136 430087 1005138
rect 429824 1005080 430026 1005136
rect 430082 1005080 430087 1005136
rect 429824 1005078 430087 1005080
rect 551356 1005136 551527 1005138
rect 551356 1005080 551466 1005136
rect 551522 1005080 551527 1005136
rect 551356 1005078 551527 1005080
rect 361389 1005075 361455 1005078
rect 430021 1005075 430087 1005078
rect 551461 1005075 551527 1005078
rect 153745 1005002 153811 1005005
rect 209221 1005002 209287 1005005
rect 313825 1005002 313891 1005005
rect 355685 1005002 355751 1005005
rect 423489 1005002 423555 1005005
rect 431217 1005002 431283 1005005
rect 507025 1005002 507091 1005005
rect 556797 1005002 556863 1005005
rect 153745 1005000 153916 1005002
rect 153745 1004944 153750 1005000
rect 153806 1004944 153916 1005000
rect 153745 1004942 153916 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 313628 1005000 313891 1005002
rect 313628 1004944 313830 1005000
rect 313886 1004944 313891 1005000
rect 313628 1004942 313891 1004944
rect 355488 1005000 355751 1005002
rect 355488 1004944 355690 1005000
rect 355746 1004944 355751 1005000
rect 355488 1004942 355751 1004944
rect 423292 1005000 423555 1005002
rect 423292 1004944 423494 1005000
rect 423550 1004944 423555 1005000
rect 423292 1004942 423555 1004944
rect 431020 1005000 431283 1005002
rect 431020 1004944 431222 1005000
rect 431278 1004944 431283 1005000
rect 431020 1004942 431283 1004944
rect 506828 1005000 507091 1005002
rect 506828 1004944 507030 1005000
rect 507086 1004944 507091 1005000
rect 506828 1004942 507091 1004944
rect 556600 1005000 556863 1005002
rect 556600 1004944 556802 1005000
rect 556858 1004944 556863 1005000
rect 556600 1004942 556863 1004944
rect 153745 1004939 153811 1004942
rect 209221 1004939 209287 1004942
rect 313825 1004939 313891 1004942
rect 355685 1004939 355751 1004942
rect 423489 1004939 423555 1004942
rect 431217 1004939 431283 1004942
rect 507025 1004939 507091 1004942
rect 556797 1004939 556863 1004942
rect 151721 1004866 151787 1004869
rect 160645 1004866 160711 1004869
rect 207565 1004866 207631 1004869
rect 151721 1004864 151892 1004866
rect 151721 1004808 151726 1004864
rect 151782 1004808 151892 1004864
rect 151721 1004806 151892 1004808
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 207460 1004864 207631 1004866
rect 207460 1004808 207570 1004864
rect 207626 1004808 207631 1004864
rect 207460 1004806 207631 1004808
rect 151721 1004803 151787 1004806
rect 160645 1004803 160711 1004806
rect 207565 1004803 207631 1004806
rect 211245 1004866 211311 1004869
rect 314653 1004866 314719 1004869
rect 362585 1004866 362651 1004869
rect 211245 1004864 211508 1004866
rect 211245 1004808 211250 1004864
rect 211306 1004808 211508 1004864
rect 211245 1004806 211508 1004808
rect 314548 1004864 314719 1004866
rect 314548 1004808 314658 1004864
rect 314714 1004808 314719 1004864
rect 314548 1004806 314719 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 211245 1004803 211311 1004806
rect 314653 1004803 314719 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 507853 1004866 507919 1004869
rect 555969 1004866 556035 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 507656 1004864 507919 1004866
rect 507656 1004808 507858 1004864
rect 507914 1004808 507919 1004864
rect 507656 1004806 507919 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 422661 1004803 422727 1004806
rect 507853 1004803 507919 1004806
rect 555969 1004803 556035 1004806
rect 154113 1004730 154179 1004733
rect 161105 1004730 161171 1004733
rect 209221 1004730 209287 1004733
rect 212533 1004730 212599 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 501321 1004730 501387 1004733
rect 557625 1004730 557691 1004733
rect 154113 1004728 154376 1004730
rect 154113 1004672 154118 1004728
rect 154174 1004672 154376 1004728
rect 154113 1004670 154376 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 212336 1004728 212599 1004730
rect 212336 1004672 212538 1004728
rect 212594 1004672 212599 1004728
rect 212336 1004670 212599 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 501124 1004728 501387 1004730
rect 501124 1004672 501326 1004728
rect 501382 1004672 501387 1004728
rect 501124 1004670 501387 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 154113 1004667 154179 1004670
rect 161105 1004667 161171 1004670
rect 209221 1004667 209287 1004670
rect 212533 1004667 212599 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 501321 1004667 501387 1004670
rect 557625 1004667 557691 1004670
rect 505369 1004594 505435 1004597
rect 505369 1004592 505632 1004594
rect 505369 1004536 505374 1004592
rect 505430 1004536 505632 1004592
rect 505369 1004534 505632 1004536
rect 505369 1004531 505435 1004534
rect 104801 1003914 104867 1003917
rect 356881 1003914 356947 1003917
rect 427169 1003914 427235 1003917
rect 505001 1003914 505067 1003917
rect 104604 1003912 104867 1003914
rect 104604 1003856 104806 1003912
rect 104862 1003856 104867 1003912
rect 104604 1003854 104867 1003856
rect 356684 1003912 356947 1003914
rect 356684 1003856 356886 1003912
rect 356942 1003856 356947 1003912
rect 356684 1003854 356947 1003856
rect 426972 1003912 427235 1003914
rect 426972 1003856 427174 1003912
rect 427230 1003856 427235 1003912
rect 426972 1003854 427235 1003856
rect 504804 1003912 505067 1003914
rect 504804 1003856 505006 1003912
rect 505062 1003856 505067 1003912
rect 504804 1003854 505067 1003856
rect 104801 1003851 104867 1003854
rect 356881 1003851 356947 1003854
rect 427169 1003851 427235 1003854
rect 505001 1003851 505067 1003854
rect 552289 1003914 552355 1003917
rect 552289 1003912 552552 1003914
rect 552289 1003856 552294 1003912
rect 552350 1003856 552552 1003912
rect 552289 1003854 552552 1003856
rect 552289 1003851 552355 1003854
rect 424317 1002826 424383 1002829
rect 424120 1002824 424383 1002826
rect 424120 1002768 424322 1002824
rect 424378 1002768 424383 1002824
rect 424120 1002766 424383 1002768
rect 424317 1002763 424383 1002766
rect 106825 1002690 106891 1002693
rect 106628 1002688 106891 1002690
rect 106628 1002632 106830 1002688
rect 106886 1002632 106891 1002688
rect 106628 1002630 106891 1002632
rect 106825 1002627 106891 1002630
rect 256141 1002690 256207 1002693
rect 261017 1002690 261083 1002693
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 260820 1002688 261083 1002690
rect 260820 1002632 261022 1002688
rect 261078 1002632 261083 1002688
rect 260820 1002630 261083 1002632
rect 256141 1002627 256207 1002630
rect 261017 1002627 261083 1002630
rect 299657 1002690 299723 1002693
rect 303245 1002690 303311 1002693
rect 306925 1002690 306991 1002693
rect 504173 1002690 504239 1002693
rect 299657 1002688 303311 1002690
rect 299657 1002632 299662 1002688
rect 299718 1002632 303250 1002688
rect 303306 1002632 303311 1002688
rect 299657 1002630 303311 1002632
rect 306728 1002688 306991 1002690
rect 306728 1002632 306930 1002688
rect 306986 1002632 306991 1002688
rect 306728 1002630 306991 1002632
rect 503976 1002688 504239 1002690
rect 503976 1002632 504178 1002688
rect 504234 1002632 504239 1002688
rect 503976 1002630 504239 1002632
rect 299657 1002627 299723 1002630
rect 303245 1002627 303311 1002630
rect 306925 1002627 306991 1002630
rect 504173 1002627 504239 1002630
rect 101489 1002554 101555 1002557
rect 108021 1002554 108087 1002557
rect 255313 1002554 255379 1002557
rect 359365 1002554 359431 1002557
rect 501689 1002554 501755 1002557
rect 101489 1002552 101752 1002554
rect 101489 1002496 101494 1002552
rect 101550 1002496 101752 1002552
rect 101489 1002494 101752 1002496
rect 107916 1002552 108087 1002554
rect 107916 1002496 108026 1002552
rect 108082 1002496 108087 1002552
rect 107916 1002494 108087 1002496
rect 255116 1002552 255379 1002554
rect 255116 1002496 255318 1002552
rect 255374 1002496 255379 1002552
rect 255116 1002494 255379 1002496
rect 359168 1002552 359431 1002554
rect 359168 1002496 359370 1002552
rect 359426 1002496 359431 1002552
rect 359168 1002494 359431 1002496
rect 501492 1002552 501755 1002554
rect 501492 1002496 501694 1002552
rect 501750 1002496 501755 1002552
rect 501492 1002494 501755 1002496
rect 101489 1002491 101555 1002494
rect 108021 1002491 108087 1002494
rect 255313 1002491 255379 1002494
rect 359365 1002491 359431 1002494
rect 501689 1002491 501755 1002494
rect 558821 1002554 558887 1002557
rect 558821 1002552 559084 1002554
rect 558821 1002496 558826 1002552
rect 558882 1002496 559084 1002552
rect 558821 1002494 559084 1002496
rect 558821 1002491 558887 1002494
rect 100293 1002418 100359 1002421
rect 103145 1002418 103211 1002421
rect 100293 1002416 100556 1002418
rect 100293 1002360 100298 1002416
rect 100354 1002360 100556 1002416
rect 100293 1002358 100556 1002360
rect 102948 1002416 103211 1002418
rect 102948 1002360 103150 1002416
rect 103206 1002360 103211 1002416
rect 102948 1002358 103211 1002360
rect 100293 1002355 100359 1002358
rect 103145 1002355 103211 1002358
rect 106825 1002418 106891 1002421
rect 150893 1002418 150959 1002421
rect 210877 1002418 210943 1002421
rect 256141 1002418 256207 1002421
rect 106825 1002416 107088 1002418
rect 106825 1002360 106830 1002416
rect 106886 1002360 107088 1002416
rect 106825 1002358 107088 1002360
rect 150893 1002416 151156 1002418
rect 150893 1002360 150898 1002416
rect 150954 1002360 151156 1002416
rect 150893 1002358 151156 1002360
rect 210877 1002416 211140 1002418
rect 210877 1002360 210882 1002416
rect 210938 1002360 211140 1002416
rect 210877 1002358 211140 1002360
rect 255944 1002416 256207 1002418
rect 255944 1002360 256146 1002416
rect 256202 1002360 256207 1002416
rect 255944 1002358 256207 1002360
rect 106825 1002355 106891 1002358
rect 150893 1002355 150959 1002358
rect 210877 1002355 210943 1002358
rect 256141 1002355 256207 1002358
rect 261017 1002418 261083 1002421
rect 357341 1002418 357407 1002421
rect 503345 1002418 503411 1002421
rect 560845 1002418 560911 1002421
rect 261017 1002416 261280 1002418
rect 261017 1002360 261022 1002416
rect 261078 1002360 261280 1002416
rect 261017 1002358 261280 1002360
rect 357144 1002416 357407 1002418
rect 357144 1002360 357346 1002416
rect 357402 1002360 357407 1002416
rect 357144 1002358 357407 1002360
rect 503148 1002416 503411 1002418
rect 503148 1002360 503350 1002416
rect 503406 1002360 503411 1002416
rect 503148 1002358 503411 1002360
rect 560740 1002416 560911 1002418
rect 560740 1002360 560850 1002416
rect 560906 1002360 560911 1002416
rect 560740 1002358 560911 1002360
rect 261017 1002355 261083 1002358
rect 357341 1002355 357407 1002358
rect 503345 1002355 503411 1002358
rect 560845 1002355 560911 1002358
rect 99097 1002282 99163 1002285
rect 101949 1002282 102015 1002285
rect 105997 1002282 106063 1002285
rect 99097 1002280 99268 1002282
rect 99097 1002224 99102 1002280
rect 99158 1002224 99268 1002280
rect 99097 1002222 99268 1002224
rect 101949 1002280 102212 1002282
rect 101949 1002224 101954 1002280
rect 102010 1002224 102212 1002280
rect 101949 1002222 102212 1002224
rect 105892 1002280 106063 1002282
rect 105892 1002224 106002 1002280
rect 106058 1002224 106063 1002280
rect 105892 1002222 106063 1002224
rect 99097 1002219 99163 1002222
rect 101949 1002219 102015 1002222
rect 105997 1002219 106063 1002222
rect 108849 1002282 108915 1002285
rect 155769 1002282 155835 1002285
rect 108849 1002280 109112 1002282
rect 108849 1002224 108854 1002280
rect 108910 1002224 109112 1002280
rect 108849 1002222 109112 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 108849 1002219 108915 1002222
rect 155769 1002219 155835 1002222
rect 156597 1002282 156663 1002285
rect 206369 1002282 206435 1002285
rect 156597 1002280 156860 1002282
rect 156597 1002224 156602 1002280
rect 156658 1002224 156860 1002280
rect 156597 1002222 156860 1002224
rect 206172 1002280 206435 1002282
rect 206172 1002224 206374 1002280
rect 206430 1002224 206435 1002280
rect 206172 1002222 206435 1002224
rect 156597 1002219 156663 1002222
rect 206369 1002219 206435 1002222
rect 254485 1002282 254551 1002285
rect 262673 1002282 262739 1002285
rect 357709 1002282 357775 1002285
rect 365069 1002282 365135 1002285
rect 428365 1002282 428431 1002285
rect 254485 1002280 254748 1002282
rect 254485 1002224 254490 1002280
rect 254546 1002224 254748 1002280
rect 254485 1002222 254748 1002224
rect 262476 1002280 262739 1002282
rect 262476 1002224 262678 1002280
rect 262734 1002224 262739 1002280
rect 262476 1002222 262739 1002224
rect 357604 1002280 357775 1002282
rect 357604 1002224 357714 1002280
rect 357770 1002224 357775 1002280
rect 357604 1002222 357775 1002224
rect 364872 1002280 365135 1002282
rect 364872 1002224 365074 1002280
rect 365130 1002224 365135 1002280
rect 364872 1002222 365135 1002224
rect 428260 1002280 428431 1002282
rect 428260 1002224 428370 1002280
rect 428426 1002224 428431 1002280
rect 428260 1002222 428431 1002224
rect 254485 1002219 254551 1002222
rect 262673 1002219 262739 1002222
rect 357709 1002219 357775 1002222
rect 365069 1002219 365135 1002222
rect 428365 1002219 428431 1002222
rect 432045 1002282 432111 1002285
rect 500493 1002282 500559 1002285
rect 509877 1002282 509943 1002285
rect 432045 1002280 432308 1002282
rect 432045 1002224 432050 1002280
rect 432106 1002224 432308 1002280
rect 432045 1002222 432308 1002224
rect 500296 1002280 500559 1002282
rect 500296 1002224 500498 1002280
rect 500554 1002224 500559 1002280
rect 500296 1002222 500559 1002224
rect 509680 1002280 509943 1002282
rect 509680 1002224 509882 1002280
rect 509938 1002224 509943 1002280
rect 509680 1002222 509943 1002224
rect 432045 1002219 432111 1002222
rect 500493 1002219 500559 1002222
rect 509877 1002219 509943 1002222
rect 554773 1002282 554839 1002285
rect 560017 1002282 560083 1002285
rect 554773 1002280 555036 1002282
rect 554773 1002224 554778 1002280
rect 554834 1002224 555036 1002280
rect 554773 1002222 555036 1002224
rect 559820 1002280 560083 1002282
rect 559820 1002224 560022 1002280
rect 560078 1002224 560083 1002280
rect 559820 1002222 560083 1002224
rect 554773 1002219 554839 1002222
rect 560017 1002219 560083 1002222
rect 100293 1002146 100359 1002149
rect 100096 1002144 100359 1002146
rect 100096 1002088 100298 1002144
rect 100354 1002088 100359 1002144
rect 100096 1002086 100359 1002088
rect 100293 1002083 100359 1002086
rect 103145 1002146 103211 1002149
rect 105629 1002146 105695 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 103145 1002144 103408 1002146
rect 103145 1002088 103150 1002144
rect 103206 1002088 103408 1002144
rect 103145 1002086 103408 1002088
rect 105432 1002144 105695 1002146
rect 105432 1002088 105634 1002144
rect 105690 1002088 105695 1002144
rect 105432 1002086 105695 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 103145 1002083 103211 1002086
rect 105629 1002083 105695 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 203517 1002146 203583 1002149
rect 206737 1002146 206803 1002149
rect 210877 1002146 210943 1002149
rect 263869 1002146 263935 1002149
rect 203517 1002144 203780 1002146
rect 203517 1002088 203522 1002144
rect 203578 1002088 203780 1002144
rect 203517 1002086 203780 1002088
rect 206540 1002144 206803 1002146
rect 206540 1002088 206742 1002144
rect 206798 1002088 206803 1002144
rect 206540 1002086 206803 1002088
rect 210680 1002144 210943 1002146
rect 210680 1002088 210882 1002144
rect 210938 1002088 210943 1002144
rect 210680 1002086 210943 1002088
rect 263764 1002144 263935 1002146
rect 263764 1002088 263874 1002144
rect 263930 1002088 263935 1002144
rect 263764 1002086 263935 1002088
rect 203517 1002083 203583 1002086
rect 206737 1002083 206803 1002086
rect 210877 1002083 210943 1002086
rect 263869 1002083 263935 1002086
rect 304901 1002146 304967 1002149
rect 360561 1002146 360627 1002149
rect 365897 1002146 365963 1002149
rect 304901 1002144 305164 1002146
rect 304901 1002088 304906 1002144
rect 304962 1002088 305164 1002144
rect 304901 1002086 305164 1002088
rect 360561 1002144 360824 1002146
rect 360561 1002088 360566 1002144
rect 360622 1002088 360824 1002144
rect 360561 1002086 360824 1002088
rect 365700 1002144 365963 1002146
rect 365700 1002088 365902 1002144
rect 365958 1002088 365963 1002144
rect 365700 1002086 365963 1002088
rect 304901 1002083 304967 1002086
rect 360561 1002083 360627 1002086
rect 365897 1002083 365963 1002086
rect 421465 1002146 421531 1002149
rect 427537 1002146 427603 1002149
rect 433333 1002146 433399 1002149
rect 421465 1002144 421636 1002146
rect 421465 1002088 421470 1002144
rect 421526 1002088 421636 1002144
rect 421465 1002086 421636 1002088
rect 427340 1002144 427603 1002146
rect 427340 1002088 427542 1002144
rect 427598 1002088 427603 1002144
rect 427340 1002086 427603 1002088
rect 433136 1002144 433399 1002146
rect 433136 1002088 433338 1002144
rect 433394 1002088 433399 1002144
rect 433136 1002086 433399 1002088
rect 421465 1002083 421531 1002086
rect 427537 1002083 427603 1002086
rect 433333 1002083 433399 1002086
rect 503345 1002146 503411 1002149
rect 510337 1002146 510403 1002149
rect 552289 1002146 552355 1002149
rect 503345 1002144 503608 1002146
rect 503345 1002088 503350 1002144
rect 503406 1002088 503608 1002144
rect 503345 1002086 503608 1002088
rect 510140 1002144 510403 1002146
rect 510140 1002088 510342 1002144
rect 510398 1002088 510403 1002144
rect 510140 1002086 510403 1002088
rect 552092 1002144 552355 1002146
rect 552092 1002088 552294 1002144
rect 552350 1002088 552355 1002144
rect 552092 1002086 552355 1002088
rect 503345 1002083 503411 1002086
rect 510337 1002083 510403 1002086
rect 552289 1002083 552355 1002086
rect 557993 1002146 558059 1002149
rect 560845 1002146 560911 1002149
rect 557993 1002144 558256 1002146
rect 557993 1002088 557998 1002144
rect 558054 1002088 558256 1002144
rect 557993 1002086 558256 1002088
rect 560845 1002144 561108 1002146
rect 560845 1002088 560850 1002144
rect 560906 1002088 561108 1002144
rect 560845 1002086 561108 1002088
rect 557993 1002083 558059 1002086
rect 560845 1002083 560911 1002086
rect 98269 1002010 98335 1002013
rect 101121 1002010 101187 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 100924 1002008 101187 1002010
rect 100924 1001952 101126 1002008
rect 101182 1001952 101187 1002008
rect 100924 1001950 101187 1001952
rect 98269 1001947 98335 1001950
rect 101121 1001947 101187 1001950
rect 102317 1002010 102383 1002013
rect 103973 1002010 104039 1002013
rect 102317 1002008 102580 1002010
rect 102317 1001952 102322 1002008
rect 102378 1001952 102580 1002008
rect 102317 1001950 102580 1001952
rect 103776 1002008 104039 1002010
rect 103776 1001952 103978 1002008
rect 104034 1001952 104039 1002008
rect 103776 1001950 104039 1001952
rect 102317 1001947 102383 1001950
rect 103973 1001947 104039 1001950
rect 105997 1002010 106063 1002013
rect 108849 1002010 108915 1002013
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 108652 1002008 108915 1002010
rect 108652 1001952 108854 1002008
rect 108910 1001952 108915 1002008
rect 108652 1001950 108915 1001952
rect 105997 1001947 106063 1001950
rect 108849 1001947 108915 1001950
rect 149237 1002010 149303 1002013
rect 154573 1002010 154639 1002013
rect 154941 1002010 155007 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 157793 1002010 157859 1002013
rect 202689 1002010 202755 1002013
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154573 1002008 154836 1002010
rect 154573 1001952 154578 1002008
rect 154634 1001952 154836 1002008
rect 154573 1001950 154836 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 155769 1002008 156032 1002010
rect 155769 1001952 155774 1002008
rect 155830 1001952 156032 1002008
rect 155769 1001950 156032 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 157596 1002008 157859 1002010
rect 157596 1001952 157798 1002008
rect 157854 1001952 157859 1002008
rect 157596 1001950 157859 1001952
rect 202492 1002008 202755 1002010
rect 202492 1001952 202694 1002008
rect 202750 1001952 202755 1002008
rect 202492 1001950 202755 1001952
rect 149237 1001947 149303 1001950
rect 154573 1001947 154639 1001950
rect 154941 1001947 155007 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 157793 1001947 157859 1001950
rect 202689 1001947 202755 1001950
rect 205541 1002010 205607 1002013
rect 207197 1002010 207263 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 207000 1002008 207263 1002010
rect 207000 1001952 207202 1002008
rect 207258 1001952 207263 1002008
rect 207000 1001950 207263 1001952
rect 205541 1001947 205607 1001950
rect 207197 1001947 207263 1001950
rect 207565 1002010 207631 1002013
rect 212073 1002010 212139 1002013
rect 263501 1002010 263567 1002013
rect 310145 1002010 310211 1002013
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 263304 1002008 263567 1002010
rect 263304 1001952 263506 1002008
rect 263562 1001952 263567 1002008
rect 263304 1001950 263567 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 207565 1001947 207631 1001950
rect 212073 1001947 212139 1001950
rect 263501 1001947 263567 1001950
rect 310145 1001947 310211 1001950
rect 354029 1002010 354095 1002013
rect 355685 1002010 355751 1002013
rect 360193 1002010 360259 1002013
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 355685 1002008 355948 1002010
rect 355685 1001952 355690 1002008
rect 355746 1001952 355948 1002008
rect 355685 1001950 355948 1001952
rect 359996 1002008 360259 1002010
rect 359996 1001952 360198 1002008
rect 360254 1001952 360259 1002008
rect 359996 1001950 360259 1001952
rect 354029 1001947 354095 1001950
rect 355685 1001947 355751 1001950
rect 360193 1001947 360259 1001950
rect 365069 1002010 365135 1002013
rect 424317 1002010 424383 1002013
rect 425145 1002010 425211 1002013
rect 425513 1002010 425579 1002013
rect 429193 1002010 429259 1002013
rect 432873 1002010 432939 1002013
rect 365069 1002008 365332 1002010
rect 365069 1001952 365074 1002008
rect 365130 1001952 365332 1002008
rect 365069 1001950 365332 1001952
rect 424317 1002008 424580 1002010
rect 424317 1001952 424322 1002008
rect 424378 1001952 424580 1002008
rect 424317 1001950 424580 1001952
rect 424948 1002008 425211 1002010
rect 424948 1001952 425150 1002008
rect 425206 1001952 425211 1002008
rect 424948 1001950 425211 1001952
rect 425316 1002008 425579 1002010
rect 425316 1001952 425518 1002008
rect 425574 1001952 425579 1002008
rect 425316 1001950 425579 1001952
rect 428996 1002008 429259 1002010
rect 428996 1001952 429198 1002008
rect 429254 1001952 429259 1002008
rect 428996 1001950 429259 1001952
rect 432676 1002008 432939 1002010
rect 432676 1001952 432878 1002008
rect 432934 1001952 432939 1002008
rect 432676 1001950 432939 1001952
rect 365069 1001947 365135 1001950
rect 424317 1001947 424383 1001950
rect 425145 1001947 425211 1001950
rect 425513 1001947 425579 1001950
rect 429193 1001947 429259 1001950
rect 432873 1001947 432939 1001950
rect 498469 1002010 498535 1002013
rect 500493 1002010 500559 1002013
rect 502149 1002010 502215 1002013
rect 502517 1002010 502583 1002013
rect 506197 1002010 506263 1002013
rect 507393 1002010 507459 1002013
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 500493 1002008 500756 1002010
rect 500493 1001952 500498 1002008
rect 500554 1001952 500756 1002008
rect 500493 1001950 500756 1001952
rect 502149 1002008 502412 1002010
rect 502149 1001952 502154 1002008
rect 502210 1001952 502412 1002008
rect 502149 1001950 502412 1001952
rect 502517 1002008 502780 1002010
rect 502517 1001952 502522 1002008
rect 502578 1001952 502780 1002008
rect 502517 1001950 502780 1001952
rect 506197 1002008 506460 1002010
rect 506197 1001952 506202 1002008
rect 506258 1001952 506460 1002008
rect 506197 1001950 506460 1001952
rect 507196 1002008 507459 1002010
rect 507196 1001952 507398 1002008
rect 507454 1001952 507459 1002008
rect 507196 1001950 507459 1001952
rect 498469 1001947 498535 1001950
rect 500493 1001947 500559 1001950
rect 502149 1001947 502215 1001950
rect 502517 1001947 502583 1001950
rect 506197 1001947 506263 1001950
rect 507393 1001947 507459 1001950
rect 554313 1002010 554379 1002013
rect 555141 1002010 555207 1002013
rect 558821 1002010 558887 1002013
rect 561673 1002010 561739 1002013
rect 554313 1002008 554576 1002010
rect 554313 1001952 554318 1002008
rect 554374 1001952 554576 1002008
rect 554313 1001950 554576 1001952
rect 555141 1002008 555404 1002010
rect 555141 1001952 555146 1002008
rect 555202 1001952 555404 1002008
rect 555141 1001950 555404 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 554313 1001947 554379 1001950
rect 555141 1001947 555207 1001950
rect 558821 1001947 558887 1001950
rect 561673 1001947 561739 1001950
rect 550265 1001194 550331 1001197
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 550265 1001131 550331 1001134
rect 258165 999154 258231 999157
rect 298461 999154 298527 999157
rect 301681 999154 301747 999157
rect 258165 999152 258428 999154
rect 258165 999096 258170 999152
rect 258226 999096 258428 999152
rect 258165 999094 258428 999096
rect 298461 999152 301747 999154
rect 298461 999096 298466 999152
rect 298522 999096 301686 999152
rect 301742 999096 301747 999152
rect 298461 999094 301747 999096
rect 258165 999091 258231 999094
rect 298461 999091 298527 999094
rect 301681 999091 301747 999094
rect 204345 998746 204411 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 204345 998683 204411 998686
rect 203885 998610 203951 998613
rect 308949 998610 309015 998613
rect 203885 998608 204148 998610
rect 203885 998552 203890 998608
rect 203946 998552 204148 998608
rect 203885 998550 204148 998552
rect 308752 998608 309015 998610
rect 308752 998552 308954 998608
rect 309010 998552 309015 998608
rect 308752 998550 309015 998552
rect 203885 998547 203951 998550
rect 308949 998547 309015 998550
rect 516685 998610 516751 998613
rect 523401 998610 523467 998613
rect 516685 998608 523467 998610
rect 516685 998552 516690 998608
rect 516746 998552 523406 998608
rect 523462 998552 523467 998608
rect 516685 998550 523467 998552
rect 516685 998547 516751 998550
rect 523401 998547 523467 998550
rect 258993 998474 259059 998477
rect 258796 998472 259059 998474
rect 258796 998416 258998 998472
rect 259054 998416 259059 998472
rect 258796 998414 259059 998416
rect 258993 998411 259059 998414
rect 298277 998474 298343 998477
rect 303245 998474 303311 998477
rect 298277 998472 303311 998474
rect 298277 998416 298282 998472
rect 298338 998416 303250 998472
rect 303306 998416 303311 998472
rect 298277 998414 303311 998416
rect 298277 998411 298343 998414
rect 303245 998411 303311 998414
rect 305269 998474 305335 998477
rect 305269 998472 305532 998474
rect 305269 998416 305274 998472
rect 305330 998416 305532 998472
rect 305269 998414 305532 998416
rect 305269 998411 305335 998414
rect 202689 998338 202755 998341
rect 307293 998338 307359 998341
rect 202689 998336 202952 998338
rect 202689 998280 202694 998336
rect 202750 998280 202952 998336
rect 202689 998278 202952 998280
rect 307293 998336 307556 998338
rect 307293 998280 307298 998336
rect 307354 998280 307556 998336
rect 307293 998278 307556 998280
rect 202689 998275 202755 998278
rect 307293 998275 307359 998278
rect 205541 998202 205607 998205
rect 205344 998200 205607 998202
rect 205344 998144 205546 998200
rect 205602 998144 205607 998200
rect 205344 998142 205607 998144
rect 205541 998139 205607 998142
rect 253657 998202 253723 998205
rect 257337 998202 257403 998205
rect 306925 998202 306991 998205
rect 458817 998202 458883 998205
rect 472433 998202 472499 998205
rect 253657 998200 253920 998202
rect 253657 998144 253662 998200
rect 253718 998144 253920 998200
rect 253657 998142 253920 998144
rect 257337 998200 257600 998202
rect 257337 998144 257342 998200
rect 257398 998144 257600 998200
rect 257337 998142 257600 998144
rect 306925 998200 307188 998202
rect 306925 998144 306930 998200
rect 306986 998144 307188 998200
rect 306925 998142 307188 998144
rect 458817 998200 472499 998202
rect 458817 998144 458822 998200
rect 458878 998144 472438 998200
rect 472494 998144 472499 998200
rect 458817 998142 472499 998144
rect 253657 998139 253723 998142
rect 257337 998139 257403 998142
rect 306925 998139 306991 998142
rect 458817 998139 458883 998142
rect 472433 998139 472499 998142
rect 201861 998066 201927 998069
rect 204713 998066 204779 998069
rect 253289 998066 253355 998069
rect 298093 998066 298159 998069
rect 303061 998066 303127 998069
rect 201861 998064 202124 998066
rect 201861 998008 201866 998064
rect 201922 998008 202124 998064
rect 201861 998006 202124 998008
rect 204713 998064 204976 998066
rect 204713 998008 204718 998064
rect 204774 998008 204976 998064
rect 204713 998006 204976 998008
rect 253289 998064 253460 998066
rect 253289 998008 253294 998064
rect 253350 998008 253460 998064
rect 253289 998006 253460 998008
rect 298093 998064 303127 998066
rect 298093 998008 298098 998064
rect 298154 998008 303066 998064
rect 303122 998008 303127 998064
rect 298093 998006 303127 998008
rect 201861 998003 201927 998006
rect 204713 998003 204779 998006
rect 253289 998003 253355 998006
rect 298093 998003 298159 998006
rect 303061 998003 303127 998006
rect 306097 998066 306163 998069
rect 308949 998066 309015 998069
rect 553117 998066 553183 998069
rect 306097 998064 306360 998066
rect 306097 998008 306102 998064
rect 306158 998008 306360 998064
rect 306097 998006 306360 998008
rect 308949 998064 309212 998066
rect 308949 998008 308954 998064
rect 309010 998008 309212 998064
rect 308949 998006 309212 998008
rect 552920 998064 553183 998066
rect 552920 998008 553122 998064
rect 553178 998008 553183 998064
rect 552920 998006 553183 998008
rect 306097 998003 306163 998006
rect 308949 998003 309015 998006
rect 553117 998003 553183 998006
rect 557165 998066 557231 998069
rect 557165 998064 557274 998066
rect 557165 998008 557170 998064
rect 557226 998008 557274 998064
rect 557165 998003 557274 998008
rect 200665 997930 200731 997933
rect 203517 997930 203583 997933
rect 252461 997930 252527 997933
rect 200665 997928 200836 997930
rect 200665 997872 200670 997928
rect 200726 997872 200836 997928
rect 200665 997870 200836 997872
rect 203320 997928 203583 997930
rect 203320 997872 203522 997928
rect 203578 997872 203583 997928
rect 203320 997870 203583 997872
rect 252264 997928 252527 997930
rect 252264 997872 252466 997928
rect 252522 997872 252527 997928
rect 252264 997870 252527 997872
rect 200665 997867 200731 997870
rect 203517 997867 203583 997870
rect 252461 997867 252527 997870
rect 256509 997930 256575 997933
rect 258993 997930 259059 997933
rect 259821 997930 259887 997933
rect 256509 997928 256772 997930
rect 256509 997872 256514 997928
rect 256570 997872 256772 997928
rect 256509 997870 256772 997872
rect 258993 997928 259164 997930
rect 258993 997872 258998 997928
rect 259054 997872 259164 997928
rect 258993 997870 259164 997872
rect 259624 997928 259887 997930
rect 259624 997872 259826 997928
rect 259882 997872 259887 997928
rect 259624 997870 259887 997872
rect 256509 997867 256575 997870
rect 258993 997867 259059 997870
rect 259821 997867 259887 997870
rect 307753 997930 307819 997933
rect 310605 997930 310671 997933
rect 307753 997928 307924 997930
rect 307753 997872 307758 997928
rect 307814 997872 307924 997928
rect 307753 997870 307924 997872
rect 310605 997928 310868 997930
rect 310605 997872 310610 997928
rect 310666 997872 310868 997928
rect 310605 997870 310868 997872
rect 307753 997867 307819 997870
rect 310605 997867 310671 997870
rect 229001 997794 229067 997797
rect 229369 997794 229435 997797
rect 229001 997792 229435 997794
rect 229001 997736 229006 997792
rect 229062 997736 229374 997792
rect 229430 997736 229435 997792
rect 229001 997734 229435 997736
rect 229001 997731 229067 997734
rect 229369 997731 229435 997734
rect 256969 997794 257035 997797
rect 258165 997794 258231 997797
rect 256969 997792 257140 997794
rect 256969 997736 256974 997792
rect 257030 997736 257140 997792
rect 256969 997734 257140 997736
rect 257968 997792 258231 997794
rect 257968 997736 258170 997792
rect 258226 997736 258231 997792
rect 257968 997734 258231 997736
rect 256969 997731 257035 997734
rect 258165 997731 258231 997734
rect 260189 997794 260255 997797
rect 261845 997794 261911 997797
rect 299289 997794 299355 997797
rect 309777 997794 309843 997797
rect 524045 997796 524111 997797
rect 524045 997794 524092 997796
rect 260189 997792 260452 997794
rect 260189 997736 260194 997792
rect 260250 997736 260452 997792
rect 260189 997734 260452 997736
rect 261845 997792 262108 997794
rect 261845 997736 261850 997792
rect 261906 997736 262108 997792
rect 261845 997734 262108 997736
rect 298142 997792 299355 997794
rect 298142 997736 299294 997792
rect 299350 997736 299355 997792
rect 298142 997734 299355 997736
rect 309580 997792 309843 997794
rect 309580 997736 309782 997792
rect 309838 997736 309843 997792
rect 309580 997734 309843 997736
rect 524000 997792 524092 997794
rect 524000 997736 524050 997792
rect 524000 997734 524092 997736
rect 260189 997731 260255 997734
rect 261845 997731 261911 997734
rect 84694 997188 84700 997252
rect 84764 997250 84770 997252
rect 93485 997250 93551 997253
rect 84764 997248 93551 997250
rect 84764 997192 93490 997248
rect 93546 997192 93551 997248
rect 84764 997190 93551 997192
rect 84764 997188 84770 997190
rect 93485 997187 93551 997190
rect 117221 997250 117287 997253
rect 144821 997250 144887 997253
rect 117221 997248 144887 997250
rect 117221 997192 117226 997248
rect 117282 997192 144826 997248
rect 144882 997192 144887 997248
rect 117221 997190 144887 997192
rect 117221 997187 117287 997190
rect 144821 997187 144887 997190
rect 170305 997250 170371 997253
rect 200205 997250 200271 997253
rect 170305 997248 200271 997250
rect 170305 997192 170310 997248
rect 170366 997192 200210 997248
rect 200266 997192 200271 997248
rect 170305 997190 200271 997192
rect 170305 997187 170371 997190
rect 200205 997187 200271 997190
rect 228817 997250 228883 997253
rect 229185 997250 229251 997253
rect 228817 997248 229251 997250
rect 228817 997192 228822 997248
rect 228878 997192 229190 997248
rect 229246 997192 229251 997248
rect 228817 997190 229251 997192
rect 228817 997187 228883 997190
rect 229185 997187 229251 997190
rect 245694 997188 245700 997252
rect 245764 997250 245770 997252
rect 250437 997250 250503 997253
rect 245764 997248 250503 997250
rect 245764 997192 250442 997248
rect 250498 997192 250503 997248
rect 245764 997190 250503 997192
rect 245764 997188 245770 997190
rect 250437 997187 250503 997190
rect 290406 997188 290412 997252
rect 290476 997250 290482 997252
rect 298142 997250 298202 997734
rect 299289 997731 299355 997734
rect 309777 997731 309843 997734
rect 524045 997732 524092 997734
rect 524156 997732 524162 997796
rect 553117 997794 553183 997797
rect 557214 997796 557274 998003
rect 553117 997792 553380 997794
rect 553117 997736 553122 997792
rect 553178 997736 553380 997792
rect 553117 997734 553380 997736
rect 524045 997731 524111 997732
rect 553117 997731 553183 997734
rect 557206 997732 557212 997796
rect 557276 997732 557282 997796
rect 290476 997190 298202 997250
rect 290476 997188 290482 997190
rect 298318 997188 298324 997252
rect 298388 997250 298394 997252
rect 299105 997250 299171 997253
rect 298388 997248 299171 997250
rect 298388 997192 299110 997248
rect 299166 997192 299171 997248
rect 298388 997190 299171 997192
rect 298388 997188 298394 997190
rect 299105 997187 299171 997190
rect 383561 997250 383627 997253
rect 390870 997250 390876 997252
rect 383561 997248 390876 997250
rect 383561 997192 383566 997248
rect 383622 997192 390876 997248
rect 383561 997190 390876 997192
rect 383561 997187 383627 997190
rect 390870 997188 390876 997190
rect 390940 997188 390946 997252
rect 439865 997250 439931 997253
rect 488901 997250 488967 997253
rect 439865 997248 488967 997250
rect 439865 997192 439870 997248
rect 439926 997192 488906 997248
rect 488962 997192 488967 997248
rect 439865 997190 488967 997192
rect 439865 997187 439931 997190
rect 488901 997187 488967 997190
rect 516685 997250 516751 997253
rect 540329 997250 540395 997253
rect 516685 997248 540395 997250
rect 516685 997192 516690 997248
rect 516746 997192 540334 997248
rect 540390 997192 540395 997248
rect 516685 997190 540395 997192
rect 516685 997187 516751 997190
rect 540329 997187 540395 997190
rect 74441 996978 74507 996981
rect 74625 996978 74691 996981
rect 74441 996976 74691 996978
rect 74441 996920 74446 996976
rect 74502 996920 74630 996976
rect 74686 996920 74691 996976
rect 74441 996918 74691 996920
rect 74441 996915 74507 996918
rect 74625 996915 74691 996918
rect 85982 996916 85988 996980
rect 86052 996978 86058 996980
rect 94497 996978 94563 996981
rect 86052 996976 94563 996978
rect 86052 996920 94502 996976
rect 94558 996920 94563 996976
rect 86052 996918 94563 996920
rect 86052 996916 86058 996918
rect 94497 996915 94563 996918
rect 116301 996978 116367 996981
rect 143993 996978 144059 996981
rect 116301 996976 144059 996978
rect 116301 996920 116306 996976
rect 116362 996920 143998 996976
rect 144054 996920 144059 996976
rect 116301 996918 144059 996920
rect 116301 996915 116367 996918
rect 143993 996915 144059 996918
rect 189022 996916 189028 996980
rect 189092 996978 189098 996980
rect 195053 996978 195119 996981
rect 189092 996976 195119 996978
rect 189092 996920 195058 996976
rect 195114 996920 195119 996976
rect 189092 996918 195119 996920
rect 189092 996916 189098 996918
rect 195053 996915 195119 996918
rect 291878 996916 291884 996980
rect 291948 996978 291954 996980
rect 299657 996978 299723 996981
rect 291948 996976 299723 996978
rect 291948 996920 299662 996976
rect 299718 996920 299723 996976
rect 291948 996918 299723 996920
rect 291948 996916 291954 996918
rect 299657 996915 299723 996918
rect 372521 996978 372587 996981
rect 399937 996978 400003 996981
rect 372521 996976 400003 996978
rect 372521 996920 372526 996976
rect 372582 996920 399942 996976
rect 399998 996920 400003 996976
rect 372521 996918 400003 996920
rect 372521 996915 372587 996918
rect 399937 996915 400003 996918
rect 439681 996978 439747 996981
rect 489085 996978 489151 996981
rect 439681 996976 489151 996978
rect 439681 996920 439686 996976
rect 439742 996920 489090 996976
rect 489146 996920 489151 996976
rect 439681 996918 489151 996920
rect 439681 996915 439747 996918
rect 489085 996915 489151 996918
rect 517053 996978 517119 996981
rect 540513 996978 540579 996981
rect 517053 996976 540579 996978
rect 517053 996920 517058 996976
rect 517114 996920 540518 996976
rect 540574 996920 540579 996976
rect 517053 996918 540579 996920
rect 517053 996915 517119 996918
rect 540513 996915 540579 996918
rect 599945 996978 600011 996981
rect 627862 996978 627868 996980
rect 599945 996976 627868 996978
rect 599945 996920 599950 996976
rect 600006 996920 627868 996976
rect 599945 996918 627868 996920
rect 599945 996915 600011 996918
rect 627862 996916 627868 996918
rect 627932 996916 627938 996980
rect 80470 996646 88074 996706
rect 80470 995757 80530 996646
rect 88014 996570 88074 996646
rect 88558 996644 88564 996708
rect 88628 996706 88634 996708
rect 94681 996706 94747 996709
rect 298318 996706 298324 996708
rect 88628 996704 94747 996706
rect 88628 996648 94686 996704
rect 94742 996648 94747 996704
rect 88628 996646 94747 996648
rect 88628 996644 88634 996646
rect 94681 996643 94747 996646
rect 282686 996646 298324 996706
rect 144821 996570 144887 996573
rect 88014 996510 88442 996570
rect 88382 996434 88442 996510
rect 142110 996568 144887 996570
rect 142110 996512 144826 996568
rect 144882 996512 144887 996568
rect 142110 996510 144887 996512
rect 93301 996434 93367 996437
rect 142110 996434 142170 996510
rect 144821 996507 144887 996510
rect 88382 996432 93367 996434
rect 88382 996376 93306 996432
rect 93362 996376 93367 996432
rect 88382 996374 93367 996376
rect 93301 996371 93367 996374
rect 140454 996374 142170 996434
rect 126237 996298 126303 996301
rect 140262 996298 140268 996300
rect 126237 996296 140268 996298
rect 126237 996240 126242 996296
rect 126298 996240 140268 996296
rect 126237 996238 140268 996240
rect 126237 996235 126303 996238
rect 140262 996236 140268 996238
rect 140332 996236 140338 996300
rect 93301 996026 93367 996029
rect 89486 996024 93367 996026
rect 89486 995968 93306 996024
rect 93362 995968 93367 996024
rect 89486 995966 93367 995968
rect 89486 995890 89546 995966
rect 93301 995963 93367 995966
rect 132350 995964 132356 996028
rect 132420 996026 132426 996028
rect 132420 995966 132970 996026
rect 132420 995964 132426 995966
rect 89302 995830 89546 995890
rect 80421 995752 80530 995757
rect 84653 995756 84719 995757
rect 84653 995754 84700 995756
rect 80421 995696 80426 995752
rect 80482 995696 80530 995752
rect 80421 995694 80530 995696
rect 84608 995752 84700 995754
rect 84608 995696 84658 995752
rect 84608 995694 84700 995696
rect 80421 995691 80487 995694
rect 84653 995692 84700 995694
rect 84764 995692 84770 995756
rect 87873 995754 87939 995757
rect 88558 995754 88564 995756
rect 87873 995752 88564 995754
rect 87873 995696 87878 995752
rect 87934 995696 88564 995752
rect 87873 995694 88564 995696
rect 84653 995691 84719 995692
rect 87873 995691 87939 995694
rect 88558 995692 88564 995694
rect 88628 995692 88634 995756
rect 88977 995754 89043 995757
rect 89302 995754 89362 995830
rect 132910 995757 132970 995966
rect 140454 995757 140514 996374
rect 192518 996372 192524 996436
rect 192588 996434 192594 996436
rect 195697 996434 195763 996437
rect 192588 996432 195763 996434
rect 192588 996376 195702 996432
rect 195758 996376 195763 996432
rect 192588 996374 195763 996376
rect 192588 996372 192594 996374
rect 195697 996371 195763 996374
rect 172329 996298 172395 996301
rect 172646 996298 172652 996300
rect 172329 996296 172652 996298
rect 172329 996240 172334 996296
rect 172390 996240 172652 996296
rect 172329 996238 172652 996240
rect 172329 996235 172395 996238
rect 172646 996236 172652 996238
rect 172716 996236 172722 996300
rect 241646 996236 241652 996300
rect 241716 996298 241722 996300
rect 251633 996298 251699 996301
rect 241716 996296 251699 996298
rect 241716 996240 251638 996296
rect 251694 996240 251699 996296
rect 241716 996238 251699 996240
rect 241716 996236 241722 996238
rect 251633 996235 251699 996238
rect 145741 996162 145807 996165
rect 88977 995752 89362 995754
rect 88977 995696 88982 995752
rect 89038 995696 89362 995752
rect 88977 995694 89362 995696
rect 89621 995754 89687 995757
rect 92657 995754 92723 995757
rect 89621 995752 92723 995754
rect 89621 995696 89626 995752
rect 89682 995696 92662 995752
rect 92718 995696 92723 995752
rect 89621 995694 92723 995696
rect 88977 995691 89043 995694
rect 89621 995691 89687 995694
rect 92657 995691 92723 995694
rect 131849 995754 131915 995757
rect 132534 995754 132540 995756
rect 131849 995752 132540 995754
rect 131849 995696 131854 995752
rect 131910 995696 132540 995752
rect 131849 995694 132540 995696
rect 131849 995691 131915 995694
rect 132534 995692 132540 995694
rect 132604 995692 132610 995756
rect 132910 995752 133019 995757
rect 132910 995696 132958 995752
rect 133014 995696 133019 995752
rect 132910 995694 133019 995696
rect 132953 995691 133019 995694
rect 140405 995752 140514 995757
rect 140405 995696 140410 995752
rect 140466 995696 140514 995752
rect 140405 995694 140514 995696
rect 140638 996160 145807 996162
rect 140638 996104 145746 996160
rect 145802 996104 145807 996160
rect 140638 996102 145807 996104
rect 140405 995691 140471 995694
rect 77937 995482 78003 995485
rect 90030 995482 90036 995484
rect 77937 995480 90036 995482
rect 77937 995424 77942 995480
rect 77998 995424 90036 995480
rect 77937 995422 90036 995424
rect 77937 995419 78003 995422
rect 90030 995420 90036 995422
rect 90100 995420 90106 995484
rect 90265 995482 90331 995485
rect 92473 995482 92539 995485
rect 90265 995480 92539 995482
rect 90265 995424 90270 995480
rect 90326 995424 92478 995480
rect 92534 995424 92539 995480
rect 90265 995422 92539 995424
rect 90265 995419 90331 995422
rect 92473 995419 92539 995422
rect 137369 995482 137435 995485
rect 140638 995482 140698 996102
rect 145741 996099 145807 996102
rect 144177 995890 144243 995893
rect 141558 995888 144243 995890
rect 141558 995832 144182 995888
rect 144238 995832 144243 995888
rect 141558 995830 144243 995832
rect 141049 995754 141115 995757
rect 141558 995754 141618 995830
rect 144177 995827 144243 995830
rect 141049 995752 141618 995754
rect 141049 995696 141054 995752
rect 141110 995696 141618 995752
rect 141049 995694 141618 995696
rect 141049 995691 141115 995694
rect 141785 995618 141851 995621
rect 147121 995618 147187 995621
rect 141785 995616 147187 995618
rect 141785 995560 141790 995616
rect 141846 995560 147126 995616
rect 147182 995560 147187 995616
rect 141785 995558 147187 995560
rect 141785 995555 141851 995558
rect 147121 995555 147187 995558
rect 155125 995618 155191 995621
rect 158486 995618 158546 996132
rect 155125 995616 158546 995618
rect 155125 995560 155130 995616
rect 155186 995560 158546 995616
rect 155125 995558 158546 995560
rect 155125 995555 155191 995558
rect 137369 995480 140698 995482
rect 137369 995424 137374 995480
rect 137430 995424 140698 995480
rect 137369 995422 140698 995424
rect 137369 995419 137435 995422
rect 132401 995348 132467 995349
rect 132350 995346 132356 995348
rect 132310 995286 132356 995346
rect 132420 995344 132467 995348
rect 132462 995288 132467 995344
rect 132350 995284 132356 995286
rect 132420 995284 132467 995288
rect 140814 995284 140820 995348
rect 140884 995346 140890 995348
rect 159222 995346 159282 996132
rect 202321 995890 202387 995893
rect 187006 995888 202387 995890
rect 187006 995832 202326 995888
rect 202382 995832 202387 995888
rect 187006 995830 202387 995832
rect 183829 995754 183895 995757
rect 187006 995754 187066 995830
rect 202321 995827 202387 995830
rect 183829 995752 187066 995754
rect 183829 995696 183834 995752
rect 183890 995696 187066 995752
rect 183829 995694 187066 995696
rect 183829 995691 183895 995694
rect 188797 995618 188863 995621
rect 189022 995618 189028 995620
rect 188797 995616 189028 995618
rect 188797 995560 188802 995616
rect 188858 995560 189028 995616
rect 188797 995558 189028 995560
rect 188797 995555 188863 995558
rect 189022 995556 189028 995558
rect 189092 995556 189098 995620
rect 190453 995618 190519 995621
rect 200757 995618 200823 995621
rect 190453 995616 200823 995618
rect 190453 995560 190458 995616
rect 190514 995560 200762 995616
rect 200818 995560 200823 995616
rect 190453 995558 200823 995560
rect 190453 995555 190519 995558
rect 200757 995555 200823 995558
rect 140884 995286 159282 995346
rect 188153 995346 188219 995349
rect 192477 995348 192543 995349
rect 190678 995346 190684 995348
rect 188153 995344 190684 995346
rect 188153 995288 188158 995344
rect 188214 995288 190684 995344
rect 188153 995286 190684 995288
rect 140884 995284 140890 995286
rect 132401 995283 132467 995284
rect 188153 995283 188219 995286
rect 190678 995284 190684 995286
rect 190748 995284 190754 995348
rect 192477 995346 192524 995348
rect 192432 995344 192524 995346
rect 192432 995288 192482 995344
rect 192432 995286 192524 995288
rect 192477 995284 192524 995286
rect 192588 995284 192594 995348
rect 192937 995346 193003 995349
rect 195881 995346 195947 995349
rect 192937 995344 195947 995346
rect 192937 995288 192942 995344
rect 192998 995288 195886 995344
rect 195942 995288 195947 995344
rect 192937 995286 195947 995288
rect 192477 995283 192543 995284
rect 192937 995283 193003 995286
rect 195881 995283 195947 995286
rect 77017 995210 77083 995213
rect 85982 995210 85988 995212
rect 77017 995208 85988 995210
rect 77017 995152 77022 995208
rect 77078 995152 85988 995208
rect 77017 995150 85988 995152
rect 77017 995147 77083 995150
rect 85982 995148 85988 995150
rect 86052 995148 86058 995212
rect 86309 995210 86375 995213
rect 93117 995210 93183 995213
rect 101397 995210 101463 995213
rect 86309 995208 93183 995210
rect 86309 995152 86314 995208
rect 86370 995152 93122 995208
rect 93178 995152 93183 995208
rect 86309 995150 93183 995152
rect 86309 995147 86375 995150
rect 93117 995147 93183 995150
rect 93810 995208 101463 995210
rect 93810 995152 101402 995208
rect 101458 995152 101463 995208
rect 93810 995150 101463 995152
rect 93810 995074 93870 995150
rect 101397 995147 101463 995150
rect 93350 995014 93870 995074
rect 124857 995074 124923 995077
rect 155125 995074 155191 995077
rect 124857 995072 155191 995074
rect 124857 995016 124862 995072
rect 124918 995016 155130 995072
rect 155186 995016 155191 995072
rect 124857 995014 155191 995016
rect 85021 994938 85087 994941
rect 92657 994938 92723 994941
rect 85021 994936 92723 994938
rect 85021 994880 85026 994936
rect 85082 994880 92662 994936
rect 92718 994880 92723 994936
rect 85021 994878 92723 994880
rect 85021 994875 85087 994878
rect 92657 994875 92723 994878
rect 90030 994604 90036 994668
rect 90100 994666 90106 994668
rect 93350 994666 93410 995014
rect 124857 995011 124923 995014
rect 155125 995011 155191 995014
rect 175917 995074 175983 995077
rect 208166 995074 208226 996132
rect 249241 996026 249307 996029
rect 241838 996024 249307 996026
rect 241838 995968 249246 996024
rect 249302 995968 249307 996024
rect 241838 995966 249307 995968
rect 239581 995754 239647 995757
rect 241838 995754 241898 995966
rect 249241 995963 249307 995966
rect 282686 995757 282746 996646
rect 298318 996644 298324 996646
rect 298388 996644 298394 996708
rect 298645 996706 298711 996709
rect 303245 996706 303311 996709
rect 298645 996704 303311 996706
rect 298645 996648 298650 996704
rect 298706 996648 303250 996704
rect 303306 996648 303311 996704
rect 298645 996646 303311 996648
rect 298645 996643 298711 996646
rect 303245 996643 303311 996646
rect 380157 996706 380223 996709
rect 383469 996706 383535 996709
rect 380157 996704 383535 996706
rect 380157 996648 380162 996704
rect 380218 996648 383474 996704
rect 383530 996648 383535 996704
rect 380157 996646 383535 996648
rect 380157 996643 380223 996646
rect 383469 996643 383535 996646
rect 489545 996706 489611 996709
rect 490097 996706 490163 996709
rect 590561 996706 590627 996709
rect 631726 996706 631732 996708
rect 489545 996704 490163 996706
rect 489545 996648 489550 996704
rect 489606 996648 490102 996704
rect 490158 996648 490163 996704
rect 489545 996646 490163 996648
rect 489545 996643 489611 996646
rect 490097 996643 490163 996646
rect 528326 996646 528570 996706
rect 472433 996570 472499 996573
rect 474774 996570 474780 996572
rect 472433 996568 474780 996570
rect 472433 996512 472438 996568
rect 472494 996512 474780 996568
rect 472433 996510 474780 996512
rect 472433 996507 472499 996510
rect 474774 996508 474780 996510
rect 474844 996508 474850 996572
rect 528134 996570 528140 996572
rect 522070 996510 528140 996570
rect 294822 996372 294828 996436
rect 294892 996434 294898 996436
rect 299381 996434 299447 996437
rect 294892 996432 299447 996434
rect 294892 996376 299386 996432
rect 299442 996376 299447 996432
rect 294892 996374 299447 996376
rect 294892 996372 294898 996374
rect 299381 996371 299447 996374
rect 372337 996434 372403 996437
rect 394918 996434 394924 996436
rect 372337 996432 394924 996434
rect 372337 996376 372342 996432
rect 372398 996376 394924 996432
rect 372337 996374 394924 996376
rect 372337 996371 372403 996374
rect 394918 996372 394924 996374
rect 394988 996372 394994 996436
rect 475878 996372 475884 996436
rect 475948 996434 475954 996436
rect 478454 996434 478460 996436
rect 475948 996374 478460 996434
rect 475948 996372 475954 996374
rect 478454 996372 478460 996374
rect 478524 996372 478530 996436
rect 494697 996434 494763 996437
rect 485638 996432 494763 996434
rect 485638 996376 494702 996432
rect 494758 996376 494763 996432
rect 485638 996374 494763 996376
rect 453205 996298 453271 996301
rect 474222 996298 474228 996300
rect 453205 996296 474228 996298
rect 453205 996240 453210 996296
rect 453266 996240 474228 996296
rect 453205 996238 474228 996240
rect 453205 996235 453271 996238
rect 474222 996236 474228 996238
rect 474292 996236 474298 996300
rect 301497 996162 301563 996165
rect 293542 996160 301563 996162
rect 293542 996104 301502 996160
rect 301558 996104 301563 996160
rect 373257 996162 373323 996165
rect 373257 996160 379530 996162
rect 293542 996102 301563 996104
rect 239581 995752 241898 995754
rect 239581 995696 239586 995752
rect 239642 995696 241898 995752
rect 239581 995694 241898 995696
rect 242065 995754 242131 995757
rect 247033 995754 247099 995757
rect 242065 995752 247099 995754
rect 242065 995696 242070 995752
rect 242126 995696 247038 995752
rect 247094 995696 247099 995752
rect 242065 995694 247099 995696
rect 282686 995752 282795 995757
rect 282686 995696 282734 995752
rect 282790 995696 282795 995752
rect 282686 995694 282795 995696
rect 239581 995691 239647 995694
rect 242065 995691 242131 995694
rect 247033 995691 247099 995694
rect 282729 995691 282795 995694
rect 290641 995754 290707 995757
rect 293542 995754 293602 996102
rect 301497 996099 301563 996102
rect 310378 995890 310438 996132
rect 296670 995830 310438 995890
rect 294781 995756 294847 995757
rect 294781 995754 294828 995756
rect 290641 995752 293602 995754
rect 290641 995696 290646 995752
rect 290702 995696 293602 995752
rect 290641 995694 293602 995696
rect 294736 995752 294828 995754
rect 294736 995696 294786 995752
rect 294736 995694 294828 995696
rect 290641 995691 290707 995694
rect 294781 995692 294828 995694
rect 294892 995692 294898 995756
rect 295057 995754 295123 995757
rect 296670 995754 296730 995830
rect 295057 995752 296730 995754
rect 295057 995696 295062 995752
rect 295118 995696 296730 995752
rect 295057 995694 296730 995696
rect 294781 995691 294847 995692
rect 295057 995691 295123 995694
rect 290457 995620 290523 995621
rect 290406 995556 290412 995620
rect 290476 995618 290523 995620
rect 301497 995618 301563 995621
rect 307017 995618 307083 995621
rect 290476 995616 290568 995618
rect 290518 995560 290568 995616
rect 290476 995558 290568 995560
rect 301497 995616 307083 995618
rect 301497 995560 301502 995616
rect 301558 995560 307022 995616
rect 307078 995560 307083 995616
rect 301497 995558 307083 995560
rect 290476 995556 290523 995558
rect 290457 995555 290523 995556
rect 301497 995555 301563 995558
rect 307017 995555 307083 995558
rect 240041 995482 240107 995485
rect 241646 995482 241652 995484
rect 240041 995480 241652 995482
rect 240041 995424 240046 995480
rect 240102 995424 241652 995480
rect 240041 995422 241652 995424
rect 240041 995419 240107 995422
rect 241646 995420 241652 995422
rect 241716 995420 241722 995484
rect 243261 995482 243327 995485
rect 246430 995482 246436 995484
rect 243261 995480 246436 995482
rect 243261 995424 243266 995480
rect 243322 995424 246436 995480
rect 243261 995422 246436 995424
rect 243261 995419 243327 995422
rect 246430 995420 246436 995422
rect 246500 995420 246506 995484
rect 280797 995346 280863 995349
rect 292297 995346 292363 995349
rect 280797 995344 292363 995346
rect 280797 995288 280802 995344
rect 280858 995288 292302 995344
rect 292358 995288 292363 995344
rect 280797 995286 292363 995288
rect 280797 995283 280863 995286
rect 292297 995283 292363 995286
rect 292481 995346 292547 995349
rect 295701 995346 295767 995349
rect 292481 995344 295767 995346
rect 292481 995288 292486 995344
rect 292542 995288 295706 995344
rect 295762 995288 295767 995344
rect 292481 995286 295767 995288
rect 292481 995283 292547 995286
rect 295701 995283 295767 995286
rect 296713 995346 296779 995349
rect 311206 995346 311266 996132
rect 296713 995344 311266 995346
rect 296713 995288 296718 995344
rect 296774 995288 311266 995344
rect 296713 995286 311266 995288
rect 296713 995283 296779 995286
rect 243905 995210 243971 995213
rect 247401 995210 247467 995213
rect 243905 995208 247467 995210
rect 243905 995152 243910 995208
rect 243966 995152 247406 995208
rect 247462 995152 247467 995208
rect 243905 995150 247467 995152
rect 243905 995147 243971 995150
rect 247401 995147 247467 995150
rect 175917 995072 208226 995074
rect 175917 995016 175922 995072
rect 175978 995016 208226 995072
rect 175917 995014 208226 995016
rect 279417 995074 279483 995077
rect 312862 995074 312922 996132
rect 373257 996104 373262 996160
rect 373318 996104 379530 996160
rect 373257 996102 379530 996104
rect 373257 996099 373323 996102
rect 379470 995754 379530 996102
rect 474414 996102 480270 996162
rect 382273 996026 382339 996029
rect 472249 996026 472315 996029
rect 474414 996026 474474 996102
rect 382273 996024 389190 996026
rect 382273 995968 382278 996024
rect 382334 995968 389190 996024
rect 382273 995966 389190 995968
rect 382273 995963 382339 995966
rect 388161 995754 388227 995757
rect 379470 995752 388227 995754
rect 379470 995696 388166 995752
rect 388222 995696 388227 995752
rect 379470 995694 388227 995696
rect 389130 995754 389190 995966
rect 472249 996024 474474 996026
rect 472249 995968 472254 996024
rect 472310 995968 474474 996024
rect 472249 995966 474474 995968
rect 472249 995963 472315 995966
rect 480210 995890 480270 996102
rect 474598 995830 476130 995890
rect 480210 995830 480546 995890
rect 415945 995754 416011 995757
rect 389130 995752 416011 995754
rect 389130 995696 415950 995752
rect 416006 995696 416011 995752
rect 389130 995694 416011 995696
rect 388161 995691 388227 995694
rect 415945 995691 416011 995694
rect 472893 995754 472959 995757
rect 473997 995754 474063 995757
rect 472893 995752 474063 995754
rect 472893 995696 472898 995752
rect 472954 995696 474002 995752
rect 474058 995696 474063 995752
rect 472893 995694 474063 995696
rect 472893 995691 472959 995694
rect 473997 995691 474063 995694
rect 474222 995692 474228 995756
rect 474292 995754 474298 995756
rect 474598 995754 474658 995830
rect 474292 995694 474658 995754
rect 476070 995754 476130 995830
rect 476941 995754 477007 995757
rect 476070 995752 477007 995754
rect 476070 995696 476946 995752
rect 477002 995696 477007 995752
rect 476070 995694 477007 995696
rect 480486 995754 480546 995830
rect 485638 995757 485698 996374
rect 494697 996371 494763 996374
rect 519813 996298 519879 996301
rect 522070 996298 522130 996510
rect 528134 996508 528140 996510
rect 528204 996508 528210 996572
rect 519813 996296 522130 996298
rect 519813 996240 519818 996296
rect 519874 996240 522130 996296
rect 519813 996238 522130 996240
rect 522297 996298 522363 996301
rect 528326 996298 528386 996646
rect 522297 996296 528386 996298
rect 522297 996240 522302 996296
rect 522358 996240 528386 996296
rect 522297 996238 528386 996240
rect 528510 996298 528570 996646
rect 590561 996704 631732 996706
rect 590561 996648 590566 996704
rect 590622 996648 631732 996704
rect 590561 996646 631732 996648
rect 590561 996643 590627 996646
rect 631726 996644 631732 996646
rect 631796 996644 631802 996708
rect 591297 996434 591363 996437
rect 599945 996434 600011 996437
rect 591297 996432 600011 996434
rect 591297 996376 591302 996432
rect 591358 996376 599950 996432
rect 600006 996376 600011 996432
rect 591297 996374 600011 996376
rect 591297 996371 591363 996374
rect 599945 996371 600011 996374
rect 618161 996434 618227 996437
rect 633934 996434 633940 996436
rect 618161 996432 633940 996434
rect 618161 996376 618166 996432
rect 618222 996376 633940 996432
rect 618161 996374 633940 996376
rect 618161 996371 618227 996374
rect 633934 996372 633940 996374
rect 634004 996372 634010 996436
rect 528510 996238 534090 996298
rect 519813 996235 519879 996238
rect 522297 996235 522363 996238
rect 480805 995754 480871 995757
rect 480486 995752 480871 995754
rect 480486 995696 480810 995752
rect 480866 995696 480871 995752
rect 480486 995694 480871 995696
rect 474292 995692 474298 995694
rect 476941 995691 477007 995694
rect 480805 995691 480871 995694
rect 485589 995752 485698 995757
rect 485589 995696 485594 995752
rect 485650 995696 485698 995752
rect 485589 995694 485698 995696
rect 485589 995691 485655 995694
rect 449157 995618 449223 995621
rect 469857 995618 469923 995621
rect 472433 995618 472499 995621
rect 474733 995620 474799 995621
rect 474733 995618 474780 995620
rect 449157 995616 466470 995618
rect 449157 995560 449162 995616
rect 449218 995560 466470 995616
rect 449157 995558 466470 995560
rect 449157 995555 449223 995558
rect 390870 995420 390876 995484
rect 390940 995482 390946 995484
rect 392393 995482 392459 995485
rect 394969 995484 395035 995485
rect 390940 995480 392459 995482
rect 390940 995424 392398 995480
rect 392454 995424 392459 995480
rect 390940 995422 392459 995424
rect 390940 995420 390946 995422
rect 392393 995419 392459 995422
rect 394918 995420 394924 995484
rect 394988 995482 395035 995484
rect 394988 995480 395080 995482
rect 395030 995424 395080 995480
rect 394988 995422 395080 995424
rect 394988 995420 395035 995422
rect 394969 995419 395035 995420
rect 375373 995346 375439 995349
rect 389357 995346 389423 995349
rect 375373 995344 389423 995346
rect 375373 995288 375378 995344
rect 375434 995288 389362 995344
rect 389418 995288 389423 995344
rect 375373 995286 389423 995288
rect 466410 995346 466470 995558
rect 469857 995616 472499 995618
rect 469857 995560 469862 995616
rect 469918 995560 472438 995616
rect 472494 995560 472499 995616
rect 469857 995558 472499 995560
rect 474688 995616 474780 995618
rect 474688 995560 474738 995616
rect 474688 995558 474780 995560
rect 469857 995555 469923 995558
rect 472433 995555 472499 995558
rect 474733 995556 474780 995558
rect 474844 995556 474850 995620
rect 478321 995618 478387 995621
rect 480253 995618 480319 995621
rect 478321 995616 480319 995618
rect 478321 995560 478326 995616
rect 478382 995560 480258 995616
rect 480314 995560 480319 995616
rect 478321 995558 480319 995560
rect 474733 995555 474799 995556
rect 478321 995555 478387 995558
rect 480253 995555 480319 995558
rect 503805 995618 503871 995621
rect 508086 995618 508146 996132
rect 503805 995616 508146 995618
rect 503805 995560 503810 995616
rect 503866 995560 508146 995616
rect 503805 995558 508146 995560
rect 503805 995555 503871 995558
rect 478229 995346 478295 995349
rect 466410 995344 478295 995346
rect 466410 995288 478234 995344
rect 478290 995288 478295 995344
rect 466410 995286 478295 995288
rect 375373 995283 375439 995286
rect 389357 995283 389423 995286
rect 478229 995283 478295 995286
rect 478454 995284 478460 995348
rect 478524 995346 478530 995348
rect 508822 995346 508882 996132
rect 523861 996026 523927 996029
rect 528870 996026 528876 996028
rect 523861 996024 528876 996026
rect 523861 995968 523866 996024
rect 523922 995968 528876 996024
rect 523861 995966 528876 995968
rect 523861 995963 523927 995966
rect 528870 995964 528876 995966
rect 528940 995964 528946 996028
rect 520917 995890 520983 995893
rect 523718 995890 523724 995892
rect 520917 995888 523724 995890
rect 520917 995832 520922 995888
rect 520978 995832 523724 995888
rect 520917 995830 523724 995832
rect 520917 995827 520983 995830
rect 523718 995828 523724 995830
rect 523788 995828 523794 995892
rect 532233 995756 532299 995757
rect 532182 995692 532188 995756
rect 532252 995754 532299 995756
rect 532252 995752 532344 995754
rect 532294 995696 532344 995752
rect 532252 995694 532344 995696
rect 532252 995692 532299 995694
rect 532233 995691 532299 995692
rect 516869 995618 516935 995621
rect 529841 995618 529907 995621
rect 516869 995616 529907 995618
rect 516869 995560 516874 995616
rect 516930 995560 529846 995616
rect 529902 995560 529907 995616
rect 516869 995558 529907 995560
rect 516869 995555 516935 995558
rect 529841 995555 529907 995558
rect 478524 995286 508882 995346
rect 522941 995346 523007 995349
rect 525333 995346 525399 995349
rect 522941 995344 525399 995346
rect 522941 995288 522946 995344
rect 523002 995288 525338 995344
rect 525394 995288 525399 995344
rect 522941 995286 525399 995288
rect 478524 995284 478530 995286
rect 522941 995283 523007 995286
rect 525333 995283 525399 995286
rect 525558 995284 525564 995348
rect 525628 995346 525634 995348
rect 525628 995286 528202 995346
rect 525628 995284 525634 995286
rect 279417 995072 312922 995074
rect 279417 995016 279422 995072
rect 279478 995016 312922 995072
rect 279417 995014 312922 995016
rect 372981 995074 373047 995077
rect 388989 995074 389055 995077
rect 372981 995072 389055 995074
rect 372981 995016 372986 995072
rect 373042 995016 388994 995072
rect 389050 995016 389055 995072
rect 372981 995014 389055 995016
rect 175917 995011 175983 995014
rect 279417 995011 279483 995014
rect 372981 995011 373047 995014
rect 388989 995011 389055 995014
rect 471237 995074 471303 995077
rect 475878 995074 475884 995076
rect 471237 995072 475884 995074
rect 471237 995016 471242 995072
rect 471298 995016 475884 995072
rect 471237 995014 475884 995016
rect 471237 995011 471303 995014
rect 475878 995012 475884 995014
rect 475948 995012 475954 995076
rect 476067 995074 476133 995077
rect 503805 995074 503871 995077
rect 476067 995072 503871 995074
rect 476067 995016 476072 995072
rect 476128 995016 503810 995072
rect 503866 995016 503871 995072
rect 476067 995014 503871 995016
rect 476067 995011 476133 995014
rect 503805 995011 503871 995014
rect 520181 995074 520247 995077
rect 523401 995074 523467 995077
rect 526069 995074 526135 995077
rect 527909 995074 527975 995077
rect 520181 995072 523234 995074
rect 520181 995016 520186 995072
rect 520242 995016 523234 995072
rect 520181 995014 523234 995016
rect 520181 995011 520247 995014
rect 132125 994802 132191 994805
rect 144361 994802 144427 994805
rect 132125 994800 144427 994802
rect 132125 994744 132130 994800
rect 132186 994744 144366 994800
rect 144422 994744 144427 994800
rect 132125 994742 144427 994744
rect 132125 994739 132191 994742
rect 144361 994739 144427 994742
rect 144545 994802 144611 994805
rect 149881 994802 149947 994805
rect 144545 994800 149947 994802
rect 144545 994744 144550 994800
rect 144606 994744 149886 994800
rect 149942 994744 149947 994800
rect 144545 994742 149947 994744
rect 144545 994739 144611 994742
rect 149881 994739 149947 994742
rect 180149 994802 180215 994805
rect 207013 994802 207079 994805
rect 180149 994800 207079 994802
rect 180149 994744 180154 994800
rect 180210 994744 207018 994800
rect 207074 994744 207079 994800
rect 180149 994742 207079 994744
rect 180149 994739 180215 994742
rect 207013 994739 207079 994742
rect 236545 994802 236611 994805
rect 251449 994802 251515 994805
rect 291837 994804 291903 994805
rect 291837 994802 291884 994804
rect 236545 994800 251515 994802
rect 236545 994744 236550 994800
rect 236606 994744 251454 994800
rect 251510 994744 251515 994800
rect 236545 994742 251515 994744
rect 291792 994800 291884 994802
rect 291792 994744 291842 994800
rect 291792 994742 291884 994744
rect 236545 994739 236611 994742
rect 251449 994739 251515 994742
rect 291837 994740 291884 994742
rect 291948 994740 291954 994804
rect 302877 994802 302943 994805
rect 292530 994800 302943 994802
rect 292530 994744 302882 994800
rect 302938 994744 302943 994800
rect 292530 994742 302943 994744
rect 291837 994739 291903 994740
rect 90100 994606 93410 994666
rect 90100 994604 90106 994606
rect 142153 994530 142219 994533
rect 157333 994530 157399 994533
rect 142153 994528 157399 994530
rect 142153 994472 142158 994528
rect 142214 994472 157338 994528
rect 157394 994472 157399 994528
rect 142153 994470 157399 994472
rect 142153 994467 142219 994470
rect 157333 994467 157399 994470
rect 187601 994530 187667 994533
rect 203333 994530 203399 994533
rect 187601 994528 203399 994530
rect 187601 994472 187606 994528
rect 187662 994472 203338 994528
rect 203394 994472 203399 994528
rect 187601 994470 203399 994472
rect 187601 994467 187667 994470
rect 203333 994467 203399 994470
rect 235257 994530 235323 994533
rect 246757 994530 246823 994533
rect 235257 994528 246823 994530
rect 235257 994472 235262 994528
rect 235318 994472 246762 994528
rect 246818 994472 246823 994528
rect 235257 994470 246823 994472
rect 235257 994467 235323 994470
rect 246757 994467 246823 994470
rect 288065 994530 288131 994533
rect 292530 994530 292590 994742
rect 302877 994739 302943 994742
rect 446397 994802 446463 994805
rect 480253 994802 480319 994805
rect 446397 994800 480319 994802
rect 446397 994744 446402 994800
rect 446458 994744 480258 994800
rect 480314 994744 480319 994800
rect 446397 994742 480319 994744
rect 523174 994802 523234 995014
rect 523401 995072 526135 995074
rect 523401 995016 523406 995072
rect 523462 995016 526074 995072
rect 526130 995016 526135 995072
rect 523401 995014 526135 995016
rect 523401 995011 523467 995014
rect 526069 995011 526135 995014
rect 526302 995072 527975 995074
rect 526302 995016 527914 995072
rect 527970 995016 527975 995072
rect 526302 995014 527975 995016
rect 528142 995074 528202 995286
rect 528318 995284 528324 995348
rect 528388 995346 528394 995348
rect 528553 995346 528619 995349
rect 528921 995348 528987 995349
rect 528388 995344 528619 995346
rect 528388 995288 528558 995344
rect 528614 995288 528619 995344
rect 528388 995286 528619 995288
rect 528388 995284 528394 995286
rect 528553 995283 528619 995286
rect 528870 995284 528876 995348
rect 528940 995346 528987 995348
rect 534030 995346 534090 996238
rect 536925 995618 536991 995621
rect 538070 995618 538076 995620
rect 536925 995616 538076 995618
rect 536925 995560 536930 995616
rect 536986 995560 538076 995616
rect 536925 995558 538076 995560
rect 536925 995555 536991 995558
rect 538070 995556 538076 995558
rect 538140 995556 538146 995620
rect 552657 995618 552723 995621
rect 557766 995618 557826 996132
rect 552657 995616 557826 995618
rect 552657 995560 552662 995616
rect 552718 995560 557826 995616
rect 552657 995558 557826 995560
rect 552657 995555 552723 995558
rect 560250 995346 560310 996132
rect 620093 996026 620159 996029
rect 623681 996026 623747 996029
rect 630622 996026 630628 996028
rect 620093 996024 621030 996026
rect 620093 995968 620098 996024
rect 620154 995968 621030 996024
rect 620093 995966 621030 995968
rect 620093 995963 620159 995966
rect 620970 995754 621030 995966
rect 623681 996024 630628 996026
rect 623681 995968 623686 996024
rect 623742 995968 630628 996024
rect 623681 995966 630628 995968
rect 623681 995963 623747 995966
rect 630622 995964 630628 995966
rect 630692 995964 630698 996028
rect 635181 995754 635247 995757
rect 620970 995752 635247 995754
rect 620970 995696 635186 995752
rect 635242 995696 635247 995752
rect 620970 995694 635247 995696
rect 635181 995691 635247 995694
rect 625521 995482 625587 995485
rect 627177 995482 627243 995485
rect 627913 995484 627979 995485
rect 625521 995480 627243 995482
rect 625521 995424 625526 995480
rect 625582 995424 627182 995480
rect 627238 995424 627243 995480
rect 625521 995422 627243 995424
rect 625521 995419 625587 995422
rect 627177 995419 627243 995422
rect 627862 995420 627868 995484
rect 627932 995482 627979 995484
rect 627932 995480 628024 995482
rect 627974 995424 628024 995480
rect 627932 995422 628024 995424
rect 627932 995420 627979 995422
rect 630622 995420 630628 995484
rect 630692 995482 630698 995484
rect 631501 995482 631567 995485
rect 633985 995484 634051 995485
rect 630692 995480 631567 995482
rect 630692 995424 631506 995480
rect 631562 995424 631567 995480
rect 630692 995422 631567 995424
rect 630692 995420 630698 995422
rect 627913 995419 627979 995420
rect 631501 995419 631567 995422
rect 633934 995420 633940 995484
rect 634004 995482 634051 995484
rect 634004 995480 634096 995482
rect 634046 995424 634096 995480
rect 634004 995422 634096 995424
rect 634004 995420 634051 995422
rect 634486 995420 634492 995484
rect 634556 995482 634562 995484
rect 634721 995482 634787 995485
rect 634556 995480 634787 995482
rect 634556 995424 634726 995480
rect 634782 995424 634787 995480
rect 634556 995422 634787 995424
rect 634556 995420 634562 995422
rect 633985 995419 634051 995420
rect 634721 995419 634787 995422
rect 528940 995344 529032 995346
rect 528982 995288 529032 995344
rect 528940 995286 529032 995288
rect 534030 995286 560310 995346
rect 631685 995348 631751 995349
rect 631685 995344 631732 995348
rect 631796 995346 631802 995348
rect 631685 995288 631690 995344
rect 528940 995284 528987 995286
rect 528921 995283 528987 995284
rect 631685 995284 631732 995288
rect 631796 995286 631842 995346
rect 631796 995284 631802 995286
rect 631685 995283 631751 995284
rect 552657 995074 552723 995077
rect 528142 995072 552723 995074
rect 528142 995016 552662 995072
rect 552718 995016 552723 995072
rect 528142 995014 552723 995016
rect 526302 994802 526362 995014
rect 527909 995011 527975 995014
rect 552657 995011 552723 995014
rect 590561 995074 590627 995077
rect 660573 995074 660639 995077
rect 590561 995072 660639 995074
rect 590561 995016 590566 995072
rect 590622 995016 660578 995072
rect 660634 995016 660639 995072
rect 590561 995014 660639 995016
rect 590561 995011 590627 995014
rect 660573 995011 660639 995014
rect 523174 994742 526362 994802
rect 526529 994802 526595 994805
rect 533705 994802 533771 994805
rect 526529 994800 533771 994802
rect 526529 994744 526534 994800
rect 526590 994744 533710 994800
rect 533766 994744 533771 994800
rect 526529 994742 533771 994744
rect 446397 994739 446463 994742
rect 480253 994739 480319 994742
rect 526529 994739 526595 994742
rect 533705 994739 533771 994742
rect 288065 994528 292590 994530
rect 288065 994472 288070 994528
rect 288126 994472 292590 994528
rect 288065 994470 292590 994472
rect 293309 994530 293375 994533
rect 298645 994530 298711 994533
rect 293309 994528 298711 994530
rect 293309 994472 293314 994528
rect 293370 994472 298650 994528
rect 298706 994472 298711 994528
rect 293309 994470 298711 994472
rect 288065 994467 288131 994470
rect 293309 994467 293375 994470
rect 298645 994467 298711 994470
rect 378041 994530 378107 994533
rect 392117 994530 392183 994533
rect 378041 994528 392183 994530
rect 378041 994472 378046 994528
rect 378102 994472 392122 994528
rect 392178 994472 392183 994528
rect 378041 994470 392183 994472
rect 378041 994467 378107 994470
rect 392117 994467 392183 994470
rect 461117 994530 461183 994533
rect 482645 994530 482711 994533
rect 461117 994528 482711 994530
rect 461117 994472 461122 994528
rect 461178 994472 482650 994528
rect 482706 994472 482711 994528
rect 461117 994470 482711 994472
rect 461117 994467 461183 994470
rect 482645 994467 482711 994470
rect 517513 994530 517579 994533
rect 533061 994530 533127 994533
rect 517513 994528 533127 994530
rect 517513 994472 517518 994528
rect 517574 994472 533066 994528
rect 533122 994472 533127 994528
rect 517513 994470 533127 994472
rect 517513 994467 517579 994470
rect 533061 994467 533127 994470
rect 86033 994394 86099 994397
rect 92841 994394 92907 994397
rect 86033 994392 92907 994394
rect 86033 994336 86038 994392
rect 86094 994336 92846 994392
rect 92902 994336 92907 994392
rect 86033 994334 92907 994336
rect 86033 994331 86099 994334
rect 92841 994331 92907 994334
rect 135897 994394 135963 994397
rect 141969 994394 142035 994397
rect 135897 994392 142035 994394
rect 135897 994336 135902 994392
rect 135958 994336 141974 994392
rect 142030 994336 142035 994392
rect 135897 994334 142035 994336
rect 135897 994331 135963 994334
rect 141969 994331 142035 994334
rect 148501 994258 148567 994261
rect 142110 994256 148567 994258
rect 142110 994200 148506 994256
rect 148562 994200 148567 994256
rect 142110 994198 148567 994200
rect 132534 994060 132540 994124
rect 132604 994122 132610 994124
rect 137553 994122 137619 994125
rect 132604 994120 137619 994122
rect 132604 994064 137558 994120
rect 137614 994064 137619 994120
rect 132604 994062 137619 994064
rect 132604 994060 132610 994062
rect 137553 994059 137619 994062
rect 137737 993986 137803 993989
rect 142110 993986 142170 994198
rect 148501 994195 148567 994198
rect 183277 994258 183343 994261
rect 208393 994258 208459 994261
rect 183277 994256 208459 994258
rect 183277 994200 183282 994256
rect 183338 994200 208398 994256
rect 208454 994200 208459 994256
rect 183277 994198 208459 994200
rect 183277 994195 183343 994198
rect 208393 994195 208459 994198
rect 240869 994258 240935 994261
rect 249057 994258 249123 994261
rect 240869 994256 249123 994258
rect 240869 994200 240874 994256
rect 240930 994200 249062 994256
rect 249118 994200 249123 994256
rect 240869 994198 249123 994200
rect 240869 994195 240935 994198
rect 249057 994195 249123 994198
rect 278630 994196 278636 994260
rect 278700 994258 278706 994260
rect 316401 994258 316467 994261
rect 278700 994256 316467 994258
rect 278700 994200 316406 994256
rect 316462 994200 316467 994256
rect 278700 994198 316467 994200
rect 278700 994196 278706 994198
rect 316401 994195 316467 994198
rect 472065 994258 472131 994261
rect 476757 994258 476823 994261
rect 472065 994256 476823 994258
rect 472065 994200 472070 994256
rect 472126 994200 476762 994256
rect 476818 994200 476823 994256
rect 472065 994198 476823 994200
rect 472065 994195 472131 994198
rect 476757 994195 476823 994198
rect 523217 994258 523283 994261
rect 526529 994258 526595 994261
rect 523217 994256 526595 994258
rect 523217 994200 523222 994256
rect 523278 994200 526534 994256
rect 526590 994200 526595 994256
rect 523217 994198 526595 994200
rect 523217 994195 523283 994198
rect 526529 994195 526595 994198
rect 137737 993984 142170 993986
rect 137737 993928 137742 993984
rect 137798 993928 142170 993984
rect 137737 993926 142170 993928
rect 142337 993986 142403 993989
rect 145557 993986 145623 993989
rect 152457 993986 152523 993989
rect 142337 993984 145623 993986
rect 142337 993928 142342 993984
rect 142398 993928 145562 993984
rect 145618 993928 145623 993984
rect 142337 993926 145623 993928
rect 137737 993923 137803 993926
rect 142337 993923 142403 993926
rect 145557 993923 145623 993926
rect 151770 993984 152523 993986
rect 151770 993928 152462 993984
rect 152518 993928 152523 993984
rect 151770 993926 152523 993928
rect 133137 993714 133203 993717
rect 139209 993714 139275 993717
rect 133137 993712 139275 993714
rect 133137 993656 133142 993712
rect 133198 993656 139214 993712
rect 139270 993656 139275 993712
rect 133137 993654 139275 993656
rect 133137 993651 133203 993654
rect 139209 993651 139275 993654
rect 139393 993714 139459 993717
rect 142153 993714 142219 993717
rect 151770 993714 151830 993926
rect 152457 993923 152523 993926
rect 190678 993924 190684 993988
rect 190748 993986 190754 993988
rect 196801 993986 196867 993989
rect 190748 993984 196867 993986
rect 190748 993928 196806 993984
rect 196862 993928 196867 993984
rect 190748 993926 196867 993928
rect 190748 993924 190754 993926
rect 196801 993923 196867 993926
rect 139393 993712 141986 993714
rect 139393 993656 139398 993712
rect 139454 993656 141986 993712
rect 139393 993654 141986 993656
rect 139393 993651 139459 993654
rect 141926 993442 141986 993654
rect 142153 993712 151830 993714
rect 142153 993656 142158 993712
rect 142214 993656 151830 993712
rect 142153 993654 151830 993656
rect 568205 993714 568271 993717
rect 641713 993714 641779 993717
rect 568205 993712 641779 993714
rect 568205 993656 568210 993712
rect 568266 993656 641718 993712
rect 641774 993656 641779 993712
rect 568205 993654 641779 993656
rect 142153 993651 142219 993654
rect 568205 993651 568271 993654
rect 641713 993651 641779 993654
rect 142337 993442 142403 993445
rect 141926 993440 142403 993442
rect 141926 993384 142342 993440
rect 142398 993384 142403 993440
rect 141926 993382 142403 993384
rect 142337 993379 142403 993382
rect 572662 990932 572668 990996
rect 572732 990994 572738 990996
rect 576301 990994 576367 990997
rect 572732 990992 576367 990994
rect 572732 990936 576306 990992
rect 576362 990936 576367 990992
rect 572732 990934 576367 990936
rect 572732 990932 572738 990934
rect 576301 990931 576367 990934
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 42149 968826 42215 968829
rect 43805 968826 43871 968829
rect 42149 968824 43871 968826
rect 42149 968768 42154 968824
rect 42210 968768 43810 968824
rect 43866 968768 43871 968824
rect 42149 968766 43871 968768
rect 42149 968763 42215 968766
rect 43805 968763 43871 968766
rect 41965 967196 42031 967197
rect 41965 967192 42012 967196
rect 42076 967194 42082 967196
rect 41965 967136 41970 967192
rect 41965 967132 42012 967136
rect 42076 967134 42122 967194
rect 42076 967132 42082 967134
rect 41965 967131 42031 967132
rect 42333 966786 42399 966789
rect 43437 966786 43503 966789
rect 42333 966784 43503 966786
rect 42333 966728 42338 966784
rect 42394 966728 43442 966784
rect 43498 966728 43503 966784
rect 42333 966726 43503 966728
rect 42333 966723 42399 966726
rect 43437 966723 43503 966726
rect 675661 966516 675727 966517
rect 675661 966512 675708 966516
rect 675772 966514 675778 966516
rect 675661 966456 675666 966512
rect 675661 966452 675708 966456
rect 675772 966454 675818 966514
rect 675772 966452 675778 966454
rect 675661 966451 675727 966452
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 42425 964746 42491 964749
rect 44633 964746 44699 964749
rect 42425 964744 44699 964746
rect 42425 964688 42430 964744
rect 42486 964688 44638 964744
rect 44694 964688 44699 964744
rect 42425 964686 44699 964688
rect 42425 964683 42491 964686
rect 44633 964683 44699 964686
rect 675293 964746 675359 964749
rect 676806 964746 676812 964748
rect 675293 964744 676812 964746
rect 675293 964688 675298 964744
rect 675354 964688 676812 964744
rect 675293 964686 676812 964688
rect 675293 964683 675359 964686
rect 676806 964684 676812 964686
rect 676876 964684 676882 964748
rect 42425 963930 42491 963933
rect 44265 963930 44331 963933
rect 42425 963928 44331 963930
rect 42425 963872 42430 963928
rect 42486 963872 44270 963928
rect 44326 963872 44331 963928
rect 42425 963870 44331 963872
rect 42425 963867 42491 963870
rect 44265 963867 44331 963870
rect 42425 963386 42491 963389
rect 43161 963386 43227 963389
rect 42425 963384 43227 963386
rect 42425 963328 42430 963384
rect 42486 963328 43166 963384
rect 43222 963328 43227 963384
rect 42425 963326 43227 963328
rect 42425 963323 42491 963326
rect 43161 963323 43227 963326
rect 675477 963388 675543 963389
rect 675477 963384 675524 963388
rect 675588 963386 675594 963388
rect 675477 963328 675482 963384
rect 675477 963324 675524 963328
rect 675588 963326 675634 963386
rect 675588 963324 675594 963326
rect 675477 963323 675543 963324
rect 42333 963114 42399 963117
rect 42793 963114 42859 963117
rect 42333 963112 42859 963114
rect 42333 963056 42338 963112
rect 42394 963056 42798 963112
rect 42854 963056 42859 963112
rect 42333 963054 42859 963056
rect 42333 963051 42399 963054
rect 42793 963051 42859 963054
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 673361 962842 673427 962845
rect 675477 962842 675543 962845
rect 673361 962840 675543 962842
rect 673361 962784 673366 962840
rect 673422 962784 675482 962840
rect 675538 962784 675543 962840
rect 673361 962782 675543 962784
rect 673361 962779 673427 962782
rect 675477 962779 675543 962782
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 41454 962100 41460 962164
rect 41524 962162 41530 962164
rect 41781 962162 41847 962165
rect 41524 962160 41847 962162
rect 41524 962104 41786 962160
rect 41842 962104 41847 962160
rect 41524 962102 41847 962104
rect 41524 962100 41530 962102
rect 41781 962099 41847 962102
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 674465 959442 674531 959445
rect 675385 959442 675451 959445
rect 674465 959440 675451 959442
rect 674465 959384 674470 959440
rect 674526 959384 675390 959440
rect 675446 959384 675451 959440
rect 674465 959382 675451 959384
rect 674465 959379 674531 959382
rect 675385 959379 675451 959382
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 674925 959170 674991 959173
rect 675518 959170 675524 959172
rect 674925 959168 675524 959170
rect 674925 959112 674930 959168
rect 674986 959112 675524 959168
rect 674925 959110 675524 959112
rect 674925 959107 674991 959110
rect 675518 959108 675524 959110
rect 675588 959108 675594 959172
rect 674649 958898 674715 958901
rect 675201 958898 675267 958901
rect 674649 958896 675267 958898
rect 674649 958840 674654 958896
rect 674710 958840 675206 958896
rect 675262 958840 675267 958896
rect 674649 958838 675267 958840
rect 674649 958835 674715 958838
rect 675201 958835 675267 958838
rect 42425 958762 42491 958765
rect 43621 958762 43687 958765
rect 42425 958760 43687 958762
rect 42425 958704 42430 958760
rect 42486 958704 43626 958760
rect 43682 958704 43687 958760
rect 42425 958702 43687 958704
rect 42425 958699 42491 958702
rect 43621 958699 43687 958702
rect 673177 958218 673243 958221
rect 675293 958218 675359 958221
rect 673177 958216 675359 958218
rect 673177 958160 673182 958216
rect 673238 958160 675298 958216
rect 675354 958160 675359 958216
rect 673177 958158 675359 958160
rect 673177 958155 673243 958158
rect 675293 958155 675359 958158
rect 42057 957946 42123 957949
rect 42558 957946 42564 957948
rect 42057 957944 42564 957946
rect 42057 957888 42062 957944
rect 42118 957888 42564 957944
rect 42057 957886 42564 957888
rect 42057 957883 42123 957886
rect 42558 957884 42564 957886
rect 42628 957884 42634 957948
rect 661677 957810 661743 957813
rect 675293 957810 675359 957813
rect 661677 957808 675359 957810
rect 661677 957752 661682 957808
rect 661738 957752 675298 957808
rect 675354 957752 675359 957808
rect 661677 957750 675359 957752
rect 661677 957747 661743 957750
rect 675293 957747 675359 957750
rect 675753 957810 675819 957813
rect 676622 957810 676628 957812
rect 675753 957808 676628 957810
rect 675753 957752 675758 957808
rect 675814 957752 676628 957808
rect 675753 957750 676628 957752
rect 675753 957747 675819 957750
rect 676622 957748 676628 957750
rect 676692 957748 676698 957812
rect 674097 957130 674163 957133
rect 675477 957130 675543 957133
rect 674097 957128 675543 957130
rect 674097 957072 674102 957128
rect 674158 957072 675482 957128
rect 675538 957072 675543 957128
rect 674097 957070 675543 957072
rect 674097 957067 674163 957070
rect 675477 957067 675543 957070
rect 675753 956450 675819 956453
rect 676990 956450 676996 956452
rect 675753 956448 676996 956450
rect 675753 956392 675758 956448
rect 675814 956392 676996 956448
rect 675753 956390 676996 956392
rect 675753 956387 675819 956390
rect 676990 956388 676996 956390
rect 677060 956388 677066 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 674833 953458 674899 953461
rect 675385 953458 675451 953461
rect 674833 953456 675451 953458
rect 674833 953400 674838 953456
rect 674894 953400 675390 953456
rect 675446 953400 675451 953456
rect 674833 953398 675451 953400
rect 674833 953395 674899 953398
rect 675385 953395 675451 953398
rect 28533 952914 28599 952917
rect 43437 952914 43503 952917
rect 28533 952912 43503 952914
rect 28533 952856 28538 952912
rect 28594 952856 43442 952912
rect 43498 952856 43503 952912
rect 28533 952854 43503 952856
rect 28533 952851 28599 952854
rect 43437 952851 43503 952854
rect 39297 952234 39363 952237
rect 41454 952234 41460 952236
rect 39297 952232 41460 952234
rect 39297 952176 39302 952232
rect 39358 952176 41460 952232
rect 39297 952174 41460 952176
rect 39297 952171 39363 952174
rect 41454 952172 41460 952174
rect 41524 952172 41530 952236
rect 672993 952234 673059 952237
rect 675477 952234 675543 952237
rect 672993 952232 675543 952234
rect 672993 952176 672998 952232
rect 673054 952176 675482 952232
rect 675538 952176 675543 952232
rect 672993 952174 675543 952176
rect 672993 952171 673059 952174
rect 675477 952171 675543 952174
rect 41597 951962 41663 951965
rect 42558 951962 42564 951964
rect 41597 951960 42564 951962
rect 41597 951904 41602 951960
rect 41658 951904 42564 951960
rect 41597 951902 42564 951904
rect 41597 951899 41663 951902
rect 42558 951900 42564 951902
rect 42628 951900 42634 951964
rect 40033 951826 40099 951829
rect 41270 951826 41276 951828
rect 40033 951824 41276 951826
rect 40033 951768 40038 951824
rect 40094 951768 41276 951824
rect 40033 951766 41276 951768
rect 40033 951763 40099 951766
rect 41270 951764 41276 951766
rect 41340 951764 41346 951828
rect 41413 951690 41479 951693
rect 42006 951690 42012 951692
rect 41413 951688 42012 951690
rect 41413 951632 41418 951688
rect 41474 951632 42012 951688
rect 41413 951630 42012 951632
rect 41413 951627 41479 951630
rect 42006 951628 42012 951630
rect 42076 951628 42082 951692
rect 675201 951554 675267 951557
rect 675845 951554 675911 951557
rect 675201 951552 675911 951554
rect 675201 951496 675206 951552
rect 675262 951496 675850 951552
rect 675906 951496 675911 951552
rect 675201 951494 675911 951496
rect 675201 951491 675267 951494
rect 675845 951491 675911 951494
rect 676806 950676 676812 950740
rect 676876 950738 676882 950740
rect 683297 950738 683363 950741
rect 676876 950736 683363 950738
rect 676876 950680 683302 950736
rect 683358 950680 683363 950736
rect 676876 950678 683363 950680
rect 676876 950676 676882 950678
rect 683297 950675 683363 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 675293 949242 675359 949245
rect 675702 949242 675708 949244
rect 675293 949240 675708 949242
rect 675293 949184 675298 949240
rect 675354 949184 675708 949240
rect 675293 949182 675708 949184
rect 675293 949179 675359 949182
rect 675702 949180 675708 949182
rect 675772 949180 675778 949244
rect 676070 948772 676076 948836
rect 676140 948834 676146 948836
rect 679617 948834 679683 948837
rect 676140 948832 679683 948834
rect 676140 948776 679622 948832
rect 679678 948776 679683 948832
rect 676140 948774 679683 948776
rect 676140 948772 676146 948774
rect 679617 948771 679683 948774
rect 667197 947338 667263 947341
rect 683481 947338 683547 947341
rect 667197 947336 683547 947338
rect 667197 947280 667202 947336
rect 667258 947280 683486 947336
rect 683542 947280 683547 947336
rect 667197 947278 683547 947280
rect 667197 947275 667263 947278
rect 683481 947275 683547 947278
rect 40534 944556 40540 944620
rect 40604 944618 40610 944620
rect 42374 944618 42380 944620
rect 40604 944558 42380 944618
rect 40604 944556 40610 944558
rect 42374 944556 42380 944558
rect 42444 944556 42450 944620
rect 41597 944346 41663 944349
rect 42190 944346 42196 944348
rect 41597 944344 42196 944346
rect 41597 944288 41602 944344
rect 41658 944288 42196 944344
rect 41597 944286 42196 944288
rect 41597 944283 41663 944286
rect 42190 944284 42196 944286
rect 42260 944284 42266 944348
rect 40718 944012 40724 944076
rect 40788 944074 40794 944076
rect 42006 944074 42012 944076
rect 40788 944014 42012 944074
rect 40788 944012 40794 944014
rect 42006 944012 42012 944014
rect 42076 944012 42082 944076
rect 40401 943802 40467 943805
rect 42241 943802 42307 943805
rect 40401 943800 42307 943802
rect 40401 943744 40406 943800
rect 40462 943744 42246 943800
rect 42302 943744 42307 943800
rect 40401 943742 42307 943744
rect 40401 943739 40467 943742
rect 42241 943739 42307 943742
rect 46289 943530 46355 943533
rect 41492 943528 46355 943530
rect 41492 943472 46294 943528
rect 46350 943472 46355 943528
rect 41492 943470 46355 943472
rect 46289 943467 46355 943470
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 28533 942714 28599 942717
rect 28533 942712 28612 942714
rect 28533 942656 28538 942712
rect 28594 942656 28612 942712
rect 28533 942654 28612 942656
rect 28533 942651 28599 942654
rect 48957 942306 49023 942309
rect 41492 942304 49023 942306
rect 41492 942248 48962 942304
rect 49018 942248 49023 942304
rect 41492 942246 49023 942248
rect 48957 942243 49023 942246
rect 35801 941898 35867 941901
rect 35788 941896 35867 941898
rect 35788 941840 35806 941896
rect 35862 941840 35867 941896
rect 35788 941838 35867 941840
rect 35801 941835 35867 941838
rect 663057 941762 663123 941765
rect 676213 941762 676279 941765
rect 663057 941760 676279 941762
rect 663057 941704 663062 941760
rect 663118 941704 676218 941760
rect 676274 941704 676279 941760
rect 663057 941702 676279 941704
rect 663057 941699 663123 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 44449 941082 44515 941085
rect 41492 941080 44515 941082
rect 41492 941024 44454 941080
rect 44510 941024 44515 941080
rect 41492 941022 44515 941024
rect 44449 941019 44515 941022
rect 50337 940674 50403 940677
rect 41492 940672 50403 940674
rect 41492 940616 50342 940672
rect 50398 940616 50403 940672
rect 41492 940614 50403 940616
rect 50337 940611 50403 940614
rect 35801 940266 35867 940269
rect 35788 940264 35867 940266
rect 35788 940208 35806 940264
rect 35862 940208 35867 940264
rect 35788 940206 35867 940208
rect 35801 940203 35867 940206
rect 51717 939858 51783 939861
rect 41492 939856 51783 939858
rect 41492 939800 51722 939856
rect 51778 939800 51783 939856
rect 41492 939798 51783 939800
rect 51717 939795 51783 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683481 939722 683547 939725
rect 683438 939720 683547 939722
rect 683438 939664 683486 939720
rect 683542 939664 683547 939720
rect 683438 939659 683547 939664
rect 683438 939556 683498 939659
rect 41822 939450 41828 939452
rect 41492 939390 41828 939450
rect 41822 939388 41828 939390
rect 41892 939388 41898 939452
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 37917 939042 37983 939045
rect 37917 939040 37996 939042
rect 37917 938984 37922 939040
rect 37978 938984 37996 939040
rect 37917 938982 37996 938984
rect 37917 938979 37983 938982
rect 669957 938770 670023 938773
rect 669957 938768 676292 938770
rect 669957 938712 669962 938768
rect 670018 938712 676292 938768
rect 669957 938710 676292 938712
rect 669957 938707 670023 938710
rect 41413 938634 41479 938637
rect 41308 938632 41479 938634
rect 41308 938576 41418 938632
rect 41474 938576 41479 938632
rect 41308 938574 41479 938576
rect 41413 938571 41479 938574
rect 36537 938464 36603 938467
rect 36494 938462 36603 938464
rect 36494 938406 36542 938462
rect 36598 938406 36603 938462
rect 36494 938401 36603 938406
rect 36494 938196 36554 938401
rect 671797 938362 671863 938365
rect 671797 938360 676292 938362
rect 671797 938304 671802 938360
rect 671858 938304 676292 938360
rect 671797 938302 676292 938304
rect 671797 938299 671863 938302
rect 672165 938090 672231 938093
rect 672165 938088 676322 938090
rect 672165 938032 672170 938088
rect 672226 938032 676322 938088
rect 672165 938030 676322 938032
rect 672165 938027 672231 938030
rect 676262 937924 676322 938030
rect 42190 937818 42196 937820
rect 41492 937758 42196 937818
rect 42190 937756 42196 937758
rect 42260 937756 42266 937820
rect 668577 937818 668643 937821
rect 672717 937818 672783 937821
rect 668577 937816 672783 937818
rect 668577 937760 668582 937816
rect 668638 937760 672722 937816
rect 672778 937760 672783 937816
rect 668577 937758 672783 937760
rect 668577 937755 668643 937758
rect 672717 937755 672783 937758
rect 671429 937546 671495 937549
rect 671429 937544 676292 937546
rect 671429 937488 671434 937544
rect 671490 937488 676292 937544
rect 671429 937486 676292 937488
rect 671429 937483 671495 937486
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 660297 937274 660363 937277
rect 672165 937274 672231 937277
rect 660297 937272 672231 937274
rect 660297 937216 660302 937272
rect 660358 937216 672170 937272
rect 672226 937216 672231 937272
rect 660297 937214 672231 937216
rect 660297 937211 660363 937214
rect 672165 937211 672231 937214
rect 672717 937274 672783 937277
rect 672717 937272 676322 937274
rect 672717 937216 672722 937272
rect 672778 937216 676322 937272
rect 672717 937214 676322 937216
rect 672717 937211 672783 937214
rect 676262 937108 676322 937214
rect 43805 937002 43871 937005
rect 41492 937000 43871 937002
rect 41492 936944 43810 937000
rect 43866 936944 43871 937000
rect 41492 936942 43871 936944
rect 43805 936939 43871 936942
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 43621 936186 43687 936189
rect 41492 936184 43687 936186
rect 41492 936128 43626 936184
rect 43682 936128 43687 936184
rect 41492 936126 43687 936128
rect 43621 936123 43687 936126
rect 42006 935778 42012 935780
rect 41492 935718 42012 935778
rect 42006 935716 42012 935718
rect 42076 935716 42082 935780
rect 42241 935778 42307 935781
rect 64462 935778 64522 936836
rect 672349 936730 672415 936733
rect 672349 936728 676292 936730
rect 672349 936672 672354 936728
rect 672410 936672 676292 936728
rect 672349 936670 676292 936672
rect 672349 936667 672415 936670
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 42241 935776 64522 935778
rect 42241 935720 42246 935776
rect 42302 935720 64522 935776
rect 42241 935718 64522 935720
rect 672533 935778 672599 935781
rect 676262 935778 676322 935884
rect 672533 935776 676322 935778
rect 672533 935720 672538 935776
rect 672594 935720 676322 935776
rect 672533 935718 676322 935720
rect 42241 935715 42307 935718
rect 672533 935715 672599 935718
rect 679617 935642 679683 935645
rect 679574 935640 679683 935642
rect 679574 935584 679622 935640
rect 679678 935584 679683 935640
rect 679574 935579 679683 935584
rect 679574 935476 679634 935579
rect 44633 935370 44699 935373
rect 41492 935368 44699 935370
rect 41492 935312 44638 935368
rect 44694 935312 44699 935368
rect 41492 935310 44699 935312
rect 44633 935307 44699 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43161 934962 43227 934965
rect 41492 934960 43227 934962
rect 41492 934904 43166 934960
rect 43222 934904 43227 934960
rect 41492 934902 43227 934904
rect 43161 934899 43227 934902
rect 675477 934690 675543 934693
rect 675477 934688 676292 934690
rect 675477 934632 675482 934688
rect 675538 934632 676292 934688
rect 675477 934630 676292 934632
rect 675477 934627 675543 934630
rect 39990 934387 40050 934524
rect 39990 934382 40099 934387
rect 39990 934326 40038 934382
rect 40094 934326 40099 934382
rect 39990 934324 40099 934326
rect 40033 934321 40099 934324
rect 675109 934282 675175 934285
rect 675109 934280 676292 934282
rect 675109 934224 675114 934280
rect 675170 934224 676292 934280
rect 675109 934222 676292 934224
rect 675109 934219 675175 934222
rect 42885 934146 42951 934149
rect 41492 934144 42951 934146
rect 41492 934088 42890 934144
rect 42946 934088 42951 934144
rect 41492 934086 42951 934088
rect 42885 934083 42951 934086
rect 674465 933874 674531 933877
rect 674465 933872 676292 933874
rect 674465 933816 674470 933872
rect 674526 933816 676292 933872
rect 674465 933814 676292 933816
rect 674465 933811 674531 933814
rect 44265 933738 44331 933741
rect 41492 933736 44331 933738
rect 41492 933680 44270 933736
rect 44326 933680 44331 933736
rect 41492 933678 44331 933680
rect 44265 933675 44331 933678
rect 672993 933466 673059 933469
rect 672993 933464 676292 933466
rect 672993 933408 672998 933464
rect 673054 933408 676292 933464
rect 672993 933406 676292 933408
rect 672993 933403 673059 933406
rect 43621 933330 43687 933333
rect 41492 933328 43687 933330
rect 41492 933272 43626 933328
rect 43682 933272 43687 933328
rect 41492 933270 43687 933272
rect 43621 933267 43687 933270
rect 674281 933058 674347 933061
rect 674281 933056 676292 933058
rect 674281 933000 674286 933056
rect 674342 933000 676292 933056
rect 674281 932998 676292 933000
rect 674281 932995 674347 932998
rect 41321 932922 41387 932925
rect 41308 932920 41387 932922
rect 27662 932484 27722 932892
rect 41308 932864 41326 932920
rect 41382 932864 41387 932920
rect 41308 932862 41387 932864
rect 41321 932859 41387 932862
rect 673361 932650 673427 932653
rect 673361 932648 676292 932650
rect 673361 932592 673366 932648
rect 673422 932592 676292 932648
rect 673361 932590 676292 932592
rect 673361 932587 673427 932590
rect 683297 932378 683363 932381
rect 683254 932376 683363 932378
rect 683254 932320 683302 932376
rect 683358 932320 683363 932376
rect 683254 932315 683363 932320
rect 683254 932212 683314 932315
rect 43805 932106 43871 932109
rect 41492 932104 43871 932106
rect 41492 932048 43810 932104
rect 43866 932048 43871 932104
rect 41492 932046 43871 932048
rect 43805 932043 43871 932046
rect 676990 931908 676996 931972
rect 677060 931908 677066 931972
rect 676998 931804 677058 931908
rect 676622 931500 676628 931564
rect 676692 931500 676698 931564
rect 676630 931396 676690 931500
rect 674649 931018 674715 931021
rect 674649 931016 676292 931018
rect 674649 930960 674654 931016
rect 674710 930960 676292 931016
rect 674649 930958 676292 930960
rect 674649 930955 674715 930958
rect 673177 930610 673243 930613
rect 673177 930608 676292 930610
rect 673177 930552 673182 930608
rect 673238 930552 676292 930608
rect 673177 930550 676292 930552
rect 673177 930547 673243 930550
rect 674097 930202 674163 930205
rect 674097 930200 676292 930202
rect 674097 930144 674102 930200
rect 674158 930144 676292 930200
rect 674097 930142 676292 930144
rect 674097 930139 674163 930142
rect 671981 929522 672047 929525
rect 676262 929522 676322 929764
rect 671981 929520 676322 929522
rect 671981 929464 671986 929520
rect 672042 929464 676322 929520
rect 671981 929462 676322 929464
rect 671981 929459 672047 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 673177 928298 673243 928301
rect 676262 928298 676322 928540
rect 673177 928296 676322 928298
rect 673177 928240 673182 928296
rect 673238 928240 676322 928296
rect 673177 928238 676322 928240
rect 673177 928235 673243 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 42241 911980 42307 911981
rect 42190 911978 42196 911980
rect 42150 911918 42196 911978
rect 42260 911976 42307 911980
rect 42302 911920 42307 911976
rect 42190 911916 42196 911918
rect 42260 911916 42307 911920
rect 42241 911915 42307 911916
rect 41781 911842 41847 911845
rect 42006 911842 42012 911844
rect 41781 911840 42012 911842
rect 41781 911784 41786 911840
rect 41842 911784 42012 911840
rect 41781 911782 42012 911784
rect 41781 911779 41847 911782
rect 42006 911780 42012 911782
rect 42076 911780 42082 911844
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 44081 892802 44147 892805
rect 55857 892802 55923 892805
rect 44081 892800 55923 892802
rect 44081 892744 44086 892800
rect 44142 892744 55862 892800
rect 55918 892744 55923 892800
rect 44081 892742 55923 892744
rect 44081 892739 44147 892742
rect 55857 892739 55923 892742
rect 44081 892530 44147 892533
rect 53281 892530 53347 892533
rect 44081 892528 53347 892530
rect 44081 892472 44086 892528
rect 44142 892472 53286 892528
rect 53342 892472 53347 892528
rect 44081 892470 53347 892472
rect 44081 892467 44147 892470
rect 53281 892467 53347 892470
rect 42931 892258 42997 892261
rect 54477 892258 54543 892261
rect 42931 892256 54543 892258
rect 42931 892200 42936 892256
rect 42992 892200 54482 892256
rect 54538 892200 54543 892256
rect 42931 892198 54543 892200
rect 42931 892195 42997 892198
rect 54477 892195 54543 892198
rect 43069 891986 43135 891989
rect 47577 891986 47643 891989
rect 43069 891984 47643 891986
rect 43069 891928 43074 891984
rect 43130 891928 47582 891984
rect 47638 891928 47643 891984
rect 43069 891926 47643 891928
rect 43069 891923 43135 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 670601 876890 670667 876893
rect 675109 876890 675175 876893
rect 670601 876888 675175 876890
rect 670601 876832 670606 876888
rect 670662 876832 675114 876888
rect 675170 876832 675175 876888
rect 670601 876830 675175 876832
rect 670601 876827 670667 876830
rect 675109 876827 675175 876830
rect 669221 876346 669287 876349
rect 675109 876346 675175 876349
rect 669221 876344 675175 876346
rect 669221 876288 669226 876344
rect 669282 876288 675114 876344
rect 675170 876288 675175 876344
rect 669221 876286 675175 876288
rect 669221 876283 669287 876286
rect 675109 876283 675175 876286
rect 675661 875938 675727 875941
rect 675886 875938 675892 875940
rect 675661 875936 675892 875938
rect 675661 875880 675666 875936
rect 675722 875880 675892 875936
rect 675661 875878 675892 875880
rect 675661 875875 675727 875878
rect 675886 875876 675892 875878
rect 675956 875876 675962 875940
rect 675753 874170 675819 874173
rect 676070 874170 676076 874172
rect 675753 874168 676076 874170
rect 675753 874112 675758 874168
rect 675814 874112 676076 874168
rect 675753 874110 676076 874112
rect 675753 874107 675819 874110
rect 676070 874108 676076 874110
rect 676140 874108 676146 874172
rect 669773 873490 669839 873493
rect 674925 873490 674991 873493
rect 669773 873488 674991 873490
rect 669773 873432 669778 873488
rect 669834 873432 674930 873488
rect 674986 873432 674991 873488
rect 669773 873430 674991 873432
rect 669773 873427 669839 873430
rect 674925 873427 674991 873430
rect 673862 873156 673868 873220
rect 673932 873218 673938 873220
rect 675109 873218 675175 873221
rect 673932 873216 675175 873218
rect 673932 873160 675114 873216
rect 675170 873160 675175 873216
rect 673932 873158 675175 873160
rect 673932 873156 673938 873158
rect 675109 873155 675175 873158
rect 668853 872266 668919 872269
rect 675109 872266 675175 872269
rect 675569 872266 675635 872269
rect 668853 872264 675175 872266
rect 668853 872208 668858 872264
rect 668914 872208 675114 872264
rect 675170 872208 675175 872264
rect 668853 872206 675175 872208
rect 668853 872203 668919 872206
rect 675109 872203 675175 872206
rect 675526 872264 675635 872266
rect 675526 872208 675574 872264
rect 675630 872208 675635 872264
rect 675526 872203 675635 872208
rect 675526 871994 675586 872203
rect 676806 871994 676812 871996
rect 675526 871934 676812 871994
rect 676806 871932 676812 871934
rect 676876 871932 676882 871996
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 672993 869410 673059 869413
rect 675109 869410 675175 869413
rect 672993 869408 675175 869410
rect 672993 869352 672998 869408
rect 673054 869352 675114 869408
rect 675170 869352 675175 869408
rect 672993 869350 675175 869352
rect 672993 869347 673059 869350
rect 675109 869347 675175 869350
rect 671153 869138 671219 869141
rect 674925 869138 674991 869141
rect 671153 869136 674991 869138
rect 671153 869080 671158 869136
rect 671214 869080 674930 869136
rect 674986 869080 674991 869136
rect 671153 869078 674991 869080
rect 671153 869075 671219 869078
rect 674925 869075 674991 869078
rect 664437 868730 664503 868733
rect 674649 868730 674715 868733
rect 664437 868728 674715 868730
rect 664437 868672 664442 868728
rect 664498 868672 674654 868728
rect 674710 868672 674715 868728
rect 664437 868670 674715 868672
rect 664437 868667 664503 868670
rect 674649 868667 674715 868670
rect 674649 868458 674715 868461
rect 675293 868458 675359 868461
rect 674649 868456 675359 868458
rect 674649 868400 674654 868456
rect 674710 868400 675298 868456
rect 675354 868400 675359 868456
rect 674649 868398 675359 868400
rect 674649 868395 674715 868398
rect 675293 868395 675359 868398
rect 669037 866690 669103 866693
rect 674925 866690 674991 866693
rect 669037 866688 674991 866690
rect 669037 866632 669042 866688
rect 669098 866632 674930 866688
rect 674986 866632 674991 866688
rect 669037 866630 674991 866632
rect 669037 866627 669103 866630
rect 674925 866627 674991 866630
rect 673913 864786 673979 864789
rect 675109 864786 675175 864789
rect 673913 864784 675175 864786
rect 673913 864728 673918 864784
rect 673974 864728 675114 864784
rect 675170 864728 675175 864784
rect 673913 864726 675175 864728
rect 673913 864723 673979 864726
rect 675109 864723 675175 864726
rect 62757 858666 62823 858669
rect 62757 858664 64492 858666
rect 62757 858608 62762 858664
rect 62818 858608 64492 858664
rect 62757 858606 64492 858608
rect 62757 858603 62823 858606
rect 651465 856354 651531 856357
rect 650164 856352 651531 856354
rect 650164 856296 651470 856352
rect 651526 856296 651531 856352
rect 650164 856294 651531 856296
rect 651465 856291 651531 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651833 843026 651899 843029
rect 650164 843024 651899 843026
rect 650164 842968 651838 843024
rect 651894 842968 651899 843024
rect 650164 842966 651899 842968
rect 651833 842963 651899 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 35801 816506 35867 816509
rect 651465 816506 651531 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 35801 816443 35867 816446
rect 651465 816443 651531 816446
rect 44909 816098 44975 816101
rect 41492 816096 44975 816098
rect 41492 816040 44914 816096
rect 44970 816040 44975 816096
rect 41492 816038 44975 816040
rect 44909 816035 44975 816038
rect 44449 815690 44515 815693
rect 41492 815688 44515 815690
rect 41492 815632 44454 815688
rect 44510 815632 44515 815688
rect 41492 815630 44515 815632
rect 44449 815627 44515 815630
rect 43069 815282 43135 815285
rect 41492 815280 43135 815282
rect 41492 815224 43074 815280
rect 43130 815224 43135 815280
rect 41492 815222 43135 815224
rect 43069 815219 43135 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 44633 814466 44699 814469
rect 41492 814464 44699 814466
rect 41492 814408 44638 814464
rect 44694 814408 44699 814464
rect 41492 814406 44699 814408
rect 44633 814403 44699 814406
rect 39982 814234 39988 814298
rect 40052 814234 40058 814298
rect 39990 814028 40050 814234
rect 45461 813650 45527 813653
rect 41492 813648 45527 813650
rect 41492 813592 45466 813648
rect 45522 813592 45527 813648
rect 41492 813590 45527 813592
rect 45461 813587 45527 813590
rect 41137 813242 41203 813245
rect 41124 813240 41203 813242
rect 41124 813184 41142 813240
rect 41198 813184 41203 813240
rect 41124 813182 41203 813184
rect 41137 813179 41203 813182
rect 41321 812834 41387 812837
rect 41308 812832 41387 812834
rect 41308 812776 41326 812832
rect 41382 812776 41387 812832
rect 41308 812774 41387 812776
rect 41321 812771 41387 812774
rect 40953 812426 41019 812429
rect 40940 812424 41019 812426
rect 40940 812368 40958 812424
rect 41014 812368 41019 812424
rect 40940 812366 41019 812368
rect 40953 812363 41019 812366
rect 41822 812018 41828 812020
rect 41492 811958 41828 812018
rect 41822 811956 41828 811958
rect 41892 811956 41898 812020
rect 39297 811610 39363 811613
rect 39284 811608 39363 811610
rect 39284 811552 39302 811608
rect 39358 811552 39363 811608
rect 39284 811550 39363 811552
rect 39297 811547 39363 811550
rect 33041 811202 33107 811205
rect 33028 811200 33107 811202
rect 33028 811144 33046 811200
rect 33102 811144 33107 811200
rect 33028 811142 33107 811144
rect 33041 811139 33107 811142
rect 45093 810794 45159 810797
rect 41492 810792 45159 810794
rect 41492 810736 45098 810792
rect 45154 810736 45159 810792
rect 41492 810734 45159 810736
rect 45093 810731 45159 810734
rect 43253 810386 43319 810389
rect 41492 810384 43319 810386
rect 41492 810328 43258 810384
rect 43314 810328 43319 810384
rect 41492 810326 43319 810328
rect 43253 810323 43319 810326
rect 45277 809978 45343 809981
rect 41492 809976 45343 809978
rect 41492 809920 45282 809976
rect 45338 809920 45343 809976
rect 41492 809918 45343 809920
rect 45277 809915 45343 809918
rect 44817 809570 44883 809573
rect 41492 809568 44883 809570
rect 41492 809512 44822 809568
rect 44878 809512 44883 809568
rect 41492 809510 44883 809512
rect 44817 809507 44883 809510
rect 41492 809102 41844 809162
rect 41784 809026 41844 809102
rect 42517 809026 42583 809029
rect 41784 809024 42583 809026
rect 41784 808968 42522 809024
rect 42578 808968 42583 809024
rect 41784 808966 42583 808968
rect 42517 808963 42583 808966
rect 42190 808754 42196 808756
rect 41492 808694 42196 808754
rect 42190 808692 42196 808694
rect 42260 808692 42266 808756
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 44173 807938 44239 807941
rect 41492 807936 44239 807938
rect 41492 807880 44178 807936
rect 44234 807880 44239 807936
rect 41492 807878 44239 807880
rect 44173 807875 44239 807878
rect 43437 807666 43503 807669
rect 41830 807664 43503 807666
rect 41830 807608 43442 807664
rect 43498 807608 43503 807664
rect 41830 807606 43503 807608
rect 41830 807530 41890 807606
rect 43437 807603 43503 807606
rect 41492 807470 41890 807530
rect 41462 806714 41522 807092
rect 42241 806714 42307 806717
rect 41462 806712 42307 806714
rect 41462 806684 42246 806712
rect 41492 806656 42246 806684
rect 42302 806656 42307 806712
rect 41492 806654 42307 806656
rect 42241 806651 42307 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43989 806306 44055 806309
rect 41492 806304 44055 806306
rect 41492 806248 43994 806304
rect 44050 806248 44055 806304
rect 41492 806246 44055 806248
rect 43989 806243 44055 806246
rect 41137 805626 41203 805629
rect 41638 805626 41644 805628
rect 41137 805624 41644 805626
rect 41137 805568 41142 805624
rect 41198 805568 41644 805624
rect 41137 805566 41644 805568
rect 41137 805563 41203 805566
rect 41638 805564 41644 805566
rect 41708 805564 41714 805628
rect 40953 805354 41019 805357
rect 41822 805354 41828 805356
rect 40953 805352 41828 805354
rect 40953 805296 40958 805352
rect 41014 805296 41828 805352
rect 40953 805294 41828 805296
rect 40953 805291 41019 805294
rect 41822 805292 41828 805294
rect 41892 805292 41898 805356
rect 40718 805020 40724 805084
rect 40788 805082 40794 805084
rect 41781 805082 41847 805085
rect 40788 805080 41847 805082
rect 40788 805024 41786 805080
rect 41842 805024 41847 805080
rect 40788 805022 41847 805024
rect 40788 805020 40794 805022
rect 41781 805019 41847 805022
rect 40534 804748 40540 804812
rect 40604 804810 40610 804812
rect 42190 804810 42196 804812
rect 40604 804750 42196 804810
rect 40604 804748 40610 804750
rect 42190 804748 42196 804750
rect 42260 804748 42266 804812
rect 40902 804340 40908 804404
rect 40972 804402 40978 804404
rect 42517 804402 42583 804405
rect 40972 804400 42583 804402
rect 40972 804344 42522 804400
rect 42578 804344 42583 804400
rect 40972 804342 42583 804344
rect 40972 804340 40978 804342
rect 42517 804339 42583 804342
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41597 801682 41663 801685
rect 42701 801682 42767 801685
rect 41597 801680 42767 801682
rect 41597 801624 41602 801680
rect 41658 801624 42706 801680
rect 42762 801624 42767 801680
rect 41597 801622 42767 801624
rect 41597 801619 41663 801622
rect 42701 801619 42767 801622
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 42517 799642 42583 799645
rect 53097 799642 53163 799645
rect 42517 799640 53163 799642
rect 42517 799584 42522 799640
rect 42578 799584 53102 799640
rect 53158 799584 53163 799640
rect 42517 799582 53163 799584
rect 42517 799579 42583 799582
rect 53097 799579 53163 799582
rect 42006 797676 42012 797740
rect 42076 797738 42082 797740
rect 44817 797738 44883 797741
rect 42076 797736 44883 797738
rect 42076 797680 44822 797736
rect 44878 797680 44883 797736
rect 42076 797678 44883 797680
rect 42076 797676 42082 797678
rect 44817 797675 44883 797678
rect 40902 796724 40908 796788
rect 40972 796786 40978 796788
rect 42517 796786 42583 796789
rect 40972 796784 42583 796786
rect 40972 796728 42522 796784
rect 42578 796728 42583 796784
rect 40972 796726 42583 796728
rect 40972 796724 40978 796726
rect 42517 796723 42583 796726
rect 44173 796378 44239 796381
rect 42198 796376 44239 796378
rect 42198 796320 44178 796376
rect 44234 796320 44239 796376
rect 42198 796318 44239 796320
rect 42198 796109 42258 796318
rect 44173 796315 44239 796318
rect 41965 796108 42031 796109
rect 41965 796106 42012 796108
rect 41920 796104 42012 796106
rect 41920 796048 41970 796104
rect 41920 796046 42012 796048
rect 41965 796044 42012 796046
rect 42076 796044 42082 796108
rect 42198 796104 42307 796109
rect 42198 796048 42246 796104
rect 42302 796048 42307 796104
rect 42198 796046 42307 796048
rect 41965 796043 42031 796044
rect 42241 796043 42307 796046
rect 40718 794956 40724 795020
rect 40788 795018 40794 795020
rect 40788 794958 42442 795018
rect 40788 794956 40794 794958
rect 42382 794341 42442 794958
rect 42382 794336 42491 794341
rect 42382 794280 42430 794336
rect 42486 794280 42491 794336
rect 42382 794278 42491 794280
rect 42425 794275 42491 794278
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 42609 792298 42675 792301
rect 45277 792298 45343 792301
rect 42609 792296 45343 792298
rect 42609 792240 42614 792296
rect 42670 792240 45282 792296
rect 45338 792240 45343 792296
rect 42609 792238 45343 792240
rect 42609 792235 42675 792238
rect 45277 792235 45343 792238
rect 42425 791754 42491 791757
rect 43253 791754 43319 791757
rect 42425 791752 43319 791754
rect 42425 791696 42430 791752
rect 42486 791696 43258 791752
rect 43314 791696 43319 791752
rect 42425 791694 43319 791696
rect 42425 791691 42491 791694
rect 43253 791691 43319 791694
rect 42149 790122 42215 790125
rect 42609 790122 42675 790125
rect 42149 790120 42675 790122
rect 42149 790064 42154 790120
rect 42210 790064 42614 790120
rect 42670 790064 42675 790120
rect 42149 790062 42675 790064
rect 42149 790059 42215 790062
rect 42609 790059 42675 790062
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 668209 789442 668275 789445
rect 675109 789442 675175 789445
rect 668209 789440 675175 789442
rect 668209 789384 668214 789440
rect 668270 789384 675114 789440
rect 675170 789384 675175 789440
rect 668209 789382 675175 789384
rect 668209 789379 668275 789382
rect 675109 789379 675175 789382
rect 41454 788564 41460 788628
rect 41524 788626 41530 788628
rect 41781 788626 41847 788629
rect 41524 788624 41847 788626
rect 41524 788568 41786 788624
rect 41842 788568 41847 788624
rect 41524 788566 41847 788568
rect 41524 788564 41530 788566
rect 41781 788563 41847 788566
rect 42701 788626 42767 788629
rect 62757 788626 62823 788629
rect 42701 788624 62823 788626
rect 42701 788568 42706 788624
rect 42762 788568 62762 788624
rect 62818 788568 62823 788624
rect 42701 788566 62823 788568
rect 42701 788563 42767 788566
rect 62757 788563 62823 788566
rect 41638 788156 41644 788220
rect 41708 788156 41714 788220
rect 41646 787946 41706 788156
rect 674465 788082 674531 788085
rect 675293 788082 675359 788085
rect 674465 788080 675359 788082
rect 674465 788024 674470 788080
rect 674526 788024 675298 788080
rect 675354 788024 675359 788080
rect 674465 788022 675359 788024
rect 674465 788019 674531 788022
rect 675293 788019 675359 788022
rect 42241 787946 42307 787949
rect 41646 787944 42307 787946
rect 41646 787888 42246 787944
rect 42302 787888 42307 787944
rect 41646 787886 42307 787888
rect 42241 787883 42307 787886
rect 42057 786450 42123 786453
rect 45185 786450 45251 786453
rect 42057 786448 45251 786450
rect 42057 786392 42062 786448
rect 42118 786392 45190 786448
rect 45246 786392 45251 786448
rect 42057 786390 45251 786392
rect 42057 786387 42123 786390
rect 45185 786387 45251 786390
rect 41781 785636 41847 785637
rect 41781 785632 41828 785636
rect 41892 785634 41898 785636
rect 41781 785576 41786 785632
rect 41781 785572 41828 785576
rect 41892 785574 41938 785634
rect 41892 785572 41898 785574
rect 41781 785571 41847 785572
rect 672809 784410 672875 784413
rect 675385 784410 675451 784413
rect 672809 784408 675451 784410
rect 672809 784352 672814 784408
rect 672870 784352 675390 784408
rect 675446 784352 675451 784408
rect 672809 784350 675451 784352
rect 672809 784347 672875 784350
rect 675385 784347 675451 784350
rect 669589 783866 669655 783869
rect 675477 783866 675543 783869
rect 669589 783864 675543 783866
rect 669589 783808 669594 783864
rect 669650 783808 675482 783864
rect 675538 783808 675543 783864
rect 669589 783806 675543 783808
rect 669589 783803 669655 783806
rect 675477 783803 675543 783806
rect 674230 782988 674236 783052
rect 674300 783050 674306 783052
rect 675385 783050 675451 783053
rect 674300 783048 675451 783050
rect 674300 782992 675390 783048
rect 675446 782992 675451 783048
rect 674300 782990 675451 782992
rect 674300 782988 674306 782990
rect 675385 782987 675451 782990
rect 670325 782506 670391 782509
rect 675477 782506 675543 782509
rect 670325 782504 675543 782506
rect 670325 782448 670330 782504
rect 670386 782448 675482 782504
rect 675538 782448 675543 782504
rect 670325 782446 675543 782448
rect 670325 782443 670391 782446
rect 675477 782443 675543 782446
rect 674833 780874 674899 780877
rect 676990 780874 676996 780876
rect 674833 780872 676996 780874
rect 674833 780816 674838 780872
rect 674894 780816 676996 780872
rect 674833 780814 676996 780816
rect 674833 780811 674899 780814
rect 676990 780812 676996 780814
rect 677060 780812 677066 780876
rect 672717 780602 672783 780605
rect 675477 780602 675543 780605
rect 672717 780600 675543 780602
rect 672717 780544 672722 780600
rect 672778 780544 675482 780600
rect 675538 780544 675543 780600
rect 672717 780542 675543 780544
rect 672717 780539 672783 780542
rect 675477 780539 675543 780542
rect 62757 780466 62823 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 62757 780403 62823 780406
rect 673729 779242 673795 779245
rect 675293 779242 675359 779245
rect 673729 779240 675359 779242
rect 673729 779184 673734 779240
rect 673790 779184 675298 779240
rect 675354 779184 675359 779240
rect 673729 779182 675359 779184
rect 673729 779179 673795 779182
rect 675293 779179 675359 779182
rect 660297 778970 660363 778973
rect 675201 778970 675267 778973
rect 660297 778968 675267 778970
rect 660297 778912 660302 778968
rect 660358 778912 675206 778968
rect 675262 778912 675267 778968
rect 660297 778910 675267 778912
rect 660297 778907 660363 778910
rect 675201 778907 675267 778910
rect 674281 778698 674347 778701
rect 675477 778698 675543 778701
rect 674281 778696 675543 778698
rect 674281 778640 674286 778696
rect 674342 778640 675482 778696
rect 675538 778640 675543 778696
rect 674281 778638 675543 778640
rect 674281 778635 674347 778638
rect 675477 778635 675543 778638
rect 666277 778426 666343 778429
rect 670785 778426 670851 778429
rect 666277 778424 670851 778426
rect 666277 778368 666282 778424
rect 666338 778368 670790 778424
rect 670846 778368 670851 778424
rect 666277 778366 670851 778368
rect 666277 778363 666343 778366
rect 670785 778363 670851 778366
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 652385 776658 652451 776661
rect 650164 776656 652451 776658
rect 650164 776600 652390 776656
rect 652446 776600 652451 776656
rect 650164 776598 652451 776600
rect 652385 776595 652451 776598
rect 670785 776522 670851 776525
rect 675477 776522 675543 776525
rect 670785 776520 675543 776522
rect 670785 776464 670790 776520
rect 670846 776464 675482 776520
rect 675538 776464 675543 776520
rect 670785 776462 675543 776464
rect 670785 776459 670851 776462
rect 675477 776459 675543 776462
rect 670141 775706 670207 775709
rect 674833 775706 674899 775709
rect 670141 775704 674899 775706
rect 670141 775648 670146 775704
rect 670202 775648 674838 775704
rect 674894 775648 674899 775704
rect 670141 775646 674899 775648
rect 670141 775643 670207 775646
rect 674833 775643 674899 775646
rect 671613 775026 671679 775029
rect 675385 775026 675451 775029
rect 671613 775024 675451 775026
rect 671613 774968 671618 775024
rect 671674 774968 675390 775024
rect 675446 774968 675451 775024
rect 671613 774966 675451 774968
rect 671613 774963 671679 774966
rect 675385 774963 675451 774966
rect 674833 774618 674899 774621
rect 675477 774618 675543 774621
rect 674833 774616 675543 774618
rect 674833 774560 674838 774616
rect 674894 774560 675482 774616
rect 675538 774560 675543 774616
rect 674833 774558 675543 774560
rect 674833 774555 674899 774558
rect 675477 774555 675543 774558
rect 41462 774346 41522 774452
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 41462 773938 41522 774044
rect 41462 773878 45570 773938
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 45001 773258 45067 773261
rect 41492 773256 45067 773258
rect 41492 773200 45006 773256
rect 45062 773200 45067 773256
rect 41492 773198 45067 773200
rect 45001 773195 45067 773198
rect 44173 772850 44239 772853
rect 41492 772848 44239 772850
rect 41492 772792 44178 772848
rect 44234 772792 44239 772848
rect 41492 772790 44239 772792
rect 45510 772850 45570 773878
rect 55857 772850 55923 772853
rect 45510 772848 55923 772850
rect 45510 772792 55862 772848
rect 55918 772792 55923 772848
rect 45510 772790 55923 772792
rect 44173 772787 44239 772790
rect 55857 772787 55923 772790
rect 43069 772442 43135 772445
rect 41492 772440 43135 772442
rect 41492 772384 43074 772440
rect 43130 772384 43135 772440
rect 41492 772382 43135 772384
rect 43069 772379 43135 772382
rect 44449 772034 44515 772037
rect 41492 772032 44515 772034
rect 41492 771976 44454 772032
rect 44510 771976 44515 772032
rect 41492 771974 44515 771976
rect 44449 771971 44515 771974
rect 673913 772034 673979 772037
rect 683205 772034 683271 772037
rect 673913 772032 683271 772034
rect 673913 771976 673918 772032
rect 673974 771976 683210 772032
rect 683266 771976 683271 772032
rect 673913 771974 683271 771976
rect 673913 771971 673979 771974
rect 683205 771971 683271 771974
rect 44633 771626 44699 771629
rect 41492 771624 44699 771626
rect 41492 771568 44638 771624
rect 44694 771568 44699 771624
rect 41492 771566 44699 771568
rect 44633 771563 44699 771566
rect 675886 771428 675892 771492
rect 675956 771490 675962 771492
rect 678237 771490 678303 771493
rect 675956 771488 678303 771490
rect 675956 771432 678242 771488
rect 678298 771432 678303 771488
rect 675956 771430 678303 771432
rect 675956 771428 675962 771430
rect 678237 771427 678303 771430
rect 44633 771218 44699 771221
rect 41492 771216 44699 771218
rect 41492 771160 44638 771216
rect 44694 771160 44699 771216
rect 41492 771158 44699 771160
rect 44633 771155 44699 771158
rect 45461 770810 45527 770813
rect 41492 770808 45527 770810
rect 41492 770752 45466 770808
rect 45522 770752 45527 770808
rect 41492 770750 45527 770752
rect 45461 770747 45527 770750
rect 674649 770674 674715 770677
rect 683389 770674 683455 770677
rect 674649 770672 683455 770674
rect 674649 770616 674654 770672
rect 674710 770616 683394 770672
rect 683450 770616 683455 770672
rect 674649 770614 683455 770616
rect 674649 770611 674715 770614
rect 683389 770611 683455 770614
rect 45001 770402 45067 770405
rect 41492 770400 45067 770402
rect 41492 770344 45006 770400
rect 45062 770344 45067 770400
rect 41492 770342 45067 770344
rect 45001 770339 45067 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 676070 768708 676076 768772
rect 676140 768770 676146 768772
rect 682377 768770 682443 768773
rect 676140 768768 682443 768770
rect 676140 768712 682382 768768
rect 682438 768712 682443 768768
rect 676140 768710 682443 768712
rect 676140 768708 676146 768710
rect 682377 768707 682443 768710
rect 35574 768229 35634 768332
rect 35574 768224 35683 768229
rect 35574 768168 35622 768224
rect 35678 768168 35683 768224
rect 35574 768166 35683 768168
rect 35617 768163 35683 768166
rect 30974 767821 31034 767924
rect 30974 767816 31083 767821
rect 35801 767818 35867 767821
rect 30974 767760 31022 767816
rect 31078 767760 31083 767816
rect 30974 767758 31083 767760
rect 31017 767755 31083 767758
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 42793 766730 42859 766733
rect 41492 766728 42859 766730
rect 41492 766672 42798 766728
rect 42854 766672 42859 766728
rect 41492 766670 42859 766672
rect 42793 766667 42859 766670
rect 674925 766594 674991 766597
rect 676121 766596 676187 766597
rect 675886 766594 675892 766596
rect 674925 766592 675892 766594
rect 674925 766536 674930 766592
rect 674986 766536 675892 766592
rect 674925 766534 675892 766536
rect 674925 766531 674991 766534
rect 675886 766532 675892 766534
rect 675956 766532 675962 766596
rect 676070 766532 676076 766596
rect 676140 766594 676187 766596
rect 676140 766592 676232 766594
rect 676182 766536 676232 766592
rect 676140 766534 676232 766536
rect 676140 766532 676187 766534
rect 676121 766531 676187 766532
rect 45185 766322 45251 766325
rect 41492 766320 45251 766322
rect 41492 766264 45190 766320
rect 45246 766264 45251 766320
rect 41492 766262 45251 766264
rect 45185 766259 45251 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 41321 765370 41387 765373
rect 42609 765370 42675 765373
rect 41321 765368 42675 765370
rect 41321 765312 41326 765368
rect 41382 765312 42614 765368
rect 42670 765312 42675 765368
rect 41321 765310 42675 765312
rect 41321 765307 41387 765310
rect 42609 765307 42675 765310
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 43345 764690 43411 764693
rect 41492 764688 43411 764690
rect 41492 764632 43350 764688
rect 43406 764632 43411 764688
rect 41492 764630 43411 764632
rect 43345 764627 43411 764630
rect 46933 764418 46999 764421
rect 41462 764416 46999 764418
rect 41462 764360 46938 764416
rect 46994 764360 46999 764416
rect 41462 764358 46999 764360
rect 41462 764252 41522 764358
rect 46933 764355 46999 764358
rect 40585 764146 40651 764149
rect 42517 764146 42583 764149
rect 40585 764144 42583 764146
rect 40585 764088 40590 764144
rect 40646 764088 42522 764144
rect 42578 764088 42583 764144
rect 40585 764086 42583 764088
rect 40585 764083 40651 764086
rect 42517 764083 42583 764086
rect 35758 763333 35818 763844
rect 40401 763738 40467 763741
rect 42333 763738 42399 763741
rect 40401 763736 42399 763738
rect 40401 763680 40406 763736
rect 40462 763680 42338 763736
rect 42394 763680 42399 763736
rect 40401 763678 42399 763680
rect 40401 763675 40467 763678
rect 42333 763675 42399 763678
rect 35758 763328 35867 763333
rect 651465 763330 651531 763333
rect 35758 763272 35806 763328
rect 35862 763272 35867 763328
rect 35758 763270 35867 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 35801 763267 35867 763270
rect 651465 763267 651531 763270
rect 43161 763058 43227 763061
rect 41492 763056 43227 763058
rect 41492 763000 43166 763056
rect 43222 763000 43227 763056
rect 41492 762998 43227 763000
rect 43161 762995 43227 762998
rect 670969 763058 671035 763061
rect 676029 763058 676095 763061
rect 670969 763056 676095 763058
rect 670969 763000 670974 763056
rect 671030 763000 676034 763056
rect 676090 763000 676095 763056
rect 670969 762998 676095 763000
rect 670969 762995 671035 762998
rect 676029 762995 676095 762998
rect 676949 761836 677015 761837
rect 676949 761832 676996 761836
rect 677060 761834 677066 761836
rect 676581 761792 676647 761793
rect 676581 761788 676628 761792
rect 676692 761790 676698 761792
rect 676581 761732 676586 761788
rect 676581 761728 676628 761732
rect 676692 761730 676738 761790
rect 676949 761776 676954 761832
rect 676949 761772 676996 761776
rect 677060 761774 677106 761834
rect 677060 761772 677066 761774
rect 676949 761771 677015 761772
rect 676692 761728 676698 761730
rect 676581 761727 676647 761728
rect 665817 761562 665883 761565
rect 665817 761560 676292 761562
rect 665817 761504 665822 761560
rect 665878 761504 676292 761560
rect 665817 761502 676292 761504
rect 665817 761499 665883 761502
rect 669270 761094 676292 761154
rect 663057 760474 663123 760477
rect 669270 760474 669330 761094
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 663057 760472 669330 760474
rect 663057 760416 663062 760472
rect 663118 760416 669330 760472
rect 663057 760414 669330 760416
rect 663057 760411 663123 760414
rect 673269 760340 673335 760341
rect 673269 760338 673316 760340
rect 673224 760336 673316 760338
rect 673224 760280 673274 760336
rect 673224 760278 673316 760280
rect 673269 760276 673316 760278
rect 673380 760276 673386 760340
rect 673502 760278 676292 760338
rect 673269 760275 673335 760276
rect 671797 760066 671863 760069
rect 673502 760066 673562 760278
rect 671797 760064 673562 760066
rect 671797 760008 671802 760064
rect 671858 760008 673562 760064
rect 671797 760006 673562 760008
rect 671797 760003 671863 760006
rect 673686 759870 676292 759930
rect 672165 759794 672231 759797
rect 673686 759794 673746 759870
rect 672165 759792 673746 759794
rect 672165 759736 672170 759792
rect 672226 759736 673746 759792
rect 672165 759734 673746 759736
rect 672165 759731 672231 759734
rect 671429 759522 671495 759525
rect 671429 759520 676292 759522
rect 671429 759464 671434 759520
rect 671490 759464 676292 759520
rect 671429 759462 676292 759464
rect 671429 759459 671495 759462
rect 36537 759114 36603 759117
rect 41638 759114 41644 759116
rect 36537 759112 41644 759114
rect 36537 759056 36542 759112
rect 36598 759056 41644 759112
rect 36537 759054 41644 759056
rect 36537 759051 36603 759054
rect 41638 759052 41644 759054
rect 41708 759052 41714 759116
rect 673361 759114 673427 759117
rect 673361 759112 676292 759114
rect 673361 759056 673366 759112
rect 673422 759056 676292 759112
rect 673361 759054 676292 759056
rect 673361 759051 673427 759054
rect 42333 758844 42399 758845
rect 42333 758840 42380 758844
rect 42444 758842 42450 758844
rect 42333 758784 42338 758840
rect 42333 758780 42380 758784
rect 42444 758782 42490 758842
rect 42444 758780 42450 758782
rect 42333 758779 42399 758780
rect 672349 758706 672415 758709
rect 672349 758704 676292 758706
rect 672349 758648 672354 758704
rect 672410 758648 676292 758704
rect 672349 758646 676292 758648
rect 672349 758643 672415 758646
rect 40585 758434 40651 758437
rect 42333 758434 42399 758437
rect 40585 758432 42399 758434
rect 40585 758376 40590 758432
rect 40646 758376 42338 758432
rect 42394 758376 42399 758432
rect 40585 758374 42399 758376
rect 40585 758371 40651 758374
rect 42333 758371 42399 758374
rect 670969 758298 671035 758301
rect 670969 758296 676292 758298
rect 670969 758240 670974 758296
rect 671030 758240 676292 758296
rect 670969 758238 676292 758240
rect 670969 758235 671035 758238
rect 672441 757890 672507 757893
rect 672441 757888 676292 757890
rect 672441 757832 672446 757888
rect 672502 757832 676292 757888
rect 672441 757830 676292 757832
rect 672441 757827 672507 757830
rect 39297 757754 39363 757757
rect 42006 757754 42012 757756
rect 39297 757752 42012 757754
rect 39297 757696 39302 757752
rect 39358 757696 42012 757752
rect 39297 757694 42012 757696
rect 39297 757691 39363 757694
rect 42006 757692 42012 757694
rect 42076 757692 42082 757756
rect 671797 757482 671863 757485
rect 671797 757480 676292 757482
rect 671797 757424 671802 757480
rect 671858 757424 676292 757480
rect 671797 757422 676292 757424
rect 671797 757419 671863 757422
rect 41781 757076 41847 757077
rect 41781 757074 41828 757076
rect 41736 757072 41828 757074
rect 41736 757016 41786 757072
rect 41736 757014 41828 757016
rect 41781 757012 41828 757014
rect 41892 757012 41898 757076
rect 678237 757074 678303 757077
rect 678237 757072 678316 757074
rect 678237 757016 678242 757072
rect 678298 757016 678316 757072
rect 678237 757014 678316 757016
rect 41781 757011 41847 757012
rect 678237 757011 678303 757014
rect 683205 756666 683271 756669
rect 683205 756664 683284 756666
rect 683205 756608 683210 756664
rect 683266 756608 683284 756664
rect 683205 756606 683284 756608
rect 683205 756603 683271 756606
rect 673862 756332 673868 756396
rect 673932 756394 673938 756396
rect 676029 756394 676095 756397
rect 673932 756392 676095 756394
rect 673932 756336 676034 756392
rect 676090 756336 676095 756392
rect 673932 756334 676095 756336
rect 673932 756332 673938 756334
rect 676029 756331 676095 756334
rect 676170 756198 676292 756258
rect 669773 756122 669839 756125
rect 676170 756122 676230 756198
rect 669773 756120 676230 756122
rect 669773 756064 669778 756120
rect 669834 756064 676230 756120
rect 669773 756062 676230 756064
rect 669773 756059 669839 756062
rect 682377 755850 682443 755853
rect 682364 755848 682443 755850
rect 682364 755792 682382 755848
rect 682438 755792 682443 755848
rect 682364 755790 682443 755792
rect 682377 755787 682443 755790
rect 41873 755444 41939 755445
rect 41822 755442 41828 755444
rect 41782 755382 41828 755442
rect 41892 755440 41939 755444
rect 41934 755384 41939 755440
rect 41822 755380 41828 755382
rect 41892 755380 41939 755384
rect 41873 755379 41939 755380
rect 669270 755382 676292 755442
rect 668853 755306 668919 755309
rect 669270 755306 669330 755382
rect 668853 755304 669330 755306
rect 668853 755248 668858 755304
rect 668914 755248 669330 755304
rect 668853 755246 669330 755248
rect 668853 755243 668919 755246
rect 676949 755034 677015 755037
rect 676949 755032 677028 755034
rect 676949 754976 676954 755032
rect 677010 754976 677028 755032
rect 676949 754974 677028 754976
rect 676949 754971 677015 754974
rect 42190 754836 42196 754900
rect 42260 754898 42266 754900
rect 45185 754898 45251 754901
rect 42260 754896 45251 754898
rect 42260 754840 45190 754896
rect 45246 754840 45251 754896
rect 42260 754838 45251 754840
rect 42260 754836 42266 754838
rect 45185 754835 45251 754838
rect 42149 754626 42215 754629
rect 42374 754626 42380 754628
rect 42149 754624 42380 754626
rect 42149 754568 42154 754624
rect 42210 754568 42380 754624
rect 42149 754566 42380 754568
rect 42149 754563 42215 754566
rect 42374 754564 42380 754566
rect 42444 754564 42450 754628
rect 670601 754626 670667 754629
rect 670601 754624 676292 754626
rect 670601 754568 670606 754624
rect 670662 754568 676292 754624
rect 670601 754566 676292 754568
rect 670601 754563 670667 754566
rect 62113 754354 62179 754357
rect 674097 754354 674163 754357
rect 675845 754354 675911 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 674097 754352 675911 754354
rect 674097 754296 674102 754352
rect 674158 754296 675850 754352
rect 675906 754296 675911 754352
rect 674097 754294 675911 754296
rect 62113 754291 62179 754294
rect 674097 754291 674163 754294
rect 675845 754291 675911 754294
rect 42057 754218 42123 754221
rect 46197 754218 46263 754221
rect 42057 754216 46263 754218
rect 42057 754160 42062 754216
rect 42118 754160 46202 754216
rect 46258 754160 46263 754216
rect 42057 754158 46263 754160
rect 42057 754155 42123 754158
rect 46197 754155 46263 754158
rect 676032 754158 676292 754218
rect 676032 754082 676092 754158
rect 669270 754022 676092 754082
rect 42333 753946 42399 753949
rect 43345 753946 43411 753949
rect 42333 753944 43411 753946
rect 42333 753888 42338 753944
rect 42394 753888 43350 753944
rect 43406 753888 43411 753944
rect 42333 753886 43411 753888
rect 42333 753883 42399 753886
rect 43345 753883 43411 753886
rect 669270 753541 669330 754022
rect 676029 753810 676095 753813
rect 676029 753808 676292 753810
rect 676029 753752 676034 753808
rect 676090 753752 676292 753808
rect 676029 753750 676292 753752
rect 676029 753747 676095 753750
rect 669221 753536 669330 753541
rect 669221 753480 669226 753536
rect 669282 753480 669330 753536
rect 669221 753478 669330 753480
rect 669221 753475 669287 753478
rect 42149 753402 42215 753405
rect 42558 753402 42564 753404
rect 42149 753400 42564 753402
rect 42149 753344 42154 753400
rect 42210 753344 42564 753400
rect 42149 753342 42564 753344
rect 42149 753339 42215 753342
rect 42558 753340 42564 753342
rect 42628 753340 42634 753404
rect 671153 753402 671219 753405
rect 671153 753400 676292 753402
rect 671153 753344 671158 753400
rect 671214 753344 676292 753400
rect 671153 753342 676292 753344
rect 671153 753339 671219 753342
rect 41965 752994 42031 752997
rect 42190 752994 42196 752996
rect 41965 752992 42196 752994
rect 41965 752936 41970 752992
rect 42026 752936 42196 752992
rect 41965 752934 42196 752936
rect 41965 752931 42031 752934
rect 42190 752932 42196 752934
rect 42260 752932 42266 752996
rect 683389 752994 683455 752997
rect 683389 752992 683468 752994
rect 683389 752936 683394 752992
rect 683450 752936 683468 752992
rect 683389 752934 683468 752936
rect 683389 752931 683455 752934
rect 676029 752586 676095 752589
rect 676029 752584 676292 752586
rect 676029 752528 676034 752584
rect 676090 752528 676292 752584
rect 676029 752526 676292 752528
rect 676029 752523 676095 752526
rect 42190 752388 42196 752452
rect 42260 752450 42266 752452
rect 42425 752450 42491 752453
rect 42260 752448 42491 752450
rect 42260 752392 42430 752448
rect 42486 752392 42491 752448
rect 42260 752390 42491 752392
rect 42260 752388 42266 752390
rect 42425 752387 42491 752390
rect 42374 752116 42380 752180
rect 42444 752178 42450 752180
rect 42885 752178 42951 752181
rect 683113 752178 683179 752181
rect 42444 752176 42951 752178
rect 42444 752120 42890 752176
rect 42946 752120 42951 752176
rect 42444 752118 42951 752120
rect 683100 752176 683179 752178
rect 683100 752120 683118 752176
rect 683174 752120 683179 752176
rect 683100 752118 683179 752120
rect 42444 752116 42450 752118
rect 42885 752115 42951 752118
rect 683113 752115 683179 752118
rect 42149 751770 42215 751773
rect 42558 751770 42564 751772
rect 42149 751768 42564 751770
rect 42149 751712 42154 751768
rect 42210 751712 42564 751768
rect 42149 751710 42564 751712
rect 42149 751707 42215 751710
rect 42558 751708 42564 751710
rect 42628 751708 42634 751772
rect 672993 751770 673059 751773
rect 672993 751768 676292 751770
rect 672993 751712 672998 751768
rect 673054 751712 676292 751768
rect 672993 751710 676292 751712
rect 672993 751707 673059 751710
rect 671153 751362 671219 751365
rect 671153 751360 676292 751362
rect 671153 751304 671158 751360
rect 671214 751304 676292 751360
rect 671153 751302 676292 751304
rect 671153 751299 671219 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 669270 750924 676660 750954
rect 669270 750894 676690 750924
rect 669037 750818 669103 750821
rect 669270 750818 669330 750894
rect 669037 750816 669330 750818
rect 669037 750760 669042 750816
rect 669098 750760 669330 750816
rect 669037 750758 669330 750760
rect 669037 750755 669103 750758
rect 676630 750516 676690 750894
rect 40718 750348 40724 750412
rect 40788 750410 40794 750412
rect 41781 750410 41847 750413
rect 40788 750408 41847 750410
rect 40788 750352 41786 750408
rect 41842 750352 41847 750408
rect 40788 750350 41847 750352
rect 40788 750348 40794 750350
rect 41781 750347 41847 750350
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 670785 750138 670851 750141
rect 670785 750136 676292 750138
rect 670785 750080 670790 750136
rect 670846 750080 676292 750136
rect 670785 750078 676292 750080
rect 670785 750075 670851 750078
rect 42149 749730 42215 749733
rect 42885 749730 42951 749733
rect 42149 749728 42951 749730
rect 42149 749672 42154 749728
rect 42210 749672 42890 749728
rect 42946 749672 42951 749728
rect 42149 749670 42951 749672
rect 42149 749667 42215 749670
rect 42885 749667 42951 749670
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 40604 749398 42074 749458
rect 40604 749396 40610 749398
rect 42014 749189 42074 749398
rect 42014 749184 42123 749189
rect 42014 749128 42062 749184
rect 42118 749128 42123 749184
rect 42014 749126 42123 749128
rect 42057 749123 42123 749126
rect 42149 746874 42215 746877
rect 42374 746874 42380 746876
rect 42149 746872 42380 746874
rect 42149 746816 42154 746872
rect 42210 746816 42380 746872
rect 42149 746814 42380 746816
rect 42149 746811 42215 746814
rect 42374 746812 42380 746814
rect 42444 746812 42450 746876
rect 42149 745516 42215 745517
rect 42149 745514 42196 745516
rect 42104 745512 42196 745514
rect 42104 745456 42154 745512
rect 42104 745454 42196 745456
rect 42149 745452 42196 745454
rect 42260 745452 42266 745516
rect 42149 745451 42215 745452
rect 41638 745180 41644 745244
rect 41708 745242 41714 745244
rect 42701 745242 42767 745245
rect 41708 745240 42767 745242
rect 41708 745184 42706 745240
rect 42762 745184 42767 745240
rect 41708 745182 42767 745184
rect 41708 745180 41714 745182
rect 42701 745179 42767 745182
rect 41454 744908 41460 744972
rect 41524 744970 41530 744972
rect 42333 744970 42399 744973
rect 41524 744968 42399 744970
rect 41524 744912 42338 744968
rect 42394 744912 42399 744968
rect 41524 744910 42399 744912
rect 41524 744908 41530 744910
rect 42333 744907 42399 744910
rect 42006 744364 42012 744428
rect 42076 744426 42082 744428
rect 42793 744426 42859 744429
rect 42076 744424 42859 744426
rect 42076 744368 42798 744424
rect 42854 744368 42859 744424
rect 42076 744366 42859 744368
rect 42076 744364 42082 744366
rect 42793 744363 42859 744366
rect 667841 743202 667907 743205
rect 675109 743202 675175 743205
rect 667841 743200 675175 743202
rect 667841 743144 667846 743200
rect 667902 743144 675114 743200
rect 675170 743144 675175 743200
rect 667841 743142 675175 743144
rect 667841 743139 667907 743142
rect 675109 743139 675175 743142
rect 62757 743066 62823 743069
rect 51030 743064 62823 743066
rect 51030 743008 62762 743064
rect 62818 743008 62823 743064
rect 51030 743006 62823 743008
rect 42885 742794 42951 742797
rect 51030 742794 51090 743006
rect 62757 743003 62823 743006
rect 42885 742792 51090 742794
rect 42885 742736 42890 742792
rect 42946 742736 51090 742792
rect 42885 742734 51090 742736
rect 42885 742731 42951 742734
rect 666461 742522 666527 742525
rect 675293 742522 675359 742525
rect 666461 742520 675359 742522
rect 666461 742464 666466 742520
rect 666522 742464 675298 742520
rect 675354 742464 675359 742520
rect 666461 742462 675359 742464
rect 666461 742459 666527 742462
rect 675293 742459 675359 742462
rect 671470 742188 671476 742252
rect 671540 742250 671546 742252
rect 675109 742250 675175 742253
rect 671540 742248 675175 742250
rect 671540 742192 675114 742248
rect 675170 742192 675175 742248
rect 671540 742190 675175 742192
rect 671540 742188 671546 742190
rect 675109 742187 675175 742190
rect 673821 741706 673887 741709
rect 675477 741706 675543 741709
rect 673821 741704 675543 741706
rect 673821 741648 673826 741704
rect 673882 741648 675482 741704
rect 675538 741648 675543 741704
rect 673821 741646 675543 741648
rect 673821 741643 673887 741646
rect 675477 741643 675543 741646
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 669221 741162 669287 741165
rect 675109 741162 675175 741165
rect 669221 741160 675175 741162
rect 669221 741104 669226 741160
rect 669282 741104 675114 741160
rect 675170 741104 675175 741160
rect 669221 741102 675175 741104
rect 669221 741099 669287 741102
rect 675109 741099 675175 741102
rect 668761 738986 668827 738989
rect 674925 738986 674991 738989
rect 668761 738984 674991 738986
rect 668761 738928 668766 738984
rect 668822 738928 674930 738984
rect 674986 738928 674991 738984
rect 668761 738926 674991 738928
rect 668761 738923 668827 738926
rect 674925 738923 674991 738926
rect 674046 738652 674052 738716
rect 674116 738714 674122 738716
rect 675385 738714 675451 738717
rect 674116 738712 675451 738714
rect 674116 738656 675390 738712
rect 675446 738656 675451 738712
rect 674116 738654 675451 738656
rect 674116 738652 674122 738654
rect 675385 738651 675451 738654
rect 674414 738108 674420 738172
rect 674484 738170 674490 738172
rect 675109 738170 675175 738173
rect 674484 738168 675175 738170
rect 674484 738112 675114 738168
rect 675170 738112 675175 738168
rect 674484 738110 675175 738112
rect 674484 738108 674490 738110
rect 675109 738107 675175 738110
rect 652017 736810 652083 736813
rect 650164 736808 652083 736810
rect 650164 736752 652022 736808
rect 652078 736752 652083 736808
rect 650164 736750 652083 736752
rect 652017 736747 652083 736750
rect 668393 735314 668459 735317
rect 674925 735314 674991 735317
rect 668393 735312 674991 735314
rect 668393 735256 668398 735312
rect 668454 735256 674930 735312
rect 674986 735256 674991 735312
rect 668393 735254 674991 735256
rect 668393 735251 668459 735254
rect 674925 735251 674991 735254
rect 671337 734906 671403 734909
rect 675109 734906 675175 734909
rect 671337 734904 675175 734906
rect 671337 734848 671342 734904
rect 671398 734848 675114 734904
rect 675170 734848 675175 734904
rect 671337 734846 675175 734848
rect 671337 734843 671403 734846
rect 675109 734843 675175 734846
rect 672349 734226 672415 734229
rect 675109 734226 675175 734229
rect 672349 734224 675175 734226
rect 672349 734168 672354 734224
rect 672410 734168 675114 734224
rect 675170 734168 675175 734224
rect 672349 734166 675175 734168
rect 672349 734163 672415 734166
rect 675109 734163 675175 734166
rect 669037 733682 669103 733685
rect 675109 733682 675175 733685
rect 669037 733680 675175 733682
rect 669037 733624 669042 733680
rect 669098 733624 675114 733680
rect 675170 733624 675175 733680
rect 669037 733622 675175 733624
rect 669037 733619 669103 733622
rect 675109 733619 675175 733622
rect 673177 733002 673243 733005
rect 675293 733002 675359 733005
rect 673177 733000 675359 733002
rect 673177 732944 673182 733000
rect 673238 732944 675298 733000
rect 675354 732944 675359 733000
rect 673177 732942 675359 732944
rect 673177 732939 673243 732942
rect 675293 732939 675359 732942
rect 671981 732868 672047 732869
rect 671981 732864 672028 732868
rect 672092 732866 672098 732868
rect 671981 732808 671986 732864
rect 671981 732804 672028 732808
rect 672092 732806 672138 732866
rect 672092 732804 672098 732806
rect 671981 732803 672047 732804
rect 669773 731506 669839 731509
rect 674925 731506 674991 731509
rect 669773 731504 674991 731506
rect 669773 731448 669778 731504
rect 669834 731448 674930 731504
rect 674986 731448 674991 731504
rect 669773 731446 674991 731448
rect 669773 731443 669839 731446
rect 674925 731443 674991 731446
rect 44817 731370 44883 731373
rect 41492 731368 44883 731370
rect 41492 731312 44822 731368
rect 44878 731312 44883 731368
rect 41492 731310 44883 731312
rect 44817 731307 44883 731310
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 670601 730554 670667 730557
rect 675293 730554 675359 730557
rect 670601 730552 675359 730554
rect 670601 730496 670606 730552
rect 670662 730496 675298 730552
rect 675354 730496 675359 730552
rect 670601 730494 675359 730496
rect 670601 730491 670667 730494
rect 675293 730491 675359 730494
rect 44173 730146 44239 730149
rect 41492 730144 44239 730146
rect 41492 730088 44178 730144
rect 44234 730088 44239 730144
rect 41492 730086 44239 730088
rect 44173 730083 44239 730086
rect 671981 730146 672047 730149
rect 675109 730146 675175 730149
rect 671981 730144 675175 730146
rect 671981 730088 671986 730144
rect 672042 730088 675114 730144
rect 675170 730088 675175 730144
rect 671981 730086 675175 730088
rect 671981 730083 672047 730086
rect 675109 730083 675175 730086
rect 675886 729948 675892 730012
rect 675956 730010 675962 730012
rect 676806 730010 676812 730012
rect 675956 729950 676812 730010
rect 675956 729948 675962 729950
rect 676806 729948 676812 729950
rect 676876 729948 676882 730012
rect 44265 729738 44331 729741
rect 41492 729736 44331 729738
rect 41492 729680 44270 729736
rect 44326 729680 44331 729736
rect 41492 729678 44331 729680
rect 44265 729675 44331 729678
rect 44449 729330 44515 729333
rect 41492 729328 44515 729330
rect 41492 729272 44454 729328
rect 44510 729272 44515 729328
rect 41492 729270 44515 729272
rect 44449 729267 44515 729270
rect 45185 728922 45251 728925
rect 41492 728920 45251 728922
rect 41492 728864 45190 728920
rect 45246 728864 45251 728920
rect 41492 728862 45251 728864
rect 45185 728859 45251 728862
rect 673310 728588 673316 728652
rect 673380 728650 673386 728652
rect 674097 728650 674163 728653
rect 673380 728648 674163 728650
rect 673380 728592 674102 728648
rect 674158 728592 674163 728648
rect 673380 728590 674163 728592
rect 673380 728588 673386 728590
rect 674097 728587 674163 728590
rect 44633 728514 44699 728517
rect 41492 728512 44699 728514
rect 41492 728456 44638 728512
rect 44694 728456 44699 728512
rect 41492 728454 44699 728456
rect 44633 728451 44699 728454
rect 672022 728452 672028 728516
rect 672092 728514 672098 728516
rect 673085 728514 673151 728517
rect 672092 728512 673151 728514
rect 672092 728456 673090 728512
rect 673146 728456 673151 728512
rect 672092 728454 673151 728456
rect 672092 728452 672098 728454
rect 673085 728451 673151 728454
rect 62757 728242 62823 728245
rect 671153 728242 671219 728245
rect 673913 728242 673979 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 671153 728240 673979 728242
rect 671153 728184 671158 728240
rect 671214 728184 673918 728240
rect 673974 728184 673979 728240
rect 671153 728182 673979 728184
rect 62757 728179 62823 728182
rect 671153 728179 671219 728182
rect 673913 728179 673979 728182
rect 44817 728106 44883 728109
rect 41492 728104 44883 728106
rect 41492 728048 44822 728104
rect 44878 728048 44883 728104
rect 41492 728046 44883 728048
rect 44817 728043 44883 728046
rect 670785 727970 670851 727973
rect 674143 727970 674209 727973
rect 670785 727968 674209 727970
rect 670785 727912 670790 727968
rect 670846 727912 674148 727968
rect 674204 727912 674209 727968
rect 670785 727910 674209 727912
rect 670785 727907 670851 727910
rect 674143 727907 674209 727910
rect 45001 727698 45067 727701
rect 41492 727696 45067 727698
rect 41492 727640 45006 727696
rect 45062 727640 45067 727696
rect 41492 727638 45067 727640
rect 45001 727635 45067 727638
rect 44633 727290 44699 727293
rect 41492 727288 44699 727290
rect 41492 727232 44638 727288
rect 44694 727232 44699 727288
rect 41492 727230 44699 727232
rect 44633 727227 44699 727230
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 674281 726882 674347 726885
rect 683113 726882 683179 726885
rect 674281 726880 683179 726882
rect 674281 726824 674286 726880
rect 674342 726824 683118 726880
rect 683174 726824 683179 726880
rect 674281 726822 683179 726824
rect 674281 726819 674347 726822
rect 683113 726819 683179 726822
rect 674557 726610 674623 726613
rect 674557 726608 678990 726610
rect 674557 726552 674562 726608
rect 674618 726552 678990 726608
rect 674557 726550 678990 726552
rect 674557 726547 674623 726550
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 678930 726474 678990 726550
rect 683389 726474 683455 726477
rect 678930 726472 683455 726474
rect 678930 726416 683394 726472
rect 683450 726416 683455 726472
rect 678930 726414 683455 726416
rect 41321 726411 41387 726414
rect 683389 726411 683455 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 680997 725794 681063 725797
rect 676140 725792 681063 725794
rect 676140 725736 681002 725792
rect 681058 725736 681063 725792
rect 676140 725734 681063 725736
rect 676140 725732 676146 725734
rect 680997 725731 681063 725734
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 672901 725522 672967 725525
rect 683573 725522 683639 725525
rect 672901 725520 683639 725522
rect 672901 725464 672906 725520
rect 672962 725464 683578 725520
rect 683634 725464 683639 725520
rect 672901 725462 683639 725464
rect 672901 725459 672967 725462
rect 683573 725459 683639 725462
rect 33777 725250 33843 725253
rect 33764 725248 33843 725250
rect 33764 725192 33782 725248
rect 33838 725192 33843 725248
rect 33764 725190 33843 725192
rect 33777 725187 33843 725190
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 31661 724434 31727 724437
rect 31661 724432 31740 724434
rect 31661 724376 31666 724432
rect 31722 724376 31740 724432
rect 31661 724374 31740 724376
rect 31661 724371 31727 724374
rect 34513 724026 34579 724029
rect 34500 724024 34579 724026
rect 34500 723968 34518 724024
rect 34574 723968 34579 724024
rect 34500 723966 34579 723968
rect 34513 723963 34579 723966
rect 673637 724026 673703 724029
rect 677317 724026 677383 724029
rect 673637 724024 677383 724026
rect 673637 723968 673642 724024
rect 673698 723968 677322 724024
rect 677378 723968 677383 724024
rect 673637 723966 677383 723968
rect 673637 723963 673703 723966
rect 677317 723963 677383 723966
rect 45001 723618 45067 723621
rect 41492 723616 45067 723618
rect 41492 723560 45006 723616
rect 45062 723560 45067 723616
rect 41492 723558 45067 723560
rect 45001 723555 45067 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 40677 723210 40743 723213
rect 40677 723208 40756 723210
rect 40677 723152 40682 723208
rect 40738 723152 40756 723208
rect 40677 723150 40756 723152
rect 40677 723147 40743 723150
rect 44173 722802 44239 722805
rect 41492 722800 44239 722802
rect 41492 722744 44178 722800
rect 44234 722744 44239 722800
rect 41492 722742 44239 722744
rect 44173 722739 44239 722742
rect 41822 722394 41828 722396
rect 41492 722334 41828 722394
rect 41822 722332 41828 722334
rect 41892 722332 41898 722396
rect 40726 721772 40786 721956
rect 40350 721708 40356 721772
rect 40420 721708 40426 721772
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 40358 721548 40418 721708
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 45553 721170 45619 721173
rect 41492 721168 45619 721170
rect 41492 721112 45558 721168
rect 45614 721112 45619 721168
rect 41492 721110 45619 721112
rect 45553 721107 45619 721110
rect 38745 720354 38811 720357
rect 38732 720352 38811 720354
rect 38732 720296 38750 720352
rect 38806 720296 38811 720352
rect 38732 720294 38811 720296
rect 38745 720291 38811 720294
rect 39852 720234 39992 720764
rect 46105 719946 46171 719949
rect 41492 719944 46171 719946
rect 41492 719888 46110 719944
rect 46166 719888 46171 719944
rect 41492 719886 46171 719888
rect 46105 719883 46171 719886
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41822 718586 41828 718588
rect 40604 718526 41828 718586
rect 40604 718524 40610 718526
rect 41822 718524 41828 718526
rect 41892 718524 41898 718588
rect 40350 716756 40356 716820
rect 40420 716818 40426 716820
rect 40902 716818 40908 716820
rect 40420 716758 40908 716818
rect 40420 716756 40426 716758
rect 40902 716756 40908 716758
rect 40972 716756 40978 716820
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 663750 716078 676292 716138
rect 658917 716002 658983 716005
rect 663750 716002 663810 716078
rect 658917 716000 663810 716002
rect 658917 715944 658922 716000
rect 658978 715944 663810 716000
rect 658917 715942 663810 715944
rect 658917 715939 658983 715942
rect 40309 715730 40375 715733
rect 42057 715730 42123 715733
rect 40309 715728 42123 715730
rect 40309 715672 40314 715728
rect 40370 715672 42062 715728
rect 42118 715672 42123 715728
rect 40309 715670 42123 715672
rect 40309 715667 40375 715670
rect 42057 715667 42123 715670
rect 669957 715730 670023 715733
rect 669957 715728 676292 715730
rect 669957 715672 669962 715728
rect 670018 715672 676292 715728
rect 669957 715670 676292 715672
rect 669957 715667 670023 715670
rect 31661 715458 31727 715461
rect 41822 715458 41828 715460
rect 31661 715456 41828 715458
rect 31661 715400 31666 715456
rect 31722 715400 41828 715456
rect 31661 715398 41828 715400
rect 31661 715395 31727 715398
rect 41822 715396 41828 715398
rect 41892 715396 41898 715460
rect 62113 715322 62179 715325
rect 672165 715322 672231 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 672165 715320 676292 715322
rect 672165 715264 672170 715320
rect 672226 715264 676292 715320
rect 672165 715262 676292 715264
rect 62113 715259 62179 715262
rect 672165 715259 672231 715262
rect 41689 715186 41755 715189
rect 42701 715186 42767 715189
rect 41689 715184 42767 715186
rect 41689 715128 41694 715184
rect 41750 715128 42706 715184
rect 42762 715128 42767 715184
rect 41689 715126 42767 715128
rect 41689 715123 41755 715126
rect 42701 715123 42767 715126
rect 672901 714914 672967 714917
rect 672901 714912 676292 714914
rect 672901 714856 672906 714912
rect 672962 714856 676292 714912
rect 672901 714854 676292 714856
rect 672901 714851 672967 714854
rect 41873 714642 41939 714645
rect 42425 714642 42491 714645
rect 41873 714640 42491 714642
rect 41873 714584 41878 714640
rect 41934 714584 42430 714640
rect 42486 714584 42491 714640
rect 41873 714582 42491 714584
rect 41873 714579 41939 714582
rect 42425 714579 42491 714582
rect 673361 714506 673427 714509
rect 673361 714504 676292 714506
rect 673361 714448 673366 714504
rect 673422 714448 676292 714504
rect 673361 714446 676292 714448
rect 673361 714443 673427 714446
rect 42057 714372 42123 714373
rect 42006 714308 42012 714372
rect 42076 714370 42123 714372
rect 42076 714368 42168 714370
rect 42118 714312 42168 714368
rect 42076 714310 42168 714312
rect 42076 714308 42123 714310
rect 42057 714307 42123 714308
rect 38745 714234 38811 714237
rect 40350 714234 40356 714236
rect 38745 714232 40356 714234
rect 38745 714176 38750 714232
rect 38806 714176 40356 714232
rect 38745 714174 40356 714176
rect 38745 714171 38811 714174
rect 40350 714172 40356 714174
rect 40420 714172 40426 714236
rect 40677 714234 40743 714237
rect 41086 714234 41092 714236
rect 40677 714232 41092 714234
rect 40677 714176 40682 714232
rect 40738 714176 41092 714232
rect 40677 714174 41092 714176
rect 40677 714171 40743 714174
rect 41086 714172 41092 714174
rect 41156 714172 41162 714236
rect 41413 714234 41479 714237
rect 41413 714232 41522 714234
rect 41413 714176 41418 714232
rect 41474 714176 41522 714232
rect 41413 714171 41522 714176
rect 41462 713554 41522 714171
rect 42701 714100 42767 714101
rect 42701 714096 42748 714100
rect 42812 714098 42818 714100
rect 671153 714098 671219 714101
rect 42701 714040 42706 714096
rect 42701 714036 42748 714040
rect 42812 714038 42858 714098
rect 671153 714096 676292 714098
rect 671153 714040 671158 714096
rect 671214 714040 676292 714096
rect 671153 714038 676292 714040
rect 42812 714036 42818 714038
rect 42701 714035 42767 714036
rect 671153 714035 671219 714038
rect 670969 713690 671035 713693
rect 670969 713688 676292 713690
rect 670969 713632 670974 713688
rect 671030 713632 676292 713688
rect 670969 713630 676292 713632
rect 670969 713627 671035 713630
rect 41781 713554 41847 713557
rect 41462 713552 41847 713554
rect 41462 713496 41786 713552
rect 41842 713496 41847 713552
rect 41462 713494 41847 713496
rect 41781 713491 41847 713494
rect 42241 713282 42307 713285
rect 42609 713282 42675 713285
rect 42241 713280 42675 713282
rect 42241 713224 42246 713280
rect 42302 713224 42614 713280
rect 42670 713224 42675 713280
rect 42241 713222 42675 713224
rect 42241 713219 42307 713222
rect 42609 713219 42675 713222
rect 670969 713282 671035 713285
rect 670969 713280 676292 713282
rect 670969 713224 670974 713280
rect 671030 713224 676292 713280
rect 670969 713222 676292 713224
rect 670969 713219 671035 713222
rect 671797 712874 671863 712877
rect 671797 712872 676292 712874
rect 671797 712816 671802 712872
rect 671858 712816 676292 712872
rect 671797 712814 676292 712816
rect 671797 712811 671863 712814
rect 673269 712466 673335 712469
rect 673269 712464 676292 712466
rect 673269 712408 673274 712464
rect 673330 712408 676292 712464
rect 673269 712406 676292 712408
rect 673269 712403 673335 712406
rect 40350 712132 40356 712196
rect 40420 712194 40426 712196
rect 41781 712194 41847 712197
rect 47577 712194 47643 712197
rect 40420 712192 41847 712194
rect 40420 712136 41786 712192
rect 41842 712136 41847 712192
rect 40420 712134 41847 712136
rect 40420 712132 40426 712134
rect 41781 712131 41847 712134
rect 42198 712192 47643 712194
rect 42198 712136 47582 712192
rect 47638 712136 47643 712192
rect 42198 712134 47643 712136
rect 42198 711109 42258 712134
rect 47577 712131 47643 712134
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 666277 711650 666343 711653
rect 666277 711648 676292 711650
rect 666277 711592 666282 711648
rect 666338 711592 676292 711648
rect 666277 711590 676292 711592
rect 666277 711587 666343 711590
rect 683389 711242 683455 711245
rect 683389 711240 683468 711242
rect 683389 711184 683394 711240
rect 683450 711184 683468 711240
rect 683389 711182 683468 711184
rect 683389 711179 683455 711182
rect 42198 711104 42307 711109
rect 42198 711048 42246 711104
rect 42302 711048 42307 711104
rect 42198 711046 42307 711048
rect 42241 711043 42307 711046
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 672625 710426 672691 710429
rect 672625 710424 676292 710426
rect 672625 710368 672630 710424
rect 672686 710368 676292 710424
rect 672625 710366 676292 710368
rect 672625 710363 672691 710366
rect 651465 710290 651531 710293
rect 650164 710288 651531 710290
rect 650164 710232 651470 710288
rect 651526 710232 651531 710288
rect 650164 710230 651531 710232
rect 651465 710227 651531 710230
rect 42701 710020 42767 710021
rect 42701 710018 42748 710020
rect 42656 710016 42748 710018
rect 42656 709960 42706 710016
rect 42656 709958 42748 709960
rect 42701 709956 42748 709958
rect 42812 709956 42818 710020
rect 670141 710018 670207 710021
rect 670141 710016 676292 710018
rect 670141 709960 670146 710016
rect 670202 709960 676292 710016
rect 670141 709958 676292 709960
rect 42701 709955 42767 709956
rect 670141 709955 670207 709958
rect 41086 709820 41092 709884
rect 41156 709882 41162 709884
rect 41781 709882 41847 709885
rect 41156 709880 41847 709882
rect 41156 709824 41786 709880
rect 41842 709824 41847 709880
rect 41156 709822 41847 709824
rect 41156 709820 41162 709822
rect 41781 709819 41847 709822
rect 668209 709610 668275 709613
rect 668209 709608 676292 709610
rect 668209 709552 668214 709608
rect 668270 709552 676292 709608
rect 668209 709550 676292 709552
rect 668209 709547 668275 709550
rect 40718 709412 40724 709476
rect 40788 709474 40794 709476
rect 40788 709414 42120 709474
rect 40788 709412 40794 709414
rect 42060 709069 42120 709414
rect 672625 709202 672691 709205
rect 672625 709200 676292 709202
rect 672625 709144 672630 709200
rect 672686 709144 676292 709200
rect 672625 709142 676292 709144
rect 672625 709139 672691 709142
rect 42057 709064 42123 709069
rect 42057 709008 42062 709064
rect 42118 709008 42123 709064
rect 42057 709003 42123 709008
rect 669589 708794 669655 708797
rect 669589 708792 676292 708794
rect 669589 708736 669594 708792
rect 669650 708736 676292 708792
rect 669589 708734 676292 708736
rect 669589 708731 669655 708734
rect 40902 708460 40908 708524
rect 40972 708522 40978 708524
rect 41781 708522 41847 708525
rect 40972 708520 41847 708522
rect 40972 708464 41786 708520
rect 41842 708464 41847 708520
rect 40972 708462 41847 708464
rect 40972 708460 40978 708462
rect 41781 708459 41847 708462
rect 683573 708386 683639 708389
rect 683573 708384 683652 708386
rect 683573 708328 683578 708384
rect 683634 708328 683652 708384
rect 683573 708326 683652 708328
rect 683573 708323 683639 708326
rect 683849 707978 683915 707981
rect 683836 707976 683915 707978
rect 683836 707920 683854 707976
rect 683910 707920 683915 707976
rect 683836 707918 683915 707920
rect 683849 707915 683915 707918
rect 42057 707842 42123 707845
rect 44173 707842 44239 707845
rect 42057 707840 44239 707842
rect 42057 707784 42062 707840
rect 42118 707784 44178 707840
rect 44234 707784 44239 707840
rect 42057 707782 44239 707784
rect 42057 707779 42123 707782
rect 44173 707779 44239 707782
rect 674230 707508 674236 707572
rect 674300 707570 674306 707572
rect 674300 707510 676292 707570
rect 674300 707508 674306 707510
rect 670325 707162 670391 707165
rect 670325 707160 676292 707162
rect 670325 707104 670330 707160
rect 670386 707104 676292 707160
rect 670325 707102 676292 707104
rect 670325 707099 670391 707102
rect 40534 706692 40540 706756
rect 40604 706754 40610 706756
rect 42241 706754 42307 706757
rect 683113 706754 683179 706757
rect 40604 706752 42307 706754
rect 40604 706696 42246 706752
rect 42302 706696 42307 706752
rect 40604 706694 42307 706696
rect 683100 706752 683179 706754
rect 683100 706696 683118 706752
rect 683174 706696 683179 706752
rect 683100 706694 683179 706696
rect 40604 706692 40610 706694
rect 42241 706691 42307 706694
rect 683113 706691 683179 706694
rect 41965 706484 42031 706485
rect 41965 706480 42012 706484
rect 42076 706482 42082 706484
rect 41965 706424 41970 706480
rect 41965 706420 42012 706424
rect 42076 706422 42122 706482
rect 42076 706420 42082 706422
rect 41965 706419 42031 706420
rect 674598 706284 674604 706348
rect 674668 706346 674674 706348
rect 674668 706286 676292 706346
rect 674668 706284 674674 706286
rect 671613 705530 671679 705533
rect 676262 705530 676322 705908
rect 671613 705528 676322 705530
rect 671613 705472 671618 705528
rect 671674 705500 676322 705528
rect 671674 705472 676292 705500
rect 671613 705470 676292 705472
rect 671613 705467 671679 705470
rect 42241 705258 42307 705261
rect 45001 705258 45067 705261
rect 42241 705256 45067 705258
rect 42241 705200 42246 705256
rect 42302 705200 45006 705256
rect 45062 705200 45067 705256
rect 42241 705198 45067 705200
rect 42241 705195 42307 705198
rect 45001 705195 45067 705198
rect 673361 705122 673427 705125
rect 673361 705120 676292 705122
rect 673361 705064 673366 705120
rect 673422 705064 676292 705120
rect 673361 705062 676292 705064
rect 673361 705059 673427 705062
rect 42241 704580 42307 704581
rect 42190 704578 42196 704580
rect 42150 704518 42196 704578
rect 42260 704576 42307 704580
rect 42302 704520 42307 704576
rect 42190 704516 42196 704518
rect 42260 704516 42307 704520
rect 42241 704515 42307 704516
rect 42149 703492 42215 703493
rect 42149 703490 42196 703492
rect 42104 703488 42196 703490
rect 42104 703432 42154 703488
rect 42104 703430 42196 703432
rect 42149 703428 42196 703430
rect 42260 703428 42266 703492
rect 42149 703427 42215 703428
rect 42057 702810 42123 702813
rect 42701 702810 42767 702813
rect 42057 702808 42767 702810
rect 42057 702752 42062 702808
rect 42118 702752 42706 702808
rect 42762 702752 42767 702808
rect 42057 702750 42767 702752
rect 42057 702747 42123 702750
rect 42701 702747 42767 702750
rect 41638 702340 41644 702404
rect 41708 702402 41714 702404
rect 42609 702402 42675 702405
rect 41708 702400 42675 702402
rect 41708 702344 42614 702400
rect 42670 702344 42675 702400
rect 41708 702342 42675 702344
rect 41708 702340 41714 702342
rect 42609 702339 42675 702342
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 669589 701178 669655 701181
rect 675109 701178 675175 701181
rect 669589 701176 675175 701178
rect 669589 701120 669594 701176
rect 669650 701120 675114 701176
rect 675170 701120 675175 701176
rect 669589 701118 675175 701120
rect 669589 701115 669655 701118
rect 675109 701115 675175 701118
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 41781 699820 41847 699821
rect 41781 699816 41828 699820
rect 41892 699818 41898 699820
rect 41781 699760 41786 699816
rect 41781 699756 41828 699760
rect 41892 699758 41938 699818
rect 41892 699756 41898 699758
rect 41781 699755 41847 699756
rect 651465 696962 651531 696965
rect 650164 696960 651531 696962
rect 650164 696904 651470 696960
rect 651526 696904 651531 696960
rect 650164 696902 651531 696904
rect 651465 696899 651531 696902
rect 670417 696962 670483 696965
rect 675109 696962 675175 696965
rect 670417 696960 675175 696962
rect 670417 696904 670422 696960
rect 670478 696904 675114 696960
rect 675170 696904 675175 696960
rect 670417 696902 675175 696904
rect 670417 696899 670483 696902
rect 675109 696899 675175 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676990 694106 676996 694108
rect 675894 694046 676996 694106
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 668393 692882 668459 692885
rect 675109 692882 675175 692885
rect 668393 692880 675175 692882
rect 668393 692824 668398 692880
rect 668454 692824 675114 692880
rect 675170 692824 675175 692880
rect 668393 692822 675175 692824
rect 668393 692819 668459 692822
rect 675109 692819 675175 692822
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 673821 690162 673887 690165
rect 675385 690162 675451 690165
rect 673821 690160 675451 690162
rect 673821 690104 673826 690160
rect 673882 690104 675390 690160
rect 675446 690104 675451 690160
rect 673821 690102 675451 690104
rect 673821 690099 673887 690102
rect 675385 690099 675451 690102
rect 674649 689618 674715 689621
rect 675293 689618 675359 689621
rect 674649 689616 675359 689618
rect 674649 689560 674654 689616
rect 674710 689560 675298 689616
rect 675354 689560 675359 689616
rect 674649 689558 675359 689560
rect 674649 689555 674715 689558
rect 675293 689555 675359 689558
rect 62757 689482 62823 689485
rect 45510 689480 62823 689482
rect 45510 689424 62762 689480
rect 62818 689424 62823 689480
rect 45510 689422 62823 689424
rect 41413 689346 41479 689349
rect 45510 689346 45570 689422
rect 62757 689419 62823 689422
rect 41413 689344 45570 689346
rect 41413 689288 41418 689344
rect 41474 689288 45570 689344
rect 41413 689286 45570 689288
rect 663057 689346 663123 689349
rect 674925 689346 674991 689349
rect 663057 689344 674991 689346
rect 663057 689288 663062 689344
rect 663118 689288 674930 689344
rect 674986 689288 674991 689344
rect 663057 689286 674991 689288
rect 41413 689283 41479 689286
rect 663057 689283 663123 689286
rect 674925 689283 674991 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 672165 689074 672231 689077
rect 675109 689074 675175 689077
rect 672165 689072 675175 689074
rect 672165 689016 672170 689072
rect 672226 689016 675114 689072
rect 675170 689016 675175 689072
rect 672165 689014 675175 689016
rect 672165 689011 672231 689014
rect 675109 689011 675175 689014
rect 667657 688938 667723 688941
rect 667657 688936 669330 688938
rect 667657 688880 667662 688936
rect 667718 688880 669330 688936
rect 667657 688878 669330 688880
rect 667657 688875 667723 688878
rect 669270 688802 669330 688878
rect 674925 688802 674991 688805
rect 669270 688800 674991 688802
rect 669270 688744 674930 688800
rect 674986 688744 674991 688800
rect 669270 688742 674991 688744
rect 674925 688739 674991 688742
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 671797 687442 671863 687445
rect 675477 687442 675543 687445
rect 671797 687440 675543 687442
rect 671797 687384 671802 687440
rect 671858 687384 675482 687440
rect 675538 687384 675543 687440
rect 671797 687382 675543 687384
rect 671797 687379 671863 687382
rect 675477 687379 675543 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 674925 687170 674991 687173
rect 675334 687170 675340 687172
rect 674925 687168 675340 687170
rect 674925 687112 674930 687168
rect 674986 687112 675340 687168
rect 674925 687110 675340 687112
rect 674925 687107 674991 687110
rect 675334 687108 675340 687110
rect 675404 687108 675410 687172
rect 44357 686898 44423 686901
rect 41492 686896 44423 686898
rect 41492 686840 44362 686896
rect 44418 686840 44423 686896
rect 41492 686838 44423 686840
rect 44357 686835 44423 686838
rect 44357 686490 44423 686493
rect 41492 686488 44423 686490
rect 41492 686432 44362 686488
rect 44418 686432 44423 686488
rect 41492 686430 44423 686432
rect 44357 686427 44423 686430
rect 45185 686082 45251 686085
rect 41492 686080 45251 686082
rect 41492 686024 45190 686080
rect 45246 686024 45251 686080
rect 41492 686022 45251 686024
rect 45185 686019 45251 686022
rect 670141 685946 670207 685949
rect 675201 685946 675267 685949
rect 670141 685944 675267 685946
rect 670141 685888 670146 685944
rect 670202 685888 675206 685944
rect 675262 685888 675267 685944
rect 670141 685886 675267 685888
rect 670141 685883 670207 685886
rect 675201 685883 675267 685886
rect 45185 685674 45251 685677
rect 41492 685672 45251 685674
rect 41492 685616 45190 685672
rect 45246 685616 45251 685672
rect 41492 685614 45251 685616
rect 45185 685611 45251 685614
rect 668209 685538 668275 685541
rect 675477 685538 675543 685541
rect 668209 685536 675543 685538
rect 668209 685480 668214 685536
rect 668270 685480 675482 685536
rect 675538 685480 675543 685536
rect 668209 685478 675543 685480
rect 668209 685475 668275 685478
rect 675477 685475 675543 685478
rect 44817 685266 44883 685269
rect 41492 685264 44883 685266
rect 41492 685208 44822 685264
rect 44878 685208 44883 685264
rect 41492 685206 44883 685208
rect 44817 685203 44883 685206
rect 44173 684858 44239 684861
rect 41492 684856 44239 684858
rect 41492 684800 44178 684856
rect 44234 684800 44239 684856
rect 41492 684798 44239 684800
rect 44173 684795 44239 684798
rect 44633 684450 44699 684453
rect 41492 684448 44699 684450
rect 41492 684392 44638 684448
rect 44694 684392 44699 684448
rect 41492 684390 44699 684392
rect 44633 684387 44699 684390
rect 45001 684042 45067 684045
rect 41492 684040 45067 684042
rect 41492 683984 45006 684040
rect 45062 683984 45067 684040
rect 41492 683982 45067 683984
rect 45001 683979 45067 683982
rect 35801 683634 35867 683637
rect 651649 683634 651715 683637
rect 35788 683632 35867 683634
rect 35788 683576 35806 683632
rect 35862 683576 35867 683632
rect 35788 683574 35867 683576
rect 650164 683632 651715 683634
rect 650164 683576 651654 683632
rect 651710 683576 651715 683632
rect 650164 683574 651715 683576
rect 35801 683571 35867 683574
rect 651649 683571 651715 683574
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35433 682818 35499 682821
rect 35420 682816 35499 682818
rect 35420 682760 35438 682816
rect 35494 682760 35499 682816
rect 35420 682758 35499 682760
rect 35433 682755 35499 682758
rect 35617 682410 35683 682413
rect 35604 682408 35683 682410
rect 35604 682352 35622 682408
rect 35678 682352 35683 682408
rect 35604 682350 35683 682352
rect 35617 682347 35683 682350
rect 673637 682410 673703 682413
rect 683205 682410 683271 682413
rect 673637 682408 683271 682410
rect 673637 682352 673642 682408
rect 673698 682352 683210 682408
rect 683266 682352 683271 682408
rect 673637 682350 683271 682352
rect 673637 682347 673703 682350
rect 683205 682347 683271 682350
rect 35801 682002 35867 682005
rect 35788 682000 35867 682002
rect 35788 681944 35806 682000
rect 35862 681944 35867 682000
rect 35788 681942 35867 681944
rect 35801 681939 35867 681942
rect 41689 681866 41755 681869
rect 42609 681866 42675 681869
rect 41689 681864 42675 681866
rect 41689 681808 41694 681864
rect 41750 681808 42614 681864
rect 42670 681808 42675 681864
rect 41689 681806 42675 681808
rect 41689 681803 41755 681806
rect 42609 681803 42675 681806
rect 32397 681594 32463 681597
rect 32397 681592 32476 681594
rect 32397 681536 32402 681592
rect 32458 681536 32476 681592
rect 32397 681534 32476 681536
rect 32397 681531 32463 681534
rect 31017 681186 31083 681189
rect 31004 681184 31083 681186
rect 31004 681128 31022 681184
rect 31078 681128 31083 681184
rect 31004 681126 31083 681128
rect 31017 681123 31083 681126
rect 674046 680988 674052 681052
rect 674116 681050 674122 681052
rect 683389 681050 683455 681053
rect 674116 681048 683455 681050
rect 674116 680992 683394 681048
rect 683450 680992 683455 681048
rect 674116 680990 683455 680992
rect 674116 680988 674122 680990
rect 683389 680987 683455 680990
rect 35617 680778 35683 680781
rect 35604 680776 35683 680778
rect 35604 680720 35622 680776
rect 35678 680720 35683 680776
rect 35604 680718 35683 680720
rect 35617 680715 35683 680718
rect 44541 680370 44607 680373
rect 41492 680368 44607 680370
rect 41492 680312 44546 680368
rect 44602 680312 44607 680368
rect 41492 680310 44607 680312
rect 44541 680307 44607 680310
rect 42885 679962 42951 679965
rect 41492 679960 42951 679962
rect 41492 679904 42890 679960
rect 42946 679904 42951 679960
rect 41492 679902 42951 679904
rect 42885 679899 42951 679902
rect 44725 679554 44791 679557
rect 41492 679552 44791 679554
rect 41492 679496 44730 679552
rect 44786 679496 44791 679552
rect 41492 679494 44791 679496
rect 44725 679491 44791 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40726 678708 40786 678928
rect 41822 678330 41828 678332
rect 41492 678270 41828 678330
rect 41822 678268 41828 678270
rect 41892 678268 41898 678332
rect 47209 677922 47275 677925
rect 41492 677920 47275 677922
rect 41492 677864 47214 677920
rect 47270 677864 47275 677920
rect 41492 677862 47275 677864
rect 47209 677859 47275 677862
rect 41781 677652 41847 677653
rect 41781 677648 41828 677652
rect 41892 677650 41898 677652
rect 41781 677592 41786 677648
rect 41781 677588 41828 677592
rect 41892 677590 41938 677650
rect 41892 677588 41898 677590
rect 41781 677587 41847 677588
rect 37230 677109 37290 677484
rect 37181 677104 37290 677109
rect 37181 677048 37186 677104
rect 37242 677076 37290 677104
rect 37242 677048 37260 677076
rect 37181 677046 37260 677048
rect 37181 677043 37247 677046
rect 45737 676698 45803 676701
rect 41492 676696 45803 676698
rect 41492 676640 45742 676696
rect 45798 676640 45803 676696
rect 41492 676638 45803 676640
rect 45737 676635 45803 676638
rect 62757 676154 62823 676157
rect 62757 676152 64492 676154
rect 62757 676096 62762 676152
rect 62818 676096 64492 676152
rect 62757 676094 64492 676096
rect 62757 676091 62823 676094
rect 40953 676018 41019 676021
rect 41454 676018 41460 676020
rect 40953 676016 41460 676018
rect 40953 675960 40958 676016
rect 41014 675960 41460 676016
rect 40953 675958 41460 675960
rect 40953 675955 41019 675958
rect 41454 675956 41460 675958
rect 41524 675956 41530 676020
rect 42006 673508 42012 673572
rect 42076 673570 42082 673572
rect 42517 673570 42583 673573
rect 42076 673568 42583 673570
rect 42076 673512 42522 673568
rect 42578 673512 42583 673568
rect 42076 673510 42583 673512
rect 42076 673508 42082 673510
rect 42517 673507 42583 673510
rect 40585 673162 40651 673165
rect 42333 673162 42399 673165
rect 40585 673160 42399 673162
rect 40585 673104 40590 673160
rect 40646 673104 42338 673160
rect 42394 673104 42399 673160
rect 40585 673102 42399 673104
rect 40585 673099 40651 673102
rect 42333 673099 42399 673102
rect 661677 673162 661743 673165
rect 676489 673162 676555 673165
rect 661677 673160 676555 673162
rect 661677 673104 661682 673160
rect 661738 673104 676494 673160
rect 676550 673104 676555 673160
rect 661677 673102 676555 673104
rect 661677 673099 661743 673102
rect 676489 673099 676555 673102
rect 39665 671938 39731 671941
rect 42333 671938 42399 671941
rect 39665 671936 42399 671938
rect 39665 671880 39670 671936
rect 39726 671880 42338 671936
rect 42394 671880 42399 671936
rect 39665 671878 42399 671880
rect 39665 671875 39731 671878
rect 42333 671875 42399 671878
rect 31017 671394 31083 671397
rect 41822 671394 41828 671396
rect 31017 671392 41828 671394
rect 31017 671336 31022 671392
rect 31078 671336 41828 671392
rect 31017 671334 41828 671336
rect 31017 671331 31083 671334
rect 41822 671332 41828 671334
rect 41892 671332 41898 671396
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 676489 671122 676555 671125
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 676446 671120 676555 671122
rect 676446 671064 676494 671120
rect 676550 671064 676555 671120
rect 667197 671059 667263 671062
rect 676446 671059 676555 671064
rect 40125 670986 40191 670989
rect 42149 670986 42215 670989
rect 40125 670984 42215 670986
rect 40125 670928 40130 670984
rect 40186 670928 42154 670984
rect 42210 670928 42215 670984
rect 676446 670956 676506 671059
rect 40125 670926 42215 670928
rect 40125 670923 40191 670926
rect 42149 670923 42215 670926
rect 668577 670578 668643 670581
rect 668577 670576 676292 670578
rect 668577 670520 668582 670576
rect 668638 670520 676292 670576
rect 668577 670518 676292 670520
rect 668577 670515 668643 670518
rect 651465 670442 651531 670445
rect 650164 670440 651531 670442
rect 650164 670384 651470 670440
rect 651526 670384 651531 670440
rect 650164 670382 651531 670384
rect 651465 670379 651531 670382
rect 671613 670306 671679 670309
rect 671613 670304 674850 670306
rect 671613 670248 671618 670304
rect 671674 670248 674850 670304
rect 671613 670246 674850 670248
rect 671613 670243 671679 670246
rect 671153 669898 671219 669901
rect 674790 669898 674850 670246
rect 675017 670170 675083 670173
rect 675017 670168 676292 670170
rect 675017 670112 675022 670168
rect 675078 670112 676292 670168
rect 675017 670110 676292 670112
rect 675017 670107 675083 670110
rect 671153 669896 674666 669898
rect 671153 669840 671158 669896
rect 671214 669840 674666 669896
rect 671153 669838 674666 669840
rect 674790 669838 676322 669898
rect 671153 669835 671219 669838
rect 672809 669490 672875 669493
rect 674606 669490 674666 669838
rect 676262 669732 676322 669838
rect 672809 669488 674482 669490
rect 672809 669432 672814 669488
rect 672870 669432 674482 669488
rect 672809 669430 674482 669432
rect 674606 669430 676322 669490
rect 672809 669427 672875 669430
rect 42190 669292 42196 669356
rect 42260 669354 42266 669356
rect 48957 669354 49023 669357
rect 42260 669352 49023 669354
rect 42260 669296 48962 669352
rect 49018 669296 49023 669352
rect 42260 669294 49023 669296
rect 42260 669292 42266 669294
rect 48957 669291 49023 669294
rect 674422 669218 674482 669430
rect 676262 669324 676322 669430
rect 675017 669218 675083 669221
rect 674422 669216 675083 669218
rect 674422 669160 675022 669216
rect 675078 669160 675083 669216
rect 674422 669158 675083 669160
rect 675017 669155 675083 669158
rect 671521 668674 671587 668677
rect 676262 668674 676322 668916
rect 671521 668672 676322 668674
rect 671521 668616 671526 668672
rect 671582 668616 676322 668672
rect 671521 668614 676322 668616
rect 671521 668611 671587 668614
rect 42057 668268 42123 668269
rect 42006 668204 42012 668268
rect 42076 668266 42123 668268
rect 670969 668266 671035 668269
rect 676262 668266 676322 668508
rect 42076 668264 42168 668266
rect 42118 668208 42168 668264
rect 42076 668206 42168 668208
rect 670969 668264 676322 668266
rect 670969 668208 670974 668264
rect 671030 668208 676322 668264
rect 670969 668206 676322 668208
rect 42076 668204 42123 668206
rect 42057 668203 42123 668204
rect 670969 668203 671035 668206
rect 671061 667994 671127 667997
rect 676262 667994 676322 668100
rect 671061 667992 676322 667994
rect 671061 667936 671066 667992
rect 671122 667936 676322 667992
rect 671061 667934 676322 667936
rect 671061 667931 671127 667934
rect 42241 667860 42307 667861
rect 42190 667796 42196 667860
rect 42260 667858 42307 667860
rect 42260 667856 42352 667858
rect 42302 667800 42352 667856
rect 42260 667798 42352 667800
rect 42260 667796 42307 667798
rect 42241 667795 42307 667796
rect 672533 667450 672599 667453
rect 676262 667450 676322 667692
rect 672533 667448 676322 667450
rect 672533 667392 672538 667448
rect 672594 667392 676322 667448
rect 672533 667390 676322 667392
rect 672533 667387 672599 667390
rect 42241 667042 42307 667045
rect 44725 667042 44791 667045
rect 676262 667042 676322 667284
rect 42241 667040 44791 667042
rect 42241 666984 42246 667040
rect 42302 666984 44730 667040
rect 44786 666984 44791 667040
rect 42241 666982 44791 666984
rect 42241 666979 42307 666982
rect 44725 666979 44791 666982
rect 674790 666982 676322 667042
rect 683205 667042 683271 667045
rect 683205 667040 683314 667042
rect 683205 666984 683210 667040
rect 683266 666984 683314 667040
rect 42057 666634 42123 666637
rect 42885 666634 42951 666637
rect 42057 666632 42951 666634
rect 42057 666576 42062 666632
rect 42118 666576 42890 666632
rect 42946 666576 42951 666632
rect 42057 666574 42951 666576
rect 42057 666571 42123 666574
rect 42885 666571 42951 666574
rect 672717 666634 672783 666637
rect 674790 666634 674850 666982
rect 683205 666979 683314 666984
rect 683254 666876 683314 666979
rect 672717 666632 674850 666634
rect 672717 666576 672722 666632
rect 672778 666576 674850 666632
rect 672717 666574 674850 666576
rect 672717 666571 672783 666574
rect 668761 666226 668827 666229
rect 674189 666226 674255 666229
rect 668761 666224 674255 666226
rect 668761 666168 668766 666224
rect 668822 666168 674194 666224
rect 674250 666168 674255 666224
rect 668761 666166 674255 666168
rect 668761 666163 668827 666166
rect 674189 666163 674255 666166
rect 674833 666226 674899 666229
rect 676262 666226 676322 666468
rect 674833 666224 676322 666226
rect 674833 666168 674838 666224
rect 674894 666168 676322 666224
rect 674833 666166 676322 666168
rect 674833 666163 674899 666166
rect 667841 665954 667907 665957
rect 676262 665954 676322 666060
rect 667841 665952 676322 665954
rect 667841 665896 667846 665952
rect 667902 665896 676322 665952
rect 667841 665894 676322 665896
rect 667841 665891 667907 665894
rect 671981 665682 672047 665685
rect 674833 665682 674899 665685
rect 671981 665680 674899 665682
rect 671981 665624 671986 665680
rect 672042 665624 674838 665680
rect 674894 665624 674899 665680
rect 671981 665622 674899 665624
rect 671981 665619 672047 665622
rect 674833 665619 674899 665622
rect 40902 665348 40908 665412
rect 40972 665410 40978 665412
rect 41781 665410 41847 665413
rect 40972 665408 41847 665410
rect 40972 665352 41786 665408
rect 41842 665352 41847 665408
rect 40972 665350 41847 665352
rect 40972 665348 40978 665350
rect 41781 665347 41847 665350
rect 666461 665410 666527 665413
rect 676262 665410 676322 665652
rect 666461 665408 676322 665410
rect 666461 665352 666466 665408
rect 666522 665352 676322 665408
rect 666461 665350 676322 665352
rect 666461 665347 666527 665350
rect 674189 665138 674255 665141
rect 676262 665138 676322 665244
rect 674189 665136 676322 665138
rect 674189 665080 674194 665136
rect 674250 665080 676322 665136
rect 674189 665078 676322 665080
rect 674189 665075 674255 665078
rect 674833 664730 674899 664733
rect 676262 664730 676322 664836
rect 674833 664728 676322 664730
rect 674833 664672 674838 664728
rect 674894 664672 676322 664728
rect 674833 664670 676322 664672
rect 674833 664667 674899 664670
rect 671470 664396 671476 664460
rect 671540 664458 671546 664460
rect 671540 664398 676292 664458
rect 671540 664396 671546 664398
rect 40718 664124 40724 664188
rect 40788 664186 40794 664188
rect 41781 664186 41847 664189
rect 40788 664184 41847 664186
rect 40788 664128 41786 664184
rect 41842 664128 41847 664184
rect 40788 664126 41847 664128
rect 40788 664124 40794 664126
rect 41781 664123 41847 664126
rect 669773 664186 669839 664189
rect 674833 664186 674899 664189
rect 669773 664184 674899 664186
rect 669773 664128 669778 664184
rect 669834 664128 674838 664184
rect 674894 664128 674899 664184
rect 669773 664126 674899 664128
rect 669773 664123 669839 664126
rect 674833 664123 674899 664126
rect 669221 663914 669287 663917
rect 676262 663914 676322 664020
rect 669221 663912 676322 663914
rect 669221 663856 669226 663912
rect 669282 663856 676322 663912
rect 669221 663854 676322 663856
rect 669221 663851 669287 663854
rect 683389 663778 683455 663781
rect 683389 663776 683498 663778
rect 683389 663720 683394 663776
rect 683450 663720 683498 663776
rect 683389 663715 683498 663720
rect 683438 663612 683498 663715
rect 42333 663372 42399 663373
rect 42333 663368 42380 663372
rect 42444 663370 42450 663372
rect 42333 663312 42338 663368
rect 42333 663308 42380 663312
rect 42444 663310 42490 663370
rect 42444 663308 42450 663310
rect 42333 663307 42399 663308
rect 62113 663098 62179 663101
rect 674833 663098 674899 663101
rect 676262 663098 676322 663204
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 674833 663096 676322 663098
rect 674833 663040 674838 663096
rect 674894 663040 676322 663096
rect 674833 663038 676322 663040
rect 62113 663035 62179 663038
rect 674833 663035 674899 663038
rect 42425 662962 42491 662965
rect 44541 662962 44607 662965
rect 42425 662960 44607 662962
rect 42425 662904 42430 662960
rect 42486 662904 44546 662960
rect 44602 662904 44607 662960
rect 42425 662902 44607 662904
rect 42425 662899 42491 662902
rect 44541 662899 44607 662902
rect 42057 662826 42123 662829
rect 41370 662824 42123 662826
rect 41370 662768 42062 662824
rect 42118 662768 42123 662824
rect 41370 662766 42123 662768
rect 40534 662628 40540 662692
rect 40604 662690 40610 662692
rect 41370 662690 41430 662766
rect 42057 662763 42123 662766
rect 672349 662826 672415 662829
rect 672349 662824 676292 662826
rect 672349 662768 672354 662824
rect 672410 662768 676292 662824
rect 672349 662766 676292 662768
rect 672349 662763 672415 662766
rect 40604 662630 41430 662690
rect 40604 662628 40610 662630
rect 669037 662554 669103 662557
rect 674833 662554 674899 662557
rect 669037 662552 674899 662554
rect 669037 662496 669042 662552
rect 669098 662496 674838 662552
rect 674894 662496 674899 662552
rect 669037 662494 674899 662496
rect 669037 662491 669103 662494
rect 674833 662491 674899 662494
rect 674414 662220 674420 662284
rect 674484 662282 674490 662284
rect 676262 662282 676322 662388
rect 674484 662222 676322 662282
rect 674484 662220 674490 662222
rect 674833 661874 674899 661877
rect 676262 661874 676322 661980
rect 674833 661872 676322 661874
rect 674833 661816 674838 661872
rect 674894 661816 676322 661872
rect 674833 661814 676322 661816
rect 674833 661811 674899 661814
rect 673085 661602 673151 661605
rect 673085 661600 676292 661602
rect 673085 661544 673090 661600
rect 673146 661544 676292 661600
rect 673085 661542 676292 661544
rect 673085 661539 673151 661542
rect 671245 661330 671311 661333
rect 674833 661330 674899 661333
rect 671245 661328 674899 661330
rect 671245 661272 671250 661328
rect 671306 661272 674838 661328
rect 674894 661272 674899 661328
rect 671245 661270 674899 661272
rect 671245 661267 671311 661270
rect 674833 661267 674899 661270
rect 671981 661058 672047 661061
rect 676262 661058 676322 661164
rect 671981 661056 676322 661058
rect 671981 661000 671986 661056
rect 672042 661000 676322 661056
rect 671981 660998 676322 661000
rect 671981 660995 672047 660998
rect 670601 660106 670667 660109
rect 676262 660106 676322 660756
rect 670601 660104 676322 660106
rect 670601 660048 670606 660104
rect 670662 660048 676322 660104
rect 670601 660046 676322 660048
rect 670601 660043 670667 660046
rect 42149 659834 42215 659837
rect 42374 659834 42380 659836
rect 42149 659832 42380 659834
rect 42149 659776 42154 659832
rect 42210 659776 42380 659832
rect 42149 659774 42380 659776
rect 42149 659771 42215 659774
rect 42374 659772 42380 659774
rect 42444 659772 42450 659836
rect 670601 659698 670667 659701
rect 676262 659698 676322 659940
rect 670601 659696 676322 659698
rect 670601 659640 670606 659696
rect 670662 659640 676322 659696
rect 670601 659638 676322 659640
rect 670601 659635 670667 659638
rect 42149 659018 42215 659021
rect 42701 659018 42767 659021
rect 42149 659016 42767 659018
rect 42149 658960 42154 659016
rect 42210 658960 42706 659016
rect 42762 658960 42767 659016
rect 42149 658958 42767 658960
rect 42149 658955 42215 658958
rect 42701 658955 42767 658958
rect 41454 658548 41460 658612
rect 41524 658610 41530 658612
rect 42609 658610 42675 658613
rect 41524 658608 42675 658610
rect 41524 658552 42614 658608
rect 42670 658552 42675 658608
rect 41524 658550 42675 658552
rect 41524 658548 41530 658550
rect 42609 658547 42675 658550
rect 41822 658276 41828 658340
rect 41892 658338 41898 658340
rect 42425 658338 42491 658341
rect 41892 658336 42491 658338
rect 41892 658280 42430 658336
rect 42486 658280 42491 658336
rect 41892 658278 42491 658280
rect 41892 658276 41898 658278
rect 42425 658275 42491 658278
rect 41638 657324 41644 657388
rect 41708 657386 41714 657388
rect 41965 657386 42031 657389
rect 41708 657384 42031 657386
rect 41708 657328 41970 657384
rect 42026 657328 42031 657384
rect 41708 657326 42031 657328
rect 41708 657324 41714 657326
rect 41965 657323 42031 657326
rect 651465 657114 651531 657117
rect 650164 657112 651531 657114
rect 650164 657056 651470 657112
rect 651526 657056 651531 657112
rect 650164 657054 651531 657056
rect 651465 657051 651531 657054
rect 62757 656162 62823 656165
rect 42566 656160 62823 656162
rect 42566 656104 62762 656160
rect 62818 656104 62823 656160
rect 42566 656102 62823 656104
rect 42566 655485 42626 656102
rect 62757 656099 62823 656102
rect 42566 655480 42675 655485
rect 42566 655424 42614 655480
rect 42670 655424 42675 655480
rect 42566 655422 42675 655424
rect 42609 655419 42675 655422
rect 669221 654258 669287 654261
rect 675385 654258 675451 654261
rect 669221 654256 675451 654258
rect 669221 654200 669226 654256
rect 669282 654200 675390 654256
rect 675446 654200 675451 654256
rect 669221 654198 675451 654200
rect 669221 654195 669287 654198
rect 675385 654195 675451 654198
rect 675334 652836 675340 652900
rect 675404 652898 675410 652900
rect 675569 652898 675635 652901
rect 675404 652896 675635 652898
rect 675404 652840 675574 652896
rect 675630 652840 675635 652896
rect 675404 652838 675635 652840
rect 675404 652836 675410 652838
rect 675569 652835 675635 652838
rect 675569 651540 675635 651541
rect 675518 651538 675524 651540
rect 675478 651478 675524 651538
rect 675588 651536 675635 651540
rect 675630 651480 675635 651536
rect 675518 651476 675524 651478
rect 675588 651476 675635 651480
rect 675569 651475 675635 651476
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674230 648892 674236 648956
rect 674300 648954 674306 648956
rect 675477 648954 675543 648957
rect 674300 648952 675543 648954
rect 674300 648896 675482 648952
rect 675538 648896 675543 648952
rect 674300 648894 675543 648896
rect 674300 648892 674306 648894
rect 675477 648891 675543 648894
rect 672993 648682 673059 648685
rect 675477 648682 675543 648685
rect 672993 648680 675543 648682
rect 672993 648624 672998 648680
rect 673054 648624 675482 648680
rect 675538 648624 675543 648680
rect 672993 648622 675543 648624
rect 672993 648619 673059 648622
rect 675477 648619 675543 648622
rect 672533 647866 672599 647869
rect 675477 647866 675543 647869
rect 672533 647864 675543 647866
rect 672533 647808 672538 647864
rect 672594 647808 675482 647864
rect 675538 647808 675543 647864
rect 672533 647806 675543 647808
rect 672533 647803 672599 647806
rect 675477 647803 675543 647806
rect 670877 647322 670943 647325
rect 675293 647322 675359 647325
rect 670877 647320 675359 647322
rect 670877 647264 670882 647320
rect 670938 647264 675298 647320
rect 675354 647264 675359 647320
rect 670877 647262 675359 647264
rect 670877 647259 670943 647262
rect 675293 647259 675359 647262
rect 674787 645826 674853 645829
rect 674966 645826 674972 645828
rect 674787 645824 674972 645826
rect 674787 645768 674792 645824
rect 674848 645768 674972 645824
rect 674787 645766 674972 645768
rect 674787 645763 674853 645766
rect 674966 645764 674972 645766
rect 675036 645764 675042 645828
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 673545 644874 673611 644877
rect 675477 644874 675543 644877
rect 673545 644872 675543 644874
rect 673545 644816 673550 644872
rect 673606 644816 675482 644872
rect 675538 644816 675543 644872
rect 673545 644814 675543 644816
rect 673545 644811 673611 644814
rect 675477 644811 675543 644814
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 35758 644504 35818 644675
rect 675753 644330 675819 644333
rect 676806 644330 676812 644332
rect 675753 644328 676812 644330
rect 675753 644272 675758 644328
rect 675814 644272 676812 644328
rect 675753 644270 676812 644272
rect 675753 644267 675819 644270
rect 676806 644268 676812 644270
rect 676876 644268 676882 644332
rect 41462 643922 41522 644096
rect 673177 644058 673243 644061
rect 675477 644058 675543 644061
rect 673177 644056 675543 644058
rect 673177 644000 673182 644056
rect 673238 644000 675482 644056
rect 675538 644000 675543 644056
rect 673177 643998 675543 644000
rect 673177 643995 673243 643998
rect 675477 643995 675543 643998
rect 41462 643862 45570 643922
rect 41462 643650 41522 643688
rect 44357 643650 44423 643653
rect 41462 643648 44423 643650
rect 41462 643592 44362 643648
rect 44418 643592 44423 643648
rect 41462 643590 44423 643592
rect 44357 643587 44423 643590
rect 44817 643378 44883 643381
rect 41462 643376 44883 643378
rect 41462 643320 44822 643376
rect 44878 643320 44883 643376
rect 41462 643318 44883 643320
rect 41462 643280 41522 643318
rect 44817 643315 44883 643318
rect 45510 643242 45570 643862
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 661677 643786 661743 643789
rect 661677 643784 663810 643786
rect 661677 643728 661682 643784
rect 661738 643728 663810 643784
rect 661677 643726 663810 643728
rect 661677 643723 661743 643726
rect 663750 643514 663810 643726
rect 675293 643514 675359 643517
rect 663750 643512 675359 643514
rect 663750 643456 675298 643512
rect 675354 643456 675359 643512
rect 663750 643454 675359 643456
rect 675293 643451 675359 643454
rect 55857 643242 55923 643245
rect 45510 643240 55923 643242
rect 45510 643184 55862 643240
rect 55918 643184 55923 643240
rect 45510 643182 55923 643184
rect 55857 643179 55923 643182
rect 667841 643242 667907 643245
rect 675150 643242 675156 643244
rect 667841 643240 675156 643242
rect 667841 643184 667846 643240
rect 667902 643184 675156 643240
rect 667841 643182 675156 643184
rect 667841 643179 667907 643182
rect 675150 643180 675156 643182
rect 675220 643180 675226 643244
rect 45185 643106 45251 643109
rect 41462 643104 45251 643106
rect 41462 643048 45190 643104
rect 45246 643048 45251 643104
rect 41462 643046 45251 643048
rect 41462 642872 41522 643046
rect 45185 643043 45251 643046
rect 44633 642562 44699 642565
rect 41462 642560 44699 642562
rect 41462 642504 44638 642560
rect 44694 642504 44699 642560
rect 41462 642502 44699 642504
rect 41462 642464 41522 642502
rect 44633 642499 44699 642502
rect 674189 642426 674255 642429
rect 674414 642426 674420 642428
rect 674189 642424 674420 642426
rect 674189 642368 674194 642424
rect 674250 642368 674420 642424
rect 674189 642366 674420 642368
rect 674189 642363 674255 642366
rect 674414 642364 674420 642366
rect 674484 642364 674490 642428
rect 44173 642290 44239 642293
rect 41462 642288 44239 642290
rect 41462 642232 44178 642288
rect 44234 642232 44239 642288
rect 41462 642230 44239 642232
rect 41462 642056 41522 642230
rect 44173 642227 44239 642230
rect 674189 641746 674255 641749
rect 675293 641746 675359 641749
rect 674189 641744 675359 641746
rect 674189 641688 674194 641744
rect 674250 641688 675298 641744
rect 675354 641688 675359 641744
rect 674189 641686 675359 641688
rect 674189 641683 674255 641686
rect 675293 641683 675359 641686
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 45001 641474 45067 641477
rect 41462 641472 45067 641474
rect 41462 641416 45006 641472
rect 45062 641416 45067 641472
rect 41462 641414 45067 641416
rect 41462 641240 41522 641414
rect 45001 641411 45067 641414
rect 675201 641340 675267 641341
rect 675150 641338 675156 641340
rect 675110 641278 675156 641338
rect 675220 641336 675267 641340
rect 675262 641280 675267 641336
rect 675150 641276 675156 641278
rect 675220 641276 675267 641280
rect 675201 641275 675267 641276
rect 41781 641202 41847 641205
rect 45369 641202 45435 641205
rect 41781 641200 45435 641202
rect 41781 641144 41786 641200
rect 41842 641144 45374 641200
rect 45430 641144 45435 641200
rect 41781 641142 45435 641144
rect 41781 641139 41847 641142
rect 45369 641139 45435 641142
rect 45185 640930 45251 640933
rect 41462 640928 45251 640930
rect 41462 640872 45190 640928
rect 45246 640872 45251 640928
rect 41462 640870 45251 640872
rect 41462 640832 41522 640870
rect 45185 640867 45251 640870
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 35390 639845 35450 640016
rect 35341 639840 35450 639845
rect 35341 639784 35346 639840
rect 35402 639784 35450 639840
rect 35341 639782 35450 639784
rect 35341 639779 35407 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 675293 639434 675359 639437
rect 675518 639434 675524 639436
rect 675293 639432 675524 639434
rect 675293 639376 675298 639432
rect 675354 639376 675524 639432
rect 675293 639374 675524 639376
rect 675293 639371 675359 639374
rect 675518 639372 675524 639374
rect 675588 639372 675594 639436
rect 35758 639200 35818 639371
rect 35758 638621 35818 638792
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 40033 638618 40099 638621
rect 41638 638618 41644 638620
rect 40033 638616 41644 638618
rect 40033 638560 40038 638616
rect 40094 638560 41644 638616
rect 40033 638558 41644 638560
rect 40033 638555 40099 638558
rect 41638 638556 41644 638558
rect 41708 638556 41714 638620
rect 669773 638618 669839 638621
rect 675477 638618 675543 638621
rect 669773 638616 675543 638618
rect 669773 638560 669778 638616
rect 669834 638560 675482 638616
rect 675538 638560 675543 638616
rect 669773 638558 675543 638560
rect 669773 638555 669839 638558
rect 675477 638555 675543 638558
rect 33734 638213 33794 638384
rect 33734 638208 33843 638213
rect 33734 638152 33782 638208
rect 33838 638152 33843 638208
rect 33734 638150 33843 638152
rect 33777 638147 33843 638150
rect 41781 638210 41847 638213
rect 47393 638210 47459 638213
rect 41781 638208 47459 638210
rect 41781 638152 41786 638208
rect 41842 638152 47398 638208
rect 47454 638152 47459 638208
rect 41781 638150 47459 638152
rect 41781 638147 41847 638150
rect 47393 638147 47459 638150
rect 41462 637802 41522 637976
rect 675334 637876 675340 637940
rect 675404 637938 675410 637940
rect 675569 637938 675635 637941
rect 675404 637936 675635 637938
rect 675404 637880 675574 637936
rect 675630 637880 675635 637936
rect 675404 637878 675635 637880
rect 675404 637876 675410 637878
rect 675569 637875 675635 637878
rect 45921 637802 45987 637805
rect 41462 637800 45987 637802
rect 41462 637744 45926 637800
rect 45982 637744 45987 637800
rect 41462 637742 45987 637744
rect 45921 637739 45987 637742
rect 674414 637740 674420 637804
rect 674484 637802 674490 637804
rect 674741 637802 674807 637805
rect 674484 637800 674807 637802
rect 674484 637744 674746 637800
rect 674802 637744 674807 637800
rect 674484 637742 674807 637744
rect 674484 637740 674490 637742
rect 674741 637739 674807 637742
rect 674966 637604 674972 637668
rect 675036 637666 675042 637668
rect 682377 637666 682443 637669
rect 675036 637664 682443 637666
rect 675036 637608 682382 637664
rect 682438 637608 682443 637664
rect 675036 637606 682443 637608
rect 675036 637604 675042 637606
rect 682377 637603 682443 637606
rect 41781 637598 41847 637601
rect 41492 637596 41847 637598
rect 41492 637540 41786 637596
rect 41842 637540 41847 637596
rect 41492 637538 41847 637540
rect 41781 637535 41847 637538
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 46289 636986 46355 636989
rect 41462 636984 46355 636986
rect 41462 636928 46294 636984
rect 46350 636928 46355 636984
rect 41462 636926 46355 636928
rect 46289 636923 46355 636926
rect 673821 636850 673887 636853
rect 683389 636850 683455 636853
rect 673821 636848 683455 636850
rect 673821 636792 673826 636848
rect 673882 636792 683394 636848
rect 683450 636792 683455 636848
rect 673821 636790 683455 636792
rect 673821 636787 673887 636790
rect 683389 636787 683455 636790
rect 41462 636578 41522 636752
rect 44265 636578 44331 636581
rect 41462 636576 44331 636578
rect 41462 636520 44270 636576
rect 44326 636520 44331 636576
rect 41462 636518 44331 636520
rect 44265 636515 44331 636518
rect 41462 636306 41522 636344
rect 42885 636306 42951 636309
rect 41462 636304 42951 636306
rect 41462 636248 42890 636304
rect 42946 636248 42951 636304
rect 41462 636246 42951 636248
rect 42885 636243 42951 636246
rect 674925 636036 674991 636037
rect 674925 636034 674972 636036
rect 674880 636032 674972 636034
rect 674880 635976 674930 636032
rect 674880 635974 674972 635976
rect 674925 635972 674972 635974
rect 675036 635972 675042 636036
rect 674925 635971 674991 635972
rect 41462 635762 41522 635936
rect 44449 635762 44515 635765
rect 41462 635760 44515 635762
rect 41462 635704 44454 635760
rect 44510 635704 44515 635760
rect 41462 635702 44515 635704
rect 44449 635699 44515 635702
rect 674925 635762 674991 635765
rect 683757 635762 683823 635765
rect 674925 635760 683823 635762
rect 674925 635704 674930 635760
rect 674986 635704 683762 635760
rect 683818 635704 683823 635760
rect 674925 635702 683823 635704
rect 674925 635699 674991 635702
rect 683757 635699 683823 635702
rect 41462 635354 41522 635528
rect 672717 635490 672783 635493
rect 683205 635490 683271 635493
rect 672717 635488 683271 635490
rect 672717 635432 672722 635488
rect 672778 635432 683210 635488
rect 683266 635432 683271 635488
rect 672717 635430 683271 635432
rect 672717 635427 672783 635430
rect 683205 635427 683271 635430
rect 45001 635354 45067 635357
rect 41462 635352 45067 635354
rect 41462 635296 45006 635352
rect 45062 635296 45067 635352
rect 41462 635294 45067 635296
rect 45001 635291 45067 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 40542 634540 40602 634712
rect 40534 634476 40540 634540
rect 40604 634476 40610 634540
rect 41462 633858 41522 634304
rect 42517 633858 42583 633861
rect 41462 633856 42583 633858
rect 41462 633800 42522 633856
rect 42578 633800 42583 633856
rect 41462 633798 42583 633800
rect 42517 633795 42583 633798
rect 41462 633450 41522 633488
rect 43345 633450 43411 633453
rect 41462 633448 43411 633450
rect 41462 633392 43350 633448
rect 43406 633392 43411 633448
rect 41462 633390 43411 633392
rect 43345 633387 43411 633390
rect 674833 631410 674899 631413
rect 675201 631410 675267 631413
rect 674833 631408 675267 631410
rect 674833 631352 674838 631408
rect 674894 631352 675206 631408
rect 675262 631352 675267 631408
rect 674833 631350 675267 631352
rect 674833 631347 674899 631350
rect 675201 631347 675267 631350
rect 675569 631410 675635 631413
rect 676070 631410 676076 631412
rect 675569 631408 676076 631410
rect 675569 631352 675574 631408
rect 675630 631352 676076 631408
rect 675569 631350 676076 631352
rect 675569 631347 675635 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 36537 630730 36603 630733
rect 41822 630730 41828 630732
rect 36537 630728 41828 630730
rect 36537 630672 36542 630728
rect 36598 630672 41828 630728
rect 36537 630670 41828 630672
rect 36537 630667 36603 630670
rect 41822 630668 41828 630670
rect 41892 630668 41898 630732
rect 651557 630594 651623 630597
rect 650164 630592 651623 630594
rect 650164 630536 651562 630592
rect 651618 630536 651623 630592
rect 650164 630534 651623 630536
rect 651557 630531 651623 630534
rect 41413 630050 41479 630053
rect 42701 630050 42767 630053
rect 41413 630048 42767 630050
rect 41413 629992 41418 630048
rect 41474 629992 42706 630048
rect 42762 629992 42767 630048
rect 41413 629990 42767 629992
rect 41413 629987 41479 629990
rect 42701 629987 42767 629990
rect 675150 629716 675156 629780
rect 675220 629778 675226 629780
rect 675385 629778 675451 629781
rect 675220 629776 675451 629778
rect 675220 629720 675390 629776
rect 675446 629720 675451 629776
rect 675220 629718 675451 629720
rect 675220 629716 675226 629718
rect 675385 629715 675451 629718
rect 674966 629444 674972 629508
rect 675036 629506 675042 629508
rect 675201 629506 675267 629509
rect 675036 629504 675267 629506
rect 675036 629448 675206 629504
rect 675262 629448 675267 629504
rect 675036 629446 675267 629448
rect 675036 629444 675042 629446
rect 675201 629443 675267 629446
rect 652017 628554 652083 628557
rect 676489 628554 676555 628557
rect 652017 628552 676555 628554
rect 652017 628496 652022 628552
rect 652078 628496 676494 628552
rect 676550 628496 676555 628552
rect 652017 628494 676555 628496
rect 652017 628491 652083 628494
rect 676489 628491 676555 628494
rect 46473 626650 46539 626653
rect 50337 626650 50403 626653
rect 46473 626648 50403 626650
rect 46473 626592 46478 626648
rect 46534 626592 50342 626648
rect 50398 626592 50403 626648
rect 46473 626590 50403 626592
rect 46473 626587 46539 626590
rect 50337 626587 50403 626590
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 42057 625834 42123 625837
rect 42517 625834 42583 625837
rect 42057 625832 42583 625834
rect 42057 625776 42062 625832
rect 42118 625776 42522 625832
rect 42578 625776 42583 625832
rect 42057 625774 42583 625776
rect 42057 625771 42123 625774
rect 42517 625771 42583 625774
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 669270 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 671613 625154 671679 625157
rect 671613 625152 676292 625154
rect 671613 625096 671618 625152
rect 671674 625096 676292 625152
rect 671613 625094 676292 625096
rect 671613 625091 671679 625094
rect 671613 624746 671679 624749
rect 671613 624744 676292 624746
rect 671613 624688 671618 624744
rect 671674 624688 676292 624744
rect 671613 624686 676292 624688
rect 671613 624683 671679 624686
rect 671429 624338 671495 624341
rect 671429 624336 676292 624338
rect 671429 624280 671434 624336
rect 671490 624280 676292 624336
rect 671429 624278 676292 624280
rect 671429 624275 671495 624278
rect 42425 624202 42491 624205
rect 46473 624202 46539 624205
rect 42425 624200 46539 624202
rect 42425 624144 42430 624200
rect 42486 624144 46478 624200
rect 46534 624144 46539 624200
rect 42425 624142 46539 624144
rect 42425 624139 42491 624142
rect 46473 624139 46539 624142
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 671245 623930 671311 623933
rect 671245 623928 676292 623930
rect 671245 623872 671250 623928
rect 671306 623872 676292 623928
rect 671245 623870 676292 623872
rect 671245 623867 671311 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42241 623794 42307 623797
rect 40788 623792 42307 623794
rect 40788 623736 42246 623792
rect 42302 623736 42307 623792
rect 40788 623734 42307 623736
rect 40788 623732 40794 623734
rect 42241 623731 42307 623734
rect 42425 623794 42491 623797
rect 42793 623794 42859 623797
rect 42425 623792 42859 623794
rect 42425 623736 42430 623792
rect 42486 623736 42798 623792
rect 42854 623736 42859 623792
rect 42425 623734 42859 623736
rect 42425 623731 42491 623734
rect 42793 623731 42859 623734
rect 671061 623522 671127 623525
rect 671061 623520 676292 623522
rect 671061 623464 671066 623520
rect 671122 623464 676292 623520
rect 671061 623462 676292 623464
rect 671061 623459 671127 623462
rect 42057 623386 42123 623389
rect 44265 623386 44331 623389
rect 42057 623384 44331 623386
rect 42057 623328 42062 623384
rect 42118 623328 44270 623384
rect 44326 623328 44331 623384
rect 42057 623326 44331 623328
rect 42057 623323 42123 623326
rect 44265 623323 44331 623326
rect 671429 623114 671495 623117
rect 671429 623112 676292 623114
rect 671429 623056 671434 623112
rect 671490 623056 676292 623112
rect 671429 623054 676292 623056
rect 671429 623051 671495 623054
rect 683205 622842 683271 622845
rect 683205 622840 683314 622842
rect 683205 622784 683210 622840
rect 683266 622784 683314 622840
rect 683205 622779 683314 622784
rect 683254 622676 683314 622779
rect 671061 622298 671127 622301
rect 671061 622296 676292 622298
rect 671061 622240 671066 622296
rect 671122 622240 676292 622296
rect 671061 622238 676292 622240
rect 671061 622235 671127 622238
rect 682377 622026 682443 622029
rect 682334 622024 682443 622026
rect 682334 621968 682382 622024
rect 682438 621968 682443 622024
rect 682334 621963 682443 621968
rect 682334 621860 682394 621963
rect 669589 621618 669655 621621
rect 676489 621618 676555 621621
rect 669589 621616 676555 621618
rect 669589 621560 669594 621616
rect 669650 621560 676494 621616
rect 676550 621560 676555 621616
rect 669589 621558 676555 621560
rect 669589 621555 669655 621558
rect 676489 621555 676555 621558
rect 667657 621210 667723 621213
rect 676262 621210 676322 621452
rect 676489 621210 676555 621213
rect 667657 621208 676322 621210
rect 667657 621152 667662 621208
rect 667718 621152 676322 621208
rect 667657 621150 676322 621152
rect 676446 621208 676555 621210
rect 676446 621152 676494 621208
rect 676550 621152 676555 621208
rect 667657 621147 667723 621150
rect 676446 621147 676555 621152
rect 676446 621044 676506 621147
rect 42057 620938 42123 620941
rect 45001 620938 45067 620941
rect 42057 620936 45067 620938
rect 42057 620880 42062 620936
rect 42118 620880 45006 620936
rect 45062 620880 45067 620936
rect 42057 620878 45067 620880
rect 42057 620875 42123 620878
rect 45001 620875 45067 620878
rect 670417 620666 670483 620669
rect 670417 620664 676292 620666
rect 670417 620608 670422 620664
rect 670478 620608 676292 620664
rect 670417 620606 676292 620608
rect 670417 620603 670483 620606
rect 670141 620394 670207 620397
rect 676489 620394 676555 620397
rect 670141 620392 676555 620394
rect 670141 620336 670146 620392
rect 670202 620336 676494 620392
rect 676550 620336 676555 620392
rect 670141 620334 676555 620336
rect 670141 620331 670207 620334
rect 676489 620331 676555 620334
rect 42241 620122 42307 620125
rect 44449 620122 44515 620125
rect 42241 620120 44515 620122
rect 42241 620064 42246 620120
rect 42302 620064 44454 620120
rect 44510 620064 44515 620120
rect 42241 620062 44515 620064
rect 42241 620059 42307 620062
rect 44449 620059 44515 620062
rect 668393 619986 668459 619989
rect 676262 619986 676322 620228
rect 676489 619986 676555 619989
rect 668393 619984 676322 619986
rect 668393 619928 668398 619984
rect 668454 619928 676322 619984
rect 668393 619926 676322 619928
rect 676446 619984 676555 619986
rect 676446 619928 676494 619984
rect 676550 619928 676555 619984
rect 668393 619923 668459 619926
rect 676446 619923 676555 619928
rect 40534 619788 40540 619852
rect 40604 619850 40610 619852
rect 42701 619850 42767 619853
rect 40604 619848 42767 619850
rect 40604 619792 42706 619848
rect 42762 619792 42767 619848
rect 676446 619820 676506 619923
rect 40604 619790 42767 619792
rect 40604 619788 40610 619790
rect 42701 619787 42767 619790
rect 42517 619578 42583 619581
rect 46289 619578 46355 619581
rect 42517 619576 46355 619578
rect 42517 619520 42522 619576
rect 42578 619520 46294 619576
rect 46350 619520 46355 619576
rect 42517 619518 46355 619520
rect 42517 619515 42583 619518
rect 46289 619515 46355 619518
rect 674649 619578 674715 619581
rect 677225 619578 677291 619581
rect 674649 619576 677291 619578
rect 674649 619520 674654 619576
rect 674710 619520 677230 619576
rect 677286 619520 677291 619576
rect 674649 619518 677291 619520
rect 674649 619515 674715 619518
rect 677225 619515 677291 619518
rect 674005 619170 674071 619173
rect 676446 619170 676506 619412
rect 674005 619168 676506 619170
rect 674005 619112 674010 619168
rect 674066 619112 676506 619168
rect 674005 619110 676506 619112
rect 674005 619107 674071 619110
rect 676990 619108 676996 619172
rect 677060 619108 677066 619172
rect 677225 619170 677291 619173
rect 683113 619170 683179 619173
rect 677225 619168 683179 619170
rect 677225 619112 677230 619168
rect 677286 619112 683118 619168
rect 683174 619112 683179 619168
rect 677225 619110 683179 619112
rect 676998 619004 677058 619108
rect 677225 619107 677291 619110
rect 683113 619107 683179 619110
rect 42517 618762 42583 618765
rect 47393 618762 47459 618765
rect 42517 618760 47459 618762
rect 42517 618704 42522 618760
rect 42578 618704 47398 618760
rect 47454 618704 47459 618760
rect 42517 618702 47459 618704
rect 42517 618699 42583 618702
rect 47393 618699 47459 618702
rect 683757 618762 683823 618765
rect 683757 618760 683866 618762
rect 683757 618704 683762 618760
rect 683818 618704 683866 618760
rect 683757 618699 683866 618704
rect 683806 618596 683866 618699
rect 671797 618218 671863 618221
rect 671797 618216 676292 618218
rect 671797 618160 671802 618216
rect 671858 618160 676292 618216
rect 671797 618158 676292 618160
rect 671797 618155 671863 618158
rect 674465 617810 674531 617813
rect 674465 617808 676292 617810
rect 674465 617752 674470 617808
rect 674526 617752 676292 617808
rect 674465 617750 676292 617752
rect 674465 617747 674531 617750
rect 683113 617538 683179 617541
rect 682886 617536 683179 617538
rect 682886 617480 683118 617536
rect 683174 617480 683179 617536
rect 682886 617478 683179 617480
rect 682886 617372 682946 617478
rect 683113 617475 683179 617478
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683389 617130 683455 617133
rect 683389 617128 683498 617130
rect 683389 617072 683394 617128
rect 683450 617072 683498 617128
rect 683389 617067 683498 617072
rect 683438 616964 683498 617067
rect 672165 616586 672231 616589
rect 672165 616584 676292 616586
rect 672165 616528 672170 616584
rect 672226 616528 676292 616584
rect 672165 616526 676292 616528
rect 672165 616523 672231 616526
rect 670417 616178 670483 616181
rect 670417 616176 676292 616178
rect 670417 616120 670422 616176
rect 670478 616120 676292 616176
rect 670417 616118 676292 616120
rect 670417 616115 670483 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 42425 616042 42491 616045
rect 41524 616040 42491 616042
rect 41524 615984 42430 616040
rect 42486 615984 42491 616040
rect 41524 615982 42491 615984
rect 41524 615980 41530 615982
rect 42425 615979 42491 615982
rect 41454 615708 41460 615772
rect 41524 615770 41530 615772
rect 41781 615770 41847 615773
rect 41524 615768 41847 615770
rect 41524 615712 41786 615768
rect 41842 615712 41847 615768
rect 41524 615710 41847 615712
rect 41524 615708 41530 615710
rect 41781 615707 41847 615710
rect 669270 615740 676660 615770
rect 669270 615710 676690 615740
rect 668209 615634 668275 615637
rect 669270 615634 669330 615710
rect 668209 615632 669330 615634
rect 668209 615576 668214 615632
rect 668270 615576 669330 615632
rect 668209 615574 669330 615576
rect 668209 615571 668275 615574
rect 676630 615332 676690 615710
rect 669589 614954 669655 614957
rect 669589 614952 676292 614954
rect 669589 614896 669594 614952
rect 669650 614896 676292 614952
rect 669589 614894 676292 614896
rect 669589 614891 669655 614894
rect 42149 613594 42215 613597
rect 45921 613594 45987 613597
rect 42149 613592 45987 613594
rect 42149 613536 42154 613592
rect 42210 613536 45926 613592
rect 45982 613536 45987 613592
rect 42149 613534 45987 613536
rect 42149 613531 42215 613534
rect 45921 613531 45987 613534
rect 41781 612780 41847 612781
rect 41781 612776 41828 612780
rect 41892 612778 41898 612780
rect 41781 612720 41786 612776
rect 41781 612716 41828 612720
rect 41892 612718 41938 612778
rect 41892 612716 41898 612718
rect 41781 612715 41847 612716
rect 43069 612370 43135 612373
rect 43713 612370 43779 612373
rect 43069 612368 43779 612370
rect 43069 612312 43074 612368
rect 43130 612312 43718 612368
rect 43774 612312 43779 612368
rect 43069 612310 43779 612312
rect 43069 612307 43135 612310
rect 43713 612307 43779 612310
rect 43345 611010 43411 611013
rect 44081 611010 44147 611013
rect 43345 611008 44147 611010
rect 43345 610952 43350 611008
rect 43406 610952 44086 611008
rect 44142 610952 44147 611008
rect 43345 610950 44147 610952
rect 43345 610947 43411 610950
rect 44081 610947 44147 610950
rect 44265 611010 44331 611013
rect 47209 611010 47275 611013
rect 44265 611008 47275 611010
rect 44265 610952 44270 611008
rect 44326 610952 47214 611008
rect 47270 610952 47275 611008
rect 44265 610950 47275 610952
rect 44265 610947 44331 610950
rect 47209 610947 47275 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 672625 608698 672691 608701
rect 674833 608698 674899 608701
rect 672625 608696 674899 608698
rect 672625 608640 672630 608696
rect 672686 608640 674838 608696
rect 674894 608640 674899 608696
rect 672625 608638 674899 608640
rect 672625 608635 672691 608638
rect 674833 608635 674899 608638
rect 675477 607884 675543 607885
rect 675477 607880 675524 607884
rect 675588 607882 675594 607884
rect 675477 607824 675482 607880
rect 675477 607820 675524 607824
rect 675588 607822 675634 607882
rect 675588 607820 675594 607822
rect 675477 607819 675543 607820
rect 672257 607338 672323 607341
rect 675293 607338 675359 607341
rect 672257 607336 675359 607338
rect 672257 607280 672262 607336
rect 672318 607280 675298 607336
rect 675354 607280 675359 607336
rect 672257 607278 675359 607280
rect 672257 607275 672323 607278
rect 675293 607275 675359 607278
rect 674833 607066 674899 607069
rect 675293 607066 675359 607069
rect 674833 607064 675359 607066
rect 674833 607008 674838 607064
rect 674894 607008 675298 607064
rect 675354 607008 675359 607064
rect 674833 607006 675359 607008
rect 674833 607003 674899 607006
rect 675293 607003 675359 607006
rect 674465 604618 674531 604621
rect 675293 604618 675359 604621
rect 674465 604616 675359 604618
rect 674465 604560 674470 604616
rect 674526 604560 675298 604616
rect 675354 604560 675359 604616
rect 674465 604558 675359 604560
rect 674465 604555 674531 604558
rect 675293 604555 675359 604558
rect 668761 604346 668827 604349
rect 675293 604346 675359 604349
rect 668761 604344 675359 604346
rect 668761 604288 668766 604344
rect 668822 604288 675298 604344
rect 675354 604288 675359 604344
rect 668761 604286 675359 604288
rect 668761 604283 668827 604286
rect 675293 604283 675359 604286
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 673913 603530 673979 603533
rect 675477 603530 675543 603533
rect 673913 603528 675543 603530
rect 673913 603472 673918 603528
rect 673974 603472 675482 603528
rect 675538 603472 675543 603528
rect 673913 603470 675543 603472
rect 673913 603467 673979 603470
rect 675477 603467 675543 603470
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675293 602986 675359 602989
rect 674484 602984 675359 602986
rect 674484 602928 675298 602984
rect 675354 602928 675359 602984
rect 674484 602926 675359 602928
rect 674484 602924 674490 602926
rect 675293 602923 675359 602926
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 48957 601354 49023 601357
rect 41492 601352 49023 601354
rect 41492 601296 48962 601352
rect 49018 601296 49023 601352
rect 41492 601294 49023 601296
rect 48957 601291 49023 601294
rect 54477 600946 54543 600949
rect 41492 600944 54543 600946
rect 41492 600888 54482 600944
rect 54538 600888 54543 600944
rect 41492 600886 54543 600888
rect 54477 600883 54543 600886
rect 44817 600538 44883 600541
rect 41492 600536 44883 600538
rect 41492 600480 44822 600536
rect 44878 600480 44883 600536
rect 41492 600478 44883 600480
rect 44817 600475 44883 600478
rect 670141 600402 670207 600405
rect 675477 600402 675543 600405
rect 670141 600400 675543 600402
rect 670141 600344 670146 600400
rect 670202 600344 675482 600400
rect 675538 600344 675543 600400
rect 670141 600342 675543 600344
rect 670141 600339 670207 600342
rect 675477 600339 675543 600342
rect 44817 600130 44883 600133
rect 41492 600128 44883 600130
rect 41492 600072 44822 600128
rect 44878 600072 44883 600128
rect 41492 600070 44883 600072
rect 44817 600067 44883 600070
rect 674966 599994 674972 599996
rect 663750 599934 674972 599994
rect 44633 599722 44699 599725
rect 41492 599720 44699 599722
rect 41492 599664 44638 599720
rect 44694 599664 44699 599720
rect 41492 599662 44699 599664
rect 44633 599659 44699 599662
rect 660297 599586 660363 599589
rect 663750 599586 663810 599934
rect 674966 599932 674972 599934
rect 675036 599932 675042 599996
rect 673453 599722 673519 599725
rect 675293 599722 675359 599725
rect 673453 599720 675359 599722
rect 673453 599664 673458 599720
rect 673514 599664 675298 599720
rect 675354 599664 675359 599720
rect 673453 599662 675359 599664
rect 673453 599659 673519 599662
rect 675293 599659 675359 599662
rect 660297 599584 663810 599586
rect 660297 599528 660302 599584
rect 660358 599528 663810 599584
rect 660297 599526 663810 599528
rect 660297 599523 660363 599526
rect 45001 599314 45067 599317
rect 41492 599312 45067 599314
rect 41492 599256 45006 599312
rect 45062 599256 45067 599312
rect 41492 599254 45067 599256
rect 45001 599251 45067 599254
rect 669037 599314 669103 599317
rect 675201 599314 675267 599317
rect 669037 599312 675267 599314
rect 669037 599256 669042 599312
rect 669098 599256 675206 599312
rect 675262 599256 675267 599312
rect 669037 599254 675267 599256
rect 669037 599251 669103 599254
rect 675201 599251 675267 599254
rect 45369 598906 45435 598909
rect 41492 598904 45435 598906
rect 41492 598848 45374 598904
rect 45430 598848 45435 598904
rect 41492 598846 45435 598848
rect 45369 598843 45435 598846
rect 44633 598498 44699 598501
rect 41492 598496 44699 598498
rect 41492 598440 44638 598496
rect 44694 598440 44699 598496
rect 41492 598438 44699 598440
rect 44633 598435 44699 598438
rect 45185 598090 45251 598093
rect 41492 598088 45251 598090
rect 41492 598032 45190 598088
rect 45246 598032 45251 598088
rect 41492 598030 45251 598032
rect 45185 598027 45251 598030
rect 62113 597954 62179 597957
rect 673729 597956 673795 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 673678 597892 673684 597956
rect 673748 597954 673795 597956
rect 673748 597952 673840 597954
rect 673790 597896 673840 597952
rect 673748 597894 673840 597896
rect 673748 597892 673795 597894
rect 673729 597891 673795 597892
rect 41492 597622 42994 597682
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 42934 597005 42994 597622
rect 673453 597410 673519 597413
rect 675385 597410 675451 597413
rect 673453 597408 675451 597410
rect 673453 597352 673458 597408
rect 673514 597352 675390 597408
rect 675446 597352 675451 597408
rect 673453 597350 675451 597352
rect 673453 597347 673519 597350
rect 675385 597347 675451 597350
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 41321 596866 41387 596869
rect 41308 596864 41387 596866
rect 41308 596808 41326 596864
rect 41382 596808 41387 596864
rect 41308 596806 41387 596808
rect 41321 596803 41387 596806
rect 674782 596804 674788 596868
rect 674852 596866 674858 596868
rect 675385 596866 675451 596869
rect 674852 596864 675451 596866
rect 674852 596808 675390 596864
rect 675446 596808 675451 596864
rect 674852 596806 675451 596808
rect 674852 596804 674858 596806
rect 675385 596803 675451 596806
rect 674005 596594 674071 596597
rect 675201 596594 675267 596597
rect 674005 596592 675267 596594
rect 674005 596536 674010 596592
rect 674066 596536 675206 596592
rect 675262 596536 675267 596592
rect 674005 596534 675267 596536
rect 674005 596531 674071 596534
rect 675201 596531 675267 596534
rect 42190 596458 42196 596460
rect 41492 596398 42196 596458
rect 42190 596396 42196 596398
rect 42260 596396 42266 596460
rect 41137 596050 41203 596053
rect 41124 596048 41203 596050
rect 41124 595992 41142 596048
rect 41198 595992 41203 596048
rect 41124 595990 41203 595992
rect 41137 595987 41203 595990
rect 33041 595642 33107 595645
rect 33028 595640 33107 595642
rect 33028 595584 33046 595640
rect 33102 595584 33107 595640
rect 33028 595582 33107 595584
rect 33041 595579 33107 595582
rect 35157 595234 35223 595237
rect 35157 595232 35236 595234
rect 35157 595176 35162 595232
rect 35218 595176 35236 595232
rect 35157 595174 35236 595176
rect 35157 595171 35223 595174
rect 40677 594826 40743 594829
rect 671061 594826 671127 594829
rect 675477 594826 675543 594829
rect 40677 594824 40756 594826
rect 40677 594768 40682 594824
rect 40738 594768 40756 594824
rect 40677 594766 40756 594768
rect 671061 594824 675543 594826
rect 671061 594768 671066 594824
rect 671122 594768 675482 594824
rect 675538 594768 675543 594824
rect 671061 594766 675543 594768
rect 40677 594763 40743 594766
rect 671061 594763 671127 594766
rect 675477 594763 675543 594766
rect 676070 594628 676076 594692
rect 676140 594690 676146 594692
rect 676990 594690 676996 594692
rect 676140 594630 676996 594690
rect 676140 594628 676146 594630
rect 676990 594628 676996 594630
rect 677060 594628 677066 594692
rect 41689 594554 41755 594557
rect 42517 594554 42583 594557
rect 41689 594552 42583 594554
rect 41689 594496 41694 594552
rect 41750 594496 42522 594552
rect 42578 594496 42583 594552
rect 41689 594494 42583 594496
rect 41689 594491 41755 594494
rect 42517 594491 42583 594494
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 42793 594010 42859 594013
rect 41492 594008 42859 594010
rect 41492 593952 42798 594008
rect 42854 593952 42859 594008
rect 41492 593950 42859 593952
rect 42793 593947 42859 593950
rect 41781 593602 41847 593605
rect 41492 593600 41847 593602
rect 41492 593544 41786 593600
rect 41842 593544 41847 593600
rect 41492 593542 41847 593544
rect 41781 593539 41847 593542
rect 668393 593602 668459 593605
rect 675477 593602 675543 593605
rect 668393 593600 675543 593602
rect 668393 593544 668398 593600
rect 668454 593544 675482 593600
rect 675538 593544 675543 593600
rect 668393 593542 675543 593544
rect 668393 593539 668459 593542
rect 675477 593539 675543 593542
rect 41781 593194 41847 593197
rect 675569 593196 675635 593197
rect 675518 593194 675524 593196
rect 41492 593192 41847 593194
rect 41492 593136 41786 593192
rect 41842 593136 41847 593192
rect 41492 593134 41847 593136
rect 675478 593134 675524 593194
rect 675588 593192 675635 593196
rect 675630 593136 675635 593192
rect 41781 593131 41847 593134
rect 675518 593132 675524 593134
rect 675588 593132 675635 593136
rect 675569 593131 675635 593132
rect 675150 592860 675156 592924
rect 675220 592922 675226 592924
rect 676029 592922 676095 592925
rect 675220 592920 676095 592922
rect 675220 592864 676034 592920
rect 676090 592864 676095 592920
rect 675220 592862 676095 592864
rect 675220 592860 675226 592862
rect 676029 592859 676095 592862
rect 41781 592786 41847 592789
rect 41492 592784 41847 592786
rect 41492 592728 41786 592784
rect 41842 592728 41847 592784
rect 41492 592726 41847 592728
rect 41781 592723 41847 592726
rect 673678 592588 673684 592652
rect 673748 592650 673754 592652
rect 683113 592650 683179 592653
rect 673748 592648 683179 592650
rect 673748 592592 683118 592648
rect 683174 592592 683179 592648
rect 673748 592590 683179 592592
rect 673748 592588 673754 592590
rect 683113 592587 683179 592590
rect 41873 592378 41939 592381
rect 41492 592376 41939 592378
rect 41492 592320 41878 592376
rect 41934 592320 41939 592376
rect 41492 592318 41939 592320
rect 41873 592315 41939 592318
rect 674741 592378 674807 592381
rect 675845 592378 675911 592381
rect 674741 592376 675911 592378
rect 674741 592320 674746 592376
rect 674802 592320 675850 592376
rect 675906 592320 675911 592376
rect 674741 592318 675911 592320
rect 674741 592315 674807 592318
rect 675845 592315 675911 592318
rect 44173 591970 44239 591973
rect 41492 591968 44239 591970
rect 41492 591912 44178 591968
rect 44234 591912 44239 591968
rect 41492 591910 44239 591912
rect 44173 591907 44239 591910
rect 43846 591562 43852 591564
rect 41492 591502 43852 591562
rect 43846 591500 43852 591502
rect 43916 591500 43922 591564
rect 674189 591290 674255 591293
rect 683389 591290 683455 591293
rect 674189 591288 683455 591290
rect 674189 591232 674194 591288
rect 674250 591232 683394 591288
rect 683450 591232 683455 591288
rect 674189 591230 683455 591232
rect 674189 591227 674255 591230
rect 683389 591227 683455 591230
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 652385 590746 652451 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 652451 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 652390 590744
rect 652446 590688 652451 590744
rect 650164 590686 652451 590688
rect 39941 590683 40007 590686
rect 652385 590683 652451 590686
rect 43437 590338 43503 590341
rect 41492 590336 43503 590338
rect 41492 590280 43442 590336
rect 43498 590280 43503 590336
rect 41492 590278 43503 590280
rect 43437 590275 43503 590278
rect 674230 589868 674236 589932
rect 674300 589930 674306 589932
rect 683665 589930 683731 589933
rect 674300 589928 683731 589930
rect 674300 589872 683670 589928
rect 683726 589872 683731 589928
rect 674300 589870 683731 589872
rect 674300 589868 674306 589870
rect 683665 589867 683731 589870
rect 40493 589660 40559 589661
rect 40493 589656 40540 589660
rect 40604 589658 40610 589660
rect 40493 589600 40498 589656
rect 40493 589596 40540 589600
rect 40604 589598 40650 589658
rect 40604 589596 40610 589598
rect 40493 589595 40559 589596
rect 40718 589460 40724 589524
rect 40788 589522 40794 589524
rect 41413 589522 41479 589525
rect 40788 589520 41479 589522
rect 40788 589464 41418 589520
rect 41474 589464 41479 589520
rect 40788 589462 41479 589464
rect 40788 589460 40794 589462
rect 41413 589459 41479 589462
rect 41873 589386 41939 589389
rect 41830 589384 41939 589386
rect 41830 589328 41878 589384
rect 41934 589328 41939 589384
rect 41830 589323 41939 589328
rect 40902 589228 40908 589292
rect 40972 589290 40978 589292
rect 41830 589290 41890 589323
rect 40972 589230 41890 589290
rect 40972 589228 40978 589230
rect 675569 586258 675635 586261
rect 676070 586258 676076 586260
rect 675569 586256 676076 586258
rect 675569 586200 675574 586256
rect 675630 586200 676076 586256
rect 675569 586198 676076 586200
rect 675569 586195 675635 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 39941 585986 40007 585989
rect 42333 585986 42399 585989
rect 39941 585984 42399 585986
rect 39941 585928 39946 585984
rect 40002 585928 42338 585984
rect 42394 585928 42399 585984
rect 39941 585926 42399 585928
rect 39941 585923 40007 585926
rect 42333 585923 42399 585926
rect 40125 584898 40191 584901
rect 42374 584898 42380 584900
rect 40125 584896 42380 584898
rect 40125 584840 40130 584896
rect 40186 584840 42380 584896
rect 40125 584838 42380 584840
rect 40125 584835 40191 584838
rect 42374 584836 42380 584838
rect 42444 584836 42450 584900
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 39389 584626 39455 584629
rect 40350 584626 40356 584628
rect 39389 584624 40356 584626
rect 39389 584568 39394 584624
rect 39450 584568 40356 584624
rect 39389 584566 40356 584568
rect 39389 584563 39455 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 40677 584626 40743 584629
rect 41822 584626 41828 584628
rect 40677 584624 41828 584626
rect 40677 584568 40682 584624
rect 40738 584568 41828 584624
rect 40677 584566 41828 584568
rect 40677 584563 40743 584566
rect 41822 584564 41828 584566
rect 41892 584564 41898 584628
rect 41781 584354 41847 584357
rect 42190 584354 42196 584356
rect 41781 584352 42196 584354
rect 41781 584296 41786 584352
rect 41842 584296 42196 584352
rect 41781 584294 42196 584296
rect 41781 584291 41847 584294
rect 42190 584292 42196 584294
rect 42260 584292 42266 584356
rect 673494 582524 673500 582588
rect 673564 582586 673570 582588
rect 673729 582586 673795 582589
rect 673564 582584 673795 582586
rect 673564 582528 673734 582584
rect 673790 582528 673795 582584
rect 673564 582526 673795 582528
rect 673564 582524 673570 582526
rect 673729 582523 673795 582526
rect 42425 582044 42491 582045
rect 42374 582042 42380 582044
rect 42334 581982 42380 582042
rect 42444 582040 42491 582044
rect 42486 581984 42491 582040
rect 42374 581980 42380 581982
rect 42444 581980 42491 581984
rect 42425 581979 42491 581980
rect 675109 581634 675175 581637
rect 675845 581634 675911 581637
rect 675109 581632 675911 581634
rect 675109 581576 675114 581632
rect 675170 581576 675850 581632
rect 675906 581576 675911 581632
rect 675109 581574 675911 581576
rect 675109 581571 675175 581574
rect 675845 581571 675911 581574
rect 40350 581300 40356 581364
rect 40420 581362 40426 581364
rect 42701 581362 42767 581365
rect 40420 581360 42767 581362
rect 40420 581304 42706 581360
rect 42762 581304 42767 581360
rect 40420 581302 42767 581304
rect 40420 581300 40426 581302
rect 42701 581299 42767 581302
rect 44173 581090 44239 581093
rect 42198 581088 44239 581090
rect 42198 581032 44178 581088
rect 44234 581032 44239 581088
rect 42198 581030 44239 581032
rect 42198 580821 42258 581030
rect 44173 581027 44239 581030
rect 669957 581090 670023 581093
rect 669957 581088 676292 581090
rect 669957 581032 669962 581088
rect 670018 581032 676292 581088
rect 669957 581030 676292 581032
rect 669957 581027 670023 581030
rect 41965 580816 42031 580821
rect 41965 580760 41970 580816
rect 42026 580760 42031 580816
rect 41965 580755 42031 580760
rect 42198 580816 42307 580821
rect 42198 580760 42246 580816
rect 42302 580760 42307 580816
rect 42198 580758 42307 580760
rect 42241 580755 42307 580758
rect 671521 580818 671587 580821
rect 675017 580818 675083 580821
rect 671521 580816 675083 580818
rect 671521 580760 671526 580816
rect 671582 580760 675022 580816
rect 675078 580760 675083 580816
rect 671521 580758 675083 580760
rect 671521 580755 671587 580758
rect 675017 580755 675083 580758
rect 41968 580546 42028 580755
rect 47577 580546 47643 580549
rect 676262 580546 676322 580652
rect 41968 580544 47643 580546
rect 41968 580488 47582 580544
rect 47638 580488 47643 580544
rect 41968 580486 47643 580488
rect 47577 580483 47643 580486
rect 674606 580486 676322 580546
rect 673545 580412 673611 580413
rect 673494 580348 673500 580412
rect 673564 580410 673611 580412
rect 673564 580408 673656 580410
rect 673606 580352 673656 580408
rect 673564 580350 673656 580352
rect 673564 580348 673611 580350
rect 673545 580347 673611 580348
rect 41965 580274 42031 580277
rect 42190 580274 42196 580276
rect 41965 580272 42196 580274
rect 41965 580216 41970 580272
rect 42026 580216 42196 580272
rect 41965 580214 42196 580216
rect 41965 580211 42031 580214
rect 42190 580212 42196 580214
rect 42260 580212 42266 580276
rect 664437 580138 664503 580141
rect 674606 580138 674666 580486
rect 676262 580138 676322 580244
rect 664437 580136 674666 580138
rect 664437 580080 664442 580136
rect 664498 580080 674666 580136
rect 664437 580078 674666 580080
rect 674790 580078 676322 580138
rect 664437 580075 664503 580078
rect 658917 579730 658983 579733
rect 674790 579730 674850 580078
rect 675017 579866 675083 579869
rect 675017 579864 676292 579866
rect 675017 579808 675022 579864
rect 675078 579808 676292 579864
rect 675017 579806 676292 579808
rect 675017 579803 675083 579806
rect 658917 579728 674850 579730
rect 658917 579672 658922 579728
rect 658978 579672 674850 579728
rect 658917 579670 674850 579672
rect 658917 579667 658983 579670
rect 671429 579322 671495 579325
rect 676262 579322 676322 579428
rect 671429 579320 676322 579322
rect 671429 579264 671434 579320
rect 671490 579264 676322 579320
rect 671429 579262 676322 579264
rect 671429 579259 671495 579262
rect 671245 578914 671311 578917
rect 676262 578914 676322 579020
rect 671245 578912 676322 578914
rect 671245 578856 671250 578912
rect 671306 578856 676322 578912
rect 671245 578854 676322 578856
rect 671245 578851 671311 578854
rect 672809 578642 672875 578645
rect 672809 578640 676292 578642
rect 672809 578584 672814 578640
rect 672870 578584 676292 578640
rect 672809 578582 676292 578584
rect 672809 578579 672875 578582
rect 675477 578370 675543 578373
rect 674606 578368 675543 578370
rect 674606 578312 675482 578368
rect 675538 578312 675543 578368
rect 674606 578310 675543 578312
rect 40718 578172 40724 578236
rect 40788 578234 40794 578236
rect 41781 578234 41847 578237
rect 40788 578232 41847 578234
rect 40788 578176 41786 578232
rect 41842 578176 41847 578232
rect 40788 578174 41847 578176
rect 40788 578172 40794 578174
rect 41781 578171 41847 578174
rect 674606 578098 674666 578310
rect 675477 578307 675543 578310
rect 676262 578098 676322 578204
rect 671110 578038 674666 578098
rect 674790 578038 676322 578098
rect 40902 577492 40908 577556
rect 40972 577554 40978 577556
rect 41781 577554 41847 577557
rect 40972 577552 41847 577554
rect 40972 577496 41786 577552
rect 41842 577496 41847 577552
rect 40972 577494 41847 577496
rect 671110 577554 671170 578038
rect 671429 577826 671495 577829
rect 671429 577824 673470 577826
rect 671429 577768 671434 577824
rect 671490 577768 673470 577824
rect 671429 577766 673470 577768
rect 671429 577763 671495 577766
rect 673410 577690 673470 577766
rect 674790 577690 674850 578038
rect 673410 577630 674850 577690
rect 675017 577690 675083 577693
rect 676262 577690 676322 577796
rect 675017 577688 676322 577690
rect 675017 577632 675022 577688
rect 675078 577632 676322 577688
rect 675017 577630 676322 577632
rect 675017 577627 675083 577630
rect 671613 577554 671679 577557
rect 671110 577552 671679 577554
rect 671110 577496 671618 577552
rect 671674 577496 671679 577552
rect 671110 577494 671679 577496
rect 40972 577492 40978 577494
rect 41781 577491 41847 577494
rect 671613 577491 671679 577494
rect 651465 577418 651531 577421
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 651465 577355 651531 577358
rect 671797 577282 671863 577285
rect 676262 577282 676322 577388
rect 671797 577280 676322 577282
rect 671797 577224 671802 577280
rect 671858 577224 676322 577280
rect 671797 577222 676322 577224
rect 671797 577219 671863 577222
rect 675477 577010 675543 577013
rect 675477 577008 676292 577010
rect 675477 576952 675482 577008
rect 675538 576952 676292 577008
rect 675477 576950 676292 576952
rect 675477 576947 675543 576950
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 671429 576874 671495 576877
rect 675017 576874 675083 576877
rect 40604 576814 42074 576874
rect 40604 576812 40610 576814
rect 42014 576605 42074 576814
rect 671429 576872 675083 576874
rect 671429 576816 671434 576872
rect 671490 576816 675022 576872
rect 675078 576816 675083 576872
rect 671429 576814 675083 576816
rect 671429 576811 671495 576814
rect 675017 576811 675083 576814
rect 42333 576738 42399 576741
rect 42701 576738 42767 576741
rect 42333 576736 42767 576738
rect 42333 576680 42338 576736
rect 42394 576680 42706 576736
rect 42762 576680 42767 576736
rect 42333 576678 42767 576680
rect 42333 576675 42399 576678
rect 42701 576675 42767 576678
rect 42014 576600 42123 576605
rect 42014 576544 42062 576600
rect 42118 576544 42123 576600
rect 42014 576542 42123 576544
rect 42057 576539 42123 576542
rect 676029 576602 676095 576605
rect 676029 576600 676292 576602
rect 676029 576544 676034 576600
rect 676090 576544 676292 576600
rect 676029 576542 676292 576544
rect 676029 576539 676095 576542
rect 667841 576058 667907 576061
rect 676262 576058 676322 576164
rect 667841 576056 676322 576058
rect 667841 576000 667846 576056
rect 667902 576000 676322 576056
rect 667841 575998 676322 576000
rect 667841 575995 667907 575998
rect 676990 575996 676996 576060
rect 677060 575996 677066 576060
rect 676998 575756 677058 575996
rect 675845 575378 675911 575381
rect 675845 575376 676292 575378
rect 675845 575320 675850 575376
rect 675906 575320 676292 575376
rect 675845 575318 676292 575320
rect 675845 575315 675911 575318
rect 670877 574834 670943 574837
rect 676262 574834 676322 574940
rect 670877 574832 676322 574834
rect 670877 574776 670882 574832
rect 670938 574776 676322 574832
rect 670877 574774 676322 574776
rect 670877 574771 670943 574774
rect 669773 574426 669839 574429
rect 676262 574426 676322 574532
rect 669773 574424 676322 574426
rect 669773 574368 669778 574424
rect 669834 574368 676322 574424
rect 669773 574366 676322 574368
rect 669773 574363 669839 574366
rect 669221 574154 669287 574157
rect 669221 574152 676292 574154
rect 669221 574096 669226 574152
rect 669282 574096 676292 574152
rect 669221 574094 676292 574096
rect 669221 574091 669287 574094
rect 683665 574018 683731 574021
rect 683622 574016 683731 574018
rect 683622 573960 683670 574016
rect 683726 573960 683731 574016
rect 683622 573955 683731 573960
rect 42149 573882 42215 573885
rect 42701 573882 42767 573885
rect 42149 573880 42767 573882
rect 42149 573824 42154 573880
rect 42210 573824 42706 573880
rect 42762 573824 42767 573880
rect 42149 573822 42767 573824
rect 42149 573819 42215 573822
rect 42701 573819 42767 573822
rect 683622 573716 683682 573955
rect 41454 573276 41460 573340
rect 41524 573338 41530 573340
rect 42609 573338 42675 573341
rect 41524 573336 42675 573338
rect 41524 573280 42614 573336
rect 42670 573280 42675 573336
rect 41524 573278 42675 573280
rect 41524 573276 41530 573278
rect 42609 573275 42675 573278
rect 672993 573202 673059 573205
rect 676262 573202 676322 573308
rect 672993 573200 676322 573202
rect 672993 573144 672998 573200
rect 673054 573144 676322 573200
rect 672993 573142 676322 573144
rect 683389 573202 683455 573205
rect 683389 573200 683498 573202
rect 683389 573144 683394 573200
rect 683450 573144 683498 573200
rect 672993 573139 673059 573142
rect 683389 573139 683498 573144
rect 683438 572900 683498 573139
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 676814 572492 676874 572732
rect 41638 572052 41644 572116
rect 41708 572114 41714 572116
rect 42517 572114 42583 572117
rect 41708 572112 42583 572114
rect 41708 572056 42522 572112
rect 42578 572056 42583 572112
rect 41708 572054 42583 572056
rect 41708 572052 41714 572054
rect 42517 572051 42583 572054
rect 672441 571978 672507 571981
rect 676262 571978 676322 572084
rect 683113 571978 683179 571981
rect 672441 571976 676322 571978
rect 672441 571920 672446 571976
rect 672502 571920 676322 571976
rect 672441 571918 676322 571920
rect 683070 571976 683179 571978
rect 683070 571920 683118 571976
rect 683174 571920 683179 571976
rect 672441 571915 672507 571918
rect 683070 571915 683179 571920
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 683070 571676 683130 571915
rect 673177 571162 673243 571165
rect 676262 571162 676322 571268
rect 673177 571160 676322 571162
rect 673177 571104 673182 571160
rect 673238 571104 676322 571160
rect 673177 571102 676322 571104
rect 673177 571099 673243 571102
rect 676262 570754 676322 570860
rect 682377 570754 682443 570757
rect 674790 570694 676322 570754
rect 682334 570752 682443 570754
rect 682334 570696 682382 570752
rect 682438 570696 682443 570752
rect 672993 570346 673059 570349
rect 674790 570346 674850 570694
rect 672993 570344 674850 570346
rect 672993 570288 672998 570344
rect 673054 570288 674850 570344
rect 672993 570286 674850 570288
rect 682334 570691 682443 570696
rect 672993 570283 673059 570286
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682334 570044 682394 570691
rect 671797 569530 671863 569533
rect 676262 569530 676322 569636
rect 671797 569528 676322 569530
rect 671797 569472 671802 569528
rect 671858 569472 676322 569528
rect 671797 569470 676322 569472
rect 671797 569467 671863 569470
rect 42333 569258 42399 569261
rect 62113 569258 62179 569261
rect 42333 569256 62179 569258
rect 42333 569200 42338 569256
rect 42394 569200 62118 569256
rect 62174 569200 62179 569256
rect 42333 569198 62179 569200
rect 42333 569195 42399 569198
rect 62113 569195 62179 569198
rect 667841 564498 667907 564501
rect 675385 564498 675451 564501
rect 667841 564496 675451 564498
rect 667841 564440 667846 564496
rect 667902 564440 675390 564496
rect 675446 564440 675451 564496
rect 667841 564438 675451 564440
rect 667841 564435 667907 564438
rect 675385 564435 675451 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675569 562732 675635 562733
rect 675518 562730 675524 562732
rect 675478 562670 675524 562730
rect 675588 562728 675635 562732
rect 675630 562672 675635 562728
rect 675518 562668 675524 562670
rect 675588 562668 675635 562672
rect 675569 562667 675635 562668
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 674833 559466 674899 559469
rect 675477 559466 675543 559469
rect 674833 559464 675543 559466
rect 674833 559408 674838 559464
rect 674894 559408 675482 559464
rect 675538 559408 675543 559464
rect 674833 559406 675543 559408
rect 674833 559403 674899 559406
rect 675477 559403 675543 559406
rect 673177 559058 673243 559061
rect 675385 559058 675451 559061
rect 673177 559056 675451 559058
rect 673177 559000 673182 559056
rect 673238 559000 675390 559056
rect 675446 559000 675451 559056
rect 673177 558998 675451 559000
rect 673177 558995 673243 558998
rect 675385 558995 675451 558998
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 50337 558514 50403 558517
rect 41492 558512 50403 558514
rect 41492 558456 50342 558512
rect 50398 558456 50403 558512
rect 41492 558454 50403 558456
rect 50337 558451 50403 558454
rect 674189 558378 674255 558381
rect 675385 558378 675451 558381
rect 674189 558376 675451 558378
rect 674189 558320 674194 558376
rect 674250 558320 675390 558376
rect 675446 558320 675451 558376
rect 674189 558318 675451 558320
rect 674189 558315 674255 558318
rect 675385 558315 675451 558318
rect 41321 558106 41387 558109
rect 41308 558104 41387 558106
rect 41308 558048 41326 558104
rect 41382 558048 41387 558104
rect 41308 558046 41387 558048
rect 41321 558043 41387 558046
rect 48957 557698 49023 557701
rect 41492 557696 49023 557698
rect 41492 557640 48962 557696
rect 49018 557640 49023 557696
rect 41492 557638 49023 557640
rect 48957 557635 49023 557638
rect 669221 557562 669287 557565
rect 675477 557562 675543 557565
rect 669221 557560 675543 557562
rect 669221 557504 669226 557560
rect 669282 557504 675482 557560
rect 675538 557504 675543 557560
rect 669221 557502 675543 557504
rect 669221 557499 669287 557502
rect 675477 557499 675543 557502
rect 675753 557562 675819 557565
rect 676254 557562 676260 557564
rect 675753 557560 676260 557562
rect 675753 557504 675758 557560
rect 675814 557504 676260 557560
rect 675753 557502 676260 557504
rect 675753 557499 675819 557502
rect 676254 557500 676260 557502
rect 676324 557500 676330 557564
rect 44817 557290 44883 557293
rect 41492 557288 44883 557290
rect 41492 557232 44822 557288
rect 44878 557232 44883 557288
rect 41492 557230 44883 557232
rect 44817 557227 44883 557230
rect 45553 556882 45619 556885
rect 41492 556880 45619 556882
rect 41492 556824 45558 556880
rect 45614 556824 45619 556880
rect 41492 556822 45619 556824
rect 45553 556819 45619 556822
rect 45001 556474 45067 556477
rect 41492 556472 45067 556474
rect 41492 556416 45006 556472
rect 45062 556416 45067 556472
rect 41492 556414 45067 556416
rect 45001 556411 45067 556414
rect 44909 556066 44975 556069
rect 41492 556064 44975 556066
rect 41492 556008 44914 556064
rect 44970 556008 44975 556064
rect 41492 556006 44975 556008
rect 44909 556003 44975 556006
rect 44633 555658 44699 555661
rect 41492 555656 44699 555658
rect 41492 555600 44638 555656
rect 44694 555600 44699 555656
rect 41492 555598 44699 555600
rect 44633 555595 44699 555598
rect 44725 555250 44791 555253
rect 41492 555248 44791 555250
rect 41492 555192 44730 555248
rect 44786 555192 44791 555248
rect 41492 555190 44791 555192
rect 44725 555187 44791 555190
rect 41321 554842 41387 554845
rect 41308 554840 41387 554842
rect 41308 554784 41326 554840
rect 41382 554784 41387 554840
rect 41308 554782 41387 554784
rect 41321 554779 41387 554782
rect 667657 554706 667723 554709
rect 675385 554706 675451 554709
rect 667657 554704 675451 554706
rect 667657 554648 667662 554704
rect 667718 554648 675390 554704
rect 675446 554648 675451 554704
rect 667657 554646 675451 554648
rect 667657 554643 667723 554646
rect 675385 554643 675451 554646
rect 44357 554434 44423 554437
rect 41492 554432 44423 554434
rect 41492 554376 44362 554432
rect 44418 554376 44423 554432
rect 41492 554374 44423 554376
rect 44357 554371 44423 554374
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 658917 554026 658983 554029
rect 669957 554026 670023 554029
rect 658917 554024 670023 554026
rect 658917 553968 658922 554024
rect 658978 553968 669962 554024
rect 670018 553968 670023 554024
rect 658917 553966 670023 553968
rect 658917 553963 658983 553966
rect 669957 553963 670023 553966
rect 675753 553890 675819 553893
rect 676806 553890 676812 553892
rect 675753 553888 676812 553890
rect 675753 553832 675758 553888
rect 675814 553832 676812 553888
rect 675753 553830 676812 553832
rect 675753 553827 675819 553830
rect 676806 553828 676812 553830
rect 676876 553828 676882 553892
rect 41278 553413 41338 553588
rect 669773 553482 669839 553485
rect 675385 553482 675451 553485
rect 669773 553480 675451 553482
rect 669773 553424 669778 553480
rect 669834 553424 675390 553480
rect 675446 553424 675451 553480
rect 669773 553422 675451 553424
rect 669773 553419 669839 553422
rect 675385 553419 675451 553422
rect 41229 553408 41338 553413
rect 41229 553352 41234 553408
rect 41290 553352 41338 553408
rect 41229 553350 41338 553352
rect 41229 553347 41295 553350
rect 41822 553210 41828 553212
rect 41492 553150 41828 553210
rect 41822 553148 41828 553150
rect 41892 553148 41898 553212
rect 41137 552802 41203 552805
rect 41124 552800 41203 552802
rect 41124 552744 41142 552800
rect 41198 552744 41203 552800
rect 41124 552742 41203 552744
rect 41137 552739 41203 552742
rect 42885 552394 42951 552397
rect 41492 552392 42951 552394
rect 41492 552336 42890 552392
rect 42946 552336 42951 552392
rect 41492 552334 42951 552336
rect 42885 552331 42951 552334
rect 670877 552122 670943 552125
rect 675385 552122 675451 552125
rect 670877 552120 675451 552122
rect 670877 552064 670882 552120
rect 670938 552064 675390 552120
rect 675446 552064 675451 552120
rect 670877 552062 675451 552064
rect 670877 552059 670943 552062
rect 675385 552059 675451 552062
rect 32397 551986 32463 551989
rect 41781 551988 41847 551989
rect 32397 551984 32476 551986
rect 32397 551928 32402 551984
rect 32458 551928 32476 551984
rect 32397 551926 32476 551928
rect 41781 551984 41828 551988
rect 41892 551986 41898 551988
rect 41781 551928 41786 551984
rect 32397 551923 32463 551926
rect 41781 551924 41828 551928
rect 41892 551926 41938 551986
rect 41892 551924 41898 551926
rect 41781 551923 41847 551924
rect 45093 551578 45159 551581
rect 41492 551576 45159 551578
rect 41492 551520 45098 551576
rect 45154 551520 45159 551576
rect 41492 551518 45159 551520
rect 45093 551515 45159 551518
rect 669957 551578 670023 551581
rect 675385 551578 675451 551581
rect 669957 551576 675451 551578
rect 669957 551520 669962 551576
rect 670018 551520 675390 551576
rect 675446 551520 675451 551576
rect 669957 551518 675451 551520
rect 669957 551515 670023 551518
rect 675385 551515 675451 551518
rect 41781 551170 41847 551173
rect 41492 551168 41847 551170
rect 41492 551112 41786 551168
rect 41842 551112 41847 551168
rect 41492 551110 41847 551112
rect 41781 551107 41847 551110
rect 651465 550898 651531 550901
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 651465 550835 651531 550838
rect 44541 550762 44607 550765
rect 41492 550760 44607 550762
rect 41492 550704 44546 550760
rect 44602 550704 44607 550760
rect 41492 550702 44607 550704
rect 44541 550699 44607 550702
rect 675201 550626 675267 550629
rect 675886 550626 675892 550628
rect 675201 550624 675892 550626
rect 675201 550568 675206 550624
rect 675262 550568 675892 550624
rect 675201 550566 675892 550568
rect 675201 550563 675267 550566
rect 675886 550564 675892 550566
rect 675956 550564 675962 550628
rect 40769 550354 40835 550357
rect 40756 550352 40835 550354
rect 40756 550296 40774 550352
rect 40830 550296 40835 550352
rect 40756 550294 40835 550296
rect 40769 550291 40835 550294
rect 675753 550354 675819 550357
rect 676990 550354 676996 550356
rect 675753 550352 676996 550354
rect 675753 550296 675758 550352
rect 675814 550296 676996 550352
rect 675753 550294 676996 550296
rect 675753 550291 675819 550294
rect 676990 550292 676996 550294
rect 677060 550292 677066 550356
rect 41873 550218 41939 550221
rect 43069 550218 43135 550221
rect 41873 550216 43135 550218
rect 41873 550160 41878 550216
rect 41934 550160 43074 550216
rect 43130 550160 43135 550216
rect 41873 550158 43135 550160
rect 41873 550155 41939 550158
rect 43069 550155 43135 550158
rect 41781 549946 41847 549949
rect 41492 549944 41847 549946
rect 41492 549888 41786 549944
rect 41842 549888 41847 549944
rect 41492 549886 41847 549888
rect 41781 549883 41847 549886
rect 41229 549538 41295 549541
rect 41229 549536 41308 549538
rect 41229 549480 41234 549536
rect 41290 549480 41308 549536
rect 41229 549478 41308 549480
rect 41229 549475 41295 549478
rect 44173 549130 44239 549133
rect 41492 549128 44239 549130
rect 41492 549072 44178 549128
rect 44234 549072 44239 549128
rect 41492 549070 44239 549072
rect 44173 549067 44239 549070
rect 45277 548722 45343 548725
rect 41492 548720 45343 548722
rect 41492 548664 45282 548720
rect 45338 548664 45343 548720
rect 41492 548662 45343 548664
rect 45277 548659 45343 548662
rect 674649 548314 674715 548317
rect 675385 548314 675451 548317
rect 674649 548312 675451 548314
rect 41278 548147 41338 548284
rect 674649 548256 674654 548312
rect 674710 548256 675390 548312
rect 675446 548256 675451 548312
rect 674649 548254 675451 548256
rect 674649 548251 674715 548254
rect 675385 548251 675451 548254
rect 31753 548144 31819 548147
rect 31710 548142 31819 548144
rect 31710 548086 31758 548142
rect 31814 548086 31819 548142
rect 31710 548081 31819 548086
rect 41229 548142 41338 548147
rect 41229 548086 41234 548142
rect 41290 548086 41338 548142
rect 41689 548178 41755 548181
rect 43621 548178 43687 548181
rect 41689 548176 43687 548178
rect 41689 548120 41694 548176
rect 41750 548120 43626 548176
rect 43682 548120 43687 548176
rect 41689 548118 43687 548120
rect 41689 548115 41755 548118
rect 43621 548115 43687 548118
rect 41229 548084 41338 548086
rect 41229 548081 41295 548084
rect 28766 547498 28826 547890
rect 31710 547498 31770 548081
rect 675937 547636 676003 547637
rect 675886 547634 675892 547636
rect 675846 547574 675892 547634
rect 675956 547632 676003 547636
rect 675998 547576 676003 547632
rect 675886 547572 675892 547574
rect 675956 547572 676003 547576
rect 676254 547572 676260 547636
rect 676324 547634 676330 547636
rect 677409 547634 677475 547637
rect 676324 547632 677475 547634
rect 676324 547576 677414 547632
rect 677470 547576 677475 547632
rect 676324 547574 677475 547576
rect 676324 547572 676330 547574
rect 675937 547571 676003 547572
rect 677409 547571 677475 547574
rect 28766 547468 31770 547498
rect 28796 547438 31770 547468
rect 43805 547090 43871 547093
rect 41492 547088 43871 547090
rect 41492 547032 43810 547088
rect 43866 547032 43871 547088
rect 41492 547030 43871 547032
rect 43805 547027 43871 547030
rect 673637 547090 673703 547093
rect 683205 547090 683271 547093
rect 673637 547088 683271 547090
rect 673637 547032 673642 547088
rect 673698 547032 683210 547088
rect 683266 547032 683271 547088
rect 673637 547030 683271 547032
rect 673637 547027 673703 547030
rect 683205 547027 683271 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 682377 546818 682443 546821
rect 676140 546816 682443 546818
rect 676140 546760 682382 546816
rect 682438 546760 682443 546816
rect 676140 546758 682443 546760
rect 676140 546756 676146 546758
rect 682377 546755 682443 546758
rect 674833 546274 674899 546277
rect 675385 546274 675451 546277
rect 674833 546272 675451 546274
rect 674833 546216 674838 546272
rect 674894 546216 675390 546272
rect 675446 546216 675451 546272
rect 674833 546214 675451 546216
rect 674833 546211 674899 546214
rect 675385 546211 675451 546214
rect 674833 546002 674899 546005
rect 675334 546002 675340 546004
rect 674833 546000 675340 546002
rect 674833 545944 674838 546000
rect 674894 545944 675340 546000
rect 674833 545942 675340 545944
rect 674833 545939 674899 545942
rect 675334 545940 675340 545942
rect 675404 545940 675410 546004
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40769 545732 40835 545733
rect 40718 545730 40724 545732
rect 40678 545670 40724 545730
rect 40788 545728 40835 545732
rect 40830 545672 40835 545728
rect 40718 545668 40724 545670
rect 40788 545668 40835 545672
rect 40769 545667 40835 545668
rect 673913 545730 673979 545733
rect 683389 545730 683455 545733
rect 673913 545728 683455 545730
rect 673913 545672 673918 545728
rect 673974 545672 683394 545728
rect 683450 545672 683455 545728
rect 673913 545670 683455 545672
rect 673913 545667 673979 545670
rect 683389 545667 683455 545670
rect 40585 545460 40651 545461
rect 40534 545458 40540 545460
rect 40494 545398 40540 545458
rect 40604 545456 40651 545460
rect 40646 545400 40651 545456
rect 40534 545396 40540 545398
rect 40604 545396 40651 545400
rect 40585 545395 40651 545396
rect 675201 545458 675267 545461
rect 675518 545458 675524 545460
rect 675201 545456 675524 545458
rect 675201 545400 675206 545456
rect 675262 545400 675524 545456
rect 675201 545398 675524 545400
rect 675201 545395 675267 545398
rect 675518 545396 675524 545398
rect 675588 545396 675594 545460
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 663057 538794 663123 538797
rect 676489 538794 676555 538797
rect 663057 538792 676555 538794
rect 663057 538736 663062 538792
rect 663118 538736 676494 538792
rect 676550 538736 676555 538792
rect 663057 538734 676555 538736
rect 663057 538731 663123 538734
rect 676489 538731 676555 538734
rect 651465 537570 651531 537573
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 651465 537507 651531 537510
rect 42517 537434 42583 537437
rect 44173 537434 44239 537437
rect 42517 537432 44239 537434
rect 42517 537376 42522 537432
rect 42578 537376 44178 537432
rect 44234 537376 44239 537432
rect 42517 537374 44239 537376
rect 42517 537371 42583 537374
rect 44173 537371 44239 537374
rect 40718 536964 40724 537028
rect 40788 537026 40794 537028
rect 41781 537026 41847 537029
rect 40788 537024 41847 537026
rect 40788 536968 41786 537024
rect 41842 536968 41847 537024
rect 40788 536966 41847 536968
rect 40788 536964 40794 536966
rect 41781 536963 41847 536966
rect 42057 537026 42123 537029
rect 45277 537026 45343 537029
rect 42057 537024 45343 537026
rect 42057 536968 42062 537024
rect 42118 536968 45282 537024
rect 45338 536968 45343 537024
rect 42057 536966 45343 536968
rect 42057 536963 42123 536966
rect 45277 536963 45343 536966
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 676489 535938 676555 535941
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 676446 535936 676555 535938
rect 676446 535880 676494 535936
rect 676550 535880 676555 535936
rect 668577 535875 668643 535878
rect 676446 535875 676555 535880
rect 676446 535704 676506 535875
rect 674005 535394 674071 535397
rect 674005 535392 676322 535394
rect 674005 535336 674010 535392
rect 674066 535336 676322 535392
rect 674005 535334 676322 535336
rect 674005 535331 674071 535334
rect 676262 535296 676322 535334
rect 40534 535196 40540 535260
rect 40604 535258 40610 535260
rect 41781 535258 41847 535261
rect 40604 535256 41847 535258
rect 40604 535200 41786 535256
rect 41842 535200 41847 535256
rect 40604 535198 41847 535200
rect 40604 535196 40610 535198
rect 41781 535195 41847 535198
rect 672349 535122 672415 535125
rect 675753 535122 675819 535125
rect 672349 535120 675819 535122
rect 672349 535064 672354 535120
rect 672410 535064 675758 535120
rect 675814 535064 675819 535120
rect 672349 535062 675819 535064
rect 672349 535059 672415 535062
rect 675753 535059 675819 535062
rect 671245 534714 671311 534717
rect 676262 534714 676322 534888
rect 671245 534712 676322 534714
rect 671245 534656 671250 534712
rect 671306 534656 676322 534712
rect 671245 534654 676322 534656
rect 671245 534651 671311 534654
rect 675753 534510 675819 534513
rect 675753 534508 676292 534510
rect 675753 534452 675758 534508
rect 675814 534452 676292 534508
rect 675753 534450 676292 534452
rect 675753 534447 675819 534450
rect 672809 534306 672875 534309
rect 672809 534304 676322 534306
rect 672809 534248 672814 534304
rect 672870 534248 676322 534304
rect 672809 534246 676322 534248
rect 672809 534243 672875 534246
rect 42885 534170 42951 534173
rect 42198 534168 42951 534170
rect 42198 534112 42890 534168
rect 42946 534112 42951 534168
rect 42198 534110 42951 534112
rect 42198 533901 42258 534110
rect 42885 534107 42951 534110
rect 667197 534170 667263 534173
rect 667197 534168 672642 534170
rect 667197 534112 667202 534168
rect 667258 534112 672642 534168
rect 667197 534110 672642 534112
rect 667197 534107 667263 534110
rect 672582 534034 672642 534110
rect 676262 534072 676322 534246
rect 674005 534034 674071 534037
rect 672582 534032 674071 534034
rect 672582 533976 674010 534032
rect 674066 533976 674071 534032
rect 672582 533974 674071 533976
rect 674005 533971 674071 533974
rect 42149 533896 42258 533901
rect 42149 533840 42154 533896
rect 42210 533840 42258 533896
rect 42149 533838 42258 533840
rect 42149 533835 42215 533838
rect 674414 533836 674420 533900
rect 674484 533898 674490 533900
rect 683573 533898 683639 533901
rect 674484 533896 683639 533898
rect 674484 533840 683578 533896
rect 683634 533840 683639 533896
rect 674484 533838 683639 533840
rect 674484 533836 674490 533838
rect 683573 533835 683639 533838
rect 674005 533490 674071 533493
rect 676262 533490 676322 533664
rect 674005 533488 676322 533490
rect 674005 533432 674010 533488
rect 674066 533432 676322 533488
rect 674005 533430 676322 533432
rect 674005 533427 674071 533430
rect 671429 533082 671495 533085
rect 676262 533082 676322 533256
rect 671429 533080 676322 533082
rect 671429 533024 671434 533080
rect 671490 533024 676322 533080
rect 671429 533022 676322 533024
rect 671429 533019 671495 533022
rect 44541 532810 44607 532813
rect 42566 532808 44607 532810
rect 42566 532752 44546 532808
rect 44602 532752 44607 532808
rect 42566 532750 44607 532752
rect 42566 532677 42626 532750
rect 44541 532747 44607 532750
rect 62113 532810 62179 532813
rect 672809 532810 672875 532813
rect 676262 532810 676322 532848
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 672809 532808 676322 532810
rect 672809 532752 672814 532808
rect 672870 532752 676322 532808
rect 672809 532750 676322 532752
rect 62113 532747 62179 532750
rect 672809 532747 672875 532750
rect 42517 532672 42626 532677
rect 42517 532616 42522 532672
rect 42578 532616 42626 532672
rect 42517 532614 42626 532616
rect 42517 532611 42583 532614
rect 674557 532266 674623 532269
rect 676262 532266 676322 532440
rect 674557 532264 676322 532266
rect 674557 532208 674562 532264
rect 674618 532208 676322 532264
rect 674557 532206 676322 532208
rect 674557 532203 674623 532206
rect 672717 531994 672783 531997
rect 676262 531994 676322 532032
rect 672717 531992 676322 531994
rect 672717 531936 672722 531992
rect 672778 531936 676322 531992
rect 672717 531934 676322 531936
rect 672717 531931 672783 531934
rect 672533 531722 672599 531725
rect 672533 531720 676322 531722
rect 672533 531664 672538 531720
rect 672594 531664 676322 531720
rect 672533 531662 676322 531664
rect 672533 531659 672599 531662
rect 676262 531624 676322 531662
rect 671613 531450 671679 531453
rect 674557 531450 674623 531453
rect 671613 531448 674623 531450
rect 671613 531392 671618 531448
rect 671674 531392 674562 531448
rect 674618 531392 674623 531448
rect 671613 531390 674623 531392
rect 671613 531387 671679 531390
rect 674557 531387 674623 531390
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 682377 531042 682443 531045
rect 682334 531040 682443 531042
rect 682334 530984 682382 531040
rect 682438 530984 682443 531040
rect 682334 530979 682443 530984
rect 682334 530808 682394 530979
rect 674373 530634 674439 530637
rect 674373 530632 676322 530634
rect 674373 530576 674378 530632
rect 674434 530576 676322 530632
rect 674373 530574 676322 530576
rect 674373 530571 674439 530574
rect 676262 530400 676322 530574
rect 41454 529892 41460 529956
rect 41524 529954 41530 529956
rect 670141 529954 670207 529957
rect 676262 529954 676322 529992
rect 41524 529894 42258 529954
rect 41524 529892 41530 529894
rect 42198 529549 42258 529894
rect 670141 529952 676322 529954
rect 670141 529896 670146 529952
rect 670202 529896 676322 529952
rect 670141 529894 676322 529896
rect 670141 529891 670207 529894
rect 42425 529818 42491 529821
rect 45093 529818 45159 529821
rect 42425 529816 45159 529818
rect 42425 529760 42430 529816
rect 42486 529760 45098 529816
rect 45154 529760 45159 529816
rect 42425 529758 45159 529760
rect 42425 529755 42491 529758
rect 45093 529755 45159 529758
rect 42198 529544 42307 529549
rect 42198 529488 42246 529544
rect 42302 529488 42307 529544
rect 42198 529486 42307 529488
rect 42241 529483 42307 529486
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 674557 529410 674623 529413
rect 676262 529410 676322 529584
rect 674557 529408 676322 529410
rect 674557 529352 674562 529408
rect 674618 529352 676322 529408
rect 674557 529350 676322 529352
rect 674557 529347 674623 529350
rect 41638 529076 41644 529140
rect 41708 529138 41714 529140
rect 42701 529138 42767 529141
rect 41708 529136 42767 529138
rect 41708 529080 42706 529136
rect 42762 529080 42767 529136
rect 41708 529078 42767 529080
rect 41708 529076 41714 529078
rect 42701 529075 42767 529078
rect 672165 529138 672231 529141
rect 676262 529138 676322 529176
rect 672165 529136 676322 529138
rect 672165 529080 672170 529136
rect 672226 529080 676322 529136
rect 672165 529078 676322 529080
rect 672165 529075 672231 529078
rect 668761 528866 668827 528869
rect 668761 528864 676322 528866
rect 668761 528808 668766 528864
rect 668822 528808 676322 528864
rect 668761 528806 676322 528808
rect 668761 528803 668827 528806
rect 676262 528768 676322 528806
rect 668393 528594 668459 528597
rect 674557 528594 674623 528597
rect 668393 528592 674623 528594
rect 668393 528536 668398 528592
rect 668454 528536 674562 528592
rect 674618 528536 674623 528592
rect 668393 528534 674623 528536
rect 668393 528531 668459 528534
rect 674557 528531 674623 528534
rect 673821 528322 673887 528325
rect 676262 528322 676322 528360
rect 673821 528320 676322 528322
rect 673821 528264 673826 528320
rect 673882 528264 676322 528320
rect 673821 528262 676322 528264
rect 673821 528259 673887 528262
rect 683205 528186 683271 528189
rect 683205 528184 683314 528186
rect 683205 528128 683210 528184
rect 683266 528128 683314 528184
rect 683205 528123 683314 528128
rect 683254 527952 683314 528123
rect 669037 527370 669103 527373
rect 676262 527370 676322 527544
rect 669037 527368 676322 527370
rect 669037 527312 669042 527368
rect 669098 527312 676322 527368
rect 669037 527310 676322 527312
rect 683573 527370 683639 527373
rect 683573 527368 683682 527370
rect 683573 527312 683578 527368
rect 683634 527312 683682 527368
rect 669037 527307 669103 527310
rect 683573 527307 683682 527312
rect 683622 527136 683682 527307
rect 673545 526962 673611 526965
rect 673545 526960 676322 526962
rect 673545 526904 673550 526960
rect 673606 526904 676322 526960
rect 673545 526902 676322 526904
rect 673545 526899 673611 526902
rect 676262 526728 676322 526902
rect 683389 526554 683455 526557
rect 683389 526552 683498 526554
rect 683389 526496 683394 526552
rect 683450 526496 683498 526552
rect 683389 526491 683498 526496
rect 683438 526320 683498 526491
rect 682886 525738 682946 525912
rect 683113 525738 683179 525741
rect 682886 525736 683179 525738
rect 682886 525680 683118 525736
rect 683174 525680 683179 525736
rect 682886 525678 683179 525680
rect 683113 525675 683179 525678
rect 671061 524922 671127 524925
rect 676262 524922 676322 525504
rect 671061 524920 676322 524922
rect 671061 524864 671066 524920
rect 671122 524864 676322 524920
rect 671061 524862 676322 524864
rect 671061 524859 671127 524862
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 675017 510234 675083 510237
rect 675845 510234 675911 510237
rect 675017 510232 675911 510234
rect 675017 510176 675022 510232
rect 675078 510176 675850 510232
rect 675906 510176 675911 510232
rect 675017 510174 675911 510176
rect 675017 510171 675083 510174
rect 675845 510171 675911 510174
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 675201 503706 675267 503709
rect 675845 503706 675911 503709
rect 675201 503704 675911 503706
rect 675201 503648 675206 503704
rect 675262 503648 675850 503704
rect 675906 503648 675911 503704
rect 675201 503646 675911 503648
rect 675201 503643 675267 503646
rect 675845 503643 675911 503646
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683573 503706 683639 503709
rect 677060 503704 683639 503706
rect 677060 503648 683578 503704
rect 683634 503648 683639 503704
rect 677060 503646 683639 503648
rect 677060 503644 677066 503646
rect 683573 503643 683639 503646
rect 676806 503372 676812 503436
rect 676876 503434 676882 503436
rect 683389 503434 683455 503437
rect 676876 503432 683455 503434
rect 676876 503376 683394 503432
rect 683450 503376 683455 503432
rect 676876 503374 683455 503376
rect 676876 503372 676882 503374
rect 683389 503371 683455 503374
rect 675017 503162 675083 503165
rect 675385 503162 675451 503165
rect 675017 503160 675451 503162
rect 675017 503104 675022 503160
rect 675078 503104 675390 503160
rect 675446 503104 675451 503160
rect 675017 503102 675451 503104
rect 675017 503099 675083 503102
rect 675385 503099 675451 503102
rect 671981 501666 672047 501669
rect 677041 501666 677107 501669
rect 671981 501664 677107 501666
rect 671981 501608 671986 501664
rect 672042 501608 677046 501664
rect 677102 501608 677107 501664
rect 671981 501606 677107 501608
rect 671981 501603 672047 501606
rect 677041 501603 677107 501606
rect 672993 500986 673059 500989
rect 675661 500986 675727 500989
rect 672993 500984 675727 500986
rect 672993 500928 672998 500984
rect 673054 500928 675666 500984
rect 675722 500928 675727 500984
rect 672993 500926 675727 500928
rect 672993 500923 673059 500926
rect 675661 500923 675727 500926
rect 652569 497722 652635 497725
rect 650164 497720 652635 497722
rect 650164 497664 652574 497720
rect 652630 497664 652635 497720
rect 650164 497662 652635 497664
rect 652569 497659 652635 497662
rect 664437 494730 664503 494733
rect 683113 494730 683179 494733
rect 664437 494728 683179 494730
rect 664437 494672 664442 494728
rect 664498 494672 683118 494728
rect 683174 494672 683179 494728
rect 664437 494670 683179 494672
rect 664437 494667 664503 494670
rect 683113 494667 683179 494670
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 665817 492146 665883 492149
rect 665817 492144 676292 492146
rect 665817 492088 665822 492144
rect 665878 492088 676292 492144
rect 665817 492086 676292 492088
rect 665817 492083 665883 492086
rect 663750 491678 676292 491738
rect 661677 491602 661743 491605
rect 663750 491602 663810 491678
rect 661677 491600 663810 491602
rect 661677 491544 661682 491600
rect 661738 491544 663810 491600
rect 661677 491542 663810 491544
rect 661677 491539 661743 491542
rect 683113 491330 683179 491333
rect 683100 491328 683179 491330
rect 683100 491272 683118 491328
rect 683174 491272 683179 491328
rect 683100 491270 683179 491272
rect 683113 491267 683179 491270
rect 672441 490922 672507 490925
rect 672441 490920 676292 490922
rect 672441 490864 672446 490920
rect 672502 490864 676292 490920
rect 672441 490862 676292 490864
rect 672441 490859 672507 490862
rect 675569 490514 675635 490517
rect 675569 490512 676292 490514
rect 675569 490456 675574 490512
rect 675630 490456 676292 490512
rect 675569 490454 676292 490456
rect 675569 490451 675635 490454
rect 674005 490106 674071 490109
rect 674005 490104 676292 490106
rect 674005 490048 674010 490104
rect 674066 490048 676292 490104
rect 674005 490046 676292 490048
rect 674005 490043 674071 490046
rect 672441 489698 672507 489701
rect 672441 489696 676292 489698
rect 672441 489640 672446 489696
rect 672502 489640 676292 489696
rect 672441 489638 676292 489640
rect 672441 489635 672507 489638
rect 672809 489290 672875 489293
rect 672809 489288 676292 489290
rect 672809 489232 672814 489288
rect 672870 489232 676292 489288
rect 672809 489230 676292 489232
rect 672809 489227 672875 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 672625 488474 672691 488477
rect 672625 488472 676292 488474
rect 672625 488416 672630 488472
rect 672686 488416 676292 488472
rect 672625 488414 676292 488416
rect 672625 488411 672691 488414
rect 672625 488066 672691 488069
rect 672625 488064 676292 488066
rect 672625 488008 672630 488064
rect 672686 488008 676292 488064
rect 672625 488006 676292 488008
rect 672625 488003 672691 488006
rect 675109 487658 675175 487661
rect 675109 487656 676292 487658
rect 675109 487600 675114 487656
rect 675170 487600 676292 487656
rect 675109 487598 676292 487600
rect 675109 487595 675175 487598
rect 683573 487250 683639 487253
rect 683573 487248 683652 487250
rect 683573 487192 683578 487248
rect 683634 487192 683652 487248
rect 683573 487190 683652 487192
rect 683573 487187 683639 487190
rect 679617 486842 679683 486845
rect 679604 486840 679683 486842
rect 679604 486784 679622 486840
rect 679678 486784 679683 486840
rect 679604 486782 679683 486784
rect 679617 486779 679683 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 669221 486026 669287 486029
rect 669221 486024 676292 486026
rect 669221 485968 669226 486024
rect 669282 485968 676292 486024
rect 669221 485966 676292 485968
rect 669221 485963 669287 485966
rect 674741 485618 674807 485621
rect 674741 485616 676292 485618
rect 674741 485560 674746 485616
rect 674802 485560 676292 485616
rect 674741 485558 676292 485560
rect 674741 485555 674807 485558
rect 667841 485210 667907 485213
rect 667841 485208 676292 485210
rect 667841 485152 667846 485208
rect 667902 485152 676292 485208
rect 667841 485150 676292 485152
rect 667841 485147 667907 485150
rect 673177 484802 673243 484805
rect 673177 484800 676292 484802
rect 673177 484744 673182 484800
rect 673238 484744 676292 484800
rect 673177 484742 676292 484744
rect 673177 484739 673243 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 674189 484394 674255 484397
rect 674189 484392 676292 484394
rect 674189 484336 674194 484392
rect 674250 484336 676292 484392
rect 674189 484334 676292 484336
rect 674189 484331 674255 484334
rect 670877 483986 670943 483989
rect 670877 483984 676292 483986
rect 670877 483928 670882 483984
rect 670938 483928 676292 483984
rect 670877 483926 676292 483928
rect 670877 483923 670943 483926
rect 683389 483578 683455 483581
rect 683389 483576 683468 483578
rect 683389 483520 683394 483576
rect 683450 483520 683468 483576
rect 683389 483518 683468 483520
rect 683389 483515 683455 483518
rect 683113 483170 683179 483173
rect 683100 483168 683179 483170
rect 683100 483112 683118 483168
rect 683174 483112 683179 483168
rect 683100 483110 683179 483112
rect 683113 483107 683179 483110
rect 667657 482762 667723 482765
rect 667657 482760 676292 482762
rect 667657 482704 667662 482760
rect 667718 482704 676292 482760
rect 667657 482702 676292 482704
rect 667657 482699 667723 482702
rect 669773 482354 669839 482357
rect 669773 482352 676292 482354
rect 669773 482296 669778 482352
rect 669834 482296 676292 482352
rect 669773 482294 676292 482296
rect 669773 482291 669839 482294
rect 675753 481946 675819 481949
rect 675753 481944 676292 481946
rect 675753 481888 675758 481944
rect 675814 481888 676292 481944
rect 675753 481886 676292 481888
rect 675753 481883 675819 481886
rect 680997 481538 681063 481541
rect 678500 481536 681063 481538
rect 678500 481508 681002 481536
rect 678470 481480 681002 481508
rect 681058 481480 681063 481536
rect 678470 481478 681063 481480
rect 678470 481100 678530 481478
rect 680997 481475 681063 481478
rect 675526 480662 676292 480722
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 675526 480045 675586 480662
rect 675477 480040 675586 480045
rect 675477 479984 675482 480040
rect 675538 479984 675586 480040
rect 675477 479982 675586 479984
rect 675477 479979 675543 479982
rect 674598 474812 674604 474876
rect 674668 474874 674674 474876
rect 676397 474874 676463 474877
rect 674668 474872 676463 474874
rect 674668 474816 676402 474872
rect 676458 474816 676463 474872
rect 674668 474814 676463 474816
rect 674668 474812 674674 474814
rect 676397 474811 676463 474814
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 673085 457058 673151 457061
rect 676121 457058 676187 457061
rect 673085 457056 676187 457058
rect 673085 457000 673090 457056
rect 673146 457000 676126 457056
rect 676182 457000 676187 457056
rect 673085 456998 676187 457000
rect 673085 456995 673151 456998
rect 676121 456995 676187 456998
rect 673821 456106 673887 456109
rect 676397 456106 676463 456109
rect 673821 456104 676463 456106
rect 673821 456048 673826 456104
rect 673882 456048 676402 456104
rect 676458 456048 676463 456104
rect 673821 456046 676463 456048
rect 673821 456043 673887 456046
rect 676397 456043 676463 456046
rect 670601 455834 670667 455837
rect 673729 455834 673795 455837
rect 670601 455832 673795 455834
rect 670601 455776 670606 455832
rect 670662 455776 673734 455832
rect 673790 455776 673795 455832
rect 670601 455774 673795 455776
rect 670601 455771 670667 455774
rect 673729 455771 673795 455774
rect 673591 455562 673657 455565
rect 675845 455562 675911 455565
rect 673591 455560 675911 455562
rect 673591 455504 673596 455560
rect 673652 455504 675850 455560
rect 675906 455504 675911 455560
rect 673591 455502 675911 455504
rect 673591 455499 673657 455502
rect 675845 455499 675911 455502
rect 670417 455290 670483 455293
rect 673381 455290 673447 455293
rect 670417 455288 673447 455290
rect 670417 455232 670422 455288
rect 670478 455232 673386 455288
rect 673442 455232 673447 455288
rect 670417 455230 673447 455232
rect 670417 455227 670483 455230
rect 673381 455227 673447 455230
rect 669589 455018 669655 455021
rect 672257 455018 672323 455021
rect 669589 455016 672323 455018
rect 669589 454960 669594 455016
rect 669650 454960 672262 455016
rect 672318 454960 672323 455016
rect 669589 454958 672323 454960
rect 669589 454955 669655 454958
rect 672257 454955 672323 454958
rect 672901 454882 672967 454885
rect 676857 454882 676923 454885
rect 672901 454880 676923 454882
rect 672901 454824 672906 454880
rect 672962 454824 676862 454880
rect 676918 454824 676923 454880
rect 672901 454822 676923 454824
rect 672901 454819 672967 454822
rect 676857 454819 676923 454822
rect 62113 454610 62179 454613
rect 673157 454610 673223 454613
rect 676029 454610 676095 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 673157 454608 676095 454610
rect 673157 454552 673162 454608
rect 673218 454552 676034 454608
rect 676090 454552 676095 454608
rect 673157 454550 676095 454552
rect 62113 454547 62179 454550
rect 673157 454547 673223 454550
rect 676029 454547 676095 454550
rect 672809 454202 672875 454205
rect 675569 454202 675635 454205
rect 672809 454200 675635 454202
rect 672809 454144 672814 454200
rect 672870 454144 675574 454200
rect 675630 454144 675635 454200
rect 672809 454142 675635 454144
rect 672809 454139 672875 454142
rect 675569 454139 675635 454142
rect 672257 453930 672323 453933
rect 674741 453930 674807 453933
rect 672257 453928 674807 453930
rect 672257 453872 672262 453928
rect 672318 453872 674746 453928
rect 674802 453872 674807 453928
rect 672257 453870 674807 453872
rect 672257 453867 672323 453870
rect 674741 453867 674807 453870
rect 674925 453930 674991 453933
rect 675334 453930 675340 453932
rect 674925 453928 675340 453930
rect 674925 453872 674930 453928
rect 674986 453872 675340 453928
rect 674925 453870 675340 453872
rect 674925 453867 674991 453870
rect 675334 453868 675340 453870
rect 675404 453868 675410 453932
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45553 429722 45619 429725
rect 41492 429720 45619 429722
rect 41492 429664 45558 429720
rect 45614 429664 45619 429720
rect 41492 429662 45619 429664
rect 45553 429659 45619 429662
rect 44541 429314 44607 429317
rect 41492 429312 44607 429314
rect 41492 429256 44546 429312
rect 44602 429256 44607 429312
rect 41492 429254 44607 429256
rect 44541 429251 44607 429254
rect 44909 428906 44975 428909
rect 41492 428904 44975 428906
rect 41492 428848 44914 428904
rect 44970 428848 44975 428904
rect 41492 428846 44975 428848
rect 44909 428843 44975 428846
rect 45001 428498 45067 428501
rect 41492 428496 45067 428498
rect 41492 428440 45006 428496
rect 45062 428440 45067 428496
rect 41492 428438 45067 428440
rect 45001 428435 45067 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44725 428090 44791 428093
rect 41492 428088 44791 428090
rect 41492 428032 44730 428088
rect 44786 428032 44791 428088
rect 41492 428030 44791 428032
rect 44725 428027 44791 428030
rect 44357 427682 44423 427685
rect 41492 427680 44423 427682
rect 41492 427624 44362 427680
rect 44418 427624 44423 427680
rect 41492 427622 44423 427624
rect 44357 427619 44423 427622
rect 44173 427274 44239 427277
rect 41492 427272 44239 427274
rect 41492 427216 44178 427272
rect 44234 427216 44239 427272
rect 41492 427214 44239 427216
rect 44173 427211 44239 427214
rect 45185 426866 45251 426869
rect 41492 426864 45251 426866
rect 41492 426808 45190 426864
rect 45246 426808 45251 426864
rect 41492 426806 45251 426808
rect 45185 426803 45251 426806
rect 46933 426458 46999 426461
rect 41492 426456 46999 426458
rect 41492 426400 46938 426456
rect 46994 426400 46999 426456
rect 41492 426398 46999 426400
rect 46933 426395 46999 426398
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 40953 425642 41019 425645
rect 40940 425640 41019 425642
rect 40940 425584 40958 425640
rect 41014 425584 41019 425640
rect 40940 425582 41019 425584
rect 40953 425579 41019 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 33685 424418 33751 424421
rect 33685 424416 33764 424418
rect 33685 424360 33690 424416
rect 33746 424360 33764 424416
rect 33685 424358 33764 424360
rect 33685 424355 33751 424358
rect 41321 424010 41387 424013
rect 41308 424008 41387 424010
rect 41308 423952 41326 424008
rect 41382 423952 41387 424008
rect 41308 423950 41387 423952
rect 41321 423947 41387 423950
rect 41781 423874 41847 423877
rect 42793 423874 42859 423877
rect 41781 423872 42859 423874
rect 41781 423816 41786 423872
rect 41842 423816 42798 423872
rect 42854 423816 42859 423872
rect 41781 423814 42859 423816
rect 41781 423811 41847 423814
rect 42793 423811 42859 423814
rect 47117 423602 47183 423605
rect 41492 423600 47183 423602
rect 41492 423544 47122 423600
rect 47178 423544 47183 423600
rect 41492 423542 47183 423544
rect 47117 423539 47183 423542
rect 45369 423194 45435 423197
rect 41492 423192 45435 423194
rect 41492 423136 45374 423192
rect 45430 423136 45435 423192
rect 41492 423134 45435 423136
rect 45369 423131 45435 423134
rect 42149 422786 42215 422789
rect 41492 422784 42215 422786
rect 41492 422728 42154 422784
rect 42210 422728 42215 422784
rect 41492 422726 42215 422728
rect 42149 422723 42215 422726
rect 41321 422378 41387 422381
rect 41308 422376 41387 422378
rect 41308 422320 41326 422376
rect 41382 422320 41387 422376
rect 41308 422318 41387 422320
rect 41321 422315 41387 422318
rect 41781 422378 41847 422381
rect 43161 422378 43227 422381
rect 41781 422376 43227 422378
rect 41781 422320 41786 422376
rect 41842 422320 43166 422376
rect 43222 422320 43227 422376
rect 41781 422318 43227 422320
rect 41781 422315 41847 422318
rect 43161 422315 43227 422318
rect 42333 421970 42399 421973
rect 41492 421968 42399 421970
rect 41492 421912 42338 421968
rect 42394 421912 42399 421968
rect 41492 421910 42399 421912
rect 42333 421907 42399 421910
rect 44173 421562 44239 421565
rect 41492 421560 44239 421562
rect 41492 421504 44178 421560
rect 44234 421504 44239 421560
rect 41492 421502 44239 421504
rect 44173 421499 44239 421502
rect 41781 421292 41847 421293
rect 41781 421290 41828 421292
rect 41736 421288 41828 421290
rect 41736 421232 41786 421288
rect 41736 421230 41828 421232
rect 41781 421228 41828 421230
rect 41892 421228 41898 421292
rect 41781 421227 41847 421228
rect 41321 421154 41387 421157
rect 41308 421152 41387 421154
rect 41308 421096 41326 421152
rect 41382 421096 41387 421152
rect 41308 421094 41387 421096
rect 41321 421091 41387 421094
rect 41781 421018 41847 421021
rect 42977 421018 43043 421021
rect 41781 421016 43043 421018
rect 41781 420960 41786 421016
rect 41842 420960 42982 421016
rect 43038 420960 43043 421016
rect 41781 420958 43043 420960
rect 41781 420955 41847 420958
rect 42977 420955 43043 420958
rect 44817 420746 44883 420749
rect 41492 420744 44883 420746
rect 41492 420688 44822 420744
rect 44878 420688 44883 420744
rect 41492 420686 44883 420688
rect 44817 420683 44883 420686
rect 41462 419930 41522 420308
rect 42517 419930 42583 419933
rect 41462 419928 42583 419930
rect 41462 419900 42522 419928
rect 41492 419872 42522 419900
rect 42578 419872 42583 419928
rect 41492 419870 42583 419872
rect 42517 419867 42583 419870
rect 43989 419522 44055 419525
rect 41492 419520 44055 419522
rect 41492 419464 43994 419520
rect 44050 419464 44055 419520
rect 41492 419462 44055 419464
rect 43989 419459 44055 419462
rect 40718 418780 40724 418844
rect 40788 418842 40794 418844
rect 42149 418842 42215 418845
rect 40788 418840 42215 418842
rect 40788 418784 42154 418840
rect 42210 418784 42215 418840
rect 40788 418782 42215 418784
rect 40788 418780 40794 418782
rect 42149 418779 42215 418782
rect 40350 418508 40356 418572
rect 40420 418570 40426 418572
rect 42333 418570 42399 418573
rect 40420 418568 42399 418570
rect 40420 418512 42338 418568
rect 42394 418512 42399 418568
rect 40420 418510 42399 418512
rect 40420 418508 40426 418510
rect 42333 418507 42399 418510
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 62941 415442 63007 415445
rect 62941 415440 64492 415442
rect 62941 415384 62946 415440
rect 63002 415384 64492 415440
rect 62941 415382 64492 415384
rect 62941 415379 63007 415382
rect 42057 411906 42123 411909
rect 42609 411906 42675 411909
rect 42057 411904 42675 411906
rect 42057 411848 42062 411904
rect 42118 411848 42614 411904
rect 42670 411848 42675 411904
rect 42057 411846 42675 411848
rect 42057 411843 42123 411846
rect 42609 411843 42675 411846
rect 660297 411906 660363 411909
rect 683297 411906 683363 411909
rect 660297 411904 683363 411906
rect 660297 411848 660302 411904
rect 660358 411848 683302 411904
rect 683358 411848 683363 411904
rect 660297 411846 683363 411848
rect 660297 411843 660363 411846
rect 683297 411843 683363 411846
rect 675334 410484 675340 410548
rect 675404 410546 675410 410548
rect 676029 410546 676095 410549
rect 675404 410544 676095 410546
rect 675404 410488 676034 410544
rect 676090 410488 676095 410544
rect 675404 410486 676095 410488
rect 675404 410484 675410 410486
rect 676029 410483 676095 410486
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 42977 407826 43043 407829
rect 42425 407824 43043 407826
rect 42425 407768 42430 407824
rect 42486 407768 42982 407824
rect 43038 407768 43043 407824
rect 42425 407766 43043 407768
rect 42425 407763 42491 407766
rect 42977 407763 43043 407766
rect 42425 407146 42491 407149
rect 43161 407146 43227 407149
rect 42425 407144 43227 407146
rect 42425 407088 42430 407144
rect 42486 407088 43166 407144
rect 43222 407088 43227 407144
rect 42425 407086 43227 407088
rect 42425 407083 42491 407086
rect 43161 407083 43227 407086
rect 42425 406874 42491 406877
rect 44173 406874 44239 406877
rect 42425 406872 44239 406874
rect 42425 406816 42430 406872
rect 42486 406816 44178 406872
rect 44234 406816 44239 406872
rect 42425 406814 44239 406816
rect 42425 406811 42491 406814
rect 44173 406811 44239 406814
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669957 403746 670023 403749
rect 676262 403746 676322 403852
rect 683297 403746 683363 403749
rect 669957 403744 676322 403746
rect 669957 403688 669962 403744
rect 670018 403688 676322 403744
rect 669957 403686 676322 403688
rect 683254 403744 683363 403746
rect 683254 403688 683302 403744
rect 683358 403688 683363 403744
rect 669957 403683 670023 403686
rect 683254 403683 683363 403688
rect 683254 403444 683314 403683
rect 683113 403338 683179 403341
rect 683070 403336 683179 403338
rect 683070 403280 683118 403336
rect 683174 403280 683179 403336
rect 683070 403275 683179 403280
rect 683070 403036 683130 403275
rect 42333 402930 42399 402933
rect 45369 402930 45435 402933
rect 42333 402928 45435 402930
rect 42333 402872 42338 402928
rect 42394 402872 45374 402928
rect 45430 402872 45435 402928
rect 42333 402870 45435 402872
rect 42333 402867 42399 402870
rect 45369 402867 45435 402870
rect 676029 402658 676095 402661
rect 676029 402656 676292 402658
rect 676029 402600 676034 402656
rect 676090 402600 676292 402656
rect 676029 402598 676292 402600
rect 676029 402595 676095 402598
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674649 402250 674715 402253
rect 674649 402248 676292 402250
rect 674649 402192 674654 402248
rect 674710 402192 676292 402248
rect 674649 402190 676292 402192
rect 674649 402187 674715 402190
rect 41454 401780 41460 401844
rect 41524 401842 41530 401844
rect 41781 401842 41847 401845
rect 41524 401840 41847 401842
rect 41524 401784 41786 401840
rect 41842 401784 41847 401840
rect 41524 401782 41847 401784
rect 41524 401780 41530 401782
rect 41781 401779 41847 401782
rect 672441 401706 672507 401709
rect 676262 401706 676322 401812
rect 672441 401704 676322 401706
rect 672441 401648 672446 401704
rect 672502 401648 676322 401704
rect 672441 401646 676322 401648
rect 672441 401643 672507 401646
rect 674189 401434 674255 401437
rect 674189 401432 676292 401434
rect 674189 401376 674194 401432
rect 674250 401376 676292 401432
rect 674189 401374 676292 401376
rect 674189 401371 674255 401374
rect 676806 401236 676812 401300
rect 676876 401236 676882 401300
rect 676814 400996 676874 401236
rect 673269 400482 673335 400485
rect 676262 400482 676322 400588
rect 673269 400480 676322 400482
rect 673269 400424 673274 400480
rect 673330 400424 676322 400480
rect 673269 400422 676322 400424
rect 673269 400419 673335 400422
rect 42425 400210 42491 400213
rect 47117 400210 47183 400213
rect 42425 400208 47183 400210
rect 42425 400152 42430 400208
rect 42486 400152 47122 400208
rect 47178 400152 47183 400208
rect 42425 400150 47183 400152
rect 42425 400147 42491 400150
rect 47117 400147 47183 400150
rect 672625 400074 672691 400077
rect 676262 400074 676322 400180
rect 672625 400072 676322 400074
rect 672625 400016 672630 400072
rect 672686 400016 676322 400072
rect 672625 400014 676322 400016
rect 672625 400011 672691 400014
rect 42425 399802 42491 399805
rect 46933 399802 46999 399805
rect 42425 399800 46999 399802
rect 42425 399744 42430 399800
rect 42486 399744 46938 399800
rect 46994 399744 46999 399800
rect 42425 399742 46999 399744
rect 42425 399739 42491 399742
rect 46933 399739 46999 399742
rect 676262 399666 676322 399772
rect 674790 399606 676322 399666
rect 41781 398852 41847 398853
rect 41781 398848 41828 398852
rect 41892 398850 41898 398852
rect 672533 398850 672599 398853
rect 674790 398850 674850 399606
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41781 398792 41786 398848
rect 41781 398788 41828 398792
rect 41892 398790 41938 398850
rect 672533 398848 674850 398850
rect 672533 398792 672538 398848
rect 672594 398792 674850 398848
rect 672533 398790 674850 398792
rect 41892 398788 41898 398790
rect 41781 398787 41847 398788
rect 672533 398787 672599 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 672717 397218 672783 397221
rect 676262 397218 676322 397324
rect 672717 397216 676322 397218
rect 672717 397160 672722 397216
rect 672778 397160 676322 397216
rect 672717 397158 676322 397160
rect 672717 397155 672783 397158
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 674373 396538 674439 396541
rect 674373 396536 676292 396538
rect 674373 396480 674378 396536
rect 674434 396480 676292 396536
rect 674373 396478 676292 396480
rect 674373 396475 674439 396478
rect 674005 396130 674071 396133
rect 674005 396128 676292 396130
rect 674005 396072 674010 396128
rect 674066 396072 676292 396128
rect 674005 396070 676292 396072
rect 674005 396067 674071 396070
rect 673821 395722 673887 395725
rect 673821 395720 676292 395722
rect 673821 395664 673826 395720
rect 673882 395664 676292 395720
rect 673821 395662 676292 395664
rect 673821 395659 673887 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 674833 394498 674899 394501
rect 674833 394496 676292 394498
rect 674833 394440 674838 394496
rect 674894 394440 676292 394496
rect 674833 394438 676292 394440
rect 674833 394435 674899 394438
rect 673085 394226 673151 394229
rect 673085 394224 676322 394226
rect 673085 394168 673090 394224
rect 673146 394168 676322 394224
rect 673085 394166 676322 394168
rect 673085 394163 673151 394166
rect 676262 394060 676322 394166
rect 672901 393954 672967 393957
rect 674833 393954 674899 393957
rect 672901 393952 674899 393954
rect 672901 393896 672906 393952
rect 672962 393896 674838 393952
rect 674894 393896 674899 393952
rect 672901 393894 674899 393896
rect 672901 393891 672967 393894
rect 674833 393891 674899 393894
rect 670601 393546 670667 393549
rect 676262 393546 676322 393652
rect 670601 393544 676322 393546
rect 670601 393488 670606 393544
rect 670662 393488 676322 393544
rect 670601 393486 676322 393488
rect 670601 393483 670667 393486
rect 683070 392733 683130 393244
rect 683021 392728 683130 392733
rect 683021 392672 683026 392728
rect 683082 392672 683130 392728
rect 683021 392670 683130 392672
rect 683021 392667 683087 392670
rect 672165 392322 672231 392325
rect 676262 392322 676322 392428
rect 672165 392320 676322 392322
rect 672165 392264 672170 392320
rect 672226 392264 676322 392320
rect 672165 392262 676322 392264
rect 672165 392259 672231 392262
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 675886 388996 675892 389060
rect 675956 389058 675962 389060
rect 683021 389058 683087 389061
rect 675956 389056 683087 389058
rect 675956 389000 683026 389056
rect 683082 389000 683087 389056
rect 675956 388998 683087 389000
rect 675956 388996 675962 388998
rect 683021 388995 683087 388998
rect 41492 387638 48330 387698
rect 41270 387562 41276 387564
rect 40910 387502 41276 387562
rect 40910 387260 40970 387502
rect 41270 387500 41276 387502
rect 41340 387500 41346 387564
rect 48270 387562 48330 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 48270 387502 51090 387562
rect 41822 387228 41828 387292
rect 41892 387290 41898 387292
rect 41892 387230 49250 387290
rect 41892 387228 41898 387230
rect 41137 387154 41203 387157
rect 41094 387152 41203 387154
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387091 41203 387096
rect 41094 386852 41154 387091
rect 41873 387018 41939 387021
rect 41873 387016 48330 387018
rect 41873 386960 41878 387016
rect 41934 386960 48330 387016
rect 41873 386958 48330 386960
rect 41873 386955 41939 386958
rect 48270 386882 48330 386958
rect 48957 386882 49023 386885
rect 48270 386880 49023 386882
rect 48270 386824 48962 386880
rect 49018 386824 49023 386880
rect 48270 386822 49023 386824
rect 48957 386819 49023 386822
rect 41321 386746 41387 386749
rect 41278 386744 41387 386746
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386683 41387 386688
rect 41505 386746 41571 386749
rect 44541 386746 44607 386749
rect 41505 386744 44607 386746
rect 41505 386688 41510 386744
rect 41566 386688 44546 386744
rect 44602 386688 44607 386744
rect 41505 386686 44607 386688
rect 41505 386683 41571 386686
rect 44541 386683 44607 386686
rect 41278 386444 41338 386683
rect 49190 386474 49250 387230
rect 51030 386746 51090 387502
rect 51717 386746 51783 386749
rect 51030 386744 51783 386746
rect 51030 386688 51722 386744
rect 51778 386688 51783 386744
rect 51030 386686 51783 386688
rect 51717 386683 51783 386686
rect 51901 386474 51967 386477
rect 49190 386472 51967 386474
rect 49190 386416 51906 386472
rect 51962 386416 51967 386472
rect 49190 386414 51967 386416
rect 51901 386411 51967 386414
rect 44633 386066 44699 386069
rect 41492 386064 44699 386066
rect 41492 386008 44638 386064
rect 44694 386008 44699 386064
rect 41492 386006 44699 386008
rect 44633 386003 44699 386006
rect 45093 385658 45159 385661
rect 41492 385656 45159 385658
rect 41492 385600 45098 385656
rect 45154 385600 45159 385656
rect 41492 385598 45159 385600
rect 45093 385595 45159 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 44357 384842 44423 384845
rect 41492 384840 44423 384842
rect 41492 384784 44362 384840
rect 44418 384784 44423 384840
rect 41492 384782 44423 384784
rect 44357 384779 44423 384782
rect 45185 384434 45251 384437
rect 41492 384432 45251 384434
rect 41492 384376 45190 384432
rect 45246 384376 45251 384432
rect 41492 384374 45251 384376
rect 45185 384371 45251 384374
rect 45369 384026 45435 384029
rect 41492 384024 45435 384026
rect 41492 383968 45374 384024
rect 45430 383968 45435 384024
rect 41492 383966 45435 383968
rect 45369 383963 45435 383966
rect 45185 383618 45251 383621
rect 41492 383616 45251 383618
rect 41492 383560 45190 383616
rect 45246 383560 45251 383616
rect 41492 383558 45251 383560
rect 45185 383555 45251 383558
rect 41278 383077 41338 383180
rect 41278 383072 41387 383077
rect 41278 383016 41326 383072
rect 41382 383016 41387 383072
rect 41278 383014 41387 383016
rect 41321 383011 41387 383014
rect 41094 382669 41154 382772
rect 41094 382664 41203 382669
rect 41094 382608 41142 382664
rect 41198 382608 41203 382664
rect 41094 382606 41203 382608
rect 41137 382603 41203 382606
rect 40174 382261 40234 382364
rect 40174 382256 40283 382261
rect 40174 382200 40222 382256
rect 40278 382200 40283 382256
rect 40174 382198 40283 382200
rect 40217 382195 40283 382198
rect 674373 382258 674439 382261
rect 675385 382258 675451 382261
rect 674373 382256 675451 382258
rect 674373 382200 674378 382256
rect 674434 382200 675390 382256
rect 675446 382200 675451 382256
rect 674373 382198 675451 382200
rect 674373 382195 674439 382198
rect 675385 382195 675451 382198
rect 39990 381853 40050 381956
rect 39990 381848 40099 381853
rect 39990 381792 40038 381848
rect 40094 381792 40099 381848
rect 39990 381790 40099 381792
rect 40033 381787 40099 381790
rect 41462 381442 41522 381548
rect 41638 381442 41644 381444
rect 41462 381382 41644 381442
rect 41638 381380 41644 381382
rect 41708 381380 41714 381444
rect 674005 381442 674071 381445
rect 675109 381442 675175 381445
rect 674005 381440 675175 381442
rect 674005 381384 674010 381440
rect 674066 381384 675114 381440
rect 675170 381384 675175 381440
rect 674005 381382 675175 381384
rect 674005 381379 674071 381382
rect 675109 381379 675175 381382
rect 41278 381037 41338 381140
rect 41278 381032 41387 381037
rect 41278 380976 41326 381032
rect 41382 380976 41387 381032
rect 41278 380974 41387 380976
rect 41321 380971 41387 380974
rect 46933 380762 46999 380765
rect 41492 380760 46999 380762
rect 41492 380704 46938 380760
rect 46994 380704 46999 380760
rect 41492 380702 46999 380704
rect 46933 380699 46999 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 45553 380354 45619 380357
rect 41492 380352 45619 380354
rect 41492 380296 45558 380352
rect 45614 380296 45619 380352
rect 41492 380294 45619 380296
rect 45553 380291 45619 380294
rect 44449 379946 44515 379949
rect 41492 379944 44515 379946
rect 41492 379888 44454 379944
rect 44510 379888 44515 379944
rect 41492 379886 44515 379888
rect 44449 379883 44515 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 41689 379402 41755 379405
rect 42977 379402 43043 379405
rect 41689 379400 43043 379402
rect 41689 379344 41694 379400
rect 41750 379344 42982 379400
rect 43038 379344 43043 379400
rect 41689 379342 43043 379344
rect 41689 379339 41755 379342
rect 42977 379339 43043 379342
rect 47117 379130 47183 379133
rect 41492 379128 47183 379130
rect 41492 379072 47122 379128
rect 47178 379072 47183 379128
rect 41492 379070 47183 379072
rect 47117 379067 47183 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 41321 378586 41387 378589
rect 42333 378586 42399 378589
rect 41321 378584 42399 378586
rect 41321 378528 41326 378584
rect 41382 378528 42338 378584
rect 42394 378528 42399 378584
rect 41321 378526 42399 378528
rect 41321 378523 41387 378526
rect 42333 378523 42399 378526
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 673453 378178 673519 378181
rect 650164 378176 673519 378178
rect 650164 378120 673458 378176
rect 673514 378120 673519 378176
rect 650164 378118 673519 378120
rect 673453 378115 673519 378118
rect 675109 378042 675175 378045
rect 676070 378042 676076 378044
rect 675109 378040 676076 378042
rect 675109 377984 675114 378040
rect 675170 377984 676076 378040
rect 675109 377982 676076 377984
rect 675109 377979 675175 377982
rect 676070 377980 676076 377982
rect 676140 377980 676146 378044
rect 672717 377906 672783 377909
rect 674782 377906 674788 377908
rect 672717 377904 674788 377906
rect 40910 377772 40970 377876
rect 672717 377848 672722 377904
rect 672778 377848 674788 377904
rect 672717 377846 674788 377848
rect 672717 377843 672783 377846
rect 674782 377844 674788 377846
rect 674852 377844 674858 377908
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 35758 376549 35818 377060
rect 40217 376954 40283 376957
rect 41454 376954 41460 376956
rect 40217 376952 41460 376954
rect 40217 376896 40222 376952
rect 40278 376896 41460 376952
rect 40217 376894 41460 376896
rect 40217 376891 40283 376894
rect 41454 376892 41460 376894
rect 41524 376892 41530 376956
rect 672901 376954 672967 376957
rect 675293 376954 675359 376957
rect 672901 376952 675359 376954
rect 672901 376896 672906 376952
rect 672962 376896 675298 376952
rect 675354 376896 675359 376952
rect 672901 376894 675359 376896
rect 672901 376891 672967 376894
rect 675293 376891 675359 376894
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 40033 376546 40099 376549
rect 42006 376546 42012 376548
rect 40033 376544 42012 376546
rect 40033 376488 40038 376544
rect 40094 376488 42012 376544
rect 40033 376486 42012 376488
rect 40033 376483 40099 376486
rect 42006 376484 42012 376486
rect 42076 376484 42082 376548
rect 62113 376274 62179 376277
rect 673085 376274 673151 376277
rect 675385 376274 675451 376277
rect 62113 376272 64492 376274
rect 28950 376141 29010 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 673085 376272 675451 376274
rect 673085 376216 673090 376272
rect 673146 376216 675390 376272
rect 675446 376216 675451 376272
rect 673085 376214 675451 376216
rect 62113 376211 62179 376214
rect 673085 376211 673151 376214
rect 675385 376211 675451 376214
rect 28901 376136 29010 376141
rect 28901 376080 28906 376136
rect 28962 376080 29010 376136
rect 28901 376078 29010 376080
rect 28901 376075 28967 376078
rect 39573 375730 39639 375733
rect 40350 375730 40356 375732
rect 39573 375728 40356 375730
rect 39573 375672 39578 375728
rect 39634 375672 40356 375728
rect 39573 375670 40356 375672
rect 39573 375667 39639 375670
rect 40350 375668 40356 375670
rect 40420 375668 40426 375732
rect 673821 375458 673887 375461
rect 675293 375458 675359 375461
rect 673821 375456 675359 375458
rect 673821 375400 673826 375456
rect 673882 375400 675298 375456
rect 675354 375400 675359 375456
rect 673821 375398 675359 375400
rect 673821 375395 673887 375398
rect 675293 375395 675359 375398
rect 675661 373010 675727 373013
rect 675886 373010 675892 373012
rect 675661 373008 675892 373010
rect 675661 372952 675666 373008
rect 675722 372952 675892 373008
rect 675661 372950 675892 372952
rect 675661 372947 675727 372950
rect 675886 372948 675892 372950
rect 675956 372948 675962 373012
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 41689 371922 41755 371925
rect 43345 371922 43411 371925
rect 41689 371920 43411 371922
rect 41689 371864 41694 371920
rect 41750 371864 43350 371920
rect 43406 371864 43411 371920
rect 41689 371862 43411 371864
rect 41689 371859 41755 371862
rect 43345 371859 43411 371862
rect 40350 368596 40356 368660
rect 40420 368658 40426 368660
rect 41781 368658 41847 368661
rect 40420 368656 41847 368658
rect 40420 368600 41786 368656
rect 41842 368600 41847 368656
rect 40420 368598 41847 368600
rect 40420 368596 40426 368598
rect 41781 368595 41847 368598
rect 42425 367026 42491 367029
rect 46197 367026 46263 367029
rect 42425 367024 46263 367026
rect 42425 366968 42430 367024
rect 42486 366968 46202 367024
rect 46258 366968 46263 367024
rect 42425 366966 46263 366968
rect 42425 366963 42491 366966
rect 46197 366963 46263 366966
rect 42425 365802 42491 365805
rect 42977 365802 43043 365805
rect 42425 365800 43043 365802
rect 42425 365744 42430 365800
rect 42486 365744 42982 365800
rect 43038 365744 43043 365800
rect 42425 365742 43043 365744
rect 42425 365739 42491 365742
rect 42977 365739 43043 365742
rect 651833 364850 651899 364853
rect 650164 364848 651899 364850
rect 650164 364792 651838 364848
rect 651894 364792 651899 364848
rect 650164 364790 651899 364792
rect 651833 364787 651899 364790
rect 40902 364244 40908 364308
rect 40972 364306 40978 364308
rect 41781 364306 41847 364309
rect 40972 364304 41847 364306
rect 40972 364248 41786 364304
rect 41842 364248 41847 364304
rect 40972 364246 41847 364248
rect 40972 364244 40978 364246
rect 41781 364243 41847 364246
rect 40718 363564 40724 363628
rect 40788 363626 40794 363628
rect 41781 363626 41847 363629
rect 40788 363624 41847 363626
rect 40788 363568 41786 363624
rect 41842 363568 41847 363624
rect 40788 363566 41847 363568
rect 40788 363564 40794 363566
rect 41781 363563 41847 363566
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 41873 362948 41939 362949
rect 41822 362946 41828 362948
rect 41782 362886 41828 362946
rect 41892 362944 41939 362948
rect 41934 362888 41939 362944
rect 41822 362884 41828 362886
rect 41892 362884 41939 362888
rect 41873 362883 41939 362884
rect 42425 361586 42491 361589
rect 47117 361586 47183 361589
rect 42425 361584 47183 361586
rect 42425 361528 42430 361584
rect 42486 361528 47122 361584
rect 47178 361528 47183 361584
rect 42425 361526 47183 361528
rect 42425 361523 42491 361526
rect 47117 361523 47183 361526
rect 667197 360906 667263 360909
rect 675845 360906 675911 360909
rect 667197 360904 675911 360906
rect 667197 360848 667202 360904
rect 667258 360848 675850 360904
rect 675906 360848 675911 360904
rect 667197 360846 675911 360848
rect 667197 360843 667263 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 42149 359954 42215 359957
rect 44449 359954 44515 359957
rect 42149 359952 44515 359954
rect 42149 359896 42154 359952
rect 42210 359896 44454 359952
rect 44510 359896 44515 359952
rect 42149 359894 44515 359896
rect 42149 359891 42215 359894
rect 44449 359891 44515 359894
rect 42057 358732 42123 358733
rect 42006 358730 42012 358732
rect 41966 358670 42012 358730
rect 42076 358728 42123 358732
rect 42118 358672 42123 358728
rect 42006 358668 42012 358670
rect 42076 358668 42123 358672
rect 42057 358667 42123 358668
rect 663750 358670 676292 358730
rect 663241 358594 663307 358597
rect 663750 358594 663810 358670
rect 663241 358592 663810 358594
rect 663241 358536 663246 358592
rect 663302 358536 663810 358592
rect 663241 358534 663810 358536
rect 663241 358531 663307 358534
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 674649 357506 674715 357509
rect 674649 357504 676292 357506
rect 674649 357448 674654 357504
rect 674710 357448 676292 357504
rect 674649 357446 676292 357448
rect 674649 357443 674715 357446
rect 42425 357370 42491 357373
rect 45553 357370 45619 357373
rect 42425 357368 45619 357370
rect 42425 357312 42430 357368
rect 42486 357312 45558 357368
rect 45614 357312 45619 357368
rect 42425 357310 45619 357312
rect 42425 357307 42491 357310
rect 45553 357307 45619 357310
rect 672717 357098 672783 357101
rect 672717 357096 676292 357098
rect 672717 357040 672722 357096
rect 672778 357040 676292 357096
rect 672717 357038 676292 357040
rect 672717 357035 672783 357038
rect 44265 356690 44331 356693
rect 45645 356690 45711 356693
rect 44265 356688 45711 356690
rect 44265 356632 44270 356688
rect 44326 356632 45650 356688
rect 45706 356632 45711 356688
rect 44265 356630 45711 356632
rect 44265 356627 44331 356630
rect 45645 356627 45711 356630
rect 674189 356690 674255 356693
rect 674189 356688 676292 356690
rect 674189 356632 674194 356688
rect 674250 356632 676292 356688
rect 674189 356630 676292 356632
rect 674189 356627 674255 356630
rect 674189 356282 674255 356285
rect 674189 356280 676292 356282
rect 674189 356224 674194 356280
rect 674250 356224 676292 356280
rect 674189 356222 676292 356224
rect 674189 356219 674255 356222
rect 42425 356146 42491 356149
rect 46933 356146 46999 356149
rect 42425 356144 46999 356146
rect 42425 356088 42430 356144
rect 42486 356088 46938 356144
rect 46994 356088 46999 356144
rect 42425 356086 46999 356088
rect 42425 356083 42491 356086
rect 46933 356083 46999 356086
rect 43345 355874 43411 355877
rect 45921 355874 45987 355877
rect 43345 355872 45987 355874
rect 43345 355816 43350 355872
rect 43406 355816 45926 355872
rect 45982 355816 45987 355872
rect 43345 355814 45987 355816
rect 43345 355811 43411 355814
rect 45921 355811 45987 355814
rect 673269 355874 673335 355877
rect 673269 355872 676292 355874
rect 673269 355816 673274 355872
rect 673330 355816 676292 355872
rect 673269 355814 676292 355816
rect 673269 355811 673335 355814
rect 41454 355676 41460 355740
rect 41524 355738 41530 355740
rect 41781 355738 41847 355741
rect 41524 355736 41847 355738
rect 41524 355680 41786 355736
rect 41842 355680 41847 355736
rect 41524 355678 41847 355680
rect 41524 355676 41530 355678
rect 41781 355675 41847 355678
rect 673269 355466 673335 355469
rect 673269 355464 676292 355466
rect 673269 355408 673274 355464
rect 673330 355408 676292 355464
rect 673269 355406 676292 355408
rect 673269 355403 673335 355406
rect 672533 355058 672599 355061
rect 672533 355056 676292 355058
rect 672533 355000 672538 355056
rect 672594 355000 676292 355056
rect 672533 354998 676292 355000
rect 672533 354995 672599 354998
rect 673085 354650 673151 354653
rect 673085 354648 676292 354650
rect 673085 354592 673090 354648
rect 673146 354592 676292 354648
rect 673085 354590 676292 354592
rect 673085 354587 673151 354590
rect 43897 354244 43963 354245
rect 43846 354180 43852 354244
rect 43916 354242 43963 354244
rect 43916 354240 44008 354242
rect 43958 354184 44008 354240
rect 43916 354182 44008 354184
rect 43916 354180 43963 354182
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 43897 354179 43963 354180
rect 44214 353772 44220 353836
rect 44284 353834 44290 353836
rect 44725 353834 44791 353837
rect 44284 353832 44791 353834
rect 44284 353776 44730 353832
rect 44786 353776 44791 353832
rect 44284 353774 44791 353776
rect 44284 353772 44290 353774
rect 44725 353771 44791 353774
rect 675702 353772 675708 353836
rect 675772 353834 675778 353836
rect 675772 353774 676292 353834
rect 675772 353772 675778 353774
rect 673637 353426 673703 353429
rect 673637 353424 676292 353426
rect 673637 353368 673642 353424
rect 673698 353368 676292 353424
rect 673637 353366 676292 353368
rect 673637 353363 673703 353366
rect 675334 352956 675340 353020
rect 675404 353018 675410 353020
rect 675404 352958 676292 353018
rect 675404 352956 675410 352958
rect 672901 352610 672967 352613
rect 672901 352608 676292 352610
rect 672901 352552 672906 352608
rect 672962 352552 676292 352608
rect 672901 352550 676292 352552
rect 672901 352547 672967 352550
rect 672533 352202 672599 352205
rect 672533 352200 676292 352202
rect 672533 352144 672538 352200
rect 672594 352144 676292 352200
rect 672533 352142 676292 352144
rect 672533 352139 672599 352142
rect 675845 351794 675911 351797
rect 675845 351792 676292 351794
rect 675845 351736 675850 351792
rect 675906 351736 676292 351792
rect 675845 351734 676292 351736
rect 675845 351731 675911 351734
rect 652385 351658 652451 351661
rect 650164 351656 652451 351658
rect 650164 351600 652390 351656
rect 652446 351600 652451 351656
rect 650164 351598 652451 351600
rect 652385 351595 652451 351598
rect 674741 351386 674807 351389
rect 674741 351384 676292 351386
rect 674741 351328 674746 351384
rect 674802 351328 676292 351384
rect 674741 351326 676292 351328
rect 674741 351323 674807 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 673821 350570 673887 350573
rect 673821 350568 676292 350570
rect 673821 350512 673826 350568
rect 673882 350512 676292 350568
rect 673821 350510 676292 350512
rect 673821 350507 673887 350510
rect 62757 350298 62823 350301
rect 675845 350300 675911 350301
rect 675845 350298 675892 350300
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 675800 350296 675892 350298
rect 675800 350240 675850 350296
rect 675800 350238 675892 350240
rect 62757 350235 62823 350238
rect 675845 350236 675892 350238
rect 675956 350236 675962 350300
rect 675845 350235 675911 350236
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 672349 349754 672415 349757
rect 672349 349752 676292 349754
rect 672349 349696 672354 349752
rect 672410 349696 676292 349752
rect 672349 349694 676292 349696
rect 672349 349691 672415 349694
rect 674005 349482 674071 349485
rect 674005 349480 676230 349482
rect 674005 349424 674010 349480
rect 674066 349424 676230 349480
rect 674005 349422 676230 349424
rect 674005 349419 674071 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 671981 348938 672047 348941
rect 671981 348936 676292 348938
rect 671981 348880 671986 348936
rect 672042 348880 676292 348936
rect 671981 348878 676292 348880
rect 671981 348875 672047 348878
rect 673862 348468 673868 348532
rect 673932 348530 673938 348532
rect 673932 348470 676292 348530
rect 673932 348468 673938 348470
rect 674557 347714 674623 347717
rect 683070 347714 683130 348092
rect 674557 347712 683130 347714
rect 674557 347656 674562 347712
rect 674618 347684 683130 347712
rect 674618 347656 683100 347684
rect 674557 347654 683100 347656
rect 674557 347651 674623 347654
rect 670417 347306 670483 347309
rect 670417 347304 676292 347306
rect 670417 347248 670422 347304
rect 670478 347248 676292 347304
rect 670417 347246 676292 347248
rect 670417 347243 670483 347246
rect 676029 346626 676095 346629
rect 676622 346626 676628 346628
rect 676029 346624 676628 346626
rect 676029 346568 676034 346624
rect 676090 346568 676628 346624
rect 676029 346566 676628 346568
rect 676029 346563 676095 346566
rect 676622 346564 676628 346566
rect 676692 346564 676698 346628
rect 62941 345674 63007 345677
rect 45510 345672 63007 345674
rect 45510 345616 62946 345672
rect 63002 345616 63007 345672
rect 45510 345614 63007 345616
rect 40217 345538 40283 345541
rect 45510 345538 45570 345614
rect 62941 345611 63007 345614
rect 40217 345536 45570 345538
rect 40217 345480 40222 345536
rect 40278 345480 45570 345536
rect 40217 345478 45570 345480
rect 40217 345475 40283 345478
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 35758 343909 35818 344148
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 35758 343904 35867 343909
rect 35758 343848 35806 343904
rect 35862 343848 35867 343904
rect 35758 343846 35867 343848
rect 35801 343843 35867 343846
rect 28582 343740 28642 343843
rect 45001 343362 45067 343365
rect 41492 343360 45067 343362
rect 41492 343304 45006 343360
rect 45062 343304 45067 343360
rect 41492 343302 45067 343304
rect 45001 343299 45067 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 44214 342682 44220 342684
rect 41462 342622 44220 342682
rect 41462 342516 41522 342622
rect 44214 342620 44220 342622
rect 44284 342620 44290 342684
rect 44398 342138 44404 342140
rect 41492 342078 44404 342138
rect 44398 342076 44404 342078
rect 44468 342076 44474 342140
rect 45369 341730 45435 341733
rect 41492 341728 45435 341730
rect 41492 341672 45374 341728
rect 45430 341672 45435 341728
rect 41492 341670 45435 341672
rect 45369 341667 45435 341670
rect 45461 341322 45527 341325
rect 41492 341320 45527 341322
rect 41492 341264 45466 341320
rect 45522 341264 45527 341320
rect 41492 341262 45527 341264
rect 45461 341259 45527 341262
rect 45185 340914 45251 340917
rect 41492 340912 45251 340914
rect 41492 340856 45190 340912
rect 45246 340856 45251 340912
rect 41492 340854 45251 340856
rect 45185 340851 45251 340854
rect 673637 340778 673703 340781
rect 675109 340778 675175 340781
rect 673637 340776 675175 340778
rect 673637 340720 673642 340776
rect 673698 340720 675114 340776
rect 675170 340720 675175 340776
rect 673637 340718 675175 340720
rect 673637 340715 673703 340718
rect 675109 340715 675175 340718
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340370 675819 340373
rect 676254 340370 676260 340372
rect 675753 340368 676260 340370
rect 675753 340312 675758 340368
rect 675814 340312 676260 340368
rect 675753 340310 676260 340312
rect 675753 340307 675819 340310
rect 676254 340308 676260 340310
rect 676324 340308 676330 340372
rect 45829 340098 45895 340101
rect 41492 340096 45895 340098
rect 41492 340040 45834 340096
rect 45890 340040 45895 340096
rect 41492 340038 45895 340040
rect 45829 340035 45895 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 675661 339418 675727 339421
rect 675886 339418 675892 339420
rect 675661 339416 675892 339418
rect 675661 339360 675666 339416
rect 675722 339360 675892 339416
rect 675661 339358 675892 339360
rect 675661 339355 675727 339358
rect 675886 339356 675892 339358
rect 675956 339356 675962 339420
rect 45645 339282 45711 339285
rect 41492 339280 45711 339282
rect 41492 339224 45650 339280
rect 45706 339224 45711 339280
rect 41492 339222 45711 339224
rect 45645 339219 45711 339222
rect 46013 338874 46079 338877
rect 41492 338872 46079 338874
rect 41492 338816 46018 338872
rect 46074 338816 46079 338872
rect 41492 338814 46079 338816
rect 46013 338811 46079 338814
rect 41462 338196 41522 338436
rect 652017 338330 652083 338333
rect 650164 338328 652083 338330
rect 650164 338272 652022 338328
rect 652078 338272 652083 338328
rect 650164 338270 652083 338272
rect 652017 338267 652083 338270
rect 41454 338132 41460 338196
rect 41524 338132 41530 338196
rect 41278 337786 41338 338028
rect 41822 337786 41828 337788
rect 41278 337726 41828 337786
rect 41822 337724 41828 337726
rect 41892 337724 41898 337788
rect 41462 337378 41522 337620
rect 42926 337378 42932 337380
rect 41462 337318 42932 337378
rect 42926 337316 42932 337318
rect 42996 337316 43002 337380
rect 62113 337242 62179 337245
rect 675385 337244 675451 337245
rect 675334 337242 675340 337244
rect 62113 337240 64492 337242
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 41278 336970 41338 337212
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 675294 337182 675340 337242
rect 675404 337240 675451 337244
rect 675446 337184 675451 337240
rect 62113 337179 62179 337182
rect 675334 337180 675340 337182
rect 675404 337180 675451 337184
rect 675385 337179 675451 337180
rect 43110 336970 43116 336972
rect 41278 336910 43116 336970
rect 43110 336908 43116 336910
rect 43180 336908 43186 336972
rect 40542 336804 40602 336908
rect 36629 336562 36695 336565
rect 41638 336562 41644 336564
rect 36629 336560 41644 336562
rect 36629 336504 36634 336560
rect 36690 336504 41644 336560
rect 36629 336502 41644 336504
rect 36629 336499 36695 336502
rect 41638 336500 41644 336502
rect 41708 336500 41714 336564
rect 675753 336562 675819 336565
rect 676438 336562 676444 336564
rect 675753 336560 676444 336562
rect 675753 336504 675758 336560
rect 675814 336504 676444 336560
rect 675753 336502 676444 336504
rect 675753 336499 675819 336502
rect 676438 336500 676444 336502
rect 676508 336500 676514 336564
rect 41462 336154 41522 336396
rect 41462 336094 43178 336154
rect 41462 335746 41522 335988
rect 42742 335746 42748 335748
rect 41462 335686 42748 335746
rect 42742 335684 42748 335686
rect 42812 335684 42818 335748
rect 40726 335340 40786 335580
rect 40718 335276 40724 335340
rect 40788 335276 40794 335340
rect 41462 334930 41522 335172
rect 41462 334870 41844 334930
rect 41278 334522 41338 334764
rect 41784 334658 41844 334870
rect 43118 334661 43178 336094
rect 672533 335882 672599 335885
rect 674782 335882 674788 335884
rect 672533 335880 674788 335882
rect 672533 335824 672538 335880
rect 672594 335824 674788 335880
rect 672533 335822 674788 335824
rect 672533 335819 672599 335822
rect 674782 335820 674788 335822
rect 674852 335820 674858 335884
rect 672349 335610 672415 335613
rect 675109 335610 675175 335613
rect 672349 335608 675175 335610
rect 672349 335552 672354 335608
rect 672410 335552 675114 335608
rect 675170 335552 675175 335608
rect 672349 335550 675175 335552
rect 672349 335547 672415 335550
rect 675109 335547 675175 335550
rect 42793 334658 42859 334661
rect 41784 334656 42859 334658
rect 41784 334600 42798 334656
rect 42854 334600 42859 334656
rect 41784 334598 42859 334600
rect 42793 334595 42859 334598
rect 43069 334656 43178 334661
rect 43069 334600 43074 334656
rect 43130 334600 43178 334656
rect 43069 334598 43178 334600
rect 43069 334595 43135 334598
rect 41597 334522 41663 334525
rect 41278 334520 41663 334522
rect 41278 334464 41602 334520
rect 41658 334464 41663 334520
rect 41278 334462 41663 334464
rect 41597 334459 41663 334462
rect 41462 334114 41522 334356
rect 42742 334324 42748 334388
rect 42812 334386 42818 334388
rect 44173 334386 44239 334389
rect 42812 334384 44239 334386
rect 42812 334328 44178 334384
rect 44234 334328 44239 334384
rect 42812 334326 44239 334328
rect 42812 334324 42818 334326
rect 44173 334323 44239 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 672901 333978 672967 333981
rect 675109 333978 675175 333981
rect 672901 333976 675175 333978
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 672901 333920 672906 333976
rect 672962 333920 675114 333976
rect 675170 333920 675175 333976
rect 672901 333918 675175 333920
rect 672901 333915 672967 333918
rect 675109 333915 675175 333918
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 41597 333706 41663 333709
rect 43253 333706 43319 333709
rect 41597 333704 43319 333706
rect 41597 333648 41602 333704
rect 41658 333648 43258 333704
rect 43314 333648 43319 333704
rect 41597 333646 43319 333648
rect 41597 333643 41663 333646
rect 43253 333643 43319 333646
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 674005 332754 674071 332757
rect 675109 332754 675175 332757
rect 674005 332752 675175 332754
rect 674005 332696 674010 332752
rect 674066 332696 675114 332752
rect 675170 332696 675175 332752
rect 674005 332694 675175 332696
rect 674005 332691 674071 332694
rect 675109 332691 675175 332694
rect 675753 332346 675819 332349
rect 676622 332346 676628 332348
rect 675753 332344 676628 332346
rect 675753 332288 675758 332344
rect 675814 332288 676628 332344
rect 675753 332286 676628 332288
rect 675753 332283 675819 332286
rect 676622 332284 676628 332286
rect 676692 332284 676698 332348
rect 673821 331122 673887 331125
rect 675293 331122 675359 331125
rect 673821 331120 675359 331122
rect 673821 331064 673826 331120
rect 673882 331064 675298 331120
rect 675354 331064 675359 331120
rect 673821 331062 675359 331064
rect 673821 331059 673887 331062
rect 675293 331059 675359 331062
rect 671981 329762 672047 329765
rect 675109 329762 675175 329765
rect 671981 329760 675175 329762
rect 671981 329704 671986 329760
rect 672042 329704 675114 329760
rect 675170 329704 675175 329760
rect 671981 329702 675175 329704
rect 671981 329699 672047 329702
rect 675109 329699 675175 329702
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 674782 326844 674788 326908
rect 674852 326906 674858 326908
rect 675385 326906 675451 326909
rect 674852 326904 675451 326906
rect 674852 326848 675390 326904
rect 675446 326848 675451 326904
rect 674852 326846 675451 326848
rect 674852 326844 674858 326846
rect 675385 326843 675451 326846
rect 41781 326772 41847 326773
rect 41781 326768 41828 326772
rect 41892 326770 41898 326772
rect 41781 326712 41786 326768
rect 41781 326708 41828 326712
rect 41892 326710 41938 326770
rect 41892 326708 41898 326710
rect 41781 326707 41847 326708
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41873 324868 41939 324869
rect 41822 324866 41828 324868
rect 41782 324806 41828 324866
rect 41892 324864 41939 324868
rect 41934 324808 41939 324864
rect 41822 324804 41828 324806
rect 41892 324804 41939 324808
rect 41873 324803 41939 324804
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 42057 322826 42123 322829
rect 43069 322826 43135 322829
rect 42057 322824 43135 322826
rect 42057 322768 42062 322824
rect 42118 322768 43074 322824
rect 43130 322768 43135 322824
rect 42057 322766 43135 322768
rect 42057 322763 42123 322766
rect 43069 322763 43135 322766
rect 42517 321466 42583 321469
rect 53097 321466 53163 321469
rect 42517 321464 53163 321466
rect 42517 321408 42522 321464
rect 42578 321408 53102 321464
rect 53158 321408 53163 321464
rect 42517 321406 53163 321408
rect 42517 321403 42583 321406
rect 53097 321403 53163 321406
rect 42241 321194 42307 321197
rect 43253 321194 43319 321197
rect 42241 321192 43319 321194
rect 42241 321136 42246 321192
rect 42302 321136 43258 321192
rect 43314 321136 43319 321192
rect 42241 321134 43319 321136
rect 42241 321131 42307 321134
rect 43253 321131 43319 321134
rect 42425 320922 42491 320925
rect 44173 320922 44239 320925
rect 42425 320920 44239 320922
rect 42425 320864 42430 320920
rect 42486 320864 44178 320920
rect 44234 320864 44239 320920
rect 42425 320862 44239 320864
rect 42425 320859 42491 320862
rect 44173 320859 44239 320862
rect 41454 319908 41460 319972
rect 41524 319970 41530 319972
rect 41781 319970 41847 319973
rect 41524 319968 41847 319970
rect 41524 319912 41786 319968
rect 41842 319912 41847 319968
rect 41524 319910 41847 319912
rect 41524 319908 41530 319910
rect 41781 319907 41847 319910
rect 40718 317460 40724 317524
rect 40788 317522 40794 317524
rect 42241 317522 42307 317525
rect 40788 317520 42307 317522
rect 40788 317464 42246 317520
rect 42302 317464 42307 317520
rect 40788 317462 42307 317464
rect 40788 317460 40794 317462
rect 42241 317459 42307 317462
rect 40534 316644 40540 316708
rect 40604 316706 40610 316708
rect 41781 316706 41847 316709
rect 40604 316704 41847 316706
rect 40604 316648 41786 316704
rect 41842 316648 41847 316704
rect 40604 316646 41847 316648
rect 40604 316644 40610 316646
rect 41781 316643 41847 316646
rect 42149 316026 42215 316029
rect 43110 316026 43116 316028
rect 42149 316024 43116 316026
rect 42149 315968 42154 316024
rect 42210 315968 43116 316024
rect 42149 315966 43116 315968
rect 42149 315963 42215 315966
rect 43110 315964 43116 315966
rect 43180 315964 43186 316028
rect 42149 315482 42215 315485
rect 46013 315482 46079 315485
rect 42149 315480 46079 315482
rect 42149 315424 42154 315480
rect 42210 315424 46018 315480
rect 46074 315424 46079 315480
rect 42149 315422 46079 315424
rect 42149 315419 42215 315422
rect 46013 315419 46079 315422
rect 665817 315482 665883 315485
rect 676029 315482 676095 315485
rect 665817 315480 676095 315482
rect 665817 315424 665822 315480
rect 665878 315424 676034 315480
rect 676090 315424 676095 315480
rect 665817 315422 676095 315424
rect 665817 315419 665883 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 45829 313714 45895 313717
rect 42149 313712 45895 313714
rect 42149 313656 42154 313712
rect 42210 313656 45834 313712
rect 45890 313656 45895 313712
rect 42149 313654 45895 313656
rect 42149 313651 42215 313654
rect 45829 313651 45895 313654
rect 663750 313654 676292 313714
rect 661677 313578 661743 313581
rect 663750 313578 663810 313654
rect 661677 313576 663810 313578
rect 661677 313520 661682 313576
rect 661738 313520 663810 313576
rect 661677 313518 663810 313520
rect 661677 313515 661743 313518
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 674649 313034 674715 313037
rect 674649 313032 675034 313034
rect 674649 312976 674654 313032
rect 674710 312976 675034 313032
rect 674649 312974 675034 312976
rect 674649 312971 674715 312974
rect 674974 312898 675034 312974
rect 674974 312838 676292 312898
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 672901 312762 672967 312765
rect 674833 312762 674899 312765
rect 672901 312760 674899 312762
rect 672901 312704 672906 312760
rect 672962 312704 674838 312760
rect 674894 312704 674899 312760
rect 672901 312702 674899 312704
rect 672901 312699 672967 312702
rect 674833 312699 674899 312702
rect 672717 312490 672783 312493
rect 672717 312488 676292 312490
rect 672717 312432 672722 312488
rect 672778 312432 676292 312488
rect 672717 312430 676292 312432
rect 672717 312427 672783 312430
rect 42149 312354 42215 312357
rect 45645 312354 45711 312357
rect 42149 312352 45711 312354
rect 42149 312296 42154 312352
rect 42210 312296 45650 312352
rect 45706 312296 45711 312352
rect 42149 312294 45711 312296
rect 42149 312291 42215 312294
rect 45645 312291 45711 312294
rect 674833 312082 674899 312085
rect 674833 312080 676292 312082
rect 674833 312024 674838 312080
rect 674894 312024 676292 312080
rect 674833 312022 676292 312024
rect 674833 312019 674899 312022
rect 668577 311946 668643 311949
rect 674649 311946 674715 311949
rect 668577 311944 674715 311946
rect 668577 311888 668582 311944
rect 668638 311888 674654 311944
rect 674710 311888 674715 311944
rect 668577 311886 674715 311888
rect 668577 311883 668643 311886
rect 674649 311883 674715 311886
rect 651465 311810 651531 311813
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 651465 311747 651531 311750
rect 674189 311674 674255 311677
rect 674189 311672 676292 311674
rect 674189 311616 674194 311672
rect 674250 311616 676292 311672
rect 674189 311614 676292 311616
rect 674189 311611 674255 311614
rect 44214 311476 44220 311540
rect 44284 311538 44290 311540
rect 44541 311538 44607 311541
rect 44284 311536 44607 311538
rect 44284 311480 44546 311536
rect 44602 311480 44607 311536
rect 44284 311478 44607 311480
rect 44284 311476 44290 311478
rect 44541 311475 44607 311478
rect 44357 311268 44423 311269
rect 44357 311266 44404 311268
rect 44312 311264 44404 311266
rect 44312 311208 44362 311264
rect 44312 311206 44404 311208
rect 44357 311204 44404 311206
rect 44468 311204 44474 311268
rect 674649 311266 674715 311269
rect 674649 311264 676292 311266
rect 674649 311208 674654 311264
rect 674710 311208 676292 311264
rect 674649 311206 676292 311208
rect 44357 311203 44423 311204
rect 674649 311203 674715 311206
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 62113 311067 62179 311070
rect 673269 310858 673335 310861
rect 673269 310856 676292 310858
rect 673269 310800 673274 310856
rect 673330 310800 676292 310856
rect 673269 310798 676292 310800
rect 673269 310795 673335 310798
rect 674281 310450 674347 310453
rect 674281 310448 676292 310450
rect 674281 310392 674286 310448
rect 674342 310392 676292 310448
rect 674281 310390 676292 310392
rect 674281 310387 674347 310390
rect 673085 310042 673151 310045
rect 673085 310040 676292 310042
rect 673085 309984 673090 310040
rect 673146 309984 676292 310040
rect 673085 309982 676292 309984
rect 673085 309979 673151 309982
rect 673085 309634 673151 309637
rect 673085 309632 676292 309634
rect 673085 309576 673090 309632
rect 673146 309576 676292 309632
rect 673085 309574 676292 309576
rect 673085 309571 673151 309574
rect 675017 309226 675083 309229
rect 675017 309224 676292 309226
rect 675017 309168 675022 309224
rect 675078 309168 676292 309224
rect 675017 309166 676292 309168
rect 675017 309163 675083 309166
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 674833 308002 674899 308005
rect 674833 308000 676292 308002
rect 674833 307944 674838 308000
rect 674894 307944 676292 308000
rect 674833 307942 676292 307944
rect 674833 307939 674899 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 675886 306716 675892 306780
rect 675956 306778 675962 306780
rect 675956 306718 676292 306778
rect 675956 306716 675962 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 675886 305900 675892 305964
rect 675956 305962 675962 305964
rect 675956 305902 676292 305962
rect 675956 305900 675962 305902
rect 674097 305554 674163 305557
rect 674097 305552 676292 305554
rect 674097 305496 674102 305552
rect 674158 305496 676292 305552
rect 674097 305494 676292 305496
rect 674097 305491 674163 305494
rect 676024 305084 676030 305148
rect 676094 305146 676100 305148
rect 676094 305086 676292 305146
rect 676094 305084 676100 305086
rect 672441 304738 672507 304741
rect 672441 304736 676292 304738
rect 672441 304680 672446 304736
rect 672502 304680 676292 304736
rect 672441 304678 676292 304680
rect 672441 304675 672507 304678
rect 672625 304330 672691 304333
rect 672625 304328 676292 304330
rect 672625 304272 672630 304328
rect 672686 304272 676292 304328
rect 672625 304270 676292 304272
rect 672625 304267 672691 304270
rect 674465 303922 674531 303925
rect 674465 303920 676292 303922
rect 674465 303864 674470 303920
rect 674526 303864 676292 303920
rect 674465 303862 676292 303864
rect 674465 303859 674531 303862
rect 673269 303514 673335 303517
rect 673269 303512 676292 303514
rect 673269 303456 673274 303512
rect 673330 303456 676292 303512
rect 673269 303454 676292 303456
rect 673269 303451 673335 303454
rect 41781 303106 41847 303109
rect 46381 303106 46447 303109
rect 41781 303104 46447 303106
rect 41781 303048 41786 303104
rect 41842 303048 46386 303104
rect 46442 303048 46447 303104
rect 41781 303046 46447 303048
rect 41781 303043 41847 303046
rect 46381 303043 46447 303046
rect 683070 302701 683130 303076
rect 683021 302696 683130 302701
rect 683021 302640 683026 302696
rect 683082 302668 683130 302696
rect 683082 302640 683100 302668
rect 683021 302638 683100 302640
rect 683021 302635 683087 302638
rect 669221 302290 669287 302293
rect 669221 302288 676292 302290
rect 669221 302232 669226 302288
rect 669282 302232 676292 302288
rect 669221 302230 676292 302232
rect 669221 302227 669287 302230
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44541 300114 44607 300117
rect 41492 300112 44607 300114
rect 41492 300056 44546 300112
rect 44602 300056 44607 300112
rect 41492 300054 44607 300056
rect 44541 300051 44607 300054
rect 44633 299706 44699 299709
rect 41492 299704 44699 299706
rect 41492 299648 44638 299704
rect 44694 299648 44699 299704
rect 41492 299646 44699 299648
rect 44633 299643 44699 299646
rect 675702 299372 675708 299436
rect 675772 299434 675778 299436
rect 683021 299434 683087 299437
rect 675772 299432 683087 299434
rect 675772 299376 683026 299432
rect 683082 299376 683087 299432
rect 675772 299374 683087 299376
rect 675772 299372 675778 299374
rect 683021 299371 683087 299374
rect 44357 299298 44423 299301
rect 41492 299296 44423 299298
rect 41492 299240 44362 299296
rect 44418 299240 44423 299296
rect 41492 299238 44423 299240
rect 44357 299235 44423 299238
rect 45185 298890 45251 298893
rect 41492 298888 45251 298890
rect 41492 298832 45190 298888
rect 45246 298832 45251 298888
rect 41492 298830 45251 298832
rect 45185 298827 45251 298830
rect 45461 298482 45527 298485
rect 652201 298482 652267 298485
rect 41492 298480 45527 298482
rect 41492 298424 45466 298480
rect 45522 298424 45527 298480
rect 41492 298422 45527 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 45461 298419 45527 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 42885 298074 42951 298077
rect 41492 298072 42951 298074
rect 41492 298016 42890 298072
rect 42946 298016 42951 298072
rect 41492 298014 42951 298016
rect 42885 298011 42951 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 675886 297332 675892 297396
rect 675956 297394 675962 297396
rect 678237 297394 678303 297397
rect 675956 297392 678303 297394
rect 675956 297336 678242 297392
rect 678298 297336 678303 297392
rect 675956 297334 678303 297336
rect 675956 297332 675962 297334
rect 678237 297331 678303 297334
rect 43253 297258 43319 297261
rect 41492 297256 43319 297258
rect 41492 297200 43258 297256
rect 43314 297200 43319 297256
rect 41492 297198 43319 297200
rect 43253 297195 43319 297198
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 675334 296788 675340 296852
rect 675404 296850 675410 296852
rect 676029 296850 676095 296853
rect 675404 296848 676095 296850
rect 675404 296792 676034 296848
rect 676090 296792 676095 296848
rect 675404 296790 676095 296792
rect 675404 296788 675410 296790
rect 676029 296787 676095 296790
rect 675518 296516 675524 296580
rect 675588 296578 675594 296580
rect 675845 296578 675911 296581
rect 675588 296576 675911 296578
rect 675588 296520 675850 296576
rect 675906 296520 675911 296576
rect 675588 296518 675911 296520
rect 675588 296516 675594 296518
rect 675845 296515 675911 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 42057 296034 42123 296037
rect 41492 296032 42123 296034
rect 41492 295976 42062 296032
rect 42118 295976 42123 296032
rect 41492 295974 42123 295976
rect 42057 295971 42123 295974
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 45001 295218 45067 295221
rect 41492 295216 45067 295218
rect 41492 295160 45006 295216
rect 45062 295160 45067 295216
rect 41492 295158 45067 295160
rect 45001 295155 45067 295158
rect 675753 295218 675819 295221
rect 676806 295218 676812 295220
rect 675753 295216 676812 295218
rect 675753 295160 675758 295216
rect 675814 295160 676812 295216
rect 675753 295158 676812 295160
rect 675753 295155 675819 295158
rect 676806 295156 676812 295158
rect 676876 295156 676882 295220
rect 37917 294810 37983 294813
rect 37917 294808 37996 294810
rect 37917 294752 37922 294808
rect 37978 294752 37996 294808
rect 37917 294750 37996 294752
rect 37917 294747 37983 294750
rect 43437 294402 43503 294405
rect 41492 294400 43503 294402
rect 41492 294344 43442 294400
rect 43498 294344 43503 294400
rect 41492 294342 43503 294344
rect 43437 294339 43503 294342
rect 44357 293994 44423 293997
rect 41492 293992 44423 293994
rect 41492 293936 44362 293992
rect 44418 293936 44423 293992
rect 41492 293934 44423 293936
rect 44357 293931 44423 293934
rect 43069 293586 43135 293589
rect 41492 293584 43135 293586
rect 41492 293528 43074 293584
rect 43130 293528 43135 293584
rect 41492 293526 43135 293528
rect 43069 293523 43135 293526
rect 43621 293178 43687 293181
rect 41492 293176 43687 293178
rect 41492 293120 43626 293176
rect 43682 293120 43687 293176
rect 41492 293118 43687 293120
rect 43621 293115 43687 293118
rect 674833 292906 674899 292909
rect 675385 292906 675451 292909
rect 674833 292904 675451 292906
rect 674833 292848 674838 292904
rect 674894 292848 675390 292904
rect 675446 292848 675451 292904
rect 674833 292846 675451 292848
rect 674833 292843 674899 292846
rect 675385 292843 675451 292846
rect 41781 292772 41847 292773
rect 41781 292768 41828 292772
rect 41892 292770 41898 292772
rect 40910 292592 40970 292740
rect 41781 292712 41786 292768
rect 41781 292708 41828 292712
rect 41892 292710 41938 292770
rect 41892 292708 41898 292710
rect 41781 292707 41847 292708
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40542 292332 40602 292528
rect 41822 292300 41828 292364
rect 41892 292362 41898 292364
rect 42057 292362 42123 292365
rect 41892 292360 42123 292362
rect 41892 292304 42062 292360
rect 42118 292304 42123 292360
rect 41892 292302 42123 292304
rect 41892 292300 41898 292302
rect 42057 292299 42123 292302
rect 675569 292092 675635 292093
rect 675518 292028 675524 292092
rect 675588 292090 675635 292092
rect 675588 292088 675680 292090
rect 675630 292032 675680 292088
rect 675588 292030 675680 292032
rect 675588 292028 675635 292030
rect 675569 292027 675635 292028
rect 43805 291954 43871 291957
rect 41492 291952 43871 291954
rect 41492 291896 43810 291952
rect 43866 291896 43871 291952
rect 41492 291894 43871 291896
rect 43805 291891 43871 291894
rect 44817 291954 44883 291957
rect 45461 291954 45527 291957
rect 44817 291952 45527 291954
rect 44817 291896 44822 291952
rect 44878 291896 45466 291952
rect 45522 291896 45527 291952
rect 44817 291894 45527 291896
rect 44817 291891 44883 291894
rect 45461 291891 45527 291894
rect 44173 291546 44239 291549
rect 41492 291544 44239 291546
rect 41492 291488 44178 291544
rect 44234 291488 44239 291544
rect 41492 291486 44239 291488
rect 44173 291483 44239 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 42241 291138 42307 291141
rect 41492 291136 42307 291138
rect 41492 291080 42246 291136
rect 42302 291080 42307 291136
rect 41492 291078 42307 291080
rect 42241 291075 42307 291078
rect 41492 290670 41890 290730
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 41830 290186 41890 290670
rect 42057 290458 42123 290461
rect 49141 290458 49207 290461
rect 42057 290456 49207 290458
rect 42057 290400 42062 290456
rect 42118 290400 49146 290456
rect 49202 290400 49207 290456
rect 42057 290398 49207 290400
rect 42057 290395 42123 290398
rect 49141 290395 49207 290398
rect 50337 290186 50403 290189
rect 41830 290184 50403 290186
rect 41830 290128 50342 290184
rect 50398 290128 50403 290184
rect 41830 290126 50403 290128
rect 50337 290123 50403 290126
rect 672441 290186 672507 290189
rect 675385 290186 675451 290189
rect 672441 290184 675451 290186
rect 672441 290128 672446 290184
rect 672502 290128 675390 290184
rect 675446 290128 675451 290184
rect 672441 290126 675451 290128
rect 672441 290123 672507 290126
rect 675385 290123 675451 290126
rect 42057 289914 42123 289917
rect 41492 289912 42123 289914
rect 41492 289856 42062 289912
rect 42118 289856 42123 289912
rect 41492 289854 42123 289856
rect 42057 289851 42123 289854
rect 42241 289914 42307 289917
rect 51717 289914 51783 289917
rect 675293 289916 675359 289917
rect 675293 289914 675340 289916
rect 42241 289912 51783 289914
rect 42241 289856 42246 289912
rect 42302 289856 51722 289912
rect 51778 289856 51783 289912
rect 42241 289854 51783 289856
rect 675248 289912 675340 289914
rect 675248 289856 675298 289912
rect 675248 289854 675340 289856
rect 42241 289851 42307 289854
rect 51717 289851 51783 289854
rect 675293 289852 675340 289854
rect 675404 289852 675410 289916
rect 675293 289851 675359 289852
rect 672625 287874 672691 287877
rect 675109 287874 675175 287877
rect 672625 287872 675175 287874
rect 672625 287816 672630 287872
rect 672686 287816 675114 287872
rect 675170 287816 675175 287872
rect 672625 287814 675175 287816
rect 672625 287811 672691 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 674465 286650 674531 286653
rect 675385 286650 675451 286653
rect 674465 286648 675451 286650
rect 674465 286592 674470 286648
rect 674526 286592 675390 286648
rect 675446 286592 675451 286648
rect 674465 286590 675451 286592
rect 674465 286587 674531 286590
rect 675385 286587 675451 286590
rect 674097 285562 674163 285565
rect 675109 285562 675175 285565
rect 674097 285560 675175 285562
rect 674097 285504 674102 285560
rect 674158 285504 675114 285560
rect 675170 285504 675175 285560
rect 674097 285502 675175 285504
rect 674097 285499 674163 285502
rect 675109 285499 675175 285502
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62941 285154 63007 285157
rect 62941 285152 64492 285154
rect 62941 285096 62946 285152
rect 63002 285096 64492 285152
rect 62941 285094 64492 285096
rect 62941 285091 63007 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282844 675727 282845
rect 675661 282840 675708 282844
rect 675772 282842 675778 282844
rect 675661 282784 675666 282840
rect 675661 282780 675708 282784
rect 675772 282782 675818 282842
rect 675772 282780 675778 282782
rect 675661 282779 675727 282780
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 675661 281210 675727 281213
rect 675886 281210 675892 281212
rect 675661 281208 675892 281210
rect 675661 281152 675666 281208
rect 675722 281152 675892 281208
rect 675661 281150 675892 281152
rect 675661 281147 675727 281150
rect 675886 281148 675892 281150
rect 675956 281148 675962 281212
rect 42149 279850 42215 279853
rect 43621 279850 43687 279853
rect 42149 279848 43687 279850
rect 42149 279792 42154 279848
rect 42210 279792 43626 279848
rect 43682 279792 43687 279848
rect 42149 279790 43687 279792
rect 42149 279787 42215 279790
rect 43621 279787 43687 279790
rect 42425 278762 42491 278765
rect 55857 278762 55923 278765
rect 42425 278760 55923 278762
rect 42425 278704 42430 278760
rect 42486 278704 55862 278760
rect 55918 278704 55923 278760
rect 42425 278702 55923 278704
rect 42425 278699 42491 278702
rect 55857 278699 55923 278702
rect 673862 278564 673868 278628
rect 673932 278564 673938 278628
rect 42425 278218 42491 278221
rect 44173 278218 44239 278221
rect 42425 278216 44239 278218
rect 42425 278160 42430 278216
rect 42486 278160 44178 278216
rect 44234 278160 44239 278216
rect 42425 278158 44239 278160
rect 42425 278155 42491 278158
rect 44173 278155 44239 278158
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 41781 277946 41847 277949
rect 40972 277944 41847 277946
rect 40972 277888 41786 277944
rect 41842 277888 41847 277944
rect 40972 277886 41847 277888
rect 40972 277884 40978 277886
rect 41781 277883 41847 277886
rect 40718 277612 40724 277676
rect 40788 277674 40794 277676
rect 42333 277674 42399 277677
rect 673870 277676 673930 278564
rect 40788 277672 42399 277674
rect 40788 277616 42338 277672
rect 42394 277616 42399 277672
rect 40788 277614 42399 277616
rect 40788 277612 40794 277614
rect 42333 277611 42399 277614
rect 673862 277612 673868 277676
rect 673932 277612 673938 277676
rect 42149 277402 42215 277405
rect 43805 277402 43871 277405
rect 42149 277400 43871 277402
rect 42149 277344 42154 277400
rect 42210 277344 43810 277400
rect 43866 277344 43871 277400
rect 42149 277342 43871 277344
rect 42149 277339 42215 277342
rect 43805 277339 43871 277342
rect 42057 276586 42123 276589
rect 45001 276586 45067 276589
rect 42057 276584 45067 276586
rect 42057 276528 42062 276584
rect 42118 276528 45006 276584
rect 45062 276528 45067 276584
rect 42057 276526 45067 276528
rect 42057 276523 42123 276526
rect 45001 276523 45067 276526
rect 671337 275362 671403 275365
rect 683297 275362 683363 275365
rect 671337 275360 683363 275362
rect 671337 275304 671342 275360
rect 671398 275304 683302 275360
rect 683358 275304 683363 275360
rect 671337 275302 683363 275304
rect 671337 275299 671403 275302
rect 683297 275299 683363 275302
rect 535729 275226 535795 275229
rect 633341 275226 633407 275229
rect 535729 275224 633407 275226
rect 535729 275168 535734 275224
rect 535790 275168 633346 275224
rect 633402 275168 633407 275224
rect 535729 275166 633407 275168
rect 535729 275163 535795 275166
rect 633341 275163 633407 275166
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 513189 274138 513255 274141
rect 602521 274138 602587 274141
rect 513189 274136 602587 274138
rect 513189 274080 513194 274136
rect 513250 274080 602526 274136
rect 602582 274080 602587 274136
rect 513189 274078 602587 274080
rect 513189 274075 513255 274078
rect 602521 274075 602587 274078
rect 533429 273866 533495 273869
rect 630949 273866 631015 273869
rect 533429 273864 631015 273866
rect 533429 273808 533434 273864
rect 533490 273808 630954 273864
rect 631010 273808 631015 273864
rect 533429 273806 631015 273808
rect 533429 273803 533495 273806
rect 630949 273803 631015 273806
rect 42057 273458 42123 273461
rect 43069 273458 43135 273461
rect 42057 273456 43135 273458
rect 42057 273400 42062 273456
rect 42118 273400 43074 273456
rect 43130 273400 43135 273456
rect 42057 273398 43135 273400
rect 42057 273395 42123 273398
rect 43069 273395 43135 273398
rect 521469 273050 521535 273053
rect 614389 273050 614455 273053
rect 521469 273048 614455 273050
rect 521469 272992 521474 273048
rect 521530 272992 614394 273048
rect 614450 272992 614455 273048
rect 521469 272990 614455 272992
rect 521469 272987 521535 272990
rect 614389 272987 614455 272990
rect 42057 272914 42123 272917
rect 44357 272914 44423 272917
rect 42057 272912 44423 272914
rect 42057 272856 42062 272912
rect 42118 272856 44362 272912
rect 44418 272856 44423 272912
rect 42057 272854 44423 272856
rect 42057 272851 42123 272854
rect 44357 272851 44423 272854
rect 533889 272778 533955 272781
rect 632145 272778 632211 272781
rect 533889 272776 632211 272778
rect 533889 272720 533894 272776
rect 533950 272720 632150 272776
rect 632206 272720 632211 272776
rect 533889 272718 632211 272720
rect 533889 272715 533955 272718
rect 632145 272715 632211 272718
rect 539317 272506 539383 272509
rect 639229 272506 639295 272509
rect 539317 272504 639295 272506
rect 539317 272448 539322 272504
rect 539378 272448 639234 272504
rect 639290 272448 639295 272504
rect 539317 272446 639295 272448
rect 539317 272443 539383 272446
rect 639229 272443 639295 272446
rect 479701 271418 479767 271421
rect 551737 271418 551803 271421
rect 479701 271416 551803 271418
rect 479701 271360 479706 271416
rect 479762 271360 551742 271416
rect 551798 271360 551803 271416
rect 479701 271358 551803 271360
rect 479701 271355 479767 271358
rect 551737 271355 551803 271358
rect 507761 271146 507827 271149
rect 593137 271146 593203 271149
rect 507761 271144 593203 271146
rect 507761 271088 507766 271144
rect 507822 271088 593142 271144
rect 593198 271088 593203 271144
rect 507761 271086 593203 271088
rect 507761 271083 507827 271086
rect 593137 271083 593203 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 42425 270466 42491 270469
rect 43437 270466 43503 270469
rect 42425 270464 43503 270466
rect 42425 270408 42430 270464
rect 42486 270408 43442 270464
rect 43498 270408 43503 270464
rect 42425 270406 43503 270408
rect 42425 270403 42491 270406
rect 43437 270403 43503 270406
rect 530945 270330 531011 270333
rect 626625 270330 626691 270333
rect 530945 270328 626691 270330
rect 530945 270272 530950 270328
rect 531006 270272 626630 270328
rect 626686 270272 626691 270328
rect 530945 270270 626691 270272
rect 530945 270267 531011 270270
rect 626625 270267 626691 270270
rect 538029 270058 538095 270061
rect 637573 270058 637639 270061
rect 538029 270056 637639 270058
rect 538029 270000 538034 270056
rect 538090 270000 637578 270056
rect 637634 270000 637639 270056
rect 538029 269998 637639 270000
rect 538029 269995 538095 269998
rect 637573 269995 637639 269998
rect 102041 269786 102107 269789
rect 161289 269786 161355 269789
rect 102041 269784 161355 269786
rect 102041 269728 102046 269784
rect 102102 269728 161294 269784
rect 161350 269728 161355 269784
rect 102041 269726 161355 269728
rect 102041 269723 102107 269726
rect 161289 269723 161355 269726
rect 468477 269786 468543 269789
rect 537661 269786 537727 269789
rect 468477 269784 537727 269786
rect 468477 269728 468482 269784
rect 468538 269728 537666 269784
rect 537722 269728 537727 269784
rect 468477 269726 537727 269728
rect 468477 269723 468543 269726
rect 537661 269723 537727 269726
rect 540513 269786 540579 269789
rect 640701 269786 640767 269789
rect 540513 269784 640767 269786
rect 540513 269728 540518 269784
rect 540574 269728 640706 269784
rect 640762 269728 640767 269784
rect 540513 269726 640767 269728
rect 540513 269723 540579 269726
rect 640701 269723 640767 269726
rect 497457 269514 497523 269517
rect 568573 269514 568639 269517
rect 497457 269512 568639 269514
rect 497457 269456 497462 269512
rect 497518 269456 568578 269512
rect 568634 269456 568639 269512
rect 497457 269454 568639 269456
rect 497457 269451 497523 269454
rect 568573 269451 568639 269454
rect 470961 269242 471027 269245
rect 539501 269242 539567 269245
rect 470961 269240 539567 269242
rect 470961 269184 470966 269240
rect 471022 269184 539506 269240
rect 539562 269184 539567 269240
rect 470961 269182 539567 269184
rect 470961 269179 471027 269182
rect 539501 269179 539567 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 676262 268562 676322 268668
rect 683297 268562 683363 268565
rect 663750 268502 676322 268562
rect 683254 268560 683363 268562
rect 683254 268504 683302 268560
rect 683358 268504 683363 268560
rect 506105 268426 506171 268429
rect 591113 268426 591179 268429
rect 506105 268424 591179 268426
rect 506105 268368 506110 268424
rect 506166 268368 591118 268424
rect 591174 268368 591179 268424
rect 506105 268366 591179 268368
rect 506105 268363 506171 268366
rect 591113 268363 591179 268366
rect 663057 268154 663123 268157
rect 663750 268154 663810 268502
rect 683254 268499 683363 268504
rect 683254 268260 683314 268499
rect 683113 268154 683179 268157
rect 663057 268152 663810 268154
rect 663057 268096 663062 268152
rect 663118 268096 663810 268152
rect 663057 268094 663810 268096
rect 683070 268152 683179 268154
rect 683070 268096 683118 268152
rect 683174 268096 683179 268152
rect 663057 268091 663123 268094
rect 683070 268091 683179 268096
rect 683070 267852 683130 268091
rect 519813 267338 519879 267341
rect 563697 267338 563763 267341
rect 519813 267336 563763 267338
rect 519813 267280 519818 267336
rect 519874 267280 563702 267336
rect 563758 267280 563763 267336
rect 519813 267278 563763 267280
rect 519813 267275 519879 267278
rect 563697 267275 563763 267278
rect 672809 267338 672875 267341
rect 676262 267338 676322 267444
rect 672809 267336 676322 267338
rect 672809 267280 672814 267336
rect 672870 267280 676322 267336
rect 672809 267278 676322 267280
rect 672809 267275 672875 267278
rect 40677 267066 40743 267069
rect 62757 267066 62823 267069
rect 40677 267064 62823 267066
rect 40677 267008 40682 267064
rect 40738 267008 62762 267064
rect 62818 267008 62823 267064
rect 40677 267006 62823 267008
rect 40677 267003 40743 267006
rect 62757 267003 62823 267006
rect 75913 267066 75979 267069
rect 138105 267066 138171 267069
rect 75913 267064 138171 267066
rect 75913 267008 75918 267064
rect 75974 267008 138110 267064
rect 138166 267008 138171 267064
rect 75913 267006 138171 267008
rect 75913 267003 75979 267006
rect 138105 267003 138171 267006
rect 484117 267066 484183 267069
rect 507945 267066 508011 267069
rect 484117 267064 508011 267066
rect 484117 267008 484122 267064
rect 484178 267008 507950 267064
rect 508006 267008 508011 267064
rect 484117 267006 508011 267008
rect 484117 267003 484183 267006
rect 507945 267003 508011 267006
rect 517145 267066 517211 267069
rect 585777 267066 585843 267069
rect 517145 267064 585843 267066
rect 517145 267008 517150 267064
rect 517206 267008 585782 267064
rect 585838 267008 585843 267064
rect 517145 267006 585843 267008
rect 517145 267003 517211 267006
rect 585777 267003 585843 267006
rect 674005 267066 674071 267069
rect 674005 267064 676292 267066
rect 674005 267008 674010 267064
rect 674066 267008 676292 267064
rect 674005 267006 676292 267008
rect 674005 267003 674071 267006
rect 674649 266658 674715 266661
rect 674649 266656 676292 266658
rect 674649 266600 674654 266656
rect 674710 266600 676292 266656
rect 674649 266598 676292 266600
rect 674649 266595 674715 266598
rect 477585 266386 477651 266389
rect 479701 266386 479767 266389
rect 477585 266384 479767 266386
rect 477585 266328 477590 266384
rect 477646 266328 479706 266384
rect 479762 266328 479767 266384
rect 477585 266326 479767 266328
rect 477585 266323 477651 266326
rect 479701 266323 479767 266326
rect 676446 266117 676506 266220
rect 674281 266114 674347 266117
rect 674281 266112 676322 266114
rect 674281 266056 674286 266112
rect 674342 266056 676322 266112
rect 674281 266054 676322 266056
rect 676446 266112 676555 266117
rect 676446 266056 676494 266112
rect 676550 266056 676555 266112
rect 676446 266054 676555 266056
rect 674281 266051 674347 266054
rect 676262 265812 676322 266054
rect 676489 266051 676555 266054
rect 672533 265706 672599 265709
rect 672533 265704 676322 265706
rect 672533 265648 672538 265704
rect 672594 265648 676322 265704
rect 672533 265646 676322 265648
rect 672533 265643 672599 265646
rect 676262 265404 676322 265646
rect 674557 265298 674623 265301
rect 676489 265298 676555 265301
rect 674557 265296 676555 265298
rect 674557 265240 674562 265296
rect 674618 265240 676494 265296
rect 676550 265240 676555 265296
rect 674557 265238 676555 265240
rect 674557 265235 674623 265238
rect 676489 265235 676555 265238
rect 673085 265026 673151 265029
rect 673085 265024 676292 265026
rect 673085 264968 673090 265024
rect 673146 264968 676292 265024
rect 673085 264966 676292 264968
rect 673085 264963 673151 264966
rect 674833 264482 674899 264485
rect 676262 264482 676322 264588
rect 674833 264480 676322 264482
rect 674833 264424 674838 264480
rect 674894 264424 676322 264480
rect 674833 264422 676322 264424
rect 674833 264419 674899 264422
rect 676446 264077 676506 264180
rect 670141 264074 670207 264077
rect 670141 264072 676322 264074
rect 670141 264016 670146 264072
rect 670202 264016 676322 264072
rect 670141 264014 676322 264016
rect 676446 264072 676555 264077
rect 676446 264016 676494 264072
rect 676550 264016 676555 264072
rect 676446 264014 676555 264016
rect 670141 264011 670207 264014
rect 672901 263802 672967 263805
rect 674833 263802 674899 263805
rect 672901 263800 674899 263802
rect 672901 263744 672906 263800
rect 672962 263744 674838 263800
rect 674894 263744 674899 263800
rect 676262 263772 676322 264014
rect 676489 264011 676555 264014
rect 672901 263742 674899 263744
rect 672901 263739 672967 263742
rect 674833 263739 674899 263742
rect 674966 263604 674972 263668
rect 675036 263666 675042 263668
rect 676489 263666 676555 263669
rect 675036 263664 676555 263666
rect 675036 263608 676494 263664
rect 676550 263608 676555 263664
rect 675036 263606 676555 263608
rect 675036 263604 675042 263606
rect 676489 263603 676555 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 676070 262380 676076 262444
rect 676140 262442 676146 262444
rect 676262 262442 676322 262548
rect 676140 262382 676322 262442
rect 676140 262380 676146 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671705 262034 671771 262037
rect 676262 262034 676322 262140
rect 671705 262032 676322 262034
rect 671705 261976 671710 262032
rect 671766 261976 676322 262032
rect 671705 261974 676322 261976
rect 671705 261971 671771 261974
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 679574 261221 679634 261324
rect 679574 261216 679683 261221
rect 679574 261160 679622 261216
rect 679678 261160 679683 261216
rect 679574 261158 679683 261160
rect 679617 261155 679683 261158
rect 673821 260946 673887 260949
rect 673821 260944 676292 260946
rect 673821 260888 673826 260944
rect 673882 260888 676292 260944
rect 673821 260886 676292 260888
rect 673821 260883 673887 260886
rect 673085 260402 673151 260405
rect 676262 260402 676322 260508
rect 673085 260400 676322 260402
rect 673085 260344 673090 260400
rect 673146 260344 676322 260400
rect 673085 260342 676322 260344
rect 673085 260339 673151 260342
rect 35801 259994 35867 259997
rect 46197 259994 46263 259997
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 35801 259992 46263 259994
rect 35801 259936 35806 259992
rect 35862 259936 46202 259992
rect 46258 259936 46263 259992
rect 35801 259934 46263 259936
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 35801 259931 35867 259934
rect 46197 259931 46263 259934
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 669957 259586 670023 259589
rect 676262 259586 676322 259692
rect 669957 259584 676322 259586
rect 669957 259528 669962 259584
rect 670018 259528 676322 259584
rect 669957 259526 676322 259528
rect 669957 259523 670023 259526
rect 671521 259178 671587 259181
rect 676262 259178 676322 259284
rect 671521 259176 676322 259178
rect 671521 259120 671526 259176
rect 671582 259120 676322 259176
rect 671521 259118 676322 259120
rect 671521 259115 671587 259118
rect 675937 258770 676003 258773
rect 676262 258770 676322 258876
rect 675937 258768 676322 258770
rect 675937 258712 675942 258768
rect 675998 258712 676322 258768
rect 675937 258710 676322 258712
rect 675937 258707 676003 258710
rect 673637 258498 673703 258501
rect 673637 258496 676292 258498
rect 673637 258440 673642 258496
rect 673698 258440 676292 258496
rect 673637 258438 676292 258440
rect 673637 258435 673703 258438
rect 35801 258362 35867 258365
rect 35758 258360 35867 258362
rect 35758 258304 35806 258360
rect 35862 258304 35867 258360
rect 35758 258299 35867 258304
rect 35758 258060 35818 258299
rect 675937 258226 676003 258229
rect 675894 258224 676003 258226
rect 675894 258168 675942 258224
rect 675998 258168 676003 258224
rect 675894 258163 676003 258168
rect 671337 257954 671403 257957
rect 675894 257954 675954 258163
rect 671337 257952 675954 257954
rect 671337 257896 671342 257952
rect 671398 257896 675954 257952
rect 671337 257894 675954 257896
rect 671337 257891 671403 257894
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 41462 257546 41522 257652
rect 53281 257546 53347 257549
rect 41462 257544 53347 257546
rect 41462 257488 53286 257544
rect 53342 257488 53347 257544
rect 41462 257486 53347 257488
rect 53281 257483 53347 257486
rect 675293 257546 675359 257549
rect 676262 257546 676322 258060
rect 675293 257544 676322 257546
rect 675293 257488 675298 257544
rect 675354 257488 676322 257544
rect 675293 257486 676322 257488
rect 675293 257483 675359 257486
rect 35758 257141 35818 257244
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 672717 257138 672783 257141
rect 676262 257138 676322 257244
rect 672717 257136 676322 257138
rect 672717 257080 672722 257136
rect 672778 257080 676322 257136
rect 672717 257078 676322 257080
rect 672717 257075 672783 257078
rect 44633 256866 44699 256869
rect 41492 256864 44699 256866
rect 41492 256808 44638 256864
rect 44694 256808 44699 256864
rect 41492 256806 44699 256808
rect 44633 256803 44699 256806
rect 671981 256730 672047 256733
rect 675293 256730 675359 256733
rect 671981 256728 675359 256730
rect 671981 256672 671986 256728
rect 672042 256672 675298 256728
rect 675354 256672 675359 256728
rect 671981 256670 675359 256672
rect 671981 256667 672047 256670
rect 675293 256667 675359 256670
rect 43621 256458 43687 256461
rect 41492 256456 43687 256458
rect 41492 256400 43626 256456
rect 43682 256400 43687 256456
rect 41492 256398 43687 256400
rect 43621 256395 43687 256398
rect 45093 256050 45159 256053
rect 41492 256048 45159 256050
rect 41492 255992 45098 256048
rect 45154 255992 45159 256048
rect 41492 255990 45159 255992
rect 45093 255987 45159 255990
rect 675201 255914 675267 255917
rect 676121 255914 676187 255917
rect 675201 255912 676187 255914
rect 675201 255856 675206 255912
rect 675262 255856 676126 255912
rect 676182 255856 676187 255912
rect 675201 255854 676187 255856
rect 675201 255851 675267 255854
rect 676121 255851 676187 255854
rect 43437 255642 43503 255645
rect 553761 255642 553827 255645
rect 41492 255640 43503 255642
rect 41492 255584 43442 255640
rect 43498 255584 43503 255640
rect 41492 255582 43503 255584
rect 552460 255640 553827 255642
rect 552460 255584 553766 255640
rect 553822 255584 553827 255640
rect 552460 255582 553827 255584
rect 43437 255579 43503 255582
rect 553761 255579 553827 255582
rect 42885 255234 42951 255237
rect 41492 255232 42951 255234
rect 41492 255176 42890 255232
rect 42946 255176 42951 255232
rect 41492 255174 42951 255176
rect 42885 255171 42951 255174
rect 42885 254826 42951 254829
rect 41492 254824 42951 254826
rect 41492 254768 42890 254824
rect 42946 254768 42951 254824
rect 41492 254766 42951 254768
rect 42885 254763 42951 254766
rect 43253 254418 43319 254421
rect 41492 254416 43319 254418
rect 41492 254360 43258 254416
rect 43314 254360 43319 254416
rect 41492 254358 43319 254360
rect 43253 254355 43319 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35758 253469 35818 253572
rect 35758 253464 35867 253469
rect 554405 253466 554471 253469
rect 35758 253408 35806 253464
rect 35862 253408 35867 253464
rect 35758 253406 35867 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35801 253403 35867 253406
rect 554405 253403 554471 253406
rect 35574 253061 35634 253164
rect 35574 253056 35683 253061
rect 35574 253000 35622 253056
rect 35678 253000 35683 253056
rect 35574 252998 35683 253000
rect 35617 252995 35683 252998
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 41321 252242 41387 252245
rect 42517 252242 42583 252245
rect 41321 252240 42583 252242
rect 41321 252184 41326 252240
rect 41382 252184 42522 252240
rect 42578 252184 42583 252240
rect 41321 252182 42583 252184
rect 41321 252179 41387 252182
rect 42517 252179 42583 252182
rect 44357 251970 44423 251973
rect 41492 251968 44423 251970
rect 41492 251912 44362 251968
rect 44418 251912 44423 251968
rect 41492 251910 44423 251912
rect 44357 251907 44423 251910
rect 675017 251834 675083 251837
rect 676029 251834 676095 251837
rect 675017 251832 676095 251834
rect 675017 251776 675022 251832
rect 675078 251776 676034 251832
rect 676090 251776 676095 251832
rect 675017 251774 676095 251776
rect 675017 251771 675083 251774
rect 676029 251771 676095 251774
rect 40542 251428 40602 251532
rect 40534 251364 40540 251428
rect 40604 251364 40610 251428
rect 553485 251290 553551 251293
rect 552460 251288 553551 251290
rect 552460 251232 553490 251288
rect 553546 251232 553551 251288
rect 552460 251230 553551 251232
rect 553485 251227 553551 251230
rect 45553 251154 45619 251157
rect 41492 251152 45619 251154
rect 41492 251096 45558 251152
rect 45614 251096 45619 251152
rect 41492 251094 45619 251096
rect 45553 251091 45619 251094
rect 45829 250746 45895 250749
rect 41492 250744 45895 250746
rect 41492 250688 45834 250744
rect 45890 250688 45895 250744
rect 41492 250686 45895 250688
rect 45829 250683 45895 250686
rect 43069 250338 43135 250341
rect 41492 250336 43135 250338
rect 41492 250280 43074 250336
rect 43130 250280 43135 250336
rect 41492 250278 43135 250280
rect 43069 250275 43135 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 673862 249596 673868 249660
rect 673932 249658 673938 249660
rect 674281 249658 674347 249661
rect 673932 249656 674347 249658
rect 673932 249600 674286 249656
rect 674342 249600 674347 249656
rect 673932 249598 674347 249600
rect 673932 249596 673938 249598
rect 674281 249595 674347 249598
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675385 249658 675451 249661
rect 674852 249656 675451 249658
rect 674852 249600 675390 249656
rect 675446 249600 675451 249656
rect 674852 249598 675451 249600
rect 674852 249596 674858 249598
rect 675385 249595 675451 249598
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 674925 249386 674991 249389
rect 676078 249386 676138 249596
rect 674925 249384 676138 249386
rect 674925 249328 674930 249384
rect 674986 249328 676138 249384
rect 674925 249326 676138 249328
rect 674925 249323 674991 249326
rect 43805 249114 43871 249117
rect 554037 249114 554103 249117
rect 41492 249112 43871 249114
rect 41492 249056 43810 249112
rect 43866 249056 43871 249112
rect 41492 249054 43871 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 43805 249051 43871 249054
rect 554037 249051 554103 249054
rect 44541 248706 44607 248709
rect 41492 248704 44607 248706
rect 41492 248648 44546 248704
rect 44602 248648 44607 248704
rect 41492 248646 44607 248648
rect 44541 248643 44607 248646
rect 45001 248298 45067 248301
rect 41492 248296 45067 248298
rect 41492 248240 45006 248296
rect 45062 248240 45067 248296
rect 41492 248238 45067 248240
rect 45001 248235 45067 248238
rect 46197 247890 46263 247893
rect 41492 247888 46263 247890
rect 41492 247832 46202 247888
rect 46258 247832 46263 247888
rect 41492 247830 46263 247832
rect 46197 247827 46263 247830
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46933 247074 46999 247077
rect 41492 247072 46999 247074
rect 41492 247016 46938 247072
rect 46994 247016 46999 247072
rect 41492 247014 46999 247016
rect 46933 247011 46999 247014
rect 553853 246938 553919 246941
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 553853 246875 553919 246878
rect 41462 246530 41522 246636
rect 50521 246530 50587 246533
rect 41462 246528 50587 246530
rect 41462 246472 50526 246528
rect 50582 246472 50587 246528
rect 41462 246470 50587 246472
rect 50521 246467 50587 246470
rect 673821 246530 673887 246533
rect 675385 246530 675451 246533
rect 673821 246528 675451 246530
rect 673821 246472 673826 246528
rect 673882 246472 675390 246528
rect 675446 246472 675451 246528
rect 673821 246470 675451 246472
rect 673821 246467 673887 246470
rect 675385 246467 675451 246470
rect 673453 246258 673519 246261
rect 674598 246258 674604 246260
rect 673453 246256 674604 246258
rect 673453 246200 673458 246256
rect 673514 246200 674604 246256
rect 673453 246198 674604 246200
rect 673453 246195 673519 246198
rect 674598 246196 674604 246198
rect 674668 246196 674674 246260
rect 669957 245850 670023 245853
rect 675385 245850 675451 245853
rect 669957 245848 675451 245850
rect 669957 245792 669962 245848
rect 670018 245792 675390 245848
rect 675446 245792 675451 245848
rect 669957 245790 675451 245792
rect 669957 245787 670023 245790
rect 675385 245787 675451 245790
rect 674925 245578 674991 245581
rect 676806 245578 676812 245580
rect 674925 245576 676812 245578
rect 674925 245520 674930 245576
rect 674986 245520 676812 245576
rect 674925 245518 676812 245520
rect 674925 245515 674991 245518
rect 676806 245516 676812 245518
rect 676876 245516 676882 245580
rect 673177 245306 673243 245309
rect 675334 245306 675340 245308
rect 673177 245304 675340 245306
rect 673177 245248 673182 245304
rect 673238 245248 675340 245304
rect 673177 245246 675340 245248
rect 673177 245243 673243 245246
rect 675334 245244 675340 245246
rect 675404 245244 675410 245308
rect 671705 245034 671771 245037
rect 675150 245034 675156 245036
rect 671705 245032 675156 245034
rect 671705 244976 671710 245032
rect 671766 244976 675156 245032
rect 671705 244974 675156 244976
rect 671705 244971 671771 244974
rect 675150 244972 675156 244974
rect 675220 244972 675226 245036
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 41689 242858 41755 242861
rect 42701 242858 42767 242861
rect 41689 242856 42767 242858
rect 41689 242800 41694 242856
rect 41750 242800 42706 242856
rect 42762 242800 42767 242856
rect 41689 242798 42767 242800
rect 41689 242795 41755 242798
rect 42701 242795 42767 242798
rect 671521 242858 671587 242861
rect 675109 242858 675175 242861
rect 671521 242856 675175 242858
rect 671521 242800 671526 242856
rect 671582 242800 675114 242856
rect 675170 242800 675175 242856
rect 671521 242798 675175 242800
rect 671521 242795 671587 242798
rect 675109 242795 675175 242798
rect 40677 242586 40743 242589
rect 43253 242586 43319 242589
rect 553669 242586 553735 242589
rect 40677 242584 43319 242586
rect 40677 242528 40682 242584
rect 40738 242528 43258 242584
rect 43314 242528 43319 242584
rect 40677 242526 43319 242528
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 40677 242523 40743 242526
rect 43253 242523 43319 242526
rect 553669 242523 553735 242526
rect 671337 241498 671403 241501
rect 675109 241498 675175 241501
rect 671337 241496 675175 241498
rect 671337 241440 671342 241496
rect 671398 241440 675114 241496
rect 675170 241440 675175 241496
rect 671337 241438 675175 241440
rect 671337 241435 671403 241438
rect 675109 241435 675175 241438
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 675385 240276 675451 240277
rect 675334 240274 675340 240276
rect 675294 240214 675340 240274
rect 675404 240272 675451 240276
rect 675446 240216 675451 240272
rect 675334 240212 675340 240214
rect 675404 240212 675451 240216
rect 675385 240211 675451 240212
rect 40534 240076 40540 240140
rect 40604 240138 40610 240140
rect 41781 240138 41847 240141
rect 40604 240136 41847 240138
rect 40604 240080 41786 240136
rect 41842 240080 41847 240136
rect 40604 240078 41847 240080
rect 40604 240076 40610 240078
rect 41781 240075 41847 240078
rect 42057 238506 42123 238509
rect 46933 238506 46999 238509
rect 42057 238504 46999 238506
rect 42057 238448 42062 238504
rect 42118 238448 46938 238504
rect 46994 238448 46999 238504
rect 42057 238446 46999 238448
rect 42057 238443 42123 238446
rect 46933 238443 46999 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 671981 238098 672047 238101
rect 675385 238098 675451 238101
rect 671981 238096 675451 238098
rect 671981 238040 671986 238096
rect 672042 238040 675390 238096
rect 675446 238040 675451 238096
rect 671981 238038 675451 238040
rect 671981 238035 672047 238038
rect 675385 238035 675451 238038
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42517 237418 42583 237421
rect 42076 237416 42583 237418
rect 42076 237360 42522 237416
rect 42578 237360 42583 237416
rect 42076 237358 42583 237360
rect 42076 237356 42082 237358
rect 42517 237355 42583 237358
rect 672717 237418 672783 237421
rect 673678 237418 673684 237420
rect 672717 237416 673684 237418
rect 672717 237360 672722 237416
rect 672778 237360 673684 237416
rect 672717 237358 673684 237360
rect 672717 237355 672783 237358
rect 673678 237356 673684 237358
rect 673748 237356 673754 237420
rect 675201 237284 675267 237285
rect 675150 237282 675156 237284
rect 675110 237222 675156 237282
rect 675220 237280 675267 237284
rect 675262 237224 675267 237280
rect 675150 237220 675156 237222
rect 675220 237220 675267 237224
rect 675201 237219 675267 237220
rect 667013 237146 667079 237149
rect 673521 237146 673587 237149
rect 667013 237144 673587 237146
rect 667013 237088 667018 237144
rect 667074 237088 673526 237144
rect 673582 237088 673587 237144
rect 667013 237086 673587 237088
rect 667013 237083 667079 237086
rect 673521 237083 673587 237086
rect 672625 236466 672691 236469
rect 673637 236466 673703 236469
rect 672625 236464 673703 236466
rect 672625 236408 672630 236464
rect 672686 236408 673642 236464
rect 673698 236408 673703 236464
rect 672625 236406 673703 236408
rect 672625 236403 672691 236406
rect 673637 236403 673703 236406
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 40718 235860 40724 235924
rect 40788 235922 40794 235924
rect 41781 235922 41847 235925
rect 40788 235920 41847 235922
rect 40788 235864 41786 235920
rect 41842 235864 41847 235920
rect 40788 235862 41847 235864
rect 40788 235860 40794 235862
rect 41781 235859 41847 235862
rect 42425 235922 42491 235925
rect 45001 235922 45067 235925
rect 42425 235920 45067 235922
rect 42425 235864 42430 235920
rect 42486 235864 45006 235920
rect 45062 235864 45067 235920
rect 42425 235862 45067 235864
rect 42425 235859 42491 235862
rect 45001 235859 45067 235862
rect 670141 235922 670207 235925
rect 675017 235922 675083 235925
rect 670141 235920 675083 235922
rect 670141 235864 670146 235920
rect 670202 235864 675022 235920
rect 675078 235864 675083 235920
rect 670141 235862 675083 235864
rect 670141 235859 670207 235862
rect 675017 235859 675083 235862
rect 674419 235106 674485 235109
rect 676806 235106 676812 235108
rect 674419 235104 676812 235106
rect 674419 235048 674424 235104
rect 674480 235048 676812 235104
rect 674419 235046 676812 235048
rect 674419 235043 674485 235046
rect 676806 235044 676812 235046
rect 676876 235044 676882 235108
rect 671889 234834 671955 234837
rect 674281 234834 674347 234837
rect 671889 234832 674347 234834
rect 671889 234776 671894 234832
rect 671950 234776 674286 234832
rect 674342 234776 674347 234832
rect 671889 234774 674347 234776
rect 671889 234771 671955 234774
rect 674281 234771 674347 234774
rect 671286 234500 671292 234564
rect 671356 234562 671362 234564
rect 672073 234562 672139 234565
rect 671356 234560 672139 234562
rect 671356 234504 672078 234560
rect 672134 234504 672139 234560
rect 671356 234502 672139 234504
rect 671356 234500 671362 234502
rect 672073 234499 672139 234502
rect 668485 234290 668551 234293
rect 671705 234290 671771 234293
rect 668485 234288 671771 234290
rect 668485 234232 668490 234288
rect 668546 234232 671710 234288
rect 671766 234232 671771 234288
rect 668485 234230 671771 234232
rect 668485 234227 668551 234230
rect 671705 234227 671771 234230
rect 42241 234154 42307 234157
rect 44541 234154 44607 234157
rect 42241 234152 44607 234154
rect 42241 234096 42246 234152
rect 42302 234096 44546 234152
rect 44602 234096 44607 234152
rect 42241 234094 44607 234096
rect 42241 234091 42307 234094
rect 44541 234091 44607 234094
rect 674529 234154 674595 234157
rect 675845 234154 675911 234157
rect 674529 234152 675911 234154
rect 674529 234096 674534 234152
rect 674590 234096 675850 234152
rect 675906 234096 675911 234152
rect 674529 234094 675911 234096
rect 674529 234091 674595 234094
rect 675845 234091 675911 234094
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683205 233882 683271 233885
rect 658917 233880 683271 233882
rect 658917 233824 658922 233880
rect 658978 233824 683210 233880
rect 683266 233824 683271 233880
rect 658917 233822 683271 233824
rect 658917 233819 658983 233822
rect 683205 233819 683271 233822
rect 670785 233610 670851 233613
rect 675109 233610 675175 233613
rect 670785 233608 675175 233610
rect 670785 233552 670790 233608
rect 670846 233552 675114 233608
rect 675170 233552 675175 233608
rect 670785 233550 675175 233552
rect 670785 233547 670851 233550
rect 675109 233547 675175 233550
rect 42149 233338 42215 233341
rect 44357 233338 44423 233341
rect 42149 233336 44423 233338
rect 42149 233280 42154 233336
rect 42210 233280 44362 233336
rect 44418 233280 44423 233336
rect 42149 233278 44423 233280
rect 42149 233275 42215 233278
rect 44357 233275 44423 233278
rect 670049 233202 670115 233205
rect 671153 233202 671219 233205
rect 670049 233200 671219 233202
rect 670049 233144 670054 233200
rect 670110 233144 671158 233200
rect 671214 233144 671219 233200
rect 670049 233142 671219 233144
rect 670049 233139 670115 233142
rect 671153 233139 671219 233142
rect 669589 232794 669655 232797
rect 673729 232794 673795 232797
rect 669589 232792 673795 232794
rect 669589 232736 669594 232792
rect 669650 232736 673734 232792
rect 673790 232736 673795 232792
rect 669589 232734 673795 232736
rect 669589 232731 669655 232734
rect 673729 232731 673795 232734
rect 42425 232522 42491 232525
rect 46013 232522 46079 232525
rect 673637 232524 673703 232525
rect 673637 232522 673684 232524
rect 42425 232520 46079 232522
rect 42425 232464 42430 232520
rect 42486 232464 46018 232520
rect 46074 232464 46079 232520
rect 42425 232462 46079 232464
rect 673592 232520 673684 232522
rect 673592 232464 673642 232520
rect 673592 232462 673684 232464
rect 42425 232459 42491 232462
rect 46013 232459 46079 232462
rect 673637 232460 673684 232462
rect 673748 232460 673754 232524
rect 673637 232459 673703 232460
rect 42425 231842 42491 231845
rect 43805 231842 43871 231845
rect 42425 231840 43871 231842
rect 42425 231784 42430 231840
rect 42486 231784 43810 231840
rect 43866 231784 43871 231840
rect 42425 231782 43871 231784
rect 42425 231779 42491 231782
rect 43805 231779 43871 231782
rect 673678 231780 673684 231844
rect 673748 231842 673754 231844
rect 674649 231842 674715 231845
rect 673748 231840 674715 231842
rect 673748 231784 674654 231840
rect 674710 231784 674715 231840
rect 673748 231782 674715 231784
rect 673748 231780 673754 231782
rect 674649 231779 674715 231782
rect 672257 231570 672323 231573
rect 673310 231570 673316 231572
rect 672257 231568 673316 231570
rect 672257 231512 672262 231568
rect 672318 231512 673316 231568
rect 672257 231510 673316 231512
rect 672257 231507 672323 231510
rect 673310 231508 673316 231510
rect 673380 231508 673386 231572
rect 674649 231570 674715 231573
rect 675845 231570 675911 231573
rect 674649 231568 675911 231570
rect 674649 231512 674654 231568
rect 674710 231512 675850 231568
rect 675906 231512 675911 231568
rect 674649 231510 675911 231512
rect 674649 231507 674715 231510
rect 675845 231507 675911 231510
rect 663793 231298 663859 231301
rect 675063 231298 675129 231301
rect 663793 231296 675129 231298
rect 663793 231240 663798 231296
rect 663854 231240 675068 231296
rect 675124 231240 675129 231296
rect 663793 231238 675129 231240
rect 663793 231235 663859 231238
rect 675063 231235 675129 231238
rect 665817 231026 665883 231029
rect 674725 231026 674791 231029
rect 665817 231024 674791 231026
rect 665817 230968 665822 231024
rect 665878 230968 674730 231024
rect 674786 230968 674791 231024
rect 665817 230966 674791 230968
rect 665817 230963 665883 230966
rect 674725 230963 674791 230966
rect 663057 230754 663123 230757
rect 674833 230754 674899 230757
rect 663057 230752 674899 230754
rect 663057 230696 663062 230752
rect 663118 230696 674838 230752
rect 674894 230696 674899 230752
rect 663057 230694 674899 230696
rect 663057 230691 663123 230694
rect 674833 230691 674899 230694
rect 675017 230754 675083 230757
rect 675845 230754 675911 230757
rect 675017 230752 675911 230754
rect 675017 230696 675022 230752
rect 675078 230696 675850 230752
rect 675906 230696 675911 230752
rect 675017 230694 675911 230696
rect 675017 230691 675083 230694
rect 675845 230691 675911 230694
rect 42149 230482 42215 230485
rect 43069 230482 43135 230485
rect 42149 230480 43135 230482
rect 42149 230424 42154 230480
rect 42210 230424 43074 230480
rect 43130 230424 43135 230480
rect 42149 230422 43135 230424
rect 42149 230419 42215 230422
rect 43069 230419 43135 230422
rect 673913 230482 673979 230485
rect 676213 230482 676279 230485
rect 673913 230480 676279 230482
rect 673913 230424 673918 230480
rect 673974 230424 676218 230480
rect 676274 230424 676279 230480
rect 673913 230422 676279 230424
rect 673913 230419 673979 230422
rect 676213 230419 676279 230422
rect 665173 230346 665239 230349
rect 665173 230344 673700 230346
rect 665173 230288 665178 230344
rect 665234 230288 673700 230344
rect 665173 230286 673700 230288
rect 665173 230283 665239 230286
rect 673640 230210 673700 230286
rect 674649 230210 674715 230213
rect 677041 230210 677107 230213
rect 673640 230174 674482 230210
rect 673640 230150 674394 230174
rect 674389 230118 674394 230150
rect 674450 230118 674482 230174
rect 674649 230208 677107 230210
rect 674649 230152 674654 230208
rect 674710 230152 677046 230208
rect 677102 230152 677107 230208
rect 674649 230150 677107 230152
rect 674649 230147 674715 230150
rect 677041 230147 677107 230150
rect 674389 230116 674482 230118
rect 674389 230113 674455 230116
rect 71037 230074 71103 230077
rect 150801 230074 150867 230077
rect 671521 230076 671587 230077
rect 71037 230072 150867 230074
rect 71037 230016 71042 230072
rect 71098 230016 150806 230072
rect 150862 230016 150867 230072
rect 71037 230014 150867 230016
rect 71037 230011 71103 230014
rect 150801 230011 150867 230014
rect 671470 230012 671476 230076
rect 671540 230074 671587 230076
rect 673453 230076 673519 230077
rect 673453 230074 673500 230076
rect 671540 230072 671632 230074
rect 671582 230016 671632 230072
rect 671540 230014 671632 230016
rect 673408 230072 673500 230074
rect 673408 230016 673458 230072
rect 673408 230014 673500 230016
rect 671540 230012 671587 230014
rect 671521 230011 671587 230012
rect 673453 230012 673500 230014
rect 673564 230012 673570 230076
rect 673453 230011 673519 230012
rect 674165 229938 674231 229941
rect 675109 229938 675175 229941
rect 674165 229936 675175 229938
rect 674165 229880 674170 229936
rect 674226 229880 675114 229936
rect 675170 229880 675175 229936
rect 674165 229878 675175 229880
rect 674165 229875 674231 229878
rect 675109 229875 675175 229878
rect 65517 229802 65583 229805
rect 148225 229802 148291 229805
rect 65517 229800 148291 229802
rect 65517 229744 65522 229800
rect 65578 229744 148230 229800
rect 148286 229744 148291 229800
rect 65517 229742 148291 229744
rect 65517 229739 65583 229742
rect 148225 229739 148291 229742
rect 639597 229802 639663 229805
rect 673821 229802 673887 229805
rect 639597 229800 673887 229802
rect 639597 229744 639602 229800
rect 639658 229744 673826 229800
rect 673882 229744 673887 229800
rect 639597 229742 673887 229744
rect 639597 229739 639663 229742
rect 673821 229739 673887 229742
rect 660941 229530 661007 229533
rect 673637 229530 673703 229533
rect 660941 229528 673703 229530
rect 660941 229472 660946 229528
rect 661002 229472 673642 229528
rect 673698 229472 673703 229528
rect 660941 229470 673703 229472
rect 660941 229467 661007 229470
rect 673637 229467 673703 229470
rect 673941 229530 674007 229533
rect 674230 229530 674236 229532
rect 673941 229528 674236 229530
rect 673941 229472 673946 229528
rect 674002 229472 674236 229528
rect 673941 229470 674236 229472
rect 673941 229467 674007 229470
rect 674230 229468 674236 229470
rect 674300 229468 674306 229532
rect 42425 229394 42491 229397
rect 45829 229394 45895 229397
rect 42425 229392 45895 229394
rect 42425 229336 42430 229392
rect 42486 229336 45834 229392
rect 45890 229336 45895 229392
rect 42425 229334 45895 229336
rect 42425 229331 42491 229334
rect 45829 229331 45895 229334
rect 673913 229258 673979 229261
rect 675109 229258 675175 229261
rect 673913 229256 675175 229258
rect 673913 229200 673918 229256
rect 673974 229200 675114 229256
rect 675170 229200 675175 229256
rect 673913 229198 675175 229200
rect 673913 229195 673979 229198
rect 675109 229195 675175 229198
rect 653397 229122 653463 229125
rect 673729 229122 673795 229125
rect 653397 229120 673795 229122
rect 653397 229064 653402 229120
rect 653458 229064 673734 229120
rect 673790 229064 673795 229120
rect 653397 229062 673795 229064
rect 653397 229059 653463 229062
rect 673729 229059 673795 229062
rect 672809 228850 672875 228853
rect 674966 228850 674972 228852
rect 672809 228848 674972 228850
rect 672809 228792 672814 228848
rect 672870 228792 674972 228848
rect 672809 228790 674972 228792
rect 672809 228787 672875 228790
rect 674966 228788 674972 228790
rect 675036 228788 675042 228852
rect 112989 228578 113055 228581
rect 184933 228578 184999 228581
rect 112989 228576 184999 228578
rect 112989 228520 112994 228576
rect 113050 228520 184938 228576
rect 184994 228520 184999 228576
rect 112989 228518 184999 228520
rect 112989 228515 113055 228518
rect 184933 228515 184999 228518
rect 672809 228578 672875 228581
rect 674782 228578 674788 228580
rect 672809 228576 674788 228578
rect 672809 228520 672814 228576
rect 672870 228520 674788 228576
rect 672809 228518 674788 228520
rect 672809 228515 672875 228518
rect 674782 228516 674788 228518
rect 674852 228516 674858 228580
rect 73705 228306 73771 228309
rect 155309 228306 155375 228309
rect 73705 228304 155375 228306
rect 73705 228248 73710 228304
rect 73766 228248 155314 228304
rect 155370 228248 155375 228304
rect 73705 228246 155375 228248
rect 73705 228243 73771 228246
rect 155309 228243 155375 228246
rect 168925 228306 168991 228309
rect 223573 228306 223639 228309
rect 168925 228304 223639 228306
rect 168925 228248 168930 228304
rect 168986 228248 223578 228304
rect 223634 228248 223639 228304
rect 168925 228246 223639 228248
rect 168925 228243 168991 228246
rect 223573 228243 223639 228246
rect 136541 227490 136607 227493
rect 202965 227490 203031 227493
rect 136541 227488 203031 227490
rect 136541 227432 136546 227488
rect 136602 227432 202970 227488
rect 203026 227432 203031 227488
rect 136541 227430 203031 227432
rect 136541 227427 136607 227430
rect 202965 227427 203031 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 89621 227218 89687 227221
rect 166901 227218 166967 227221
rect 89621 227216 166967 227218
rect 89621 227160 89626 227216
rect 89682 227160 166906 227216
rect 166962 227160 166967 227216
rect 89621 227158 166967 227160
rect 89621 227155 89687 227158
rect 166901 227155 166967 227158
rect 672349 227082 672415 227085
rect 674833 227082 674899 227085
rect 672349 227080 674899 227082
rect 672349 227024 672354 227080
rect 672410 227024 674838 227080
rect 674894 227024 674899 227080
rect 672349 227022 674899 227024
rect 672349 227019 672415 227022
rect 674833 227019 674899 227022
rect 79961 226946 80027 226949
rect 160461 226946 160527 226949
rect 79961 226944 160527 226946
rect 79961 226888 79966 226944
rect 80022 226888 160466 226944
rect 160522 226888 160527 226944
rect 79961 226886 160527 226888
rect 79961 226883 80027 226886
rect 160461 226883 160527 226886
rect 671889 226946 671955 226949
rect 671889 226944 672274 226946
rect 671889 226888 671894 226944
rect 671950 226888 672274 226944
rect 671889 226886 672274 226888
rect 671889 226883 671955 226886
rect 672214 226810 672274 226886
rect 673177 226812 673243 226813
rect 672942 226810 672948 226812
rect 672214 226750 672948 226810
rect 672942 226748 672948 226750
rect 673012 226748 673018 226812
rect 673126 226748 673132 226812
rect 673196 226810 673243 226812
rect 673196 226808 673288 226810
rect 673238 226752 673288 226808
rect 673196 226750 673288 226752
rect 673196 226748 673243 226750
rect 673177 226747 673243 226748
rect 42149 226674 42215 226677
rect 45553 226674 45619 226677
rect 42149 226672 45619 226674
rect 42149 226616 42154 226672
rect 42210 226616 45558 226672
rect 45614 226616 45619 226672
rect 42149 226614 45619 226616
rect 42149 226611 42215 226614
rect 45553 226611 45619 226614
rect 658917 226674 658983 226677
rect 671813 226674 671879 226677
rect 658917 226672 671879 226674
rect 658917 226616 658922 226672
rect 658978 226616 671818 226672
rect 671874 226616 671879 226672
rect 658917 226614 671879 226616
rect 658917 226611 658983 226614
rect 671813 226611 671879 226614
rect 672373 226538 672439 226541
rect 674465 226538 674531 226541
rect 672373 226536 674531 226538
rect 672373 226480 672378 226536
rect 672434 226480 674470 226536
rect 674526 226480 674531 226536
rect 672373 226478 674531 226480
rect 672373 226475 672439 226478
rect 674465 226475 674531 226478
rect 654777 226402 654843 226405
rect 671935 226402 672001 226405
rect 654777 226400 672001 226402
rect 654777 226344 654782 226400
rect 654838 226344 671940 226400
rect 671996 226344 672001 226400
rect 654777 226342 672001 226344
rect 654777 226339 654843 226342
rect 671935 226339 672001 226342
rect 673913 226266 673979 226269
rect 676397 226266 676463 226269
rect 673913 226264 676463 226266
rect 673913 226208 673918 226264
rect 673974 226208 676402 226264
rect 676458 226208 676463 226264
rect 673913 226206 676463 226208
rect 673913 226203 673979 226206
rect 676397 226203 676463 226206
rect 125225 226130 125291 226133
rect 196525 226130 196591 226133
rect 125225 226128 196591 226130
rect 125225 226072 125230 226128
rect 125286 226072 196530 226128
rect 196586 226072 196591 226128
rect 125225 226070 196591 226072
rect 125225 226067 125291 226070
rect 196525 226067 196591 226070
rect 672027 226130 672093 226133
rect 673453 226130 673519 226133
rect 672027 226128 673519 226130
rect 672027 226072 672032 226128
rect 672088 226072 673458 226128
rect 673514 226072 673519 226128
rect 672027 226070 673519 226072
rect 672027 226067 672093 226070
rect 673453 226067 673519 226070
rect 89437 225858 89503 225861
rect 168189 225858 168255 225861
rect 671705 225860 671771 225861
rect 671654 225858 671660 225860
rect 89437 225856 168255 225858
rect 89437 225800 89442 225856
rect 89498 225800 168194 225856
rect 168250 225800 168255 225856
rect 89437 225798 168255 225800
rect 671614 225798 671660 225858
rect 671724 225856 671771 225860
rect 671766 225800 671771 225856
rect 89437 225795 89503 225798
rect 168189 225795 168255 225798
rect 671654 225796 671660 225798
rect 671724 225796 671771 225800
rect 672942 225796 672948 225860
rect 673012 225858 673018 225860
rect 675017 225858 675083 225861
rect 673012 225856 675083 225858
rect 673012 225800 675022 225856
rect 675078 225800 675083 225856
rect 673012 225798 675083 225800
rect 673012 225796 673018 225798
rect 671705 225795 671771 225796
rect 675017 225795 675083 225798
rect 42425 225722 42491 225725
rect 43253 225722 43319 225725
rect 669405 225722 669471 225725
rect 42425 225720 43319 225722
rect 42425 225664 42430 225720
rect 42486 225664 43258 225720
rect 43314 225664 43319 225720
rect 42425 225662 43319 225664
rect 42425 225659 42491 225662
rect 43253 225659 43319 225662
rect 659610 225720 669471 225722
rect 659610 225664 669410 225720
rect 669466 225664 669471 225720
rect 659610 225662 669471 225664
rect 82721 225586 82787 225589
rect 163037 225586 163103 225589
rect 82721 225584 163103 225586
rect 82721 225528 82726 225584
rect 82782 225528 163042 225584
rect 163098 225528 163103 225584
rect 82721 225526 163103 225528
rect 82721 225523 82787 225526
rect 163037 225523 163103 225526
rect 650637 225586 650703 225589
rect 659610 225586 659670 225662
rect 669405 225659 669471 225662
rect 671813 225722 671879 225725
rect 672758 225722 672764 225724
rect 671813 225720 672764 225722
rect 671813 225664 671818 225720
rect 671874 225664 672764 225720
rect 671813 225662 672764 225664
rect 671813 225659 671879 225662
rect 672758 225660 672764 225662
rect 672828 225660 672834 225724
rect 673913 225588 673979 225589
rect 650637 225584 659670 225586
rect 650637 225528 650642 225584
rect 650698 225528 659670 225584
rect 650637 225526 659670 225528
rect 650637 225523 650703 225526
rect 673862 225524 673868 225588
rect 673932 225586 673979 225588
rect 673932 225584 674024 225586
rect 673974 225528 674024 225584
rect 673932 225526 674024 225528
rect 673932 225524 673979 225526
rect 673913 225523 673979 225524
rect 670734 225388 670740 225452
rect 670804 225450 670810 225452
rect 670969 225450 671035 225453
rect 670804 225448 671035 225450
rect 670804 225392 670974 225448
rect 671030 225392 671035 225448
rect 670804 225390 671035 225392
rect 670804 225388 670810 225390
rect 670969 225387 671035 225390
rect 671981 225450 672047 225453
rect 673729 225450 673795 225453
rect 671981 225448 673795 225450
rect 671981 225392 671986 225448
rect 672042 225392 673734 225448
rect 673790 225392 673795 225448
rect 671981 225390 673795 225392
rect 671981 225387 672047 225390
rect 673729 225387 673795 225390
rect 655605 225314 655671 225317
rect 669313 225314 669379 225317
rect 655605 225312 669379 225314
rect 655605 225256 655610 225312
rect 655666 225256 669318 225312
rect 669374 225256 669379 225312
rect 655605 225254 669379 225256
rect 655605 225251 655671 225254
rect 669313 225251 669379 225254
rect 671589 225178 671655 225181
rect 669454 225176 671655 225178
rect 669454 225120 671594 225176
rect 671650 225120 671655 225176
rect 669454 225118 671655 225120
rect 661677 225042 661743 225045
rect 669454 225042 669514 225118
rect 671589 225115 671655 225118
rect 671981 225178 672047 225181
rect 675661 225178 675727 225181
rect 671981 225176 675727 225178
rect 671981 225120 671986 225176
rect 672042 225120 675666 225176
rect 675722 225120 675727 225176
rect 671981 225118 675727 225120
rect 671981 225115 672047 225118
rect 675661 225115 675727 225118
rect 661677 225040 669514 225042
rect 661677 224984 661682 225040
rect 661738 224984 669514 225040
rect 661677 224982 669514 224984
rect 661677 224979 661743 224982
rect 72417 224770 72483 224773
rect 152733 224770 152799 224773
rect 72417 224768 152799 224770
rect 72417 224712 72422 224768
rect 72478 224712 152738 224768
rect 152794 224712 152799 224768
rect 72417 224710 152799 224712
rect 72417 224707 72483 224710
rect 152733 224707 152799 224710
rect 670969 224770 671035 224773
rect 672073 224770 672139 224773
rect 670969 224768 672139 224770
rect 670969 224712 670974 224768
rect 671030 224712 672078 224768
rect 672134 224712 672139 224768
rect 670969 224710 672139 224712
rect 670969 224707 671035 224710
rect 672073 224707 672139 224710
rect 185209 224634 185275 224637
rect 186221 224634 186287 224637
rect 185209 224632 186287 224634
rect 185209 224576 185214 224632
rect 185270 224576 186226 224632
rect 186282 224576 186287 224632
rect 185209 224574 186287 224576
rect 185209 224571 185275 224574
rect 186221 224571 186287 224574
rect 672717 224634 672783 224637
rect 673269 224634 673335 224637
rect 672717 224632 673335 224634
rect 672717 224576 672722 224632
rect 672778 224576 673274 224632
rect 673330 224576 673335 224632
rect 672717 224574 673335 224576
rect 672717 224571 672783 224574
rect 673269 224571 673335 224574
rect 41689 224498 41755 224501
rect 62941 224498 63007 224501
rect 41689 224496 63007 224498
rect 41689 224440 41694 224496
rect 41750 224440 62946 224496
rect 63002 224440 63007 224496
rect 41689 224438 63007 224440
rect 41689 224435 41755 224438
rect 62941 224435 63007 224438
rect 66897 224498 66963 224501
rect 149789 224498 149855 224501
rect 176561 224498 176627 224501
rect 66897 224496 149855 224498
rect 66897 224440 66902 224496
rect 66958 224440 149794 224496
rect 149850 224440 149855 224496
rect 66897 224438 149855 224440
rect 66897 224435 66963 224438
rect 149789 224435 149855 224438
rect 161430 224496 176627 224498
rect 161430 224440 176566 224496
rect 176622 224440 176627 224496
rect 161430 224438 176627 224440
rect 58985 224226 59051 224229
rect 145005 224226 145071 224229
rect 58985 224224 145071 224226
rect 58985 224168 58990 224224
rect 59046 224168 145010 224224
rect 145066 224168 145071 224224
rect 58985 224166 145071 224168
rect 58985 224163 59051 224166
rect 145005 224163 145071 224166
rect 146937 224226 147003 224229
rect 161430 224226 161490 224438
rect 176561 224435 176627 224438
rect 671654 224300 671660 224364
rect 671724 224362 671730 224364
rect 675477 224362 675543 224365
rect 671724 224360 675543 224362
rect 671724 224304 675482 224360
rect 675538 224304 675543 224360
rect 671724 224302 675543 224304
rect 671724 224300 671730 224302
rect 675477 224299 675543 224302
rect 146937 224224 161490 224226
rect 146937 224168 146942 224224
rect 146998 224168 161490 224224
rect 146937 224166 161490 224168
rect 175917 224226 175983 224229
rect 204897 224226 204963 224229
rect 175917 224224 204963 224226
rect 175917 224168 175922 224224
rect 175978 224168 204902 224224
rect 204958 224168 204963 224224
rect 175917 224166 204963 224168
rect 146937 224163 147003 224166
rect 175917 224163 175983 224166
rect 204897 224163 204963 224166
rect 658181 224226 658247 224229
rect 670923 224226 670989 224229
rect 658181 224224 670989 224226
rect 658181 224168 658186 224224
rect 658242 224168 670928 224224
rect 670984 224168 670989 224224
rect 658181 224166 670989 224168
rect 658181 224163 658247 224166
rect 670923 224163 670989 224166
rect 671613 224092 671679 224093
rect 671613 224088 671660 224092
rect 671724 224090 671730 224092
rect 672901 224090 672967 224093
rect 673126 224090 673132 224092
rect 671613 224032 671618 224088
rect 671613 224028 671660 224032
rect 671724 224030 671770 224090
rect 672901 224088 673132 224090
rect 672901 224032 672906 224088
rect 672962 224032 673132 224088
rect 672901 224030 673132 224032
rect 671724 224028 671730 224030
rect 671613 224027 671679 224028
rect 672901 224027 672967 224030
rect 673126 224028 673132 224030
rect 673196 224028 673202 224092
rect 656893 223954 656959 223957
rect 666829 223954 666895 223957
rect 670785 223956 670851 223957
rect 656893 223952 666895 223954
rect 656893 223896 656898 223952
rect 656954 223896 666834 223952
rect 666890 223896 666895 223952
rect 656893 223894 666895 223896
rect 656893 223891 656959 223894
rect 666829 223891 666895 223894
rect 670734 223892 670740 223956
rect 670804 223954 670851 223956
rect 672717 223956 672783 223957
rect 672717 223954 672764 223956
rect 670804 223952 670896 223954
rect 670846 223896 670896 223952
rect 670804 223894 670896 223896
rect 672672 223952 672764 223954
rect 672672 223896 672722 223952
rect 672672 223894 672764 223896
rect 670804 223892 670851 223894
rect 670785 223891 670851 223892
rect 672717 223892 672764 223894
rect 672828 223892 672834 223956
rect 672717 223891 672783 223892
rect 674598 223756 674604 223820
rect 674668 223818 674674 223820
rect 674668 223758 676322 223818
rect 674668 223756 674674 223758
rect 656157 223682 656223 223685
rect 669405 223682 669471 223685
rect 656157 223680 669471 223682
rect 656157 223624 656162 223680
rect 656218 223624 669410 223680
rect 669466 223624 669471 223680
rect 656157 223622 669471 223624
rect 656157 223619 656223 223622
rect 669405 223619 669471 223622
rect 673913 223682 673979 223685
rect 674465 223682 674531 223685
rect 673913 223680 674531 223682
rect 673913 223624 673918 223680
rect 673974 223624 674470 223680
rect 674526 223624 674531 223680
rect 673913 223622 674531 223624
rect 673913 223619 673979 223622
rect 674465 223619 674531 223622
rect 676262 223516 676322 223758
rect 92105 223410 92171 223413
rect 170765 223410 170831 223413
rect 92105 223408 170831 223410
rect 92105 223352 92110 223408
rect 92166 223352 170770 223408
rect 170826 223352 170831 223408
rect 92105 223350 170831 223352
rect 92105 223347 92171 223350
rect 170765 223347 170831 223350
rect 71405 223138 71471 223141
rect 152089 223138 152155 223141
rect 71405 223136 152155 223138
rect 71405 223080 71410 223136
rect 71466 223080 152094 223136
rect 152150 223080 152155 223136
rect 71405 223078 152155 223080
rect 71405 223075 71471 223078
rect 152089 223075 152155 223078
rect 657537 223138 657603 223141
rect 667933 223138 667999 223141
rect 657537 223136 667999 223138
rect 657537 223080 657542 223136
rect 657598 223080 667938 223136
rect 667994 223080 667999 223136
rect 657537 223078 667999 223080
rect 657537 223075 657603 223078
rect 667933 223075 667999 223078
rect 683205 223138 683271 223141
rect 683205 223136 683284 223138
rect 683205 223080 683210 223136
rect 683266 223080 683284 223136
rect 683205 223078 683284 223080
rect 683205 223075 683271 223078
rect 28533 222866 28599 222869
rect 54477 222866 54543 222869
rect 28533 222864 54543 222866
rect 28533 222808 28538 222864
rect 28594 222808 54482 222864
rect 54538 222808 54543 222864
rect 28533 222806 54543 222808
rect 28533 222803 28599 222806
rect 54477 222803 54543 222806
rect 64781 222866 64847 222869
rect 146661 222866 146727 222869
rect 64781 222864 146727 222866
rect 64781 222808 64786 222864
rect 64842 222808 146666 222864
rect 146722 222808 146727 222864
rect 64781 222806 146727 222808
rect 64781 222803 64847 222806
rect 146661 222803 146727 222806
rect 150893 222866 150959 222869
rect 213913 222866 213979 222869
rect 150893 222864 213979 222866
rect 150893 222808 150898 222864
rect 150954 222808 213918 222864
rect 213974 222808 213979 222864
rect 150893 222806 213979 222808
rect 150893 222803 150959 222806
rect 213913 222803 213979 222806
rect 652385 222866 652451 222869
rect 674230 222866 674236 222868
rect 652385 222864 674236 222866
rect 652385 222808 652390 222864
rect 652446 222808 674236 222864
rect 652385 222806 674236 222808
rect 652385 222803 652451 222806
rect 674230 222804 674236 222806
rect 674300 222804 674306 222868
rect 674465 222730 674531 222733
rect 675886 222730 675892 222732
rect 674465 222728 675892 222730
rect 674465 222672 674470 222728
rect 674526 222672 675892 222728
rect 674465 222670 675892 222672
rect 674465 222667 674531 222670
rect 675886 222668 675892 222670
rect 675956 222668 675962 222732
rect 683665 222730 683731 222733
rect 683652 222728 683731 222730
rect 683652 222672 683670 222728
rect 683726 222672 683731 222728
rect 683652 222670 683731 222672
rect 683665 222667 683731 222670
rect 563329 222322 563395 222325
rect 571885 222322 571951 222325
rect 563329 222320 571951 222322
rect 563329 222264 563334 222320
rect 563390 222264 571890 222320
rect 571946 222264 571951 222320
rect 563329 222262 571951 222264
rect 563329 222259 563395 222262
rect 571885 222259 571951 222262
rect 674281 222322 674347 222325
rect 674281 222320 676292 222322
rect 674281 222264 674286 222320
rect 674342 222264 676292 222320
rect 674281 222262 676292 222264
rect 674281 222259 674347 222262
rect 108665 222050 108731 222053
rect 183645 222050 183711 222053
rect 108665 222048 183711 222050
rect 108665 221992 108670 222048
rect 108726 221992 183650 222048
rect 183706 221992 183711 222048
rect 108665 221990 183711 221992
rect 108665 221987 108731 221990
rect 183645 221987 183711 221990
rect 513557 222050 513623 222053
rect 599485 222050 599551 222053
rect 513557 222048 599551 222050
rect 513557 221992 513562 222048
rect 513618 221992 599490 222048
rect 599546 221992 599551 222048
rect 513557 221990 599551 221992
rect 513557 221987 513623 221990
rect 599485 221987 599551 221990
rect 660757 222050 660823 222053
rect 667933 222050 667999 222053
rect 660757 222048 667999 222050
rect 660757 221992 660762 222048
rect 660818 221992 667938 222048
rect 667994 221992 667999 222048
rect 660757 221990 667999 221992
rect 660757 221987 660823 221990
rect 667933 221987 667999 221990
rect 672441 221916 672507 221917
rect 672390 221914 672396 221916
rect 672350 221854 672396 221914
rect 672460 221912 672507 221916
rect 672502 221856 672507 221912
rect 672390 221852 672396 221854
rect 672460 221852 672507 221856
rect 672441 221851 672507 221852
rect 673361 221914 673427 221917
rect 673361 221912 676292 221914
rect 673361 221856 673366 221912
rect 673422 221856 676292 221912
rect 673361 221854 676292 221856
rect 673361 221851 673427 221854
rect 97717 221778 97783 221781
rect 172697 221778 172763 221781
rect 97717 221776 172763 221778
rect 97717 221720 97722 221776
rect 97778 221720 172702 221776
rect 172758 221720 172763 221776
rect 97717 221718 172763 221720
rect 97717 221715 97783 221718
rect 172697 221715 172763 221718
rect 530853 221778 530919 221781
rect 603349 221778 603415 221781
rect 530853 221776 603415 221778
rect 530853 221720 530858 221776
rect 530914 221720 603354 221776
rect 603410 221720 603415 221776
rect 530853 221718 603415 221720
rect 530853 221715 530919 221718
rect 603349 221715 603415 221718
rect 664161 221778 664227 221781
rect 664161 221776 671652 221778
rect 664161 221720 664166 221776
rect 664222 221720 671652 221776
rect 664161 221718 671652 221720
rect 664161 221715 664227 221718
rect 671592 221642 671652 221718
rect 674833 221642 674899 221645
rect 671592 221640 674899 221642
rect 671592 221584 674838 221640
rect 674894 221584 674899 221640
rect 671592 221582 674899 221584
rect 674833 221579 674899 221582
rect 95417 221506 95483 221509
rect 172973 221506 173039 221509
rect 95417 221504 173039 221506
rect 95417 221448 95422 221504
rect 95478 221448 172978 221504
rect 173034 221448 173039 221504
rect 95417 221446 173039 221448
rect 95417 221443 95483 221446
rect 172973 221443 173039 221446
rect 521009 221506 521075 221509
rect 600313 221506 600379 221509
rect 521009 221504 600379 221506
rect 521009 221448 521014 221504
rect 521070 221448 600318 221504
rect 600374 221448 600379 221504
rect 521009 221446 600379 221448
rect 521009 221443 521075 221446
rect 600313 221443 600379 221446
rect 653029 221506 653095 221509
rect 671429 221506 671495 221509
rect 679801 221506 679867 221509
rect 653029 221504 671495 221506
rect 653029 221448 653034 221504
rect 653090 221448 671434 221504
rect 671490 221448 671495 221504
rect 653029 221446 671495 221448
rect 679788 221504 679867 221506
rect 679788 221448 679806 221504
rect 679862 221448 679867 221504
rect 679788 221446 679867 221448
rect 653029 221443 653095 221446
rect 671429 221443 671495 221446
rect 679801 221443 679867 221446
rect 171041 221234 171107 221237
rect 229553 221234 229619 221237
rect 171041 221232 229619 221234
rect 171041 221176 171046 221232
rect 171102 221176 229558 221232
rect 229614 221176 229619 221232
rect 171041 221174 229619 221176
rect 171041 221171 171107 221174
rect 229553 221171 229619 221174
rect 515765 221234 515831 221237
rect 600773 221234 600839 221237
rect 515765 221232 600839 221234
rect 515765 221176 515770 221232
rect 515826 221176 600778 221232
rect 600834 221176 600839 221232
rect 515765 221174 600839 221176
rect 515765 221171 515831 221174
rect 600773 221171 600839 221174
rect 671889 221234 671955 221237
rect 671889 221232 675034 221234
rect 671889 221176 671894 221232
rect 671950 221176 675034 221232
rect 671889 221174 675034 221176
rect 671889 221171 671955 221174
rect 674974 221098 675034 221174
rect 674974 221038 676292 221098
rect 517513 220962 517579 220965
rect 518525 220962 518591 220965
rect 600589 220962 600655 220965
rect 517513 220960 600655 220962
rect 517513 220904 517518 220960
rect 517574 220904 518530 220960
rect 518586 220904 600594 220960
rect 600650 220904 600655 220960
rect 517513 220902 600655 220904
rect 517513 220899 517579 220902
rect 518525 220899 518591 220902
rect 600589 220899 600655 220902
rect 667933 220962 667999 220965
rect 672901 220962 672967 220965
rect 673126 220962 673132 220964
rect 667933 220960 672642 220962
rect 667933 220904 667938 220960
rect 667994 220904 672642 220960
rect 667933 220902 672642 220904
rect 667933 220899 667999 220902
rect 147581 220690 147647 220693
rect 211337 220690 211403 220693
rect 672582 220690 672642 220902
rect 672901 220960 673132 220962
rect 672901 220904 672906 220960
rect 672962 220904 673132 220960
rect 672901 220902 673132 220904
rect 672901 220899 672967 220902
rect 673126 220900 673132 220902
rect 673196 220900 673202 220964
rect 674782 220962 674788 220964
rect 673318 220902 674788 220962
rect 673318 220690 673378 220902
rect 674782 220900 674788 220902
rect 674852 220900 674858 220964
rect 679617 220690 679683 220693
rect 147581 220688 211403 220690
rect 147581 220632 147586 220688
rect 147642 220632 211342 220688
rect 211398 220632 211403 220688
rect 147581 220630 211403 220632
rect 147581 220627 147647 220630
rect 211337 220627 211403 220630
rect 663750 220630 669330 220690
rect 672582 220630 673378 220690
rect 679604 220688 679683 220690
rect 679604 220632 679622 220688
rect 679678 220632 679683 220688
rect 679604 220630 679683 220632
rect 522573 220554 522639 220557
rect 618805 220554 618871 220557
rect 522573 220552 618871 220554
rect 522573 220496 522578 220552
rect 522634 220496 618810 220552
rect 618866 220496 618871 220552
rect 522573 220494 618871 220496
rect 522573 220491 522639 220494
rect 618805 220491 618871 220494
rect 124397 220418 124463 220421
rect 193305 220418 193371 220421
rect 124397 220416 193371 220418
rect 124397 220360 124402 220416
rect 124458 220360 193310 220416
rect 193366 220360 193371 220416
rect 124397 220358 193371 220360
rect 124397 220355 124463 220358
rect 193305 220355 193371 220358
rect 646129 220418 646195 220421
rect 663750 220418 663810 220630
rect 646129 220416 663810 220418
rect 646129 220360 646134 220416
rect 646190 220360 663810 220416
rect 646129 220358 663810 220360
rect 669270 220418 669330 220630
rect 679617 220627 679683 220630
rect 675017 220554 675083 220557
rect 673502 220552 675083 220554
rect 673502 220496 675022 220552
rect 675078 220496 675083 220552
rect 673502 220494 675083 220496
rect 673502 220418 673562 220494
rect 675017 220491 675083 220494
rect 669270 220358 673562 220418
rect 646129 220355 646195 220358
rect 527541 220282 527607 220285
rect 619633 220282 619699 220285
rect 527541 220280 619699 220282
rect 527541 220224 527546 220280
rect 527602 220224 619638 220280
rect 619694 220224 619699 220280
rect 527541 220222 619699 220224
rect 527541 220219 527607 220222
rect 619633 220219 619699 220222
rect 674649 220282 674715 220285
rect 674649 220280 676292 220282
rect 674649 220224 674654 220280
rect 674710 220224 676292 220280
rect 674649 220222 676292 220224
rect 674649 220219 674715 220222
rect 117773 220146 117839 220149
rect 187877 220146 187943 220149
rect 117773 220144 187943 220146
rect 117773 220088 117778 220144
rect 117834 220088 187882 220144
rect 187938 220088 187943 220144
rect 117773 220086 187943 220088
rect 117773 220083 117839 220086
rect 187877 220083 187943 220086
rect 637573 220146 637639 220149
rect 674046 220146 674052 220148
rect 637573 220144 674052 220146
rect 637573 220088 637578 220144
rect 637634 220088 674052 220144
rect 637573 220086 674052 220088
rect 637573 220083 637639 220086
rect 674046 220084 674052 220086
rect 674116 220084 674122 220148
rect 524965 220010 525031 220013
rect 530025 220010 530091 220013
rect 620461 220010 620527 220013
rect 524965 220008 529122 220010
rect 524965 219952 524970 220008
rect 525026 219952 529122 220008
rect 524965 219950 529122 219952
rect 524965 219947 525031 219950
rect 518893 219740 518959 219741
rect 518893 219736 518940 219740
rect 519004 219738 519010 219740
rect 528461 219738 528527 219741
rect 528870 219738 528876 219740
rect 518893 219680 518898 219736
rect 518893 219676 518940 219680
rect 519004 219678 519050 219738
rect 528461 219736 528876 219738
rect 528461 219680 528466 219736
rect 528522 219680 528876 219736
rect 528461 219678 528876 219680
rect 519004 219676 519010 219678
rect 518893 219675 518959 219676
rect 528461 219675 528527 219678
rect 528870 219676 528876 219678
rect 528940 219676 528946 219740
rect 529062 219738 529122 219950
rect 530025 220008 620527 220010
rect 530025 219952 530030 220008
rect 530086 219952 620466 220008
rect 620522 219952 620527 220008
rect 530025 219950 620527 219952
rect 530025 219947 530091 219950
rect 620461 219947 620527 219950
rect 648613 219874 648679 219877
rect 673545 219874 673611 219877
rect 648613 219872 673611 219874
rect 648613 219816 648618 219872
rect 648674 219816 673550 219872
rect 673606 219816 673611 219872
rect 648613 219814 673611 219816
rect 648613 219811 648679 219814
rect 673545 219811 673611 219814
rect 675109 219874 675175 219877
rect 676029 219874 676095 219877
rect 675109 219872 676095 219874
rect 675109 219816 675114 219872
rect 675170 219816 676034 219872
rect 676090 219816 676095 219872
rect 675109 219814 676095 219816
rect 675109 219811 675175 219814
rect 676029 219811 676095 219814
rect 683389 219874 683455 219877
rect 683389 219872 683468 219874
rect 683389 219816 683394 219872
rect 683450 219816 683468 219872
rect 683389 219814 683468 219816
rect 683389 219811 683455 219814
rect 619817 219738 619883 219741
rect 529062 219736 619883 219738
rect 529062 219680 619822 219736
rect 619878 219680 619883 219736
rect 529062 219678 619883 219680
rect 619817 219675 619883 219678
rect 491937 219466 492003 219469
rect 553117 219466 553183 219469
rect 562358 219466 562364 219468
rect 491937 219464 553183 219466
rect 491937 219408 491942 219464
rect 491998 219408 553122 219464
rect 553178 219408 553183 219464
rect 491937 219406 553183 219408
rect 491937 219403 492003 219406
rect 553117 219403 553183 219406
rect 554086 219406 562364 219466
rect 554086 219330 554146 219406
rect 562358 219404 562364 219406
rect 562428 219404 562434 219468
rect 562734 219466 563070 219500
rect 562550 219440 563070 219466
rect 562550 219406 562794 219440
rect 563010 219432 563070 219440
rect 553902 219270 554146 219330
rect 494697 219194 494763 219197
rect 505093 219194 505159 219197
rect 494697 219192 505159 219194
rect 494697 219136 494702 219192
rect 494758 219136 505098 219192
rect 505154 219136 505159 219192
rect 494697 219134 505159 219136
rect 494697 219131 494763 219134
rect 505093 219131 505159 219134
rect 505277 219194 505343 219197
rect 533889 219194 533955 219197
rect 534073 219194 534139 219197
rect 505277 219192 533722 219194
rect 505277 219136 505282 219192
rect 505338 219163 533722 219192
rect 533889 219192 534139 219194
rect 505338 219158 533771 219163
rect 505338 219136 533710 219158
rect 505277 219134 533710 219136
rect 505277 219131 505343 219134
rect 533662 219102 533710 219134
rect 533766 219102 533771 219158
rect 533889 219136 533894 219192
rect 533950 219136 534078 219192
rect 534134 219136 534139 219192
rect 533889 219134 534139 219136
rect 533889 219131 533955 219134
rect 534073 219131 534139 219134
rect 534257 219194 534323 219197
rect 553902 219194 553962 219270
rect 534257 219192 553962 219194
rect 534257 219136 534262 219192
rect 534318 219136 553962 219192
rect 534257 219134 553962 219136
rect 554221 219194 554287 219197
rect 562550 219194 562610 219406
rect 563010 219372 563346 219432
rect 563462 219404 563468 219468
rect 563532 219466 563538 219468
rect 571926 219466 571932 219468
rect 563532 219406 571932 219466
rect 563532 219404 563538 219406
rect 571926 219404 571932 219406
rect 571996 219404 572002 219468
rect 594149 219466 594215 219469
rect 621289 219466 621355 219469
rect 572486 219406 591682 219466
rect 554221 219192 562610 219194
rect 554221 219136 554226 219192
rect 554282 219136 562610 219192
rect 554221 219134 562610 219136
rect 563286 219194 563346 219372
rect 572486 219330 572546 219406
rect 572118 219270 572546 219330
rect 572118 219194 572178 219270
rect 563286 219134 572178 219194
rect 534257 219131 534323 219134
rect 554221 219131 554287 219134
rect 572846 219132 572852 219196
rect 572916 219194 572922 219196
rect 591389 219194 591455 219197
rect 572916 219192 591455 219194
rect 572916 219136 591394 219192
rect 591450 219136 591455 219192
rect 572916 219134 591455 219136
rect 591622 219194 591682 219406
rect 594149 219464 621355 219466
rect 594149 219408 594154 219464
rect 594210 219408 621294 219464
rect 621350 219408 621355 219464
rect 594149 219406 621355 219408
rect 594149 219403 594215 219406
rect 621289 219403 621355 219406
rect 673545 219466 673611 219469
rect 673545 219464 676292 219466
rect 673545 219408 673550 219464
rect 673606 219408 676292 219464
rect 673545 219406 676292 219408
rect 673545 219403 673611 219406
rect 595161 219194 595227 219197
rect 591622 219192 595227 219194
rect 591622 219136 595166 219192
rect 595222 219136 595227 219192
rect 591622 219134 595227 219136
rect 572916 219132 572922 219134
rect 591389 219131 591455 219134
rect 595161 219131 595227 219134
rect 651281 219194 651347 219197
rect 672717 219194 672783 219197
rect 651281 219192 672783 219194
rect 651281 219136 651286 219192
rect 651342 219136 672722 219192
rect 672778 219136 672783 219192
rect 651281 219134 672783 219136
rect 651281 219131 651347 219134
rect 672717 219131 672783 219134
rect 533662 219100 533771 219102
rect 533705 219097 533771 219100
rect 675518 218996 675524 219060
rect 675588 219058 675594 219060
rect 675588 218998 676292 219058
rect 675588 218996 675594 218998
rect 493685 218922 493751 218925
rect 499205 218922 499271 218925
rect 493685 218920 499271 218922
rect 493685 218864 493690 218920
rect 493746 218864 499210 218920
rect 499266 218864 499271 218920
rect 493685 218862 499271 218864
rect 493685 218859 493751 218862
rect 499205 218859 499271 218862
rect 499430 218860 499436 218924
rect 499500 218922 499506 218924
rect 567837 218922 567903 218925
rect 499500 218920 567903 218922
rect 499500 218864 567842 218920
rect 567898 218864 567903 218920
rect 499500 218862 567903 218864
rect 499500 218860 499506 218862
rect 567837 218859 567903 218862
rect 568297 218922 568363 218925
rect 572478 218922 572484 218924
rect 568297 218920 572484 218922
rect 568297 218864 568302 218920
rect 568358 218864 572484 218920
rect 568297 218862 572484 218864
rect 568297 218859 568363 218862
rect 572478 218860 572484 218862
rect 572548 218860 572554 218924
rect 572713 218922 572779 218925
rect 641161 218922 641227 218925
rect 675109 218922 675175 218925
rect 572713 218920 611370 218922
rect 572713 218864 572718 218920
rect 572774 218864 611370 218920
rect 572713 218862 611370 218864
rect 572713 218859 572779 218862
rect 77201 218650 77267 218653
rect 157701 218650 157767 218653
rect 77201 218648 157767 218650
rect 77201 218592 77206 218648
rect 77262 218592 157706 218648
rect 157762 218592 157767 218648
rect 77201 218590 157767 218592
rect 77201 218587 77267 218590
rect 157701 218587 157767 218590
rect 159817 218650 159883 218653
rect 200757 218650 200823 218653
rect 159817 218648 200823 218650
rect 159817 218592 159822 218648
rect 159878 218592 200762 218648
rect 200818 218592 200823 218648
rect 159817 218590 200823 218592
rect 159817 218587 159883 218590
rect 200757 218587 200823 218590
rect 490281 218650 490347 218653
rect 496670 218650 496676 218652
rect 490281 218648 496676 218650
rect 490281 218592 490286 218648
rect 490342 218592 496676 218648
rect 490281 218590 496676 218592
rect 490281 218587 490347 218590
rect 496670 218588 496676 218590
rect 496740 218588 496746 218652
rect 496997 218650 497063 218653
rect 497549 218650 497615 218653
rect 602061 218650 602127 218653
rect 496997 218648 602127 218650
rect 496997 218592 497002 218648
rect 497058 218592 497554 218648
rect 497610 218592 602066 218648
rect 602122 218592 602127 218648
rect 496997 218590 602127 218592
rect 611310 218650 611370 218862
rect 641161 218920 675175 218922
rect 641161 218864 641166 218920
rect 641222 218864 675114 218920
rect 675170 218864 675175 218920
rect 641161 218862 675175 218864
rect 641161 218859 641227 218862
rect 675109 218859 675175 218862
rect 630673 218650 630739 218653
rect 611310 218648 630739 218650
rect 611310 218592 630678 218648
rect 630734 218592 630739 218648
rect 611310 218590 630739 218592
rect 496997 218587 497063 218590
rect 497549 218587 497615 218590
rect 602061 218587 602127 218590
rect 630673 218587 630739 218590
rect 666318 218588 666324 218652
rect 666388 218650 666394 218652
rect 666388 218590 676292 218650
rect 666388 218588 666394 218590
rect 487797 218378 487863 218381
rect 499573 218378 499639 218381
rect 487797 218376 499639 218378
rect 487797 218320 487802 218376
rect 487858 218320 499578 218376
rect 499634 218320 499639 218376
rect 487797 218318 499639 218320
rect 487797 218315 487863 218318
rect 499573 218315 499639 218318
rect 499757 218378 499823 218381
rect 567653 218378 567719 218381
rect 499757 218376 567719 218378
rect 499757 218320 499762 218376
rect 499818 218320 567658 218376
rect 567714 218320 567719 218376
rect 499757 218318 567719 218320
rect 499757 218315 499823 218318
rect 567653 218315 567719 218318
rect 567837 218378 567903 218381
rect 572437 218378 572503 218381
rect 567837 218376 572503 218378
rect 567837 218320 567842 218376
rect 567898 218320 572442 218376
rect 572498 218320 572503 218376
rect 567837 218318 572503 218320
rect 567837 218315 567903 218318
rect 572437 218315 572503 218318
rect 572621 218378 572687 218381
rect 612733 218378 612799 218381
rect 572621 218376 612799 218378
rect 572621 218320 572626 218376
rect 572682 218320 612738 218376
rect 612794 218320 612799 218376
rect 572621 218318 612799 218320
rect 572621 218315 572687 218318
rect 612733 218315 612799 218318
rect 643829 218378 643895 218381
rect 673177 218378 673243 218381
rect 643829 218376 673243 218378
rect 643829 218320 643834 218376
rect 643890 218320 673182 218376
rect 673238 218320 673243 218376
rect 643829 218318 673243 218320
rect 643829 218315 643895 218318
rect 673177 218315 673243 218318
rect 676024 218180 676030 218244
rect 676094 218242 676100 218244
rect 676094 218182 676292 218242
rect 676094 218180 676100 218182
rect 484577 218106 484643 218109
rect 485037 218106 485103 218109
rect 518893 218106 518959 218109
rect 484577 218104 518959 218106
rect 484577 218048 484582 218104
rect 484638 218048 485042 218104
rect 485098 218048 518898 218104
rect 518954 218048 518959 218104
rect 484577 218046 518959 218048
rect 484577 218043 484643 218046
rect 485037 218043 485103 218046
rect 518893 218043 518959 218046
rect 519077 218106 519143 218109
rect 524413 218106 524479 218109
rect 519077 218104 524479 218106
rect 519077 218048 519082 218104
rect 519138 218048 524418 218104
rect 524474 218048 524479 218104
rect 519077 218046 524479 218048
rect 519077 218043 519143 218046
rect 524413 218043 524479 218046
rect 524597 218106 524663 218109
rect 572989 218106 573055 218109
rect 524597 218104 573055 218106
rect 524597 218048 524602 218104
rect 524658 218048 572994 218104
rect 573050 218048 573055 218104
rect 524597 218046 573055 218048
rect 524597 218043 524663 218046
rect 572989 218043 573055 218046
rect 573214 218044 573220 218108
rect 573284 218106 573290 218108
rect 582097 218106 582163 218109
rect 573284 218104 582163 218106
rect 573284 218048 582102 218104
rect 582158 218048 582163 218104
rect 573284 218046 582163 218048
rect 573284 218044 573290 218046
rect 582097 218043 582163 218046
rect 582281 218106 582347 218109
rect 627729 218106 627795 218109
rect 675201 218106 675267 218109
rect 582281 218104 627795 218106
rect 582281 218048 582286 218104
rect 582342 218048 627734 218104
rect 627790 218048 627795 218104
rect 582281 218046 627795 218048
rect 582281 218043 582347 218046
rect 627729 218043 627795 218046
rect 672376 218104 675267 218106
rect 672376 218048 675206 218104
rect 675262 218048 675267 218104
rect 672376 218046 675267 218048
rect 672376 217970 672436 218046
rect 675201 218043 675267 218046
rect 669270 217910 672436 217970
rect 499205 217834 499271 217837
rect 499757 217834 499823 217837
rect 499205 217832 499823 217834
rect 499205 217776 499210 217832
rect 499266 217776 499762 217832
rect 499818 217776 499823 217832
rect 499205 217774 499823 217776
rect 499205 217771 499271 217774
rect 499757 217771 499823 217774
rect 507761 217834 507827 217837
rect 510981 217834 511047 217837
rect 514937 217834 515003 217837
rect 507761 217832 509434 217834
rect 507761 217776 507766 217832
rect 507822 217776 509434 217832
rect 507761 217774 509434 217776
rect 507761 217771 507827 217774
rect 501045 217564 501111 217565
rect 501045 217562 501092 217564
rect 501000 217560 501092 217562
rect 501000 217504 501050 217560
rect 501000 217502 501092 217504
rect 501045 217500 501092 217502
rect 501156 217500 501162 217564
rect 502977 217562 503043 217565
rect 503345 217564 503411 217565
rect 503294 217562 503300 217564
rect 502977 217560 503300 217562
rect 503364 217562 503411 217564
rect 503621 217564 503687 217565
rect 503621 217562 503668 217564
rect 503364 217560 503456 217562
rect 502977 217504 502982 217560
rect 503038 217504 503300 217560
rect 503406 217504 503456 217560
rect 502977 217502 503300 217504
rect 501045 217499 501111 217500
rect 502977 217499 503043 217502
rect 503294 217500 503300 217502
rect 503364 217502 503456 217504
rect 503576 217560 503668 217562
rect 503576 217504 503626 217560
rect 503576 217502 503668 217504
rect 503364 217500 503411 217502
rect 503345 217499 503411 217500
rect 503621 217500 503668 217502
rect 503732 217500 503738 217564
rect 505461 217562 505527 217565
rect 506105 217564 506171 217565
rect 506054 217562 506060 217564
rect 505461 217560 506060 217562
rect 506124 217562 506171 217564
rect 508681 217562 508747 217565
rect 509182 217562 509188 217564
rect 506124 217560 506216 217562
rect 505461 217504 505466 217560
rect 505522 217504 506060 217560
rect 506166 217504 506216 217560
rect 505461 217502 506060 217504
rect 503621 217499 503687 217500
rect 505461 217499 505527 217502
rect 506054 217500 506060 217502
rect 506124 217502 506216 217504
rect 508681 217560 509188 217562
rect 508681 217504 508686 217560
rect 508742 217504 509188 217560
rect 508681 217502 509188 217504
rect 506124 217500 506171 217502
rect 506105 217499 506171 217500
rect 508681 217499 508747 217502
rect 509182 217500 509188 217502
rect 509252 217500 509258 217564
rect 509374 217562 509434 217774
rect 510981 217832 515003 217834
rect 510981 217776 510986 217832
rect 511042 217776 514942 217832
rect 514998 217776 515003 217832
rect 510981 217774 515003 217776
rect 510981 217771 511047 217774
rect 514937 217771 515003 217774
rect 515121 217834 515187 217837
rect 518341 217834 518407 217837
rect 515121 217832 518407 217834
rect 515121 217776 515126 217832
rect 515182 217776 518346 217832
rect 518402 217776 518407 217832
rect 515121 217774 518407 217776
rect 515121 217771 515187 217774
rect 518341 217771 518407 217774
rect 518709 217834 518775 217837
rect 591849 217834 591915 217837
rect 518709 217832 591915 217834
rect 518709 217776 518714 217832
rect 518770 217776 591854 217832
rect 591910 217776 591915 217832
rect 518709 217774 591915 217776
rect 518709 217771 518775 217774
rect 591849 217771 591915 217774
rect 592166 217772 592172 217836
rect 592236 217834 592242 217836
rect 597553 217834 597619 217837
rect 592236 217832 597619 217834
rect 592236 217776 597558 217832
rect 597614 217776 597619 217832
rect 592236 217774 597619 217776
rect 592236 217772 592242 217774
rect 597553 217771 597619 217774
rect 644933 217834 644999 217837
rect 669270 217834 669330 217910
rect 644933 217832 669330 217834
rect 644933 217776 644938 217832
rect 644994 217776 669330 217832
rect 644933 217774 669330 217776
rect 674833 217834 674899 217837
rect 674833 217832 676292 217834
rect 674833 217776 674838 217832
rect 674894 217776 676292 217832
rect 674833 217774 676292 217776
rect 644933 217771 644999 217774
rect 674833 217771 674899 217774
rect 674598 217698 674604 217700
rect 669454 217638 674604 217698
rect 518893 217562 518959 217565
rect 509374 217560 518959 217562
rect 509374 217504 518898 217560
rect 518954 217504 518959 217560
rect 509374 217502 518959 217504
rect 518893 217499 518959 217502
rect 519077 217562 519143 217565
rect 563053 217562 563119 217565
rect 519077 217560 563119 217562
rect 519077 217504 519082 217560
rect 519138 217504 563058 217560
rect 563114 217504 563119 217560
rect 519077 217502 563119 217504
rect 519077 217499 519143 217502
rect 563053 217499 563119 217502
rect 563237 217562 563303 217565
rect 572253 217562 572319 217565
rect 563237 217560 572319 217562
rect 563237 217504 563242 217560
rect 563298 217504 572258 217560
rect 572314 217504 572319 217560
rect 563237 217502 572319 217504
rect 563237 217499 563303 217502
rect 572253 217499 572319 217502
rect 572897 217562 572963 217565
rect 582097 217562 582163 217565
rect 572897 217560 582163 217562
rect 572897 217504 572902 217560
rect 572958 217504 582102 217560
rect 582158 217504 582163 217560
rect 572897 217502 582163 217504
rect 572897 217499 572963 217502
rect 582097 217499 582163 217502
rect 582281 217562 582347 217565
rect 606753 217562 606819 217565
rect 617793 217562 617859 217565
rect 582281 217560 606586 217562
rect 582281 217504 582286 217560
rect 582342 217504 606586 217560
rect 582281 217502 606586 217504
rect 582281 217499 582347 217502
rect 495249 217290 495315 217293
rect 582373 217290 582439 217293
rect 591798 217290 591804 217292
rect 495249 217288 582439 217290
rect 495249 217232 495254 217288
rect 495310 217232 582378 217288
rect 582434 217232 582439 217288
rect 495249 217230 582439 217232
rect 495249 217227 495315 217230
rect 582373 217227 582439 217230
rect 582790 217230 591804 217290
rect 489085 217154 489151 217157
rect 582790 217154 582850 217230
rect 591798 217228 591804 217230
rect 591868 217228 591874 217292
rect 606526 217290 606586 217502
rect 606753 217560 617859 217562
rect 606753 217504 606758 217560
rect 606814 217504 617798 217560
rect 617854 217504 617859 217560
rect 606753 217502 617859 217504
rect 606753 217499 606819 217502
rect 617793 217499 617859 217502
rect 639965 217562 640031 217565
rect 669454 217562 669514 217638
rect 674598 217636 674604 217638
rect 674668 217636 674674 217700
rect 639965 217560 669514 217562
rect 639965 217504 639970 217560
rect 640026 217504 669514 217560
rect 639965 217502 669514 217504
rect 639965 217499 640031 217502
rect 674465 217426 674531 217429
rect 674465 217424 676292 217426
rect 674465 217368 674470 217424
rect 674526 217368 676292 217424
rect 674465 217366 676292 217368
rect 674465 217363 674531 217366
rect 617241 217290 617307 217293
rect 591990 217230 601710 217290
rect 606526 217288 617307 217290
rect 606526 217232 617246 217288
rect 617302 217232 617307 217288
rect 606526 217230 617307 217232
rect 489085 217152 491218 217154
rect 489085 217096 489090 217152
rect 489146 217096 491218 217152
rect 489085 217094 491218 217096
rect 489085 217091 489151 217094
rect 491158 216746 491218 217094
rect 582606 217094 582850 217154
rect 503294 216956 503300 217020
rect 503364 217018 503370 217020
rect 582606 217018 582666 217094
rect 503364 216958 582666 217018
rect 582925 217018 582991 217021
rect 586646 217018 586652 217020
rect 582925 217016 586652 217018
rect 582925 216960 582930 217016
rect 582986 216960 586652 217016
rect 582925 216958 586652 216960
rect 503364 216956 503370 216958
rect 582925 216955 582991 216958
rect 586646 216956 586652 216958
rect 586716 216956 586722 217020
rect 586881 217018 586947 217021
rect 591990 217018 592050 217230
rect 586881 217016 592050 217018
rect 586881 216960 586886 217016
rect 586942 216960 592050 217016
rect 586881 216958 592050 216960
rect 592217 217018 592283 217021
rect 595713 217018 595779 217021
rect 592217 217016 595779 217018
rect 592217 216960 592222 217016
rect 592278 216960 595718 217016
rect 595774 216960 595779 217016
rect 592217 216958 595779 216960
rect 601650 217018 601710 217230
rect 617241 217227 617307 217230
rect 656525 217290 656591 217293
rect 672073 217290 672139 217293
rect 656525 217288 672139 217290
rect 656525 217232 656530 217288
rect 656586 217232 672078 217288
rect 672134 217232 672139 217288
rect 656525 217230 672139 217232
rect 656525 217227 656591 217230
rect 672073 217227 672139 217230
rect 606753 217018 606819 217021
rect 601650 217016 606819 217018
rect 601650 216960 606758 217016
rect 606814 216960 606819 217016
rect 601650 216958 606819 216960
rect 586881 216955 586947 216958
rect 592217 216955 592283 216958
rect 595713 216955 595779 216958
rect 606753 216955 606819 216958
rect 675886 216956 675892 217020
rect 675956 217018 675962 217020
rect 675956 216958 676292 217018
rect 675956 216956 675962 216958
rect 594793 216746 594859 216749
rect 491158 216744 594859 216746
rect 491158 216688 594798 216744
rect 594854 216688 594859 216744
rect 491158 216686 594859 216688
rect 594793 216683 594859 216686
rect 594977 216746 595043 216749
rect 599025 216746 599091 216749
rect 594977 216744 599091 216746
rect 594977 216688 594982 216744
rect 595038 216688 599030 216744
rect 599086 216688 599091 216744
rect 594977 216686 599091 216688
rect 594977 216683 595043 216686
rect 599025 216683 599091 216686
rect 669405 216610 669471 216613
rect 669405 216608 676292 216610
rect 669405 216552 669410 216608
rect 669466 216552 676292 216608
rect 669405 216550 676292 216552
rect 669405 216547 669471 216550
rect 518934 216412 518940 216476
rect 519004 216474 519010 216476
rect 528686 216474 528692 216476
rect 519004 216414 528692 216474
rect 519004 216412 519010 216414
rect 528686 216412 528692 216414
rect 528756 216412 528762 216476
rect 528870 216412 528876 216476
rect 528940 216474 528946 216476
rect 618345 216474 618411 216477
rect 528940 216472 618411 216474
rect 528940 216416 618350 216472
rect 618406 216416 618411 216472
rect 528940 216414 618411 216416
rect 528940 216412 528946 216414
rect 618345 216411 618411 216414
rect 503662 216140 503668 216204
rect 503732 216202 503738 216204
rect 596357 216202 596423 216205
rect 503732 216200 596423 216202
rect 503732 216144 596362 216200
rect 596418 216144 596423 216200
rect 503732 216142 596423 216144
rect 503732 216140 503738 216142
rect 596357 216139 596423 216142
rect 646589 216202 646655 216205
rect 675201 216202 675267 216205
rect 646589 216200 669330 216202
rect 646589 216144 646594 216200
rect 646650 216144 669330 216200
rect 646589 216142 669330 216144
rect 646589 216139 646655 216142
rect 501086 215868 501092 215932
rect 501156 215930 501162 215932
rect 582373 215930 582439 215933
rect 501156 215928 582439 215930
rect 501156 215872 582378 215928
rect 582434 215872 582439 215928
rect 501156 215870 582439 215872
rect 501156 215868 501162 215870
rect 582373 215867 582439 215870
rect 582557 215930 582623 215933
rect 611721 215930 611787 215933
rect 582557 215928 611787 215930
rect 582557 215872 582562 215928
rect 582618 215872 611726 215928
rect 611782 215872 611787 215928
rect 582557 215870 611787 215872
rect 582557 215867 582623 215870
rect 611721 215867 611787 215870
rect 643001 215930 643067 215933
rect 669270 215930 669330 216142
rect 675201 216200 676292 216202
rect 675201 216144 675206 216200
rect 675262 216144 676292 216200
rect 675201 216142 676292 216144
rect 675201 216139 675267 216142
rect 675661 215930 675727 215933
rect 643001 215928 663810 215930
rect 643001 215872 643006 215928
rect 643062 215872 663810 215928
rect 643001 215870 663810 215872
rect 669270 215928 675727 215930
rect 669270 215872 675666 215928
rect 675722 215872 675727 215928
rect 669270 215870 675727 215872
rect 643001 215867 643067 215870
rect 509182 215596 509188 215660
rect 509252 215658 509258 215660
rect 594609 215658 594675 215661
rect 597921 215658 597987 215661
rect 509252 215656 594675 215658
rect 509252 215600 594614 215656
rect 594670 215600 594675 215656
rect 509252 215598 594675 215600
rect 509252 215596 509258 215598
rect 594609 215595 594675 215598
rect 594934 215656 597987 215658
rect 594934 215600 597926 215656
rect 597982 215600 597987 215656
rect 594934 215598 597987 215600
rect 506054 215324 506060 215388
rect 506124 215386 506130 215388
rect 594934 215386 594994 215598
rect 597921 215595 597987 215598
rect 506124 215326 594994 215386
rect 663750 215386 663810 215870
rect 675661 215867 675727 215870
rect 676170 215734 676292 215794
rect 667974 215596 667980 215660
rect 668044 215658 668050 215660
rect 669221 215658 669287 215661
rect 668044 215656 669287 215658
rect 668044 215600 669226 215656
rect 669282 215600 669287 215656
rect 668044 215598 669287 215600
rect 668044 215596 668050 215598
rect 669221 215595 669287 215598
rect 669446 215596 669452 215660
rect 669516 215658 669522 215660
rect 676170 215658 676230 215734
rect 669516 215598 676230 215658
rect 669516 215596 669522 215598
rect 675017 215386 675083 215389
rect 663750 215384 675083 215386
rect 663750 215328 675022 215384
rect 675078 215328 675083 215384
rect 663750 215326 675083 215328
rect 506124 215324 506130 215326
rect 675017 215323 675083 215326
rect 675702 215324 675708 215388
rect 675772 215386 675778 215388
rect 675772 215326 676292 215386
rect 675772 215324 675778 215326
rect 528686 215052 528692 215116
rect 528756 215114 528762 215116
rect 577037 215114 577103 215117
rect 528756 215112 577103 215114
rect 528756 215056 577042 215112
rect 577098 215056 577103 215112
rect 528756 215054 577103 215056
rect 528756 215052 528762 215054
rect 577037 215051 577103 215054
rect 586646 215052 586652 215116
rect 586716 215114 586722 215116
rect 596081 215114 596147 215117
rect 586716 215112 596147 215114
rect 586716 215056 596086 215112
rect 596142 215056 596147 215112
rect 586716 215054 596147 215056
rect 586716 215052 586722 215054
rect 596081 215051 596147 215054
rect 662045 215114 662111 215117
rect 676029 215114 676095 215117
rect 662045 215112 676095 215114
rect 662045 215056 662050 215112
rect 662106 215056 676034 215112
rect 676090 215056 676095 215112
rect 676254 215086 676260 215150
rect 676324 215086 676330 215150
rect 662045 215054 676095 215056
rect 662045 215051 662111 215054
rect 676029 215051 676095 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 676262 214948 676322 215086
rect 41492 214918 44883 214920
rect 44817 214915 44883 214918
rect 659285 214842 659351 214845
rect 675661 214842 675727 214845
rect 659285 214840 675727 214842
rect 659285 214784 659290 214840
rect 659346 214784 675666 214840
rect 675722 214784 675727 214840
rect 659285 214782 675727 214784
rect 659285 214779 659351 214782
rect 675661 214779 675727 214782
rect 650453 214570 650519 214573
rect 669221 214570 669287 214573
rect 669446 214570 669452 214572
rect 650453 214568 663810 214570
rect 35758 214301 35818 214540
rect 650453 214512 650458 214568
rect 650514 214512 663810 214568
rect 650453 214510 663810 214512
rect 669176 214568 669452 214570
rect 669176 214512 669226 214568
rect 669282 214512 669452 214568
rect 669176 214510 669452 214512
rect 650453 214507 650519 214510
rect 28533 214298 28599 214301
rect 28533 214296 28642 214298
rect 28533 214240 28538 214296
rect 28594 214240 28642 214296
rect 28533 214235 28642 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 28582 214132 28642 214235
rect 575982 214026 576042 214404
rect 663750 214298 663810 214510
rect 669221 214507 669287 214510
rect 669446 214508 669452 214510
rect 669516 214508 669522 214572
rect 669681 214570 669747 214573
rect 676029 214570 676095 214573
rect 669681 214568 674114 214570
rect 669681 214512 669686 214568
rect 669742 214512 674114 214568
rect 669681 214510 674114 214512
rect 669681 214507 669747 214510
rect 673729 214298 673795 214301
rect 663750 214296 673795 214298
rect 663750 214240 673734 214296
rect 673790 214240 673795 214296
rect 663750 214238 673795 214240
rect 673729 214235 673795 214238
rect 674054 214162 674114 214510
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 674054 214102 676292 214162
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 669446 213964 669452 214028
rect 669516 214026 669522 214028
rect 670601 214026 670667 214029
rect 669516 214024 670667 214026
rect 669516 213968 670606 214024
rect 670662 213968 670667 214024
rect 669516 213966 670667 213968
rect 669516 213964 669522 213966
rect 670601 213963 670667 213966
rect 672533 214028 672599 214029
rect 672533 214024 672580 214028
rect 672644 214026 672650 214028
rect 672533 213968 672538 214024
rect 672533 213964 672580 213968
rect 672644 213966 672690 214026
rect 672644 213964 672650 213966
rect 672533 213963 672599 213964
rect 43621 213754 43687 213757
rect 41492 213752 43687 213754
rect 41492 213696 43626 213752
rect 43682 213696 43687 213752
rect 41492 213694 43687 213696
rect 43621 213691 43687 213694
rect 664805 213754 664871 213757
rect 672073 213754 672139 213757
rect 664805 213752 671906 213754
rect 664805 213696 664810 213752
rect 664866 213696 671906 213752
rect 664805 213694 671906 213696
rect 664805 213691 664871 213694
rect 661493 213482 661559 213485
rect 671846 213482 671906 213694
rect 672073 213752 676292 213754
rect 672073 213696 672078 213752
rect 672134 213696 676292 213752
rect 672073 213694 676292 213696
rect 672073 213691 672139 213694
rect 676029 213482 676095 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 671846 213480 676095 213482
rect 671846 213424 676034 213480
rect 676090 213424 676095 213480
rect 671846 213422 676095 213424
rect 661493 213419 661559 213422
rect 47945 213346 48011 213349
rect 41492 213344 48011 213346
rect 41492 213288 47950 213344
rect 48006 213288 48011 213344
rect 41492 213286 48011 213288
rect 47945 213283 48011 213286
rect 647141 213210 647207 213213
rect 669270 213210 669330 213422
rect 676029 213419 676095 213422
rect 683297 213346 683363 213349
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 683297 213283 683363 213286
rect 676029 213210 676095 213213
rect 647141 213208 663810 213210
rect 647141 213152 647146 213208
rect 647202 213152 663810 213208
rect 647141 213150 663810 213152
rect 669270 213208 676095 213210
rect 669270 213152 676034 213208
rect 676090 213152 676095 213208
rect 669270 213150 676095 213152
rect 647141 213147 647207 213150
rect 43437 212938 43503 212941
rect 41492 212936 43503 212938
rect 41492 212880 43442 212936
rect 43498 212880 43503 212936
rect 41492 212878 43503 212880
rect 663750 212938 663810 213150
rect 676029 213147 676095 213150
rect 673913 212938 673979 212941
rect 663750 212936 673979 212938
rect 663750 212880 673918 212936
rect 673974 212880 673979 212936
rect 663750 212878 673979 212880
rect 43437 212875 43503 212878
rect 673913 212875 673979 212878
rect 683070 212533 683130 212908
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 35574 212261 35634 212500
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 683113 212467 683179 212470
rect 35574 212256 35683 212261
rect 35574 212200 35622 212256
rect 35678 212200 35683 212256
rect 35574 212198 35683 212200
rect 35617 212195 35683 212198
rect 42885 212122 42951 212125
rect 41492 212120 42951 212122
rect 41492 212064 42890 212120
rect 42946 212064 42951 212120
rect 41492 212062 42951 212064
rect 42885 212059 42951 212062
rect 575982 211714 576042 212228
rect 674046 212060 674052 212124
rect 674116 212122 674122 212124
rect 674116 212062 676292 212122
rect 674116 212060 674122 212062
rect 578233 211714 578299 211717
rect 575982 211712 578299 211714
rect 35758 211445 35818 211684
rect 575982 211656 578238 211712
rect 578294 211656 578299 211712
rect 575982 211654 578299 211656
rect 578233 211651 578299 211654
rect 35758 211440 35867 211445
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211382 35867 211384
rect 35801 211379 35867 211382
rect 670601 211442 670667 211445
rect 670601 211440 678990 211442
rect 670601 211384 670606 211440
rect 670662 211384 678990 211440
rect 670601 211382 678990 211384
rect 670601 211379 670667 211382
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 44173 211243 44239 211246
rect 669630 211108 669636 211172
rect 669700 211170 669706 211172
rect 670417 211170 670483 211173
rect 669700 211168 670483 211170
rect 669700 211112 670422 211168
rect 670478 211112 670483 211168
rect 669700 211110 670483 211112
rect 669700 211108 669706 211110
rect 670417 211107 670483 211110
rect 673729 211170 673795 211173
rect 676765 211170 676831 211173
rect 673729 211168 676831 211170
rect 673729 211112 673734 211168
rect 673790 211112 676770 211168
rect 676826 211112 676831 211168
rect 673729 211110 676831 211112
rect 673729 211107 673795 211110
rect 676765 211107 676831 211110
rect 676949 211172 677015 211173
rect 676949 211168 676996 211172
rect 677060 211170 677066 211172
rect 678930 211170 678990 211382
rect 683113 211170 683179 211173
rect 676949 211112 676954 211168
rect 676949 211108 676996 211112
rect 677060 211110 677106 211170
rect 678930 211168 683179 211170
rect 678930 211112 683118 211168
rect 683174 211112 683179 211168
rect 678930 211110 683179 211112
rect 677060 211108 677066 211110
rect 676949 211107 677015 211108
rect 683113 211107 683179 211110
rect 48129 210898 48195 210901
rect 41492 210896 48195 210898
rect 41492 210840 48134 210896
rect 48190 210840 48195 210896
rect 41492 210838 48195 210840
rect 48129 210835 48195 210838
rect 44173 210490 44239 210493
rect 41492 210488 44239 210490
rect 41492 210432 44178 210488
rect 44234 210432 44239 210488
rect 41492 210430 44239 210432
rect 44173 210427 44239 210430
rect 672809 210354 672875 210357
rect 683297 210354 683363 210357
rect 672809 210352 683363 210354
rect 672809 210296 672814 210352
rect 672870 210296 683302 210352
rect 683358 210296 683363 210352
rect 672809 210294 683363 210296
rect 672809 210291 672875 210294
rect 683297 210291 683363 210294
rect 35758 209813 35818 210052
rect 35758 209808 35867 209813
rect 35758 209752 35806 209808
rect 35862 209752 35867 209808
rect 35758 209750 35867 209752
rect 575982 209810 576042 210052
rect 579245 209810 579311 209813
rect 575982 209808 579311 209810
rect 575982 209752 579250 209808
rect 579306 209752 579311 209808
rect 575982 209750 579311 209752
rect 35801 209747 35867 209750
rect 579245 209747 579311 209750
rect 42793 209674 42859 209677
rect 41492 209672 42859 209674
rect 41492 209616 42798 209672
rect 42854 209616 42859 209672
rect 41492 209614 42859 209616
rect 42793 209611 42859 209614
rect 673913 209674 673979 209677
rect 677869 209674 677935 209677
rect 673913 209672 677935 209674
rect 673913 209616 673918 209672
rect 673974 209616 677874 209672
rect 677930 209616 677935 209672
rect 673913 209614 677935 209616
rect 673913 209611 673979 209614
rect 677869 209611 677935 209614
rect 41462 208996 41522 209236
rect 41454 208932 41460 208996
rect 41524 208932 41530 208996
rect 41689 208994 41755 208997
rect 49601 208994 49667 208997
rect 41689 208992 49667 208994
rect 41689 208936 41694 208992
rect 41750 208936 49606 208992
rect 49662 208936 49667 208992
rect 41689 208934 49667 208936
rect 41689 208931 41755 208934
rect 49601 208931 49667 208934
rect 41278 208586 41338 208828
rect 44541 208586 44607 208589
rect 41278 208584 44607 208586
rect 41278 208528 44546 208584
rect 44602 208528 44607 208584
rect 41278 208526 44607 208528
rect 44541 208523 44607 208526
rect 40542 208180 40602 208420
rect 40534 208116 40540 208180
rect 40604 208116 40610 208180
rect 43253 208042 43319 208045
rect 41492 208040 43319 208042
rect 41492 207984 43258 208040
rect 43314 207984 43319 208040
rect 41492 207982 43319 207984
rect 43253 207979 43319 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40910 207364 40970 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40902 207300 40908 207364
rect 40972 207300 40978 207364
rect 675477 207362 675543 207365
rect 666878 207360 675543 207362
rect 666878 207304 675482 207360
rect 675538 207304 675543 207360
rect 666878 207302 675543 207304
rect 666878 207294 666938 207302
rect 675477 207299 675543 207302
rect 666356 207234 666938 207294
rect 40726 206956 40786 207196
rect 40718 206892 40724 206956
rect 40788 206892 40794 206956
rect 43621 206818 43687 206821
rect 41492 206816 43687 206818
rect 41492 206760 43626 206816
rect 43682 206760 43687 206816
rect 41492 206758 43687 206760
rect 43621 206755 43687 206758
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 44357 206002 44423 206005
rect 41492 206000 44423 206002
rect 41492 205944 44362 206000
rect 44418 205944 44423 206000
rect 41492 205942 44423 205944
rect 44357 205939 44423 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 41321 205730 41387 205733
rect 42006 205730 42012 205732
rect 41321 205728 42012 205730
rect 41321 205672 41326 205728
rect 41382 205672 42012 205728
rect 41321 205670 42012 205672
rect 41321 205667 41387 205670
rect 42006 205668 42012 205670
rect 42076 205668 42082 205732
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 669262 205668 669268 205732
rect 669332 205730 669338 205732
rect 669630 205730 669636 205732
rect 669332 205670 669636 205730
rect 669332 205668 669338 205670
rect 669630 205668 669636 205670
rect 669700 205668 669706 205732
rect 675753 205594 675819 205597
rect 676438 205594 676444 205596
rect 675753 205592 676444 205594
rect 41462 205322 41522 205564
rect 675753 205536 675758 205592
rect 675814 205536 676444 205592
rect 675753 205534 676444 205536
rect 675753 205531 675819 205534
rect 676438 205532 676444 205534
rect 676508 205532 676514 205596
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 43805 205322 43871 205325
rect 41462 205320 43871 205322
rect 41462 205264 43810 205320
rect 43866 205264 43871 205320
rect 41462 205262 43871 205264
rect 43805 205259 43871 205262
rect 41462 204914 41522 205156
rect 43989 204914 44055 204917
rect 41462 204912 44055 204914
rect 41462 204856 43994 204912
rect 44050 204856 44055 204912
rect 41462 204854 44055 204856
rect 43989 204851 44055 204854
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 41462 204506 41522 204748
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 44817 204506 44883 204509
rect 41462 204504 44883 204506
rect 41462 204448 44822 204504
rect 44878 204448 44883 204504
rect 41462 204446 44883 204448
rect 44817 204443 44883 204446
rect 41094 204101 41154 204340
rect 675477 204236 675543 204237
rect 675477 204232 675524 204236
rect 675588 204234 675594 204236
rect 675477 204176 675482 204232
rect 675477 204172 675524 204176
rect 675588 204174 675634 204234
rect 675588 204172 675594 204174
rect 675477 204171 675543 204172
rect 41094 204096 41203 204101
rect 41094 204040 41142 204096
rect 41198 204040 41203 204096
rect 41094 204038 41203 204040
rect 41137 204035 41203 204038
rect 666356 203970 666938 204030
rect 666878 203962 666938 203970
rect 673729 203962 673795 203965
rect 666878 203960 673795 203962
rect 41278 203693 41338 203932
rect 666878 203904 673734 203960
rect 673790 203904 673795 203960
rect 666878 203902 673795 203904
rect 673729 203899 673795 203902
rect 41278 203688 41387 203693
rect 41278 203632 41326 203688
rect 41382 203632 41387 203688
rect 41278 203630 41387 203632
rect 41321 203627 41387 203630
rect 46381 203554 46447 203557
rect 41492 203552 46447 203554
rect 41492 203496 46386 203552
rect 46442 203496 46447 203552
rect 41492 203494 46447 203496
rect 46381 203491 46447 203494
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 669313 202602 669379 202605
rect 675477 202602 675543 202605
rect 669313 202600 675543 202602
rect 669313 202544 669318 202600
rect 669374 202544 675482 202600
rect 675538 202544 675543 202600
rect 669313 202542 675543 202544
rect 669313 202539 669379 202542
rect 675477 202539 675543 202542
rect 668025 202466 668091 202469
rect 666694 202464 668091 202466
rect 666694 202408 668030 202464
rect 668086 202408 668091 202464
rect 666694 202406 668091 202408
rect 666694 202398 666754 202406
rect 668025 202403 668091 202406
rect 666356 202338 666754 202398
rect 41321 202194 41387 202197
rect 41822 202194 41828 202196
rect 41321 202192 41828 202194
rect 41321 202136 41326 202192
rect 41382 202136 41828 202192
rect 41321 202134 41828 202136
rect 41321 202131 41387 202134
rect 41822 202132 41828 202134
rect 41892 202132 41898 202196
rect 674833 202058 674899 202061
rect 675477 202058 675543 202061
rect 674833 202056 675543 202058
rect 674833 202000 674838 202056
rect 674894 202000 675482 202056
rect 675538 202000 675543 202056
rect 674833 201998 675543 202000
rect 674833 201995 674899 201998
rect 675477 201995 675543 201998
rect 669221 201650 669287 201653
rect 675109 201650 675175 201653
rect 669221 201648 675175 201650
rect 669221 201592 669226 201648
rect 669282 201592 675114 201648
rect 675170 201592 675175 201648
rect 669221 201590 675175 201592
rect 669221 201587 669287 201590
rect 675109 201587 675175 201590
rect 41873 201514 41939 201517
rect 49417 201514 49483 201517
rect 41873 201512 49483 201514
rect 41873 201456 41878 201512
rect 41934 201456 49422 201512
rect 49478 201456 49483 201512
rect 41873 201454 49483 201456
rect 41873 201451 41939 201454
rect 49417 201451 49483 201454
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 575982 200834 576042 201348
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672073 200834 672139 200837
rect 674925 200834 674991 200837
rect 672073 200832 674991 200834
rect 672073 200776 672078 200832
rect 672134 200776 674930 200832
rect 674986 200776 674991 200832
rect 672073 200774 674991 200776
rect 672073 200771 672139 200774
rect 674925 200771 674991 200774
rect 41137 200698 41203 200701
rect 43437 200698 43503 200701
rect 41137 200696 43503 200698
rect 41137 200640 41142 200696
rect 41198 200640 43442 200696
rect 43498 200640 43503 200696
rect 41137 200638 43503 200640
rect 41137 200635 41203 200638
rect 43437 200635 43503 200638
rect 675753 200698 675819 200701
rect 676806 200698 676812 200700
rect 675753 200696 676812 200698
rect 675753 200640 675758 200696
rect 675814 200640 676812 200696
rect 675753 200638 676812 200640
rect 675753 200635 675819 200638
rect 676806 200636 676812 200638
rect 676876 200636 676882 200700
rect 669681 200562 669747 200565
rect 675293 200562 675359 200565
rect 669681 200560 675359 200562
rect 669681 200504 669686 200560
rect 669742 200504 675298 200560
rect 675354 200504 675359 200560
rect 669681 200502 675359 200504
rect 669681 200499 669747 200502
rect 675293 200499 675359 200502
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 667933 199202 667999 199205
rect 666694 199200 667999 199202
rect 575982 198930 576042 199172
rect 666694 199144 667938 199200
rect 667994 199144 667999 199200
rect 666694 199142 667999 199144
rect 666694 199134 666754 199142
rect 667933 199139 667999 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 668117 198794 668183 198797
rect 672257 198794 672323 198797
rect 668117 198792 672323 198794
rect 668117 198736 668122 198792
rect 668178 198736 672262 198792
rect 672318 198736 672323 198792
rect 668117 198734 672323 198736
rect 668117 198731 668183 198734
rect 672257 198731 672323 198734
rect 590377 198250 590443 198253
rect 674465 198250 674531 198253
rect 675477 198250 675543 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 674465 198248 675543 198250
rect 674465 198192 674470 198248
rect 674526 198192 675482 198248
rect 675538 198192 675543 198248
rect 674465 198190 675543 198192
rect 590377 198187 590443 198190
rect 674465 198187 674531 198190
rect 675477 198187 675543 198190
rect 666356 197442 666938 197502
rect 666878 197434 666938 197442
rect 673913 197434 673979 197437
rect 666878 197432 673979 197434
rect 666878 197376 673918 197432
rect 673974 197376 673979 197432
rect 666878 197374 673979 197376
rect 673913 197371 673979 197374
rect 40534 197100 40540 197164
rect 40604 197162 40610 197164
rect 41781 197162 41847 197165
rect 40604 197160 41847 197162
rect 40604 197104 41786 197160
rect 41842 197104 41847 197160
rect 40604 197102 41847 197104
rect 40604 197100 40610 197102
rect 41781 197099 41847 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49601 196482 49667 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49601 196480 52164 196482
rect 49601 196424 49606 196480
rect 49662 196424 52164 196480
rect 49601 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49601 196419 49667 196422
rect 578509 196419 578575 196422
rect 669262 196012 669268 196076
rect 669332 196074 669338 196076
rect 669630 196074 669636 196076
rect 669332 196014 669636 196074
rect 669332 196012 669338 196014
rect 669630 196012 669636 196014
rect 669700 196012 669706 196076
rect 41781 195804 41847 195805
rect 41781 195800 41828 195804
rect 41892 195802 41898 195804
rect 41781 195744 41786 195800
rect 41781 195740 41828 195744
rect 41892 195742 41938 195802
rect 41892 195740 41898 195742
rect 41781 195739 41847 195740
rect 40902 195332 40908 195396
rect 40972 195394 40978 195396
rect 42241 195394 42307 195397
rect 40972 195392 42307 195394
rect 40972 195336 42246 195392
rect 42302 195336 42307 195392
rect 40972 195334 42307 195336
rect 40972 195332 40978 195334
rect 42241 195331 42307 195334
rect 675661 195258 675727 195261
rect 675886 195258 675892 195260
rect 675661 195256 675892 195258
rect 675661 195200 675666 195256
rect 675722 195200 675892 195256
rect 675661 195198 675892 195200
rect 675661 195195 675727 195198
rect 675886 195196 675892 195198
rect 675956 195196 675962 195260
rect 41965 195124 42031 195125
rect 41965 195120 42012 195124
rect 42076 195122 42082 195124
rect 41965 195064 41970 195120
rect 41965 195060 42012 195064
rect 42076 195062 42122 195122
rect 42076 195060 42082 195062
rect 41965 195059 42031 195060
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 48129 194442 48195 194445
rect 48129 194440 52164 194442
rect 48129 194384 48134 194440
rect 48190 194384 52164 194440
rect 48129 194382 52164 194384
rect 48129 194379 48195 194382
rect 667933 194306 667999 194309
rect 666694 194304 667999 194306
rect 666694 194248 667938 194304
rect 667994 194248 667999 194304
rect 666694 194246 667999 194248
rect 666694 194238 666754 194246
rect 667933 194243 667999 194246
rect 666356 194178 666754 194238
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42006 193156 42012 193220
rect 42076 193218 42082 193220
rect 42241 193218 42307 193221
rect 42076 193216 42307 193218
rect 42076 193160 42246 193216
rect 42302 193160 42307 193216
rect 42076 193158 42307 193160
rect 42076 193156 42082 193158
rect 42241 193155 42307 193158
rect 42425 193218 42491 193221
rect 43621 193218 43687 193221
rect 42425 193216 43687 193218
rect 42425 193160 42430 193216
rect 42486 193160 43626 193216
rect 43682 193160 43687 193216
rect 42425 193158 43687 193160
rect 42425 193155 42491 193158
rect 43621 193155 43687 193158
rect 668945 192674 669011 192677
rect 666694 192672 669011 192674
rect 49417 192402 49483 192405
rect 49417 192400 52164 192402
rect 49417 192344 49422 192400
rect 49478 192344 52164 192400
rect 49417 192342 52164 192344
rect 49417 192339 49483 192342
rect 575982 192266 576042 192644
rect 666694 192616 668950 192672
rect 669006 192616 669011 192672
rect 666694 192614 669011 192616
rect 666694 192606 666754 192614
rect 668945 192611 669011 192614
rect 666356 192546 666754 192606
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 43989 191722 44055 191725
rect 42333 191720 44055 191722
rect 42333 191664 42338 191720
rect 42394 191664 43994 191720
rect 44050 191664 44055 191720
rect 42333 191662 44055 191664
rect 42333 191659 42399 191662
rect 43989 191659 44055 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43805 190498 43871 190501
rect 42425 190496 43871 190498
rect 42425 190440 42430 190496
rect 42486 190440 43810 190496
rect 43866 190440 43871 190496
rect 42425 190438 43871 190440
rect 42425 190435 42491 190438
rect 43805 190435 43871 190438
rect 47945 190498 48011 190501
rect 47945 190496 52164 190498
rect 47945 190440 47950 190496
rect 48006 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47945 190438 52164 190440
rect 47945 190435 48011 190438
rect 670601 190362 670667 190365
rect 675293 190362 675359 190365
rect 670601 190360 675359 190362
rect 670601 190304 670606 190360
rect 670662 190304 675298 190360
rect 675354 190304 675359 190360
rect 670601 190302 675359 190304
rect 670601 190299 670667 190302
rect 675293 190299 675359 190302
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 44541 189954 44607 189957
rect 42425 189952 44607 189954
rect 42425 189896 42430 189952
rect 42486 189896 44546 189952
rect 44602 189896 44607 189952
rect 42425 189894 44607 189896
rect 42425 189891 42491 189894
rect 44541 189891 44607 189894
rect 666502 189756 666508 189820
rect 666572 189818 666578 189820
rect 675109 189818 675175 189821
rect 666572 189816 675175 189818
rect 666572 189760 675114 189816
rect 675170 189760 675175 189816
rect 666572 189758 675175 189760
rect 666572 189756 666578 189758
rect 675109 189755 675175 189758
rect 667933 189410 667999 189413
rect 666694 189408 667999 189410
rect 666694 189352 667938 189408
rect 667994 189352 667999 189408
rect 666694 189350 667999 189352
rect 666694 189342 666754 189350
rect 667933 189347 667999 189350
rect 666356 189282 666754 189342
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 666356 187650 666754 187710
rect 42425 187642 42491 187645
rect 44357 187642 44423 187645
rect 42425 187640 44423 187642
rect 42425 187584 42430 187640
rect 42486 187584 44362 187640
rect 44418 187584 44423 187640
rect 42425 187582 44423 187584
rect 666694 187642 666754 187650
rect 668117 187642 668183 187645
rect 666694 187640 668183 187642
rect 666694 187584 668122 187640
rect 668178 187584 668183 187640
rect 666694 187582 668183 187584
rect 42425 187579 42491 187582
rect 44357 187579 44423 187582
rect 668117 187579 668183 187582
rect 41454 187172 41460 187236
rect 41524 187234 41530 187236
rect 41781 187234 41847 187237
rect 41524 187232 41847 187234
rect 41524 187176 41786 187232
rect 41842 187176 41847 187232
rect 41524 187174 41847 187176
rect 41524 187172 41530 187174
rect 41781 187171 41847 187174
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 42057 186420 42123 186421
rect 42006 186418 42012 186420
rect 41966 186358 42012 186418
rect 42076 186416 42123 186420
rect 42118 186360 42123 186416
rect 42006 186356 42012 186358
rect 42076 186356 42123 186360
rect 42057 186355 42123 186356
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 42149 185876 42215 185877
rect 42149 185874 42196 185876
rect 42104 185872 42196 185874
rect 42104 185816 42154 185872
rect 42104 185814 42196 185816
rect 42149 185812 42196 185814
rect 42260 185812 42266 185876
rect 42149 185811 42215 185812
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 42425 184922 42491 184925
rect 44173 184922 44239 184925
rect 42425 184920 44239 184922
rect 42425 184864 42430 184920
rect 42486 184864 44178 184920
rect 44234 184864 44239 184920
rect 42425 184862 44239 184864
rect 42425 184859 42491 184862
rect 44173 184859 44239 184862
rect 668117 184922 668183 184925
rect 672441 184922 672507 184925
rect 668117 184920 672507 184922
rect 668117 184864 668122 184920
rect 668178 184864 672446 184920
rect 672502 184864 672507 184920
rect 668117 184862 672507 184864
rect 668117 184859 668183 184862
rect 672441 184859 672507 184862
rect 669221 184514 669287 184517
rect 666694 184512 669287 184514
rect 666694 184456 669226 184512
rect 669282 184456 669287 184512
rect 666694 184454 669287 184456
rect 666694 184446 666754 184454
rect 669221 184451 669287 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 672073 183562 672139 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672073 183560 672948 183562
rect 672073 183504 672078 183560
rect 672134 183504 672948 183560
rect 672073 183502 672948 183504
rect 589457 183499 589523 183502
rect 672073 183499 672139 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 43253 183154 43319 183157
rect 42425 183152 43319 183154
rect 42425 183096 42430 183152
rect 42486 183096 43258 183152
rect 43314 183096 43319 183152
rect 42425 183094 43319 183096
rect 42425 183091 42491 183094
rect 43253 183091 43319 183094
rect 668301 182882 668367 182885
rect 666694 182880 668367 182882
rect 666694 182824 668306 182880
rect 668362 182824 668367 182880
rect 666694 182822 668367 182824
rect 666694 182814 666754 182822
rect 668301 182819 668367 182822
rect 666356 182754 666754 182814
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667381 181386 667447 181389
rect 675845 181386 675911 181389
rect 667381 181384 675911 181386
rect 667381 181328 667386 181384
rect 667442 181328 675850 181384
rect 675906 181328 675911 181384
rect 667381 181326 675911 181328
rect 667381 181323 667447 181326
rect 675845 181323 675911 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 666356 179490 666938 179550
rect 666878 179482 666938 179490
rect 674281 179482 674347 179485
rect 666878 179480 674347 179482
rect 666878 179424 674286 179480
rect 674342 179424 674347 179480
rect 666878 179422 674347 179424
rect 674281 179419 674347 179422
rect 667749 178802 667815 178805
rect 676029 178802 676095 178805
rect 667749 178800 676095 178802
rect 667749 178744 667754 178800
rect 667810 178744 676034 178800
rect 676090 178744 676095 178800
rect 667749 178742 676095 178744
rect 667749 178739 667815 178742
rect 676029 178739 676095 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 666645 178530 666711 178533
rect 666645 178528 676292 178530
rect 666645 178472 666650 178528
rect 666706 178472 676292 178528
rect 666645 178470 676292 178472
rect 666645 178467 666711 178470
rect 675845 178122 675911 178125
rect 675845 178120 676292 178122
rect 675845 178064 675850 178120
rect 675906 178064 676292 178120
rect 675845 178062 676292 178064
rect 675845 178059 675911 178062
rect 672993 177986 673059 177989
rect 666694 177984 673059 177986
rect 666694 177928 672998 177984
rect 673054 177928 673059 177984
rect 666694 177926 673059 177928
rect 666694 177918 666754 177926
rect 672993 177923 673059 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 676029 177714 676095 177717
rect 676029 177712 676292 177714
rect 676029 177656 676034 177712
rect 676090 177656 676292 177712
rect 676029 177654 676292 177656
rect 676029 177651 676095 177654
rect 673361 177306 673427 177309
rect 673361 177304 676292 177306
rect 673361 177248 673366 177304
rect 673422 177248 676292 177304
rect 673361 177246 676292 177248
rect 673361 177243 673427 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673361 176898 673427 176901
rect 673361 176896 676292 176898
rect 673361 176840 673366 176896
rect 673422 176840 676292 176896
rect 673361 176838 676292 176840
rect 673361 176835 673427 176838
rect 671889 176490 671955 176493
rect 671889 176488 676292 176490
rect 671889 176432 671894 176488
rect 671950 176432 676292 176488
rect 671889 176430 676292 176432
rect 671889 176427 671955 176430
rect 673177 176082 673243 176085
rect 673177 176080 676292 176082
rect 673177 176024 673182 176080
rect 673238 176024 676292 176080
rect 673177 176022 676292 176024
rect 673177 176019 673243 176022
rect 674649 175674 674715 175677
rect 674649 175672 676292 175674
rect 674649 175616 674654 175672
rect 674710 175616 676292 175672
rect 674649 175614 676292 175616
rect 674649 175611 674715 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674649 175266 674715 175269
rect 674649 175264 676292 175266
rect 575982 175130 576042 175236
rect 674649 175208 674654 175264
rect 674710 175208 676292 175264
rect 674649 175206 676292 175208
rect 674649 175203 674715 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 673545 174858 673611 174861
rect 673545 174856 676292 174858
rect 673545 174800 673550 174856
rect 673606 174800 676292 174856
rect 673545 174798 676292 174800
rect 673545 174795 673611 174798
rect 667933 174722 667999 174725
rect 666694 174720 667999 174722
rect 666694 174664 667938 174720
rect 667994 174664 667999 174720
rect 666694 174662 667999 174664
rect 666694 174654 666754 174662
rect 667933 174659 667999 174662
rect 666356 174594 666754 174654
rect 674373 174450 674439 174453
rect 674373 174448 676292 174450
rect 674373 174392 674378 174448
rect 674434 174392 676292 174448
rect 674373 174390 676292 174392
rect 674373 174387 674439 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 671705 173090 671771 173093
rect 666694 173088 671771 173090
rect 666694 173032 671710 173088
rect 671766 173032 671771 173088
rect 666694 173030 671771 173032
rect 666694 173022 666754 173030
rect 671705 173027 671771 173030
rect 666356 172962 666754 173022
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 670601 172002 670667 172005
rect 670601 172000 676292 172002
rect 670601 171944 670606 172000
rect 670662 171944 676292 172000
rect 670601 171942 676292 171944
rect 670601 171939 670667 171942
rect 680997 171594 681063 171597
rect 680997 171592 681076 171594
rect 680997 171536 681002 171592
rect 681058 171536 681076 171592
rect 680997 171534 681076 171536
rect 680997 171531 681063 171534
rect 675017 171186 675083 171189
rect 675017 171184 676292 171186
rect 675017 171128 675022 171184
rect 675078 171128 676292 171184
rect 675017 171126 676292 171128
rect 675017 171123 675083 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 675702 170308 675708 170372
rect 675772 170370 675778 170372
rect 675772 170310 676292 170370
rect 675772 170308 675778 170310
rect 671889 169962 671955 169965
rect 671889 169960 676292 169962
rect 671889 169904 671894 169960
rect 671950 169904 676292 169960
rect 671889 169902 676292 169904
rect 671889 169899 671955 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 667933 169690 667999 169693
rect 666694 169688 667999 169690
rect 666694 169632 667938 169688
rect 667994 169632 667999 169688
rect 666694 169630 667999 169632
rect 667933 169627 667999 169630
rect 669773 169554 669839 169557
rect 669773 169552 676292 169554
rect 669773 169496 669778 169552
rect 669834 169496 676292 169552
rect 669773 169494 676292 169496
rect 669773 169491 669839 169494
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672993 169146 673059 169149
rect 672993 169144 676292 169146
rect 672993 169088 672998 169144
rect 673054 169088 676292 169144
rect 672993 169086 676292 169088
rect 672993 169083 673059 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673913 168738 673979 168741
rect 673913 168736 676292 168738
rect 673913 168680 673918 168736
rect 673974 168680 676292 168736
rect 673913 168678 676292 168680
rect 673913 168675 673979 168678
rect 670141 168330 670207 168333
rect 670141 168328 676292 168330
rect 670141 168272 670146 168328
rect 670202 168272 676292 168328
rect 670141 168270 676292 168272
rect 670141 168267 670207 168270
rect 668117 168194 668183 168197
rect 666694 168192 668183 168194
rect 666694 168136 668122 168192
rect 668178 168136 668183 168192
rect 666694 168134 668183 168136
rect 666694 168126 666754 168134
rect 668117 168131 668183 168134
rect 666356 168066 666754 168126
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675886 167452 675892 167516
rect 675956 167514 675962 167516
rect 675956 167454 676292 167514
rect 675956 167452 675962 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 669129 167106 669195 167109
rect 669630 167106 669636 167108
rect 669129 167104 669636 167106
rect 669129 167048 669134 167104
rect 669190 167048 669636 167104
rect 669129 167046 669636 167048
rect 669129 167043 669195 167046
rect 669630 167044 669636 167046
rect 669700 167044 669706 167108
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 671705 166970 671771 166973
rect 676170 166970 676230 167046
rect 671705 166968 676230 166970
rect 671705 166912 671710 166968
rect 671766 166912 676230 166968
rect 671705 166910 676230 166912
rect 671705 166907 671771 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 670325 165610 670391 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 670325 165608 676095 165610
rect 670325 165552 670330 165608
rect 670386 165552 676034 165608
rect 676090 165552 676095 165608
rect 670325 165550 676095 165552
rect 589457 165547 589523 165550
rect 670325 165547 670391 165550
rect 676029 165547 676095 165550
rect 669497 164930 669563 164933
rect 666694 164928 669563 164930
rect 666694 164872 669502 164928
rect 669558 164872 669563 164928
rect 666694 164870 669563 164872
rect 666694 164862 666754 164870
rect 669497 164867 669563 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668945 163298 669011 163301
rect 666694 163296 669011 163298
rect 666694 163240 668950 163296
rect 669006 163240 669011 163296
rect 666694 163238 669011 163240
rect 666694 163230 666754 163238
rect 668945 163235 669011 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675201 161394 675267 161397
rect 675845 161394 675911 161397
rect 675201 161392 675911 161394
rect 675201 161336 675206 161392
rect 675262 161336 675850 161392
rect 675906 161336 675911 161392
rect 675201 161334 675911 161336
rect 675201 161331 675267 161334
rect 675845 161331 675911 161334
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 667013 160034 667079 160037
rect 666694 160032 667079 160034
rect 575982 159898 576042 160004
rect 666694 159976 667018 160032
rect 667074 159976 667079 160032
rect 666694 159974 667079 159976
rect 666694 159966 666754 159974
rect 667013 159971 667079 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 675753 159354 675819 159357
rect 676438 159354 676444 159356
rect 675753 159352 676444 159354
rect 675753 159296 675758 159352
rect 675814 159296 676444 159352
rect 675753 159294 676444 159296
rect 675753 159291 675819 159294
rect 676438 159292 676444 159294
rect 676508 159292 676514 159356
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 671521 158402 671587 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 671587 158402
rect 666694 158344 671526 158400
rect 671582 158344 671587 158400
rect 666694 158342 671587 158344
rect 666694 158334 666754 158342
rect 671521 158339 671587 158342
rect 666356 158274 666754 158334
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 666356 155010 666938 155070
rect 666878 154594 666938 155010
rect 669773 154866 669839 154869
rect 675109 154866 675175 154869
rect 669773 154864 675175 154866
rect 669773 154808 669778 154864
rect 669834 154808 675114 154864
rect 675170 154808 675175 154864
rect 669773 154806 675175 154808
rect 669773 154803 669839 154806
rect 675109 154803 675175 154806
rect 674097 154594 674163 154597
rect 666878 154592 674163 154594
rect 666878 154536 674102 154592
rect 674158 154536 674163 154592
rect 666878 154534 674163 154536
rect 674097 154531 674163 154534
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 668761 153506 668827 153509
rect 666694 153504 668827 153506
rect 666694 153448 668766 153504
rect 668822 153448 668827 153504
rect 666694 153446 668827 153448
rect 666694 153438 666754 153446
rect 668761 153443 668827 153446
rect 666356 153378 666754 153438
rect 668761 153098 668827 153101
rect 672625 153098 672691 153101
rect 668761 153096 672691 153098
rect 668761 153040 668766 153096
rect 668822 153040 672630 153096
rect 672686 153040 672691 153096
rect 668761 153038 672691 153040
rect 668761 153035 668827 153038
rect 672625 153035 672691 153038
rect 589457 152554 589523 152557
rect 672993 152554 673059 152557
rect 675477 152554 675543 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 672993 152552 675543 152554
rect 672993 152496 672998 152552
rect 673054 152496 675482 152552
rect 675538 152496 675543 152552
rect 672993 152494 675543 152496
rect 589457 152491 589523 152494
rect 672993 152491 673059 152494
rect 675477 152491 675543 152494
rect 671889 151874 671955 151877
rect 675477 151874 675543 151877
rect 671889 151872 675543 151874
rect 671889 151816 671894 151872
rect 671950 151816 675482 151872
rect 675538 151816 675543 151872
rect 671889 151814 675543 151816
rect 671889 151811 671955 151814
rect 675477 151811 675543 151814
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675293 151602 675359 151605
rect 676254 151602 676260 151604
rect 675293 151600 676260 151602
rect 675293 151544 675298 151600
rect 675354 151544 676260 151600
rect 675293 151542 676260 151544
rect 675293 151539 675359 151542
rect 676254 151540 676260 151542
rect 676324 151540 676330 151604
rect 673913 151058 673979 151061
rect 675109 151058 675175 151061
rect 673913 151056 675175 151058
rect 673913 151000 673918 151056
rect 673974 151000 675114 151056
rect 675170 151000 675175 151056
rect 673913 150998 675175 151000
rect 673913 150995 673979 150998
rect 675109 150995 675175 150998
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 675661 150380 675727 150381
rect 675661 150376 675708 150380
rect 675772 150378 675778 150380
rect 675661 150320 675666 150376
rect 675661 150316 675708 150320
rect 675772 150318 675818 150378
rect 675772 150316 675778 150318
rect 675661 150315 675727 150316
rect 668301 150242 668367 150245
rect 666694 150240 668367 150242
rect 666694 150184 668306 150240
rect 668362 150184 668367 150240
rect 666694 150182 668367 150184
rect 666694 150174 666754 150182
rect 668301 150179 668367 150182
rect 666356 150114 666754 150174
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 670601 149018 670667 149021
rect 675293 149018 675359 149021
rect 670601 149016 675359 149018
rect 670601 148960 670606 149016
rect 670662 148960 675298 149016
rect 675354 148960 675359 149016
rect 670601 148958 675359 148960
rect 670601 148955 670667 148958
rect 675293 148955 675359 148958
rect 668485 148610 668551 148613
rect 666694 148608 668551 148610
rect 666694 148552 668490 148608
rect 668546 148552 668551 148608
rect 666694 148550 668551 148552
rect 666694 148542 666754 148550
rect 668485 148547 668551 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 675661 147658 675727 147661
rect 675886 147658 675892 147660
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 675661 147656 675892 147658
rect 675661 147600 675666 147656
rect 675722 147600 675892 147656
rect 675661 147598 675892 147600
rect 588537 147595 588603 147598
rect 675661 147595 675727 147598
rect 675886 147596 675892 147598
rect 675956 147596 675962 147660
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 671286 145346 671292 145348
rect 666694 145286 671292 145346
rect 666694 145278 666754 145286
rect 671286 145284 671292 145286
rect 671356 145284 671362 145348
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579521 144666 579587 144669
rect 575982 144664 579587 144666
rect 575982 144608 579526 144664
rect 579582 144608 579587 144664
rect 575982 144606 579587 144608
rect 579521 144603 579587 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669129 143714 669195 143717
rect 666694 143712 669195 143714
rect 666694 143656 669134 143712
rect 669190 143656 669195 143712
rect 666694 143654 669195 143656
rect 666694 143646 666754 143654
rect 669129 143651 669195 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 669037 142218 669103 142221
rect 673678 142218 673684 142220
rect 669037 142216 673684 142218
rect 669037 142160 669042 142216
rect 669098 142160 673684 142216
rect 669037 142158 673684 142160
rect 669037 142155 669103 142158
rect 673678 142156 673684 142158
rect 673748 142156 673754 142220
rect 667197 141402 667263 141405
rect 683297 141402 683363 141405
rect 667197 141400 683363 141402
rect 667197 141344 667202 141400
rect 667258 141344 683302 141400
rect 683358 141344 683363 141400
rect 667197 141342 683363 141344
rect 667197 141339 667263 141342
rect 683297 141339 683363 141342
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 672073 140450 672139 140453
rect 666694 140448 672139 140450
rect 666694 140392 672078 140448
rect 672134 140392 672139 140448
rect 666694 140390 672139 140392
rect 666694 140382 666754 140390
rect 672073 140387 672139 140390
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 669037 138818 669103 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 669103 138818
rect 666694 138760 669042 138816
rect 669098 138760 669103 138816
rect 666694 138758 669103 138760
rect 666694 138750 666754 138758
rect 669037 138755 669103 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 667933 137458 667999 137461
rect 669446 137458 669452 137460
rect 667933 137456 669452 137458
rect 667933 137400 667938 137456
rect 667994 137400 669452 137456
rect 667933 137398 669452 137400
rect 667933 137395 667999 137398
rect 669446 137396 669452 137398
rect 669516 137396 669522 137460
rect 579245 136642 579311 136645
rect 575798 136640 579311 136642
rect 575798 136584 579250 136640
rect 579306 136584 579311 136640
rect 575798 136582 579311 136584
rect 575798 136068 575858 136582
rect 579245 136579 579311 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 667565 135962 667631 135965
rect 683113 135962 683179 135965
rect 667565 135960 683179 135962
rect 667565 135904 667570 135960
rect 667626 135904 683118 135960
rect 683174 135904 683179 135960
rect 667565 135902 683179 135904
rect 667565 135899 667631 135902
rect 683113 135899 683179 135902
rect 667933 135554 667999 135557
rect 666694 135552 667999 135554
rect 666694 135496 667938 135552
rect 667994 135496 667999 135552
rect 666694 135494 667999 135496
rect 666694 135486 666754 135494
rect 667933 135491 667999 135494
rect 666356 135426 666754 135486
rect 590285 134602 590351 134605
rect 590285 134600 592572 134602
rect 590285 134544 590290 134600
rect 590346 134544 592572 134600
rect 590285 134542 592572 134544
rect 590285 134539 590351 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 673126 133922 673132 133924
rect 667982 133862 673132 133922
rect 666356 133794 666938 133854
rect 666878 133650 666938 133794
rect 667982 133650 668042 133862
rect 673126 133860 673132 133862
rect 673196 133860 673202 133924
rect 666878 133590 668042 133650
rect 666829 133106 666895 133109
rect 676262 133106 676322 133348
rect 683297 133106 683363 133109
rect 666829 133104 676322 133106
rect 666829 133048 666834 133104
rect 666890 133048 676322 133104
rect 666829 133046 676322 133048
rect 683254 133104 683363 133106
rect 683254 133048 683302 133104
rect 683358 133048 683363 133104
rect 666829 133043 666895 133046
rect 683254 133043 683363 133048
rect 588721 132970 588787 132973
rect 588721 132968 592572 132970
rect 588721 132912 588726 132968
rect 588782 132912 592572 132968
rect 683254 132940 683314 133043
rect 588721 132910 592572 132912
rect 588721 132907 588787 132910
rect 683113 132698 683179 132701
rect 683070 132696 683179 132698
rect 683070 132640 683118 132696
rect 683174 132640 683179 132696
rect 683070 132635 683179 132640
rect 683070 132532 683130 132635
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673361 132154 673427 132157
rect 673361 132152 676292 132154
rect 673361 132096 673366 132152
rect 673422 132096 676292 132152
rect 673361 132094 676292 132096
rect 673361 132091 673427 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 673177 131338 673243 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 673177 131336 676292 131338
rect 673177 131280 673182 131336
rect 673238 131280 676292 131336
rect 673177 131278 676292 131280
rect 589457 131275 589523 131278
rect 673177 131275 673243 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130658 667980 130660
rect 666694 130598 667980 130658
rect 666694 130590 666754 130598
rect 667974 130596 667980 130598
rect 668044 130596 668050 130660
rect 666356 130530 666754 130590
rect 674649 130522 674715 130525
rect 674649 130520 676292 130522
rect 674649 130464 674654 130520
rect 674710 130464 676292 130520
rect 674649 130462 676292 130464
rect 674649 130459 674715 130462
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 579061 129706 579127 129709
rect 575798 129704 579127 129706
rect 575798 129648 579066 129704
rect 579122 129648 579127 129704
rect 575798 129646 579127 129648
rect 575798 129540 575858 129646
rect 579061 129643 579127 129646
rect 589641 129706 589707 129709
rect 674373 129706 674439 129709
rect 589641 129704 592572 129706
rect 589641 129648 589646 129704
rect 589702 129648 592572 129704
rect 589641 129646 592572 129648
rect 674373 129704 676292 129706
rect 674373 129648 674378 129704
rect 674434 129648 676292 129704
rect 674373 129646 676292 129648
rect 589641 129643 589707 129646
rect 674373 129643 674439 129646
rect 674097 129298 674163 129301
rect 674097 129296 676292 129298
rect 674097 129240 674102 129296
rect 674158 129240 676292 129296
rect 674097 129238 676292 129240
rect 674097 129235 674163 129238
rect 666356 128898 666938 128958
rect 666878 128482 666938 128898
rect 676630 128620 676690 128860
rect 676622 128556 676628 128620
rect 676692 128556 676698 128620
rect 673494 128482 673500 128484
rect 666878 128422 673500 128482
rect 673494 128420 673500 128422
rect 673564 128420 673570 128484
rect 674281 128346 674347 128349
rect 676029 128346 676095 128349
rect 674281 128344 676095 128346
rect 674281 128288 674286 128344
rect 674342 128288 676034 128344
rect 676090 128288 676095 128344
rect 674281 128286 676095 128288
rect 674281 128283 674347 128286
rect 676029 128283 676095 128286
rect 679574 128213 679634 128452
rect 668945 128210 669011 128213
rect 674046 128210 674052 128212
rect 668945 128208 674052 128210
rect 668945 128152 668950 128208
rect 669006 128152 674052 128208
rect 668945 128150 674052 128152
rect 668945 128147 669011 128150
rect 674046 128148 674052 128150
rect 674116 128148 674122 128212
rect 679574 128208 679683 128213
rect 679574 128152 679622 128208
rect 679678 128152 679683 128208
rect 679574 128150 679683 128152
rect 679617 128147 679683 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 678286 127805 678346 128044
rect 579153 127802 579219 127805
rect 575798 127800 579219 127802
rect 575798 127744 579158 127800
rect 579214 127744 579219 127800
rect 575798 127742 579219 127744
rect 575798 127364 575858 127742
rect 579153 127739 579219 127742
rect 678237 127800 678346 127805
rect 678237 127744 678242 127800
rect 678298 127744 678346 127800
rect 678237 127742 678346 127744
rect 678237 127739 678303 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 676262 126989 676322 127228
rect 676213 126984 676322 126989
rect 676213 126928 676218 126984
rect 676274 126928 676322 126984
rect 676213 126926 676322 126928
rect 676213 126923 676279 126926
rect 676446 126580 676506 126820
rect 676438 126516 676444 126580
rect 676508 126516 676514 126580
rect 590101 126442 590167 126445
rect 675017 126442 675083 126445
rect 590101 126440 592572 126442
rect 590101 126384 590106 126440
rect 590162 126384 592572 126440
rect 590101 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 590101 126379 590167 126382
rect 675017 126379 675083 126382
rect 674649 126034 674715 126037
rect 674649 126032 676292 126034
rect 674649 125976 674654 126032
rect 674710 125976 676292 126032
rect 674649 125974 676292 125976
rect 674649 125971 674715 125974
rect 668761 125762 668827 125765
rect 666694 125760 668827 125762
rect 666694 125704 668766 125760
rect 668822 125704 668827 125760
rect 666694 125702 668827 125704
rect 666694 125694 666754 125702
rect 668761 125699 668827 125702
rect 666356 125634 666754 125694
rect 672349 125626 672415 125629
rect 672349 125624 676292 125626
rect 672349 125568 672354 125624
rect 672410 125568 676292 125624
rect 672349 125566 676292 125568
rect 672349 125563 672415 125566
rect 579521 125354 579587 125357
rect 575798 125352 579587 125354
rect 575798 125296 579526 125352
rect 579582 125296 579587 125352
rect 575798 125294 579587 125296
rect 575798 125188 575858 125294
rect 579521 125291 579587 125294
rect 673913 125218 673979 125221
rect 673913 125216 676292 125218
rect 673913 125160 673918 125216
rect 673974 125160 676292 125216
rect 673913 125158 676292 125160
rect 673913 125155 673979 125158
rect 675886 124884 675892 124948
rect 675956 124946 675962 124948
rect 676213 124946 676279 124949
rect 675956 124944 676279 124946
rect 675956 124888 676218 124944
rect 676274 124888 676279 124944
rect 675956 124886 676279 124888
rect 675956 124884 675962 124886
rect 676213 124883 676279 124886
rect 589917 124810 589983 124813
rect 589917 124808 592572 124810
rect 589917 124752 589922 124808
rect 589978 124752 592572 124808
rect 589917 124750 592572 124752
rect 589917 124747 589983 124750
rect 676814 124540 676874 124780
rect 676806 124476 676812 124540
rect 676876 124476 676882 124540
rect 673177 124402 673243 124405
rect 673177 124400 676292 124402
rect 673177 124344 673182 124400
rect 673238 124344 676292 124400
rect 673177 124342 676292 124344
rect 673177 124339 673243 124342
rect 672809 124130 672875 124133
rect 666694 124128 672875 124130
rect 666694 124072 672814 124128
rect 672870 124072 672875 124128
rect 666694 124070 672875 124072
rect 666694 124062 666754 124070
rect 672809 124067 672875 124070
rect 666356 124002 666754 124062
rect 673361 123722 673427 123725
rect 676262 123722 676322 123964
rect 673361 123720 676322 123722
rect 673361 123664 673366 123720
rect 673422 123664 676322 123720
rect 673361 123662 676322 123664
rect 673361 123659 673427 123662
rect 578325 123586 578391 123589
rect 575798 123584 578391 123586
rect 575798 123528 578330 123584
rect 578386 123528 578391 123584
rect 575798 123526 578391 123528
rect 575798 123012 575858 123526
rect 578325 123523 578391 123526
rect 676630 123317 676690 123556
rect 676630 123312 676739 123317
rect 676630 123256 676678 123312
rect 676734 123256 676739 123312
rect 676630 123254 676739 123256
rect 676673 123251 676739 123254
rect 589457 123178 589523 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 589457 123115 589523 123118
rect 676262 122906 676322 123148
rect 673134 122846 676322 122906
rect 672942 122708 672948 122772
rect 673012 122770 673018 122772
rect 673134 122770 673194 122846
rect 673012 122710 673194 122770
rect 673012 122708 673018 122710
rect 672717 122498 672783 122501
rect 676262 122498 676322 122740
rect 672717 122496 676322 122498
rect 672717 122440 672722 122496
rect 672778 122440 676322 122496
rect 672717 122438 676322 122440
rect 672717 122435 672783 122438
rect 669221 122226 669287 122229
rect 672942 122226 672948 122228
rect 669221 122224 672948 122226
rect 669221 122168 669226 122224
rect 669282 122168 672948 122224
rect 669221 122166 672948 122168
rect 669221 122163 669287 122166
rect 672942 122164 672948 122166
rect 673012 122164 673018 122228
rect 676070 122028 676076 122092
rect 676140 122090 676146 122092
rect 676262 122090 676322 122332
rect 676140 122030 676322 122090
rect 676140 122028 676146 122030
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 579521 121138 579587 121141
rect 575798 121136 579587 121138
rect 575798 121080 579526 121136
rect 579582 121080 579587 121136
rect 575798 121078 579587 121080
rect 575798 120836 575858 121078
rect 579521 121075 579587 121078
rect 668945 120866 669011 120869
rect 666694 120864 669011 120866
rect 666694 120808 668950 120864
rect 669006 120808 669011 120864
rect 666694 120806 669011 120808
rect 666694 120798 666754 120806
rect 668945 120803 669011 120806
rect 666356 120738 666754 120798
rect 675894 120730 675954 121622
rect 673410 120670 675954 120730
rect 668577 120594 668643 120597
rect 673410 120594 673470 120670
rect 668577 120592 673470 120594
rect 668577 120536 668582 120592
rect 668638 120536 673470 120592
rect 668577 120534 673470 120536
rect 668577 120531 668643 120534
rect 674465 120050 674531 120053
rect 676673 120050 676739 120053
rect 674465 120048 676739 120050
rect 674465 119992 674470 120048
rect 674526 119992 676678 120048
rect 676734 119992 676739 120048
rect 674465 119990 676739 119992
rect 674465 119987 674531 119990
rect 676673 119987 676739 119990
rect 589457 119914 589523 119917
rect 589457 119912 592572 119914
rect 589457 119856 589462 119912
rect 589518 119856 592572 119912
rect 589457 119854 592572 119856
rect 589457 119851 589523 119854
rect 667933 119234 667999 119237
rect 666694 119232 667999 119234
rect 666694 119176 667938 119232
rect 667994 119176 667999 119232
rect 666694 119174 667999 119176
rect 666694 119166 666754 119174
rect 667933 119171 667999 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 578693 118418 578759 118421
rect 575982 118416 578759 118418
rect 575982 118360 578698 118416
rect 578754 118360 578759 118416
rect 575982 118358 578759 118360
rect 578693 118355 578759 118358
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 676438 117948 676444 118012
rect 676508 118010 676514 118012
rect 676806 118010 676812 118012
rect 676508 117950 676812 118010
rect 676508 117948 676514 117950
rect 676806 117948 676812 117950
rect 676876 117948 676882 118012
rect 668025 117602 668091 117605
rect 666694 117600 668091 117602
rect 666694 117544 668030 117600
rect 668086 117544 668091 117600
rect 666694 117542 668091 117544
rect 666694 117534 666754 117542
rect 668025 117539 668091 117542
rect 666356 117474 666754 117534
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 679617 117330 679683 117333
rect 675772 117328 679683 117330
rect 675772 117272 679622 117328
rect 679678 117272 679683 117328
rect 675772 117270 679683 117272
rect 675772 117268 675778 117270
rect 679617 117267 679683 117270
rect 578693 116922 578759 116925
rect 575798 116920 578759 116922
rect 575798 116864 578698 116920
rect 578754 116864 578759 116920
rect 575798 116862 578759 116864
rect 575798 116484 575858 116862
rect 578693 116859 578759 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 671705 115834 671771 115837
rect 666694 115832 671771 115834
rect 666694 115776 671710 115832
rect 671766 115776 671771 115832
rect 666694 115774 671771 115776
rect 671705 115771 671771 115774
rect 590377 115018 590443 115021
rect 590377 115016 592572 115018
rect 590377 114960 590382 115016
rect 590438 114960 592572 115016
rect 590377 114958 592572 114960
rect 590377 114955 590443 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669221 114338 669287 114341
rect 666694 114336 669287 114338
rect 666694 114280 669226 114336
rect 669282 114280 669287 114336
rect 666694 114278 669287 114280
rect 666694 114270 666754 114278
rect 669221 114275 669287 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 675293 113114 675359 113117
rect 676622 113114 676628 113116
rect 675293 113112 676628 113114
rect 675293 113056 675298 113112
rect 675354 113056 676628 113112
rect 675293 113054 676628 113056
rect 675293 113051 675359 113054
rect 676622 113052 676628 113054
rect 676692 113052 676698 113116
rect 672717 112706 672783 112709
rect 666694 112704 672783 112706
rect 666694 112648 672722 112704
rect 672778 112648 672783 112704
rect 666694 112646 672783 112648
rect 666694 112638 666754 112646
rect 672717 112643 672783 112646
rect 666356 112578 666754 112638
rect 579153 112570 579219 112573
rect 575798 112568 579219 112570
rect 575798 112512 579158 112568
rect 579214 112512 579219 112568
rect 575798 112510 579219 112512
rect 575798 112132 575858 112510
rect 579153 112507 579219 112510
rect 589365 111754 589431 111757
rect 589365 111752 592572 111754
rect 589365 111696 589370 111752
rect 589426 111696 592572 111752
rect 589365 111694 592572 111696
rect 589365 111691 589431 111694
rect 672349 111346 672415 111349
rect 675385 111346 675451 111349
rect 672349 111344 675451 111346
rect 672349 111288 672354 111344
rect 672410 111288 675390 111344
rect 675446 111288 675451 111344
rect 672349 111286 675451 111288
rect 672349 111283 672415 111286
rect 675385 111283 675451 111286
rect 668577 111074 668643 111077
rect 674097 111074 674163 111077
rect 666694 111072 668643 111074
rect 666694 111016 668582 111072
rect 668638 111016 668643 111072
rect 666694 111014 668643 111016
rect 666694 111006 666754 111014
rect 668577 111011 668643 111014
rect 673410 111072 674163 111074
rect 673410 111016 674102 111072
rect 674158 111016 674163 111072
rect 673410 111014 674163 111016
rect 666356 110946 666754 111006
rect 668117 110802 668183 110805
rect 673410 110802 673470 111014
rect 674097 111011 674163 111014
rect 668117 110800 673470 110802
rect 668117 110744 668122 110800
rect 668178 110744 673470 110800
rect 668117 110742 673470 110744
rect 668117 110739 668183 110742
rect 578877 110394 578943 110397
rect 575798 110392 578943 110394
rect 575798 110336 578882 110392
rect 578938 110336 578943 110392
rect 575798 110334 578943 110336
rect 575798 109956 575858 110334
rect 578877 110331 578943 110334
rect 673177 110394 673243 110397
rect 675109 110394 675175 110397
rect 673177 110392 675175 110394
rect 673177 110336 673182 110392
rect 673238 110336 675114 110392
rect 675170 110336 675175 110392
rect 673177 110334 675175 110336
rect 673177 110331 673243 110334
rect 675109 110331 675175 110334
rect 590101 110122 590167 110125
rect 590101 110120 592572 110122
rect 590101 110064 590106 110120
rect 590162 110064 592572 110120
rect 590101 110062 592572 110064
rect 590101 110059 590167 110062
rect 666356 109314 666754 109374
rect 666694 109306 666754 109314
rect 668393 109306 668459 109309
rect 666694 109304 668459 109306
rect 666694 109248 668398 109304
rect 668454 109248 668459 109304
rect 666694 109246 668459 109248
rect 668393 109243 668459 109246
rect 675201 109034 675267 109037
rect 676438 109034 676444 109036
rect 675201 109032 676444 109034
rect 675201 108976 675206 109032
rect 675262 108976 676444 109032
rect 675201 108974 676444 108976
rect 675201 108971 675267 108974
rect 676438 108972 676444 108974
rect 676508 108972 676514 109036
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578877 108354 578943 108357
rect 575798 108352 578943 108354
rect 575798 108296 578882 108352
rect 578938 108296 578943 108352
rect 575798 108294 578943 108296
rect 575798 107780 575858 108294
rect 578877 108291 578943 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 671521 107810 671587 107813
rect 666694 107808 671587 107810
rect 666694 107752 671526 107808
rect 671582 107752 671587 107808
rect 666694 107750 671587 107752
rect 666694 107742 666754 107750
rect 671521 107747 671587 107750
rect 666356 107682 666754 107742
rect 589641 106858 589707 106861
rect 673361 106858 673427 106861
rect 675477 106858 675543 106861
rect 589641 106856 592572 106858
rect 589641 106800 589646 106856
rect 589702 106800 592572 106856
rect 589641 106798 592572 106800
rect 673361 106856 675543 106858
rect 673361 106800 673366 106856
rect 673422 106800 675482 106856
rect 675538 106800 675543 106856
rect 673361 106798 675543 106800
rect 589641 106795 589707 106798
rect 673361 106795 673427 106798
rect 675477 106795 675543 106798
rect 666829 106110 666895 106113
rect 666356 106108 666895 106110
rect 666356 106052 666834 106108
rect 666890 106052 666895 106108
rect 666356 106050 666895 106052
rect 666829 106047 666895 106050
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 673913 104682 673979 104685
rect 675109 104682 675175 104685
rect 673913 104680 675175 104682
rect 673913 104624 673918 104680
rect 673974 104624 675114 104680
rect 675170 104624 675175 104680
rect 673913 104622 675175 104624
rect 673913 104619 673979 104622
rect 675109 104619 675175 104622
rect 666356 104418 666754 104478
rect 666694 104410 666754 104418
rect 668117 104410 668183 104413
rect 666694 104408 668183 104410
rect 666694 104352 668122 104408
rect 668178 104352 668183 104408
rect 666694 104350 668183 104352
rect 668117 104347 668183 104350
rect 590285 103594 590351 103597
rect 590285 103592 592572 103594
rect 590285 103536 590290 103592
rect 590346 103536 592572 103592
rect 590285 103534 592572 103536
rect 590285 103531 590351 103534
rect 575982 103322 576042 103428
rect 578325 103322 578391 103325
rect 575982 103320 578391 103322
rect 575982 103264 578330 103320
rect 578386 103264 578391 103320
rect 575982 103262 578391 103264
rect 578325 103259 578391 103262
rect 675661 103188 675727 103189
rect 675661 103184 675708 103188
rect 675772 103186 675778 103188
rect 675661 103128 675666 103184
rect 675661 103124 675708 103128
rect 675772 103126 675818 103186
rect 675772 103124 675778 103126
rect 675661 103123 675727 103124
rect 666356 102786 666938 102846
rect 666878 102778 666938 102786
rect 667933 102778 667999 102781
rect 666878 102776 673470 102778
rect 666878 102720 667938 102776
rect 667994 102720 673470 102776
rect 666878 102718 673470 102720
rect 667933 102715 667999 102718
rect 673410 102370 673470 102718
rect 675753 102506 675819 102509
rect 676070 102506 676076 102508
rect 675753 102504 676076 102506
rect 675753 102448 675758 102504
rect 675814 102448 676076 102504
rect 675753 102446 676076 102448
rect 675753 102443 675819 102446
rect 676070 102444 676076 102446
rect 676140 102444 676146 102508
rect 674281 102370 674347 102373
rect 673410 102368 674347 102370
rect 673410 102312 674286 102368
rect 674342 102312 674347 102368
rect 673410 102310 674347 102312
rect 674281 102307 674347 102310
rect 589917 101962 589983 101965
rect 589917 101960 592572 101962
rect 589917 101904 589922 101960
rect 589978 101904 592572 101960
rect 589917 101902 592572 101904
rect 589917 101899 589983 101902
rect 578509 101690 578575 101693
rect 575798 101688 578575 101690
rect 575798 101632 578514 101688
rect 578570 101632 578575 101688
rect 575798 101630 578575 101632
rect 575798 101252 575858 101630
rect 578509 101627 578575 101630
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 579153 99242 579219 99245
rect 575798 99240 579219 99242
rect 575798 99184 579158 99240
rect 579214 99184 579219 99240
rect 575798 99182 579219 99184
rect 575798 99076 575858 99182
rect 579153 99179 579219 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 635549 96386 635615 96389
rect 647417 96386 647483 96389
rect 635549 96384 647483 96386
rect 635549 96328 635554 96384
rect 635610 96328 647422 96384
rect 647478 96328 647483 96384
rect 635549 96326 647483 96328
rect 635549 96323 635615 96326
rect 647417 96323 647483 96326
rect 634670 96052 634676 96116
rect 634740 96114 634746 96116
rect 635733 96114 635799 96117
rect 634740 96112 635799 96114
rect 634740 96056 635738 96112
rect 635794 96056 635799 96112
rect 634740 96054 635799 96056
rect 634740 96052 634746 96054
rect 635733 96051 635799 96054
rect 641989 96114 642055 96117
rect 647182 96114 647188 96116
rect 641989 96112 647188 96114
rect 641989 96056 641994 96112
rect 642050 96056 647188 96112
rect 641989 96054 647188 96056
rect 641989 96051 642055 96054
rect 647182 96052 647188 96054
rect 647252 96052 647258 96116
rect 611997 95842 612063 95845
rect 668117 95842 668183 95845
rect 611997 95840 668183 95842
rect 611997 95784 612002 95840
rect 612058 95784 668122 95840
rect 668178 95784 668183 95840
rect 611997 95782 668183 95784
rect 611997 95779 612063 95782
rect 668117 95779 668183 95782
rect 579521 95026 579587 95029
rect 575798 95024 579587 95026
rect 575798 94968 579526 95024
rect 579582 94968 579587 95024
rect 575798 94966 579587 94968
rect 575798 94724 575858 94966
rect 579521 94963 579587 94966
rect 647141 95026 647207 95029
rect 647141 95024 647434 95026
rect 647141 94968 647146 95024
rect 647202 94968 647434 95024
rect 647141 94966 647434 94968
rect 647141 94963 647207 94966
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94966
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 655053 94210 655119 94213
rect 655053 94208 656788 94210
rect 655053 94152 655058 94208
rect 655114 94152 656788 94208
rect 655053 94150 656788 94152
rect 655053 94147 655119 94150
rect 625981 93666 626047 93669
rect 625981 93664 628268 93666
rect 625981 93608 625986 93664
rect 626042 93608 628268 93664
rect 625981 93606 628268 93608
rect 625981 93603 626047 93606
rect 655421 93394 655487 93397
rect 665357 93394 665423 93397
rect 655421 93392 656788 93394
rect 655421 93336 655426 93392
rect 655482 93336 656788 93392
rect 655421 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 655421 93331 655487 93334
rect 665357 93331 665423 93334
rect 579153 93122 579219 93125
rect 575798 93120 579219 93122
rect 575798 93064 579158 93120
rect 579214 93064 579219 93120
rect 575798 93062 579219 93064
rect 575798 92548 575858 93062
rect 579153 93059 579219 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626441 92850 626507 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 626441 92787 626507 92790
rect 656758 92548 656818 93062
rect 663701 92850 663767 92853
rect 663382 92848 663767 92850
rect 663382 92792 663706 92848
rect 663762 92792 663767 92848
rect 663382 92790 663767 92792
rect 663382 92548 663442 92790
rect 663701 92787 663767 92790
rect 625797 92034 625863 92037
rect 648613 92034 648679 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648679 92034
rect 648140 91976 648618 92032
rect 648674 91976 648679 92032
rect 648140 91974 648679 91976
rect 625797 91971 625863 91974
rect 648613 91971 648679 91974
rect 664529 91762 664595 91765
rect 663596 91760 664595 91762
rect 663596 91704 664534 91760
rect 664590 91704 664595 91760
rect 663596 91702 664595 91704
rect 664529 91699 664595 91702
rect 654685 91490 654751 91493
rect 654685 91488 656788 91490
rect 654685 91432 654690 91488
rect 654746 91432 656788 91488
rect 654685 91430 656788 91432
rect 654685 91427 654751 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 578509 90946 578575 90949
rect 575798 90944 578575 90946
rect 575798 90888 578514 90944
rect 578570 90888 578575 90944
rect 575798 90886 578575 90888
rect 575798 90372 575858 90886
rect 578509 90883 578575 90886
rect 655421 90674 655487 90677
rect 664161 90674 664227 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 664227 90674
rect 663596 90616 664166 90672
rect 664222 90616 664227 90672
rect 663596 90614 664227 90616
rect 655421 90611 655487 90614
rect 664161 90611 664227 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664345 89858 664411 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664411 89858
rect 663596 89800 664350 89856
rect 664406 89800 664411 89856
rect 663596 89798 664411 89800
rect 655789 89795 655855 89798
rect 664345 89795 664411 89798
rect 626257 89586 626323 89589
rect 650269 89586 650335 89589
rect 626257 89584 628268 89586
rect 626257 89528 626262 89584
rect 626318 89528 628268 89584
rect 626257 89526 628268 89528
rect 648140 89584 650335 89586
rect 648140 89528 650274 89584
rect 650330 89528 650335 89584
rect 648140 89526 650335 89528
rect 626257 89523 626323 89526
rect 650269 89523 650335 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 626441 88770 626507 88773
rect 626441 88768 628268 88770
rect 626441 88712 626446 88768
rect 626502 88712 628268 88768
rect 626441 88710 628268 88712
rect 626441 88707 626507 88710
rect 575982 88090 576042 88196
rect 578509 88090 578575 88093
rect 575982 88088 578575 88090
rect 575982 88032 578514 88088
rect 578570 88032 578575 88088
rect 575982 88030 578575 88032
rect 578509 88027 578575 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 625613 87138 625679 87141
rect 650545 87138 650611 87141
rect 625613 87136 628268 87138
rect 625613 87080 625618 87136
rect 625674 87080 628268 87136
rect 625613 87078 628268 87080
rect 648140 87136 650611 87138
rect 648140 87080 650550 87136
rect 650606 87080 650611 87136
rect 648140 87078 650611 87080
rect 625613 87075 625679 87078
rect 650545 87075 650611 87078
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 649993 84690 650059 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 650059 84690
rect 648140 84632 649998 84688
rect 650054 84632 650059 84688
rect 648140 84630 650059 84632
rect 625245 84627 625311 84630
rect 649993 84627 650059 84630
rect 579521 84010 579587 84013
rect 575798 84008 579587 84010
rect 575798 83952 579526 84008
rect 579582 83952 579587 84008
rect 575798 83950 579587 83952
rect 575798 83844 575858 83950
rect 579521 83947 579587 83950
rect 626441 83874 626507 83877
rect 626441 83872 628268 83874
rect 626441 83816 626446 83872
rect 626502 83816 628268 83872
rect 626441 83814 628268 83816
rect 626441 83811 626507 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 578509 82242 578575 82245
rect 648889 82242 648955 82245
rect 575798 82240 578575 82242
rect 575798 82184 578514 82240
rect 578570 82184 578575 82240
rect 648140 82240 648955 82242
rect 575798 82182 578575 82184
rect 575798 81668 575858 82182
rect 578509 82179 578575 82182
rect 628790 81698 628850 82212
rect 648140 82184 648894 82240
rect 648950 82184 648955 82240
rect 648140 82182 648955 82184
rect 648889 82179 648955 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 579337 80066 579403 80069
rect 575798 80064 579403 80066
rect 575798 80008 579342 80064
rect 579398 80008 579403 80064
rect 575798 80006 579403 80008
rect 575798 79492 575858 80006
rect 579337 80003 579403 80006
rect 578509 77890 578575 77893
rect 575798 77888 578575 77890
rect 575798 77832 578514 77888
rect 578570 77832 578575 77888
rect 575798 77830 578575 77832
rect 575798 77316 575858 77830
rect 578509 77827 578575 77830
rect 580441 77890 580507 77893
rect 637062 77890 637068 77892
rect 580441 77888 637068 77890
rect 580441 77832 580446 77888
rect 580502 77832 637068 77888
rect 580441 77830 637068 77832
rect 580441 77827 580507 77830
rect 637062 77828 637068 77830
rect 637132 77890 637138 77892
rect 639597 77890 639663 77893
rect 637132 77888 639663 77890
rect 637132 77832 639602 77888
rect 639658 77832 639663 77888
rect 637132 77830 639663 77832
rect 637132 77828 637138 77830
rect 639597 77827 639663 77830
rect 633893 77618 633959 77621
rect 634670 77618 634676 77620
rect 633893 77616 634676 77618
rect 633893 77560 633898 77616
rect 633954 77560 634676 77616
rect 633893 77558 634676 77560
rect 633893 77555 633959 77558
rect 634670 77556 634676 77558
rect 634740 77556 634746 77620
rect 625981 75986 626047 75989
rect 633893 75986 633959 75989
rect 625981 75984 633959 75986
rect 625981 75928 625986 75984
rect 626042 75928 633898 75984
rect 633954 75928 633959 75984
rect 625981 75926 633959 75928
rect 625981 75923 626047 75926
rect 633893 75923 633959 75926
rect 579061 75714 579127 75717
rect 575798 75712 579127 75714
rect 575798 75656 579066 75712
rect 579122 75656 579127 75712
rect 575798 75654 579127 75656
rect 575798 75140 575858 75654
rect 579061 75651 579127 75654
rect 646313 74218 646379 74221
rect 646270 74216 646379 74218
rect 646270 74160 646318 74216
rect 646374 74160 646379 74216
rect 646270 74155 646379 74160
rect 646270 73848 646330 74155
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 646497 71770 646563 71773
rect 646454 71768 646563 71770
rect 646454 71712 646502 71768
rect 646558 71712 646563 71768
rect 646454 71707 646563 71712
rect 646454 71400 646514 71707
rect 578509 71226 578575 71229
rect 575798 71224 578575 71226
rect 575798 71168 578514 71224
rect 578570 71168 578575 71224
rect 575798 71166 578575 71168
rect 575798 70788 575858 71166
rect 578509 71163 578575 71166
rect 646129 69186 646195 69189
rect 646086 69184 646195 69186
rect 646086 69128 646134 69184
rect 646190 69128 646195 69184
rect 646086 69123 646195 69128
rect 646086 68952 646146 69123
rect 575468 66342 575802 68636
rect 648705 67146 648771 67149
rect 646638 67144 648771 67146
rect 646638 67088 648710 67144
rect 648766 67088 648771 67144
rect 646638 67086 648771 67088
rect 646638 66504 646698 67086
rect 648705 67083 648771 67086
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 647233 64426 647299 64429
rect 646638 64424 647299 64426
rect 646638 64368 647238 64424
rect 647294 64368 647299 64424
rect 646638 64366 647299 64368
rect 646638 64056 646698 64366
rect 647233 64363 647299 64366
rect 648889 62114 648955 62117
rect 646638 62112 648955 62114
rect 575982 61842 576042 62084
rect 646638 62056 648894 62112
rect 648950 62056 648955 62112
rect 646638 62054 648955 62056
rect 579521 61842 579587 61845
rect 575982 61840 579587 61842
rect 575982 61784 579526 61840
rect 579582 61784 579587 61840
rect 575982 61782 579587 61784
rect 579521 61779 579587 61782
rect 646638 61608 646698 62054
rect 648889 62051 648955 62054
rect 579521 60346 579587 60349
rect 575798 60344 579587 60346
rect 575798 60288 579526 60344
rect 579582 60288 579587 60344
rect 575798 60286 579587 60288
rect 575798 59908 575858 60286
rect 579521 60283 579587 60286
rect 646129 59394 646195 59397
rect 646086 59392 646195 59394
rect 646086 59336 646134 59392
rect 646190 59336 646195 59392
rect 646086 59331 646195 59336
rect 646086 59160 646146 59331
rect 579337 57898 579403 57901
rect 575798 57896 579403 57898
rect 575798 57840 579342 57896
rect 579398 57840 579403 57896
rect 575798 57838 579403 57840
rect 575798 57732 575858 57838
rect 579337 57835 579403 57838
rect 647417 57354 647483 57357
rect 646638 57352 647483 57354
rect 646638 57296 647422 57352
rect 647478 57296 647483 57352
rect 646638 57294 647483 57296
rect 646638 56712 646698 57294
rect 647417 57291 647483 57294
rect 578509 56130 578575 56133
rect 575798 56128 578575 56130
rect 575798 56072 578514 56128
rect 578570 56072 578575 56128
rect 575798 56070 578575 56072
rect 575798 55556 575858 56070
rect 578509 56067 578575 56070
rect 574737 55042 574803 55045
rect 459510 55040 574803 55042
rect 459510 54984 574742 55040
rect 574798 54984 574803 55040
rect 459510 54982 574803 54984
rect 459510 53685 459570 54982
rect 574737 54979 574803 54982
rect 462630 54708 462636 54772
rect 462700 54770 462706 54772
rect 584397 54770 584463 54773
rect 462700 54768 584463 54770
rect 462700 54712 584402 54768
rect 584458 54712 584463 54768
rect 462700 54710 584463 54712
rect 462700 54708 462706 54710
rect 584397 54707 584463 54710
rect 581637 54498 581703 54501
rect 459878 54496 581703 54498
rect 459878 54440 581642 54496
rect 581698 54440 581703 54496
rect 459878 54438 581703 54440
rect 459878 53685 459938 54438
rect 581637 54435 581703 54438
rect 575473 54226 575539 54229
rect 460798 54224 575539 54226
rect 460798 54168 575478 54224
rect 575534 54168 575539 54224
rect 460798 54166 575539 54168
rect 460798 53685 460858 54166
rect 575473 54163 575539 54166
rect 577681 53954 577747 53957
rect 461718 53952 577747 53954
rect 461718 53896 577686 53952
rect 577742 53896 577747 53952
rect 461718 53894 577747 53896
rect 461718 53685 461778 53894
rect 577681 53891 577747 53894
rect 459461 53680 459570 53685
rect 459461 53624 459466 53680
rect 459522 53624 459570 53680
rect 459461 53622 459570 53624
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459461 53619 459527 53622
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 462589 53619 462655 53620
rect 194358 48860 194364 48924
rect 194428 48922 194434 48924
rect 308029 48922 308095 48925
rect 194428 48920 308095 48922
rect 194428 48864 308034 48920
rect 308090 48864 308095 48920
rect 194428 48862 308095 48864
rect 194428 48860 194434 48862
rect 308029 48859 308095 48862
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 662413 48514 662479 48517
rect 662094 48512 662479 48514
rect 661480 48456 662418 48512
rect 662474 48456 662479 48512
rect 661480 48454 662479 48456
rect 661480 48452 662154 48454
rect 662413 48451 662479 48454
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661585 47791 661651 47794
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47789 661651 47791
rect 661388 47733 661590 47789
rect 661646 47733 661651 47789
rect 661388 47731 661651 47733
rect 661585 47728 661651 47731
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662597 47426 662663 47429
rect 661388 47424 662663 47426
rect 661388 47368 662602 47424
rect 662658 47368 662663 47424
rect 661388 47366 662663 47368
rect 662597 47363 662663 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 463693 44436 463759 44437
rect 463693 44432 463740 44436
rect 463804 44434 463810 44436
rect 463693 44376 463698 44432
rect 463693 44372 463740 44376
rect 463804 44374 463850 44434
rect 463804 44372 463810 44374
rect 463693 44371 463759 44372
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 464102 44236 464108 44300
rect 464172 44298 464178 44300
rect 464337 44298 464403 44301
rect 464172 44296 464403 44298
rect 464172 44240 464342 44296
rect 464398 44240 464403 44296
rect 464172 44238 464403 44240
rect 464172 44236 464178 44238
rect 464337 44235 464403 44238
rect 307293 44162 307359 44165
rect 463877 44162 463943 44165
rect 307293 44160 463943 44162
rect 307293 44104 307298 44160
rect 307354 44104 463882 44160
rect 463938 44104 463943 44160
rect 307293 44102 463943 44104
rect 307293 44099 307359 44102
rect 463877 44099 463943 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 419717 43890 419783 43893
rect 440182 43890 440188 43892
rect 419717 43888 440188 43890
rect 419717 43832 419722 43888
rect 419778 43832 440188 43888
rect 419717 43830 440188 43832
rect 419717 43827 419783 43830
rect 440182 43828 440188 43830
rect 440252 43828 440258 43892
rect 440918 43828 440924 43892
rect 440988 43890 440994 43892
rect 456057 43890 456123 43893
rect 461945 43890 462011 43893
rect 440988 43888 456123 43890
rect 440988 43832 456062 43888
rect 456118 43832 456123 43888
rect 440988 43830 456123 43832
rect 440988 43828 440994 43830
rect 456057 43827 456123 43830
rect 460890 43888 462011 43890
rect 460890 43832 461950 43888
rect 462006 43832 462011 43888
rect 460890 43830 462011 43832
rect 415393 43618 415459 43621
rect 439589 43618 439655 43621
rect 415393 43616 439655 43618
rect 415393 43560 415398 43616
rect 415454 43560 439594 43616
rect 439650 43560 439655 43616
rect 415393 43558 439655 43560
rect 415393 43555 415459 43558
rect 439589 43555 439655 43558
rect 441613 43618 441679 43621
rect 460890 43618 460950 43830
rect 461945 43827 462011 43830
rect 462681 43890 462747 43893
rect 465809 43890 465875 43893
rect 462681 43888 465875 43890
rect 462681 43832 462686 43888
rect 462742 43832 465814 43888
rect 465870 43832 465875 43888
rect 462681 43830 465875 43832
rect 462681 43827 462747 43830
rect 465809 43827 465875 43830
rect 441613 43616 460950 43618
rect 441613 43560 441618 43616
rect 441674 43560 460950 43616
rect 441613 43558 460950 43560
rect 461761 43618 461827 43621
rect 463693 43618 463759 43621
rect 461761 43616 463759 43618
rect 461761 43560 461766 43616
rect 461822 43560 463698 43616
rect 463754 43560 463759 43616
rect 461761 43558 463759 43560
rect 441613 43555 441679 43558
rect 461761 43555 461827 43558
rect 463693 43555 463759 43558
rect 456057 43346 456123 43349
rect 462865 43346 462931 43349
rect 456057 43344 462931 43346
rect 456057 43288 456062 43344
rect 456118 43288 462870 43344
rect 462926 43288 462931 43344
rect 456057 43286 462931 43288
rect 456057 43283 456123 43286
rect 462865 43283 462931 43286
rect 460749 43074 460815 43077
rect 460749 43072 470610 43074
rect 460749 43016 460754 43072
rect 460810 43016 470610 43072
rect 460749 43014 470610 43016
rect 460749 43011 460815 43014
rect 470550 42938 470610 43014
rect 470550 42878 471162 42938
rect 471102 42805 471162 42878
rect 471102 42800 471211 42805
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 471102 42744 471150 42800
rect 471206 42744 471211 42800
rect 471102 42742 471211 42744
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 471145 42739 471211 42742
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 460933 42394 460999 42397
rect 451230 42392 460999 42394
rect 451230 42336 460938 42392
rect 460994 42336 460999 42392
rect 451230 42334 460999 42336
rect 416681 42258 416747 42261
rect 446397 42258 446463 42261
rect 451230 42258 451290 42334
rect 460933 42331 460999 42334
rect 416681 42256 427830 42258
rect 416681 42200 416686 42256
rect 416742 42200 427830 42256
rect 416681 42198 427830 42200
rect 416681 42195 416747 42198
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 194317 42059 194383 42060
rect 361941 41852 362007 41853
rect 361941 41848 361988 41852
rect 362052 41850 362058 41852
rect 365161 41850 365227 41853
rect 365478 41850 365484 41852
rect 361941 41792 361946 41848
rect 361941 41788 361988 41792
rect 362052 41790 362098 41850
rect 365161 41848 365484 41850
rect 365161 41792 365166 41848
rect 365222 41792 365484 41848
rect 365161 41790 365484 41792
rect 362052 41788 362058 41790
rect 361941 41787 362007 41788
rect 365161 41787 365227 41790
rect 365478 41788 365484 41790
rect 365548 41788 365554 41852
rect 403014 41788 403020 41852
rect 403084 41850 403090 41852
rect 421966 41850 421972 41852
rect 403084 41790 421972 41850
rect 403084 41788 403090 41790
rect 421966 41788 421972 41790
rect 422036 41788 422042 41852
rect 427770 41578 427830 42198
rect 446397 42256 451290 42258
rect 446397 42200 446402 42256
rect 446458 42200 451290 42256
rect 446397 42198 451290 42200
rect 446397 42195 446463 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 464102 41850 464108 41852
rect 441908 41790 464108 41850
rect 441908 41788 441914 41790
rect 464102 41788 464108 41790
rect 464172 41788 464178 41852
rect 446397 41578 446463 41581
rect 427770 41576 446463 41578
rect 427770 41520 446402 41576
rect 446458 41520 446463 41576
rect 427770 41518 446463 41520
rect 446397 41515 446463 41518
rect 141693 40492 141759 40493
rect 141693 40488 141740 40492
rect 141804 40490 141810 40492
rect 141693 40432 141698 40488
rect 141693 40428 141740 40432
rect 141804 40430 141850 40490
rect 141804 40428 141810 40430
rect 141693 40427 141759 40428
<< via3 >>
rect 524092 997792 524156 997796
rect 524092 997736 524106 997792
rect 524106 997736 524156 997792
rect 84700 997188 84764 997252
rect 245700 997188 245764 997252
rect 290412 997188 290476 997252
rect 524092 997732 524156 997736
rect 557212 997732 557276 997796
rect 298324 997188 298388 997252
rect 390876 997188 390940 997252
rect 85988 996916 86052 996980
rect 189028 996916 189092 996980
rect 291884 996916 291948 996980
rect 627868 996916 627932 996980
rect 88564 996644 88628 996708
rect 140268 996236 140332 996300
rect 132356 995964 132420 996028
rect 84700 995752 84764 995756
rect 84700 995696 84714 995752
rect 84714 995696 84764 995752
rect 84700 995692 84764 995696
rect 88564 995692 88628 995756
rect 192524 996372 192588 996436
rect 172652 996236 172716 996300
rect 241652 996236 241716 996300
rect 132540 995692 132604 995756
rect 90036 995420 90100 995484
rect 132356 995344 132420 995348
rect 132356 995288 132406 995344
rect 132406 995288 132420 995344
rect 132356 995284 132420 995288
rect 140820 995284 140884 995348
rect 189028 995556 189092 995620
rect 190684 995284 190748 995348
rect 192524 995344 192588 995348
rect 192524 995288 192538 995344
rect 192538 995288 192588 995344
rect 192524 995284 192588 995288
rect 85988 995148 86052 995212
rect 90036 994604 90100 994668
rect 298324 996644 298388 996708
rect 474780 996508 474844 996572
rect 294828 996372 294892 996436
rect 394924 996372 394988 996436
rect 475884 996372 475948 996436
rect 478460 996372 478524 996436
rect 474228 996236 474292 996300
rect 294828 995752 294892 995756
rect 294828 995696 294842 995752
rect 294842 995696 294892 995752
rect 294828 995692 294892 995696
rect 290412 995616 290476 995620
rect 290412 995560 290462 995616
rect 290462 995560 290476 995616
rect 290412 995556 290476 995560
rect 241652 995420 241716 995484
rect 246436 995420 246500 995484
rect 474228 995692 474292 995756
rect 528140 996508 528204 996572
rect 631732 996644 631796 996708
rect 633940 996372 634004 996436
rect 390876 995420 390940 995484
rect 394924 995480 394988 995484
rect 394924 995424 394974 995480
rect 394974 995424 394988 995480
rect 394924 995420 394988 995424
rect 474780 995616 474844 995620
rect 474780 995560 474794 995616
rect 474794 995560 474844 995616
rect 474780 995556 474844 995560
rect 478460 995284 478524 995348
rect 528876 995964 528940 996028
rect 523724 995828 523788 995892
rect 532188 995752 532252 995756
rect 532188 995696 532238 995752
rect 532238 995696 532252 995752
rect 532188 995692 532252 995696
rect 525564 995284 525628 995348
rect 475884 995012 475948 995076
rect 291884 994800 291948 994804
rect 291884 994744 291898 994800
rect 291898 994744 291948 994800
rect 291884 994740 291948 994744
rect 528324 995284 528388 995348
rect 528876 995344 528940 995348
rect 538076 995556 538140 995620
rect 630628 995964 630692 996028
rect 627868 995480 627932 995484
rect 627868 995424 627918 995480
rect 627918 995424 627932 995480
rect 627868 995420 627932 995424
rect 630628 995420 630692 995484
rect 633940 995480 634004 995484
rect 633940 995424 633990 995480
rect 633990 995424 634004 995480
rect 633940 995420 634004 995424
rect 634492 995420 634556 995484
rect 528876 995288 528926 995344
rect 528926 995288 528940 995344
rect 528876 995284 528940 995288
rect 631732 995344 631796 995348
rect 631732 995288 631746 995344
rect 631746 995288 631796 995344
rect 631732 995284 631796 995288
rect 132540 994060 132604 994124
rect 278636 994196 278700 994260
rect 190684 993924 190748 993988
rect 572668 990932 572732 990996
rect 42012 967192 42076 967196
rect 42012 967136 42026 967192
rect 42026 967136 42076 967192
rect 42012 967132 42076 967136
rect 675708 966512 675772 966516
rect 675708 966456 675722 966512
rect 675722 966456 675772 966512
rect 675708 966452 675772 966456
rect 676076 965092 676140 965156
rect 676812 964684 676876 964748
rect 675524 963384 675588 963388
rect 675524 963328 675538 963384
rect 675538 963328 675588 963384
rect 675524 963324 675588 963328
rect 41460 962100 41524 962164
rect 41276 959788 41340 959852
rect 40540 959108 40604 959172
rect 675524 959108 675588 959172
rect 42564 957884 42628 957948
rect 676628 957748 676692 957812
rect 676996 956388 677060 956452
rect 40724 955436 40788 955500
rect 41460 952172 41524 952236
rect 42564 951900 42628 951964
rect 41276 951764 41340 951828
rect 42012 951628 42076 951692
rect 676812 950676 676876 950740
rect 675708 949180 675772 949244
rect 676076 948772 676140 948836
rect 40540 944556 40604 944620
rect 42380 944556 42444 944620
rect 42196 944284 42260 944348
rect 40724 944012 40788 944076
rect 42012 944012 42076 944076
rect 41828 939388 41892 939452
rect 42196 937756 42260 937820
rect 41828 936532 41892 936596
rect 42012 935716 42076 935780
rect 676996 931908 677060 931972
rect 676628 931500 676692 931564
rect 42196 911976 42260 911980
rect 42196 911920 42246 911976
rect 42246 911920 42260 911976
rect 42196 911916 42260 911920
rect 42012 911780 42076 911844
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 675892 875876 675956 875940
rect 676076 874108 676140 874172
rect 673868 873156 673932 873220
rect 676812 871932 676876 871996
rect 39988 814234 40052 814298
rect 41828 811956 41892 812020
rect 42196 808692 42260 808756
rect 41644 805564 41708 805628
rect 41828 805292 41892 805356
rect 40724 805020 40788 805084
rect 40540 804748 40604 804812
rect 42196 804748 42260 804812
rect 40908 804340 40972 804404
rect 42012 797676 42076 797740
rect 40908 796724 40972 796788
rect 42012 796104 42076 796108
rect 42012 796048 42026 796104
rect 42026 796048 42076 796104
rect 42012 796044 42076 796048
rect 40724 794956 40788 795020
rect 40540 792508 40604 792572
rect 41460 788564 41524 788628
rect 41644 788156 41708 788220
rect 41828 785632 41892 785636
rect 41828 785576 41842 785632
rect 41842 785576 41892 785632
rect 41828 785572 41892 785576
rect 674236 782988 674300 783052
rect 676996 780812 677060 780876
rect 675892 771428 675956 771492
rect 41460 769796 41524 769860
rect 676076 768708 676140 768772
rect 675892 766532 675956 766596
rect 676076 766592 676140 766596
rect 676076 766536 676126 766592
rect 676126 766536 676140 766592
rect 676076 766532 676140 766536
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 40724 764900 40788 764964
rect 676996 761832 677060 761836
rect 676628 761788 676692 761792
rect 676628 761732 676642 761788
rect 676642 761732 676692 761788
rect 676628 761728 676692 761732
rect 676996 761776 677010 761832
rect 677010 761776 677060 761832
rect 676996 761772 677060 761776
rect 673316 760336 673380 760340
rect 673316 760280 673330 760336
rect 673330 760280 673380 760336
rect 673316 760276 673380 760280
rect 41644 759052 41708 759116
rect 42380 758840 42444 758844
rect 42380 758784 42394 758840
rect 42394 758784 42444 758840
rect 42380 758780 42444 758784
rect 42012 757692 42076 757756
rect 41828 757072 41892 757076
rect 41828 757016 41842 757072
rect 41842 757016 41892 757072
rect 41828 757012 41892 757016
rect 673868 756332 673932 756396
rect 41828 755440 41892 755444
rect 41828 755384 41878 755440
rect 41878 755384 41892 755440
rect 41828 755380 41892 755384
rect 42196 754836 42260 754900
rect 42380 754564 42444 754628
rect 42564 753340 42628 753404
rect 42196 752932 42260 752996
rect 42196 752388 42260 752452
rect 42380 752116 42444 752180
rect 42564 751708 42628 751772
rect 40908 751028 40972 751092
rect 40724 750348 40788 750412
rect 40540 749396 40604 749460
rect 42380 746812 42444 746876
rect 42196 745512 42260 745516
rect 42196 745456 42210 745512
rect 42210 745456 42260 745512
rect 42196 745452 42260 745456
rect 41644 745180 41708 745244
rect 41460 744908 41524 744972
rect 42012 744364 42076 744428
rect 671476 742188 671540 742252
rect 674052 738652 674116 738716
rect 674420 738108 674484 738172
rect 672028 732864 672092 732868
rect 672028 732808 672042 732864
rect 672042 732808 672092 732864
rect 672028 732804 672092 732808
rect 675892 729948 675956 730012
rect 676812 729948 676876 730012
rect 673316 728588 673380 728652
rect 672028 728452 672092 728516
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 41828 722332 41892 722396
rect 40356 721708 40420 721772
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 718524 40604 718588
rect 41828 718524 41892 718588
rect 40356 716756 40420 716820
rect 40908 716756 40972 716820
rect 41828 715396 41892 715460
rect 42012 714368 42076 714372
rect 42012 714312 42062 714368
rect 42062 714312 42076 714368
rect 42012 714308 42076 714312
rect 40356 714172 40420 714236
rect 41092 714172 41156 714236
rect 42748 714096 42812 714100
rect 42748 714040 42762 714096
rect 42762 714040 42812 714096
rect 42748 714036 42812 714040
rect 40356 712132 40420 712196
rect 675892 711996 675956 712060
rect 42748 710016 42812 710020
rect 42748 709960 42762 710016
rect 42762 709960 42812 710016
rect 42748 709956 42812 709960
rect 41092 709820 41156 709884
rect 40724 709412 40788 709476
rect 40908 708460 40972 708524
rect 674236 707508 674300 707572
rect 40540 706692 40604 706756
rect 42012 706480 42076 706484
rect 42012 706424 42026 706480
rect 42026 706424 42076 706480
rect 42012 706420 42076 706424
rect 674604 706284 674668 706348
rect 42196 704576 42260 704580
rect 42196 704520 42246 704576
rect 42246 704520 42260 704576
rect 42196 704516 42260 704520
rect 42196 703488 42260 703492
rect 42196 703432 42210 703488
rect 42210 703432 42260 703488
rect 42196 703428 42260 703432
rect 41644 702340 41708 702404
rect 41460 700436 41524 700500
rect 41828 699816 41892 699820
rect 41828 699760 41842 699816
rect 41842 699760 41892 699816
rect 41828 699756 41892 699760
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676996 694044 677060 694108
rect 675340 687108 675404 687172
rect 674052 680988 674116 681052
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 41828 678268 41892 678332
rect 41828 677648 41892 677652
rect 41828 677592 41842 677648
rect 41842 677592 41892 677648
rect 41828 677588 41892 677592
rect 41460 675956 41524 676020
rect 42012 673508 42076 673572
rect 41828 671332 41892 671396
rect 42196 669292 42260 669356
rect 42012 668264 42076 668268
rect 42012 668208 42062 668264
rect 42062 668208 42076 668264
rect 42012 668204 42076 668208
rect 42196 667856 42260 667860
rect 42196 667800 42246 667856
rect 42246 667800 42260 667856
rect 42196 667796 42260 667800
rect 40908 665348 40972 665412
rect 671476 664396 671540 664460
rect 40724 664124 40788 664188
rect 42380 663368 42444 663372
rect 42380 663312 42394 663368
rect 42394 663312 42444 663368
rect 42380 663308 42444 663312
rect 40540 662628 40604 662692
rect 674420 662220 674484 662284
rect 42380 659772 42444 659836
rect 41460 658548 41524 658612
rect 41828 658276 41892 658340
rect 41644 657324 41708 657388
rect 675340 652836 675404 652900
rect 675524 651536 675588 651540
rect 675524 651480 675574 651536
rect 675574 651480 675588 651536
rect 675524 651476 675588 651480
rect 674236 648892 674300 648956
rect 674972 645764 675036 645828
rect 676812 644268 676876 644332
rect 675156 643180 675220 643244
rect 674420 642364 674484 642428
rect 675156 641336 675220 641340
rect 675156 641280 675206 641336
rect 675206 641280 675220 641336
rect 675156 641276 675220 641280
rect 41460 640596 41524 640660
rect 675524 639372 675588 639436
rect 41644 638556 41708 638620
rect 675340 637876 675404 637940
rect 674420 637740 674484 637804
rect 674972 637604 675036 637668
rect 674972 636032 675036 636036
rect 674972 635976 674986 636032
rect 674986 635976 675036 636032
rect 674972 635972 675036 635976
rect 40724 634884 40788 634948
rect 40540 634476 40604 634540
rect 676076 631348 676140 631412
rect 41828 630668 41892 630732
rect 675156 629716 675220 629780
rect 674972 629444 675036 629508
rect 40724 623732 40788 623796
rect 40540 619788 40604 619852
rect 676996 619108 677060 619172
rect 41460 615980 41524 616044
rect 41460 615708 41524 615772
rect 41828 612776 41892 612780
rect 41828 612720 41842 612776
rect 41842 612720 41892 612776
rect 41828 612716 41892 612720
rect 675524 607880 675588 607884
rect 675524 607824 675538 607880
rect 675538 607824 675588 607880
rect 675524 607820 675588 607824
rect 674420 602924 674484 602988
rect 674972 599932 675036 599996
rect 673684 597952 673748 597956
rect 673684 597896 673734 597952
rect 673734 597896 673748 597952
rect 673684 597892 673748 597896
rect 42012 597212 42076 597276
rect 674788 596804 674852 596868
rect 42196 596396 42260 596460
rect 676076 594628 676140 594692
rect 676996 594628 677060 594692
rect 675524 593192 675588 593196
rect 675524 593136 675574 593192
rect 675574 593136 675588 593192
rect 675524 593132 675588 593136
rect 675156 592860 675220 592924
rect 673684 592588 673748 592652
rect 43852 591500 43916 591564
rect 674236 589868 674300 589932
rect 40540 589656 40604 589660
rect 40540 589600 40554 589656
rect 40554 589600 40604 589656
rect 40540 589596 40604 589600
rect 40724 589460 40788 589524
rect 40908 589228 40972 589292
rect 676076 586196 676140 586260
rect 42380 584836 42444 584900
rect 40356 584564 40420 584628
rect 41828 584564 41892 584628
rect 42196 584292 42260 584356
rect 673500 582524 673564 582588
rect 42380 582040 42444 582044
rect 42380 581984 42430 582040
rect 42430 581984 42444 582040
rect 42380 581980 42444 581984
rect 40356 581300 40420 581364
rect 673500 580408 673564 580412
rect 673500 580352 673550 580408
rect 673550 580352 673564 580408
rect 673500 580348 673564 580352
rect 42196 580212 42260 580276
rect 40724 578172 40788 578236
rect 40908 577492 40972 577556
rect 40540 576812 40604 576876
rect 676996 575996 677060 576060
rect 41460 573276 41524 573340
rect 676812 572732 676876 572796
rect 41644 572052 41708 572116
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675524 562728 675588 562732
rect 675524 562672 675574 562728
rect 675574 562672 675588 562728
rect 675524 562668 675588 562672
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676260 557500 676324 557564
rect 41828 553964 41892 554028
rect 676812 553828 676876 553892
rect 41828 553148 41892 553212
rect 41828 551984 41892 551988
rect 41828 551928 41842 551984
rect 41842 551928 41892 551984
rect 41828 551924 41892 551928
rect 675892 550564 675956 550628
rect 676996 550292 677060 550356
rect 675892 547632 675956 547636
rect 675892 547576 675942 547632
rect 675942 547576 675956 547632
rect 675892 547572 675956 547576
rect 676260 547572 676324 547636
rect 676076 546756 676140 546820
rect 675340 545940 675404 546004
rect 40724 545728 40788 545732
rect 40724 545672 40774 545728
rect 40774 545672 40788 545728
rect 40724 545668 40788 545672
rect 40540 545456 40604 545460
rect 40540 545400 40590 545456
rect 40590 545400 40604 545456
rect 40540 545396 40604 545400
rect 675524 545396 675588 545460
rect 40724 536964 40788 537028
rect 40540 535196 40604 535260
rect 674420 533836 674484 533900
rect 41460 529892 41524 529956
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 41644 529076 41708 529140
rect 676996 503644 677060 503708
rect 676812 503372 676876 503436
rect 675892 488820 675956 488884
rect 674604 474812 674668 474876
rect 675340 453868 675404 453932
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 41828 421288 41892 421292
rect 41828 421232 41842 421288
rect 41842 421232 41892 421288
rect 41828 421228 41892 421232
rect 40724 418780 40788 418844
rect 40356 418508 40420 418572
rect 675340 410484 675404 410548
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 41460 401780 41524 401844
rect 676812 401236 676876 401300
rect 41828 398848 41892 398852
rect 41828 398792 41842 398848
rect 41842 398792 41892 398848
rect 41828 398788 41892 398792
rect 676076 398788 676140 398852
rect 676628 396748 676692 396812
rect 676260 395116 676324 395180
rect 676444 394708 676508 394772
rect 675892 388996 675956 389060
rect 41276 387500 41340 387564
rect 675708 387636 675772 387700
rect 41828 387228 41892 387292
rect 676628 384916 676692 384980
rect 41644 381380 41708 381444
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 676076 377980 676140 378044
rect 674788 377844 674852 377908
rect 40908 377708 40972 377772
rect 676260 377300 676324 377364
rect 41460 376892 41524 376956
rect 42012 376484 42076 376548
rect 40356 375668 40420 375732
rect 675892 372948 675956 373012
rect 674788 372540 674852 372604
rect 40356 368596 40420 368660
rect 40908 364244 40972 364308
rect 40724 363564 40788 363628
rect 41828 362944 41892 362948
rect 41828 362888 41878 362944
rect 41878 362888 41892 362944
rect 41828 362884 41892 362888
rect 40540 360028 40604 360092
rect 42012 358728 42076 358732
rect 42012 358672 42062 358728
rect 42062 358672 42076 358728
rect 42012 358668 42076 358672
rect 41460 355676 41524 355740
rect 43852 354240 43916 354244
rect 43852 354184 43902 354240
rect 43902 354184 43916 354240
rect 43852 354180 43916 354184
rect 675524 354180 675588 354244
rect 44220 353772 44284 353836
rect 675708 353772 675772 353836
rect 675340 352956 675404 353020
rect 675892 350916 675956 350980
rect 675892 350296 675956 350300
rect 675892 350240 675906 350296
rect 675906 350240 675956 350296
rect 675892 350236 675956 350240
rect 673868 348468 673932 348532
rect 676628 346564 676692 346628
rect 44404 342892 44468 342956
rect 44220 342620 44284 342684
rect 44404 342076 44468 342140
rect 43668 340444 43732 340508
rect 676260 340308 676324 340372
rect 675892 339356 675956 339420
rect 41460 338132 41524 338196
rect 41828 337724 41892 337788
rect 42932 337316 42996 337380
rect 40540 336908 40604 336972
rect 675340 337240 675404 337244
rect 675340 337184 675390 337240
rect 675390 337184 675404 337240
rect 675340 337180 675404 337184
rect 43116 336908 43180 336972
rect 41644 336500 41708 336564
rect 676444 336500 676508 336564
rect 42748 335684 42812 335748
rect 40724 335276 40788 335340
rect 674788 335820 674852 335884
rect 42748 334324 42812 334388
rect 40908 333644 40972 333708
rect 676628 332284 676692 332348
rect 676076 328340 676140 328404
rect 674788 326844 674852 326908
rect 41828 326768 41892 326772
rect 41828 326712 41842 326768
rect 41842 326712 41892 326768
rect 41828 326708 41892 326712
rect 40908 325348 40972 325412
rect 41828 324864 41892 324868
rect 41828 324808 41878 324864
rect 41878 324808 41892 324864
rect 41828 324804 41892 324808
rect 41460 319908 41524 319972
rect 40724 317460 40788 317524
rect 40540 316644 40604 316708
rect 43116 315964 43180 316028
rect 42932 312700 42996 312764
rect 44220 311476 44284 311540
rect 44404 311264 44468 311268
rect 44404 311208 44418 311264
rect 44418 311208 44468 311264
rect 44404 311204 44468 311208
rect 675708 308756 675772 308820
rect 675892 306716 675956 306780
rect 675892 305900 675956 305964
rect 676030 305084 676094 305148
rect 675708 299372 675772 299436
rect 43668 297604 43732 297668
rect 675892 297332 675956 297396
rect 675340 296788 675404 296852
rect 675524 296516 675588 296580
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676812 295156 676876 295220
rect 41828 292768 41892 292772
rect 41828 292712 41842 292768
rect 41842 292712 41892 292768
rect 41828 292708 41892 292712
rect 40540 292528 40604 292592
rect 40908 292528 40972 292592
rect 41828 292300 41892 292364
rect 675524 292088 675588 292092
rect 675524 292032 675574 292088
rect 675574 292032 675588 292088
rect 675524 292028 675588 292032
rect 676444 291484 676508 291548
rect 675340 289912 675404 289916
rect 675340 289856 675354 289912
rect 675354 289856 675404 289912
rect 675340 289852 675404 289856
rect 676260 286996 676324 287060
rect 676076 283596 676140 283660
rect 675708 282840 675772 282844
rect 675708 282784 675722 282840
rect 675722 282784 675772 282840
rect 675708 282780 675772 282784
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 675892 281148 675956 281212
rect 673868 278564 673932 278628
rect 40908 277884 40972 277948
rect 40724 277612 40788 277676
rect 673868 277612 673932 277676
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 674972 263604 675036 263668
rect 676076 262380 676140 262444
rect 676996 261564 677060 261628
rect 676812 259932 676876 259996
rect 40540 251364 40604 251428
rect 676996 250276 677060 250340
rect 40724 249732 40788 249796
rect 673868 249596 673932 249660
rect 674788 249596 674852 249660
rect 676076 249596 676140 249660
rect 674604 246196 674668 246260
rect 676812 245516 676876 245580
rect 675340 245244 675404 245308
rect 675156 244972 675220 245036
rect 675340 240272 675404 240276
rect 675340 240216 675390 240272
rect 675390 240216 675404 240272
rect 675340 240212 675404 240216
rect 40540 240076 40604 240140
rect 42012 237356 42076 237420
rect 673684 237356 673748 237420
rect 675156 237280 675220 237284
rect 675156 237224 675206 237280
rect 675206 237224 675220 237280
rect 675156 237220 675220 237224
rect 40724 235860 40788 235924
rect 676812 235044 676876 235108
rect 671292 234500 671356 234564
rect 673684 232520 673748 232524
rect 673684 232464 673698 232520
rect 673698 232464 673748 232520
rect 673684 232460 673748 232464
rect 673684 231780 673748 231844
rect 673316 231508 673380 231572
rect 671476 230072 671540 230076
rect 671476 230016 671526 230072
rect 671526 230016 671540 230072
rect 671476 230012 671540 230016
rect 673500 230072 673564 230076
rect 673500 230016 673514 230072
rect 673514 230016 673564 230072
rect 673500 230012 673564 230016
rect 674236 229468 674300 229532
rect 674972 228788 675036 228852
rect 674788 228516 674852 228580
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 672948 226748 673012 226812
rect 673132 226808 673196 226812
rect 673132 226752 673182 226808
rect 673182 226752 673196 226808
rect 673132 226748 673196 226752
rect 671660 225856 671724 225860
rect 671660 225800 671710 225856
rect 671710 225800 671724 225856
rect 671660 225796 671724 225800
rect 672948 225796 673012 225860
rect 672764 225660 672828 225724
rect 673868 225584 673932 225588
rect 673868 225528 673918 225584
rect 673918 225528 673932 225584
rect 673868 225524 673932 225528
rect 670740 225388 670804 225452
rect 671660 224300 671724 224364
rect 671660 224088 671724 224092
rect 671660 224032 671674 224088
rect 671674 224032 671724 224088
rect 671660 224028 671724 224032
rect 673132 224028 673196 224092
rect 670740 223952 670804 223956
rect 670740 223896 670790 223952
rect 670790 223896 670804 223952
rect 670740 223892 670804 223896
rect 672764 223952 672828 223956
rect 672764 223896 672778 223952
rect 672778 223896 672828 223952
rect 672764 223892 672828 223896
rect 674604 223756 674668 223820
rect 674236 222804 674300 222868
rect 675892 222668 675956 222732
rect 672396 221912 672460 221916
rect 672396 221856 672446 221912
rect 672446 221856 672460 221912
rect 672396 221852 672460 221856
rect 673132 220900 673196 220964
rect 674788 220900 674852 220964
rect 674052 220084 674116 220148
rect 518940 219736 519004 219740
rect 518940 219680 518954 219736
rect 518954 219680 519004 219736
rect 518940 219676 519004 219680
rect 528876 219676 528940 219740
rect 562364 219404 562428 219468
rect 563468 219404 563532 219468
rect 571932 219404 571996 219468
rect 572852 219132 572916 219196
rect 675524 218996 675588 219060
rect 499436 218860 499500 218924
rect 572484 218860 572548 218924
rect 496676 218588 496740 218652
rect 666324 218588 666388 218652
rect 676030 218180 676094 218244
rect 573220 218044 573284 218108
rect 501092 217560 501156 217564
rect 501092 217504 501106 217560
rect 501106 217504 501156 217560
rect 501092 217500 501156 217504
rect 503300 217560 503364 217564
rect 503300 217504 503350 217560
rect 503350 217504 503364 217560
rect 503300 217500 503364 217504
rect 503668 217560 503732 217564
rect 503668 217504 503682 217560
rect 503682 217504 503732 217560
rect 503668 217500 503732 217504
rect 506060 217560 506124 217564
rect 506060 217504 506110 217560
rect 506110 217504 506124 217560
rect 506060 217500 506124 217504
rect 509188 217500 509252 217564
rect 592172 217772 592236 217836
rect 591804 217228 591868 217292
rect 674604 217636 674668 217700
rect 503300 216956 503364 217020
rect 586652 216956 586716 217020
rect 675892 216956 675956 217020
rect 518940 216412 519004 216476
rect 528692 216412 528756 216476
rect 528876 216412 528940 216476
rect 503668 216140 503732 216204
rect 501092 215868 501156 215932
rect 509188 215596 509252 215660
rect 506060 215324 506124 215388
rect 667980 215596 668044 215660
rect 669452 215596 669516 215660
rect 675708 215324 675772 215388
rect 528692 215052 528756 215116
rect 586652 215052 586716 215116
rect 676260 215086 676324 215150
rect 669452 214508 669516 214572
rect 669452 213964 669516 214028
rect 672580 214024 672644 214028
rect 672580 213968 672594 214024
rect 672594 213968 672644 214024
rect 672580 213964 672644 213968
rect 674052 212060 674116 212124
rect 669636 211108 669700 211172
rect 676996 211168 677060 211172
rect 676996 211112 677010 211168
rect 677010 211112 677060 211168
rect 676996 211108 677060 211112
rect 41460 208932 41524 208996
rect 40540 208116 40604 208180
rect 40908 207300 40972 207364
rect 40724 206892 40788 206956
rect 42012 205668 42076 205732
rect 669268 205668 669332 205732
rect 669636 205668 669700 205732
rect 676444 205532 676508 205596
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 675524 204232 675588 204236
rect 675524 204176 675538 204232
rect 675538 204176 675588 204232
rect 675524 204172 675588 204176
rect 41828 202132 41892 202196
rect 676812 200636 676876 200700
rect 40540 197100 40604 197164
rect 676260 197100 676324 197164
rect 669268 196012 669332 196076
rect 669636 196012 669700 196076
rect 41828 195800 41892 195804
rect 41828 195744 41842 195800
rect 41842 195744 41892 195800
rect 41828 195740 41892 195744
rect 40908 195332 40972 195396
rect 675892 195196 675956 195260
rect 42012 195120 42076 195124
rect 42012 195064 42026 195120
rect 42026 195064 42076 195120
rect 42012 195060 42076 195064
rect 42012 193156 42076 193220
rect 676076 191524 676140 191588
rect 666508 189756 666572 189820
rect 41460 187172 41524 187236
rect 42012 186416 42076 186420
rect 42012 186360 42062 186416
rect 42062 186360 42076 186416
rect 42012 186356 42076 186360
rect 42196 185872 42260 185876
rect 42196 185816 42210 185872
rect 42210 185816 42260 185872
rect 42196 185812 42260 185816
rect 672948 183500 673012 183564
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675708 170308 675772 170372
rect 675892 167452 675956 167516
rect 669636 167044 669700 167108
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 676444 159292 676508 159356
rect 676628 156300 676692 156364
rect 676260 151540 676324 151604
rect 675708 150376 675772 150380
rect 675708 150320 675722 150376
rect 675722 150320 675772 150376
rect 675708 150316 675772 150320
rect 676076 148412 676140 148476
rect 675892 147596 675956 147660
rect 671292 145284 671356 145348
rect 673684 142156 673748 142220
rect 669452 137396 669516 137460
rect 673132 133860 673196 133924
rect 667980 130596 668044 130660
rect 676628 128556 676692 128620
rect 673500 128420 673564 128484
rect 674052 128148 674116 128212
rect 676444 126516 676508 126580
rect 675892 124884 675956 124948
rect 676812 124476 676876 124540
rect 672948 122708 673012 122772
rect 672948 122164 673012 122228
rect 676076 122028 676140 122092
rect 676444 117948 676508 118012
rect 676812 117948 676876 118012
rect 675708 117268 675772 117332
rect 676628 113052 676692 113116
rect 676444 108972 676508 109036
rect 675892 108020 675956 108084
rect 675708 103184 675772 103188
rect 675708 103128 675722 103184
rect 675722 103128 675772 103184
rect 675708 103124 675772 103128
rect 676076 102444 676140 102508
rect 676260 101356 676324 101420
rect 637252 96868 637316 96932
rect 634676 96052 634740 96116
rect 647188 96052 647252 96116
rect 650316 93060 650380 93124
rect 637068 77828 637132 77892
rect 634676 77556 634740 77620
rect 462636 54708 462700 54772
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 194364 48860 194428 48924
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 463740 44432 463804 44436
rect 463740 44376 463754 44432
rect 463754 44376 463804 44432
rect 463740 44372 463804 44376
rect 141740 43964 141804 44028
rect 464108 44236 464172 44300
rect 440188 43828 440252 43892
rect 440924 43828 440988 43892
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 361988 41848 362052 41852
rect 361988 41792 362002 41848
rect 362002 41792 362052 41848
rect 361988 41788 362052 41792
rect 365484 41788 365548 41852
rect 403020 41788 403084 41852
rect 421972 41788 422036 41852
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 464108 41788 464172 41852
rect 141740 40488 141804 40492
rect 141740 40432 141754 40488
rect 141754 40432 141804 40488
rect 141740 40428 141804 40432
<< metal4 >>
rect 524091 997796 524157 997797
rect 524091 997732 524092 997796
rect 524156 997732 524157 997796
rect 524091 997731 524157 997732
rect 557211 997796 557277 997797
rect 557211 997732 557212 997796
rect 557276 997732 557277 997796
rect 557211 997731 557277 997732
rect 524094 997338 524154 997731
rect 557214 997338 557274 997731
rect 84699 997252 84765 997253
rect 84699 997188 84700 997252
rect 84764 997188 84765 997252
rect 84699 997187 84765 997188
rect 84702 995757 84762 997187
rect 290411 997252 290477 997253
rect 290411 997188 290412 997252
rect 290476 997188 290477 997252
rect 290411 997187 290477 997188
rect 298323 997252 298389 997253
rect 298323 997188 298324 997252
rect 298388 997188 298389 997252
rect 298323 997187 298389 997188
rect 390875 997252 390941 997253
rect 390875 997188 390876 997252
rect 390940 997188 390941 997252
rect 390875 997187 390941 997188
rect 85987 996980 86053 996981
rect 85987 996916 85988 996980
rect 86052 996916 86053 996980
rect 85987 996915 86053 996916
rect 84699 995756 84765 995757
rect 84699 995692 84700 995756
rect 84764 995692 84765 995756
rect 84699 995691 84765 995692
rect 85990 995213 86050 996915
rect 88563 996708 88629 996709
rect 88563 996644 88564 996708
rect 88628 996644 88629 996708
rect 88563 996643 88629 996644
rect 88566 995757 88626 996643
rect 172654 996301 172714 997102
rect 189027 996980 189093 996981
rect 189027 996916 189028 996980
rect 189092 996916 189093 996980
rect 189027 996915 189093 996916
rect 140267 996300 140333 996301
rect 140267 996236 140268 996300
rect 140332 996236 140333 996300
rect 140267 996235 140333 996236
rect 172651 996300 172717 996301
rect 172651 996236 172652 996300
rect 172716 996236 172717 996300
rect 172651 996235 172717 996236
rect 132355 996028 132421 996029
rect 132355 995964 132356 996028
rect 132420 995964 132421 996028
rect 132355 995963 132421 995964
rect 88563 995756 88629 995757
rect 88563 995692 88564 995756
rect 88628 995692 88629 995756
rect 88563 995691 88629 995692
rect 90035 995484 90101 995485
rect 90035 995420 90036 995484
rect 90100 995420 90101 995484
rect 90035 995419 90101 995420
rect 85987 995212 86053 995213
rect 85987 995148 85988 995212
rect 86052 995148 86053 995212
rect 85987 995147 86053 995148
rect 90038 994669 90098 995419
rect 132358 995349 132418 995963
rect 140270 995890 140330 996235
rect 140270 995830 140882 995890
rect 132539 995756 132605 995757
rect 132539 995692 132540 995756
rect 132604 995692 132605 995756
rect 132539 995691 132605 995692
rect 132355 995348 132421 995349
rect 132355 995284 132356 995348
rect 132420 995284 132421 995348
rect 132355 995283 132421 995284
rect 90035 994668 90101 994669
rect 90035 994604 90036 994668
rect 90100 994604 90101 994668
rect 90035 994603 90101 994604
rect 132542 994125 132602 995691
rect 140822 995349 140882 995830
rect 189030 995621 189090 996915
rect 192523 996436 192589 996437
rect 192523 996372 192524 996436
rect 192588 996372 192589 996436
rect 192523 996371 192589 996372
rect 189027 995620 189093 995621
rect 189027 995556 189028 995620
rect 189092 995556 189093 995620
rect 189027 995555 189093 995556
rect 192526 995349 192586 996371
rect 241651 996300 241717 996301
rect 241651 996236 241652 996300
rect 241716 996236 241717 996300
rect 241651 996235 241717 996236
rect 241654 995485 241714 996235
rect 246438 995485 246498 997102
rect 241651 995484 241717 995485
rect 241651 995420 241652 995484
rect 241716 995420 241717 995484
rect 241651 995419 241717 995420
rect 246435 995484 246501 995485
rect 246435 995420 246436 995484
rect 246500 995420 246501 995484
rect 246435 995419 246501 995420
rect 140819 995348 140885 995349
rect 140819 995284 140820 995348
rect 140884 995284 140885 995348
rect 140819 995283 140885 995284
rect 190683 995348 190749 995349
rect 190683 995284 190684 995348
rect 190748 995284 190749 995348
rect 190683 995283 190749 995284
rect 192523 995348 192589 995349
rect 192523 995284 192524 995348
rect 192588 995284 192589 995348
rect 192523 995283 192589 995284
rect 132539 994124 132605 994125
rect 132539 994060 132540 994124
rect 132604 994060 132605 994124
rect 132539 994059 132605 994060
rect 190686 993989 190746 995283
rect 278638 994261 278698 997102
rect 290414 995621 290474 997187
rect 291883 996980 291949 996981
rect 291883 996916 291884 996980
rect 291948 996916 291949 996980
rect 291883 996915 291949 996916
rect 290411 995620 290477 995621
rect 290411 995556 290412 995620
rect 290476 995556 290477 995620
rect 290411 995555 290477 995556
rect 291886 994805 291946 996915
rect 298326 996709 298386 997187
rect 298323 996708 298389 996709
rect 298323 996644 298324 996708
rect 298388 996644 298389 996708
rect 298323 996643 298389 996644
rect 294827 996436 294893 996437
rect 294827 996372 294828 996436
rect 294892 996372 294893 996436
rect 294827 996371 294893 996372
rect 294830 995757 294890 996371
rect 294827 995756 294893 995757
rect 294827 995692 294828 995756
rect 294892 995692 294893 995756
rect 294827 995691 294893 995692
rect 390878 995485 390938 997187
rect 474779 996572 474845 996573
rect 474779 996508 474780 996572
rect 474844 996508 474845 996572
rect 474779 996507 474845 996508
rect 528139 996572 528205 996573
rect 528139 996508 528140 996572
rect 528204 996508 528205 996572
rect 528139 996507 528205 996508
rect 394923 996436 394989 996437
rect 394923 996372 394924 996436
rect 394988 996372 394989 996436
rect 394923 996371 394989 996372
rect 394926 995485 394986 996371
rect 474227 996300 474293 996301
rect 474227 996236 474228 996300
rect 474292 996236 474293 996300
rect 474227 996235 474293 996236
rect 474230 995757 474290 996235
rect 474227 995756 474293 995757
rect 474227 995692 474228 995756
rect 474292 995692 474293 995756
rect 474227 995691 474293 995692
rect 474782 995621 474842 996507
rect 475883 996436 475949 996437
rect 475883 996372 475884 996436
rect 475948 996372 475949 996436
rect 475883 996371 475949 996372
rect 478459 996436 478525 996437
rect 478459 996372 478460 996436
rect 478524 996372 478525 996436
rect 478459 996371 478525 996372
rect 474779 995620 474845 995621
rect 474779 995556 474780 995620
rect 474844 995556 474845 995620
rect 474779 995555 474845 995556
rect 390875 995484 390941 995485
rect 390875 995420 390876 995484
rect 390940 995420 390941 995484
rect 390875 995419 390941 995420
rect 394923 995484 394989 995485
rect 394923 995420 394924 995484
rect 394988 995420 394989 995484
rect 394923 995419 394989 995420
rect 475886 995077 475946 996371
rect 478462 995349 478522 996371
rect 523723 995892 523789 995893
rect 523723 995828 523724 995892
rect 523788 995828 523789 995892
rect 523723 995827 523789 995828
rect 478459 995348 478525 995349
rect 478459 995284 478460 995348
rect 478524 995284 478525 995348
rect 523726 995346 523786 995827
rect 525563 995348 525629 995349
rect 525563 995346 525564 995348
rect 523726 995286 525564 995346
rect 478459 995283 478525 995284
rect 525563 995284 525564 995286
rect 525628 995284 525629 995348
rect 528142 995346 528202 996507
rect 528875 996028 528941 996029
rect 528875 995964 528876 996028
rect 528940 995964 528941 996028
rect 528875 995963 528941 995964
rect 528878 995349 528938 995963
rect 532190 995757 532250 997102
rect 627867 996980 627933 996981
rect 627867 996916 627868 996980
rect 627932 996916 627933 996980
rect 627867 996915 627933 996916
rect 532187 995756 532253 995757
rect 532187 995692 532188 995756
rect 532252 995692 532253 995756
rect 532187 995691 532253 995692
rect 538075 995620 538141 995621
rect 538075 995556 538076 995620
rect 538140 995556 538141 995620
rect 538075 995555 538141 995556
rect 528323 995348 528389 995349
rect 528323 995346 528324 995348
rect 528142 995286 528324 995346
rect 525563 995283 525629 995284
rect 528323 995284 528324 995286
rect 528388 995284 528389 995348
rect 528323 995283 528389 995284
rect 528875 995348 528941 995349
rect 528875 995284 528876 995348
rect 528940 995284 528941 995348
rect 528875 995283 528941 995284
rect 475883 995076 475949 995077
rect 475883 995012 475884 995076
rect 475948 995012 475949 995076
rect 475883 995011 475949 995012
rect 291883 994804 291949 994805
rect 291883 994740 291884 994804
rect 291948 994740 291949 994804
rect 291883 994739 291949 994740
rect 278635 994260 278701 994261
rect 278635 994196 278636 994260
rect 278700 994196 278701 994260
rect 278635 994195 278701 994196
rect 190683 993988 190749 993989
rect 190683 993924 190684 993988
rect 190748 993924 190749 993988
rect 190683 993923 190749 993924
rect 538078 993258 538138 995555
rect 627870 995485 627930 996915
rect 631731 996708 631797 996709
rect 631731 996644 631732 996708
rect 631796 996644 631797 996708
rect 631731 996643 631797 996644
rect 630627 996028 630693 996029
rect 630627 995964 630628 996028
rect 630692 995964 630693 996028
rect 630627 995963 630693 995964
rect 630630 995485 630690 995963
rect 627867 995484 627933 995485
rect 627867 995420 627868 995484
rect 627932 995420 627933 995484
rect 627867 995419 627933 995420
rect 630627 995484 630693 995485
rect 630627 995420 630628 995484
rect 630692 995420 630693 995484
rect 630627 995419 630693 995420
rect 631734 995349 631794 996643
rect 633939 996436 634005 996437
rect 633939 996372 633940 996436
rect 634004 996372 634005 996436
rect 633939 996371 634005 996372
rect 633942 995485 634002 996371
rect 634494 995485 634554 997102
rect 633939 995484 634005 995485
rect 633939 995420 633940 995484
rect 634004 995420 634005 995484
rect 633939 995419 634005 995420
rect 634491 995484 634557 995485
rect 634491 995420 634492 995484
rect 634556 995420 634557 995484
rect 634491 995419 634557 995420
rect 631731 995348 631797 995349
rect 631731 995284 631732 995348
rect 631796 995284 631797 995348
rect 631731 995283 631797 995284
rect 572670 990997 572730 993022
rect 572667 990996 572733 990997
rect 572667 990932 572668 990996
rect 572732 990932 572733 990996
rect 572667 990931 572733 990932
rect 42011 967196 42077 967197
rect 42011 967132 42012 967196
rect 42076 967132 42077 967196
rect 42011 967131 42077 967132
rect 41459 962164 41525 962165
rect 41459 962100 41460 962164
rect 41524 962100 41525 962164
rect 41459 962099 41525 962100
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 944621 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 40539 944620 40605 944621
rect 40539 944556 40540 944620
rect 40604 944556 40605 944620
rect 40539 944555 40605 944556
rect 40726 944077 40786 955435
rect 41278 951829 41338 959787
rect 41462 952237 41522 962099
rect 41459 952236 41525 952237
rect 41459 952172 41460 952236
rect 41524 952172 41525 952236
rect 41459 952171 41525 952172
rect 41275 951828 41341 951829
rect 41275 951764 41276 951828
rect 41340 951764 41341 951828
rect 41275 951763 41341 951764
rect 42014 951693 42074 967131
rect 675707 966516 675773 966517
rect 675707 966452 675708 966516
rect 675772 966452 675773 966516
rect 675707 966451 675773 966452
rect 675523 963388 675589 963389
rect 675523 963324 675524 963388
rect 675588 963324 675589 963388
rect 675523 963323 675589 963324
rect 675526 959173 675586 963323
rect 675523 959172 675589 959173
rect 675523 959108 675524 959172
rect 675588 959108 675589 959172
rect 675523 959107 675589 959108
rect 42563 957948 42629 957949
rect 42563 957884 42564 957948
rect 42628 957884 42629 957948
rect 42563 957883 42629 957884
rect 42566 951965 42626 957883
rect 42563 951964 42629 951965
rect 42563 951900 42564 951964
rect 42628 951900 42629 951964
rect 42563 951899 42629 951900
rect 42011 951692 42077 951693
rect 42011 951628 42012 951692
rect 42076 951628 42077 951692
rect 42011 951627 42077 951628
rect 675710 949245 675770 966451
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675707 949244 675773 949245
rect 675707 949180 675708 949244
rect 675772 949180 675773 949244
rect 675707 949179 675773 949180
rect 676078 948837 676138 965091
rect 676811 964748 676877 964749
rect 676811 964684 676812 964748
rect 676876 964684 676877 964748
rect 676811 964683 676877 964684
rect 676627 957812 676693 957813
rect 676627 957748 676628 957812
rect 676692 957748 676693 957812
rect 676627 957747 676693 957748
rect 676075 948836 676141 948837
rect 676075 948772 676076 948836
rect 676140 948772 676141 948836
rect 676075 948771 676141 948772
rect 42379 944620 42445 944621
rect 42379 944556 42380 944620
rect 42444 944556 42445 944620
rect 42379 944555 42445 944556
rect 42195 944348 42261 944349
rect 42195 944284 42196 944348
rect 42260 944284 42261 944348
rect 42195 944283 42261 944284
rect 40723 944076 40789 944077
rect 40723 944012 40724 944076
rect 40788 944012 40789 944076
rect 40723 944011 40789 944012
rect 42011 944076 42077 944077
rect 42011 944012 42012 944076
rect 42076 944012 42077 944076
rect 42011 944011 42077 944012
rect 41827 939452 41893 939453
rect 41827 939450 41828 939452
rect 41094 939390 41828 939450
rect 41094 935670 41154 939390
rect 41827 939388 41828 939390
rect 41892 939388 41893 939452
rect 41827 939387 41893 939388
rect 42014 937050 42074 944011
rect 42198 937821 42258 944283
rect 42195 937820 42261 937821
rect 42195 937756 42196 937820
rect 42260 937756 42261 937820
rect 42195 937755 42261 937756
rect 41830 936990 42074 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 42011 935780 42077 935781
rect 42011 935716 42012 935780
rect 42076 935778 42077 935780
rect 42382 935778 42442 944555
rect 42076 935718 42442 935778
rect 42076 935716 42077 935718
rect 42011 935715 42077 935716
rect 39990 935610 41154 935670
rect 39990 814299 40050 935610
rect 676630 931565 676690 957747
rect 676814 950741 676874 964683
rect 676995 956452 677061 956453
rect 676995 956388 676996 956452
rect 677060 956388 677061 956452
rect 676995 956387 677061 956388
rect 676811 950740 676877 950741
rect 676811 950676 676812 950740
rect 676876 950676 676877 950740
rect 676811 950675 676877 950676
rect 676998 931973 677058 956387
rect 676995 931972 677061 931973
rect 676995 931908 676996 931972
rect 677060 931908 677061 931972
rect 676995 931907 677061 931908
rect 676627 931564 676693 931565
rect 676627 931500 676628 931564
rect 676692 931500 676693 931564
rect 676627 931499 676693 931500
rect 42195 911980 42261 911981
rect 42195 911916 42196 911980
rect 42260 911916 42261 911980
rect 42195 911915 42261 911916
rect 42011 911844 42077 911845
rect 42011 911780 42012 911844
rect 42076 911780 42077 911844
rect 42011 911779 42077 911780
rect 42014 885461 42074 911779
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911915
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 675891 875940 675957 875941
rect 675891 875876 675892 875940
rect 675956 875876 675957 875940
rect 675891 875875 675957 875876
rect 673867 873220 673933 873221
rect 673867 873156 673868 873220
rect 673932 873156 673933 873220
rect 673867 873155 673933 873156
rect 39987 814298 40053 814299
rect 39987 814234 39988 814298
rect 40052 814234 40053 814298
rect 39987 814233 40053 814234
rect 41827 812020 41893 812021
rect 41827 811956 41828 812020
rect 41892 811956 41893 812020
rect 41827 811955 41893 811956
rect 41830 811610 41890 811955
rect 41462 811550 41890 811610
rect 40723 805084 40789 805085
rect 40723 805020 40724 805084
rect 40788 805020 40789 805084
rect 40723 805019 40789 805020
rect 40539 804812 40605 804813
rect 40539 804748 40540 804812
rect 40604 804748 40605 804812
rect 40539 804747 40605 804748
rect 40542 792573 40602 804747
rect 40726 795021 40786 805019
rect 40907 804404 40973 804405
rect 40907 804340 40908 804404
rect 40972 804340 40973 804404
rect 40907 804339 40973 804340
rect 40910 796789 40970 804339
rect 40907 796788 40973 796789
rect 40907 796724 40908 796788
rect 40972 796724 40973 796788
rect 40907 796723 40973 796724
rect 40723 795020 40789 795021
rect 40723 794956 40724 795020
rect 40788 794956 40789 795020
rect 40723 794955 40789 794956
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 788629 41522 811550
rect 42195 808756 42261 808757
rect 42195 808692 42196 808756
rect 42260 808692 42261 808756
rect 42195 808691 42261 808692
rect 41643 805628 41709 805629
rect 41643 805564 41644 805628
rect 41708 805564 41709 805628
rect 41643 805563 41709 805564
rect 41459 788628 41525 788629
rect 41459 788564 41460 788628
rect 41524 788564 41525 788628
rect 41459 788563 41525 788564
rect 41646 788221 41706 805563
rect 41827 805356 41893 805357
rect 41827 805292 41828 805356
rect 41892 805292 41893 805356
rect 41827 805291 41893 805292
rect 41643 788220 41709 788221
rect 41643 788156 41644 788220
rect 41708 788156 41709 788220
rect 41643 788155 41709 788156
rect 41830 785637 41890 805291
rect 42198 804813 42258 808691
rect 42195 804812 42261 804813
rect 42195 804748 42196 804812
rect 42260 804748 42261 804812
rect 42195 804747 42261 804748
rect 42011 797740 42077 797741
rect 42011 797676 42012 797740
rect 42076 797676 42077 797740
rect 42011 797675 42077 797676
rect 42014 796109 42074 797675
rect 42011 796108 42077 796109
rect 42011 796044 42012 796108
rect 42076 796044 42077 796108
rect 42011 796043 42077 796044
rect 41827 785636 41893 785637
rect 41827 785572 41828 785636
rect 41892 785572 41893 785636
rect 41827 785571 41893 785572
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750413 40786 764899
rect 40910 751093 40970 765715
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40723 750412 40789 750413
rect 40723 750348 40724 750412
rect 40788 750348 40789 750412
rect 40723 750347 40789 750348
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 744973 41522 769795
rect 673315 760340 673381 760341
rect 673315 760276 673316 760340
rect 673380 760276 673381 760340
rect 673315 760275 673381 760276
rect 41643 759116 41709 759117
rect 41643 759052 41644 759116
rect 41708 759052 41709 759116
rect 41643 759051 41709 759052
rect 41646 745245 41706 759051
rect 42379 758844 42445 758845
rect 42379 758780 42380 758844
rect 42444 758780 42445 758844
rect 42379 758779 42445 758780
rect 42011 757756 42077 757757
rect 42011 757692 42012 757756
rect 42076 757692 42077 757756
rect 42011 757691 42077 757692
rect 41827 757076 41893 757077
rect 41827 757012 41828 757076
rect 41892 757012 41893 757076
rect 41827 757011 41893 757012
rect 41830 755445 41890 757011
rect 41827 755444 41893 755445
rect 41827 755380 41828 755444
rect 41892 755380 41893 755444
rect 41827 755379 41893 755380
rect 41643 745244 41709 745245
rect 41643 745180 41644 745244
rect 41708 745180 41709 745244
rect 41643 745179 41709 745180
rect 41459 744972 41525 744973
rect 41459 744908 41460 744972
rect 41524 744908 41525 744972
rect 41459 744907 41525 744908
rect 42014 744429 42074 757691
rect 42195 754900 42261 754901
rect 42195 754836 42196 754900
rect 42260 754836 42261 754900
rect 42195 754835 42261 754836
rect 42198 752997 42258 754835
rect 42382 754629 42442 758779
rect 42379 754628 42445 754629
rect 42379 754564 42380 754628
rect 42444 754564 42445 754628
rect 42379 754563 42445 754564
rect 42563 753404 42629 753405
rect 42563 753340 42564 753404
rect 42628 753340 42629 753404
rect 42563 753339 42629 753340
rect 42195 752996 42261 752997
rect 42195 752932 42196 752996
rect 42260 752932 42261 752996
rect 42195 752931 42261 752932
rect 42195 752452 42261 752453
rect 42195 752388 42196 752452
rect 42260 752388 42261 752452
rect 42195 752387 42261 752388
rect 42198 745517 42258 752387
rect 42379 752180 42445 752181
rect 42379 752116 42380 752180
rect 42444 752116 42445 752180
rect 42379 752115 42445 752116
rect 42382 746877 42442 752115
rect 42566 751773 42626 753339
rect 42563 751772 42629 751773
rect 42563 751708 42564 751772
rect 42628 751708 42629 751772
rect 42563 751707 42629 751708
rect 42379 746876 42445 746877
rect 42379 746812 42380 746876
rect 42444 746812 42445 746876
rect 42379 746811 42445 746812
rect 42195 745516 42261 745517
rect 42195 745452 42196 745516
rect 42260 745452 42261 745516
rect 42195 745451 42261 745452
rect 42011 744428 42077 744429
rect 42011 744364 42012 744428
rect 42076 744364 42077 744428
rect 42011 744363 42077 744364
rect 671475 742252 671541 742253
rect 671475 742188 671476 742252
rect 671540 742188 671541 742252
rect 671475 742187 671541 742188
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40355 721772 40421 721773
rect 40355 721708 40356 721772
rect 40420 721708 40421 721772
rect 40355 721707 40421 721708
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40358 716821 40418 721707
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40355 716820 40421 716821
rect 40355 716756 40356 716820
rect 40420 716756 40421 716820
rect 40355 716755 40421 716756
rect 40355 714236 40421 714237
rect 40355 714172 40356 714236
rect 40420 714172 40421 714236
rect 40355 714171 40421 714172
rect 40358 712197 40418 714171
rect 40355 712196 40421 712197
rect 40355 712132 40356 712196
rect 40420 712132 40421 712196
rect 40355 712131 40421 712132
rect 40542 706757 40602 718523
rect 40726 709477 40786 721707
rect 40907 716820 40973 716821
rect 40907 716756 40908 716820
rect 40972 716756 40973 716820
rect 40907 716755 40973 716756
rect 40723 709476 40789 709477
rect 40723 709412 40724 709476
rect 40788 709412 40789 709476
rect 40723 709411 40789 709412
rect 40910 708525 40970 716755
rect 41091 714236 41157 714237
rect 41091 714172 41092 714236
rect 41156 714172 41157 714236
rect 41091 714171 41157 714172
rect 41094 709885 41154 714171
rect 41091 709884 41157 709885
rect 41091 709820 41092 709884
rect 41156 709820 41157 709884
rect 41091 709819 41157 709820
rect 40907 708524 40973 708525
rect 40907 708460 40908 708524
rect 40972 708460 40973 708524
rect 40907 708459 40973 708460
rect 40539 706756 40605 706757
rect 40539 706692 40540 706756
rect 40604 706692 40605 706756
rect 40539 706691 40605 706692
rect 41462 700501 41522 726550
rect 41827 722396 41893 722397
rect 41827 722332 41828 722396
rect 41892 722332 41893 722396
rect 41827 722331 41893 722332
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41646 702405 41706 721707
rect 41830 718589 41890 722331
rect 41827 718588 41893 718589
rect 41827 718524 41828 718588
rect 41892 718524 41893 718588
rect 41827 718523 41893 718524
rect 41827 715460 41893 715461
rect 41827 715396 41828 715460
rect 41892 715396 41893 715460
rect 41827 715395 41893 715396
rect 41643 702404 41709 702405
rect 41643 702340 41644 702404
rect 41708 702340 41709 702404
rect 41643 702339 41709 702340
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 41830 699821 41890 715395
rect 42011 714372 42077 714373
rect 42011 714308 42012 714372
rect 42076 714308 42077 714372
rect 42011 714307 42077 714308
rect 42014 706485 42074 714307
rect 42747 714100 42813 714101
rect 42747 714036 42748 714100
rect 42812 714036 42813 714100
rect 42747 714035 42813 714036
rect 42750 710021 42810 714035
rect 42747 710020 42813 710021
rect 42747 709956 42748 710020
rect 42812 709956 42813 710020
rect 42747 709955 42813 709956
rect 42011 706484 42077 706485
rect 42011 706420 42012 706484
rect 42076 706420 42077 706484
rect 42011 706419 42077 706420
rect 42195 704580 42261 704581
rect 42195 704516 42196 704580
rect 42260 704516 42261 704580
rect 42195 704515 42261 704516
rect 42198 703493 42258 704515
rect 42195 703492 42261 703493
rect 42195 703428 42196 703492
rect 42260 703428 42261 703492
rect 42195 703427 42261 703428
rect 41827 699820 41893 699821
rect 41827 699756 41828 699820
rect 41892 699756 41893 699820
rect 41827 699755 41893 699756
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40910 678930 41890 678990
rect 40542 662693 40602 678927
rect 40726 664189 40786 678927
rect 40910 665413 40970 678930
rect 41830 678333 41890 678930
rect 41827 678332 41893 678333
rect 41827 678268 41828 678332
rect 41892 678268 41893 678332
rect 41827 678267 41893 678268
rect 41827 677652 41893 677653
rect 41827 677588 41828 677652
rect 41892 677588 41893 677652
rect 41827 677587 41893 677588
rect 41830 676230 41890 677587
rect 41646 676170 41890 676230
rect 41459 676020 41525 676021
rect 41459 675956 41460 676020
rect 41524 675956 41525 676020
rect 41459 675955 41525 675956
rect 40907 665412 40973 665413
rect 40907 665348 40908 665412
rect 40972 665348 40973 665412
rect 40907 665347 40973 665348
rect 40723 664188 40789 664189
rect 40723 664124 40724 664188
rect 40788 664124 40789 664188
rect 40723 664123 40789 664124
rect 40539 662692 40605 662693
rect 40539 662628 40540 662692
rect 40604 662628 40605 662692
rect 40539 662627 40605 662628
rect 41462 658613 41522 675955
rect 41459 658612 41525 658613
rect 41459 658548 41460 658612
rect 41524 658548 41525 658612
rect 41459 658547 41525 658548
rect 41646 657389 41706 676170
rect 42011 673572 42077 673573
rect 42011 673508 42012 673572
rect 42076 673508 42077 673572
rect 42011 673507 42077 673508
rect 41827 671396 41893 671397
rect 41827 671332 41828 671396
rect 41892 671332 41893 671396
rect 41827 671331 41893 671332
rect 41830 658341 41890 671331
rect 42014 668269 42074 673507
rect 42195 669356 42261 669357
rect 42195 669292 42196 669356
rect 42260 669292 42261 669356
rect 42195 669291 42261 669292
rect 42011 668268 42077 668269
rect 42011 668204 42012 668268
rect 42076 668204 42077 668268
rect 42011 668203 42077 668204
rect 42198 667861 42258 669291
rect 42195 667860 42261 667861
rect 42195 667796 42196 667860
rect 42260 667796 42261 667860
rect 42195 667795 42261 667796
rect 671478 664461 671538 742187
rect 672027 732868 672093 732869
rect 672027 732804 672028 732868
rect 672092 732804 672093 732868
rect 672027 732803 672093 732804
rect 672030 728517 672090 732803
rect 673318 728653 673378 760275
rect 673870 756397 673930 873155
rect 674235 783052 674301 783053
rect 674235 782988 674236 783052
rect 674300 782988 674301 783052
rect 674235 782987 674301 782988
rect 673867 756396 673933 756397
rect 673867 756332 673868 756396
rect 673932 756332 673933 756396
rect 673867 756331 673933 756332
rect 674051 738716 674117 738717
rect 674051 738652 674052 738716
rect 674116 738652 674117 738716
rect 674051 738651 674117 738652
rect 673315 728652 673381 728653
rect 673315 728588 673316 728652
rect 673380 728588 673381 728652
rect 673315 728587 673381 728588
rect 672027 728516 672093 728517
rect 672027 728452 672028 728516
rect 672092 728452 672093 728516
rect 672027 728451 672093 728452
rect 674054 681053 674114 738651
rect 674238 707573 674298 782987
rect 675894 771493 675954 875875
rect 676075 874172 676141 874173
rect 676075 874108 676076 874172
rect 676140 874108 676141 874172
rect 676075 874107 676141 874108
rect 675891 771492 675957 771493
rect 675891 771428 675892 771492
rect 675956 771428 675957 771492
rect 675891 771427 675957 771428
rect 676078 768773 676138 874107
rect 676811 871996 676877 871997
rect 676811 871932 676812 871996
rect 676876 871932 676877 871996
rect 676811 871931 676877 871932
rect 676075 768772 676141 768773
rect 676075 768708 676076 768772
rect 676140 768708 676141 768772
rect 676075 768707 676141 768708
rect 675891 766596 675957 766597
rect 675891 766532 675892 766596
rect 675956 766532 675957 766596
rect 675891 766531 675957 766532
rect 676075 766596 676141 766597
rect 676075 766532 676076 766596
rect 676140 766532 676141 766596
rect 676075 766531 676141 766532
rect 674419 738172 674485 738173
rect 674419 738108 674420 738172
rect 674484 738108 674485 738172
rect 674419 738107 674485 738108
rect 674235 707572 674301 707573
rect 674235 707508 674236 707572
rect 674300 707508 674301 707572
rect 674235 707507 674301 707508
rect 674051 681052 674117 681053
rect 674051 680988 674052 681052
rect 674116 680988 674117 681052
rect 674051 680987 674117 680988
rect 671475 664460 671541 664461
rect 671475 664396 671476 664460
rect 671540 664396 671541 664460
rect 671475 664395 671541 664396
rect 42379 663372 42445 663373
rect 42379 663308 42380 663372
rect 42444 663308 42445 663372
rect 42379 663307 42445 663308
rect 42382 659837 42442 663307
rect 674422 662285 674482 738107
rect 675894 730013 675954 766531
rect 675891 730012 675957 730013
rect 675891 729948 675892 730012
rect 675956 729948 675957 730012
rect 675891 729947 675957 729948
rect 676078 725797 676138 766531
rect 676627 761792 676693 761793
rect 676627 761728 676628 761792
rect 676692 761790 676693 761792
rect 676814 761790 676874 871931
rect 676995 780876 677061 780877
rect 676995 780812 676996 780876
rect 677060 780812 677061 780876
rect 676995 780811 677061 780812
rect 676998 761837 677058 780811
rect 676692 761730 676874 761790
rect 676995 761836 677061 761837
rect 676995 761772 676996 761836
rect 677060 761772 677061 761836
rect 676995 761771 677061 761772
rect 676692 761728 676693 761730
rect 676627 761727 676693 761728
rect 676811 730012 676877 730013
rect 676811 729948 676812 730012
rect 676876 729948 676877 730012
rect 676811 729947 676877 729948
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712110 676874 729947
rect 675894 712061 676874 712110
rect 675891 712060 676874 712061
rect 675891 711996 675892 712060
rect 675956 712050 676874 712060
rect 675956 711996 675957 712050
rect 675891 711995 675957 711996
rect 674603 706348 674669 706349
rect 674603 706284 674604 706348
rect 674668 706284 674669 706348
rect 674603 706283 674669 706284
rect 674419 662284 674485 662285
rect 674419 662220 674420 662284
rect 674484 662220 674485 662284
rect 674419 662219 674485 662220
rect 42379 659836 42445 659837
rect 42379 659772 42380 659836
rect 42444 659772 42445 659836
rect 42379 659771 42445 659772
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41643 657388 41709 657389
rect 41643 657324 41644 657388
rect 41708 657324 41709 657388
rect 41643 657323 41709 657324
rect 674235 648956 674301 648957
rect 674235 648892 674236 648956
rect 674300 648892 674301 648956
rect 674235 648891 674301 648892
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40539 634540 40605 634541
rect 40539 634476 40540 634540
rect 40604 634476 40605 634540
rect 40539 634475 40605 634476
rect 40542 619853 40602 634475
rect 40726 623797 40786 634883
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 619852 40605 619853
rect 40539 619788 40540 619852
rect 40604 619788 40605 619852
rect 40539 619787 40605 619788
rect 41462 616045 41522 640595
rect 41643 638620 41709 638621
rect 41643 638556 41644 638620
rect 41708 638556 41709 638620
rect 41643 638555 41709 638556
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41459 615772 41525 615773
rect 41459 615708 41460 615772
rect 41524 615770 41525 615772
rect 41646 615770 41706 638555
rect 41827 630732 41893 630733
rect 41827 630668 41828 630732
rect 41892 630668 41893 630732
rect 41827 630667 41893 630668
rect 41524 615710 41706 615770
rect 41524 615708 41525 615710
rect 41459 615707 41525 615708
rect 41830 612781 41890 630667
rect 41827 612780 41893 612781
rect 41827 612716 41828 612780
rect 41892 612716 41893 612780
rect 41827 612715 41893 612716
rect 673683 597956 673749 597957
rect 673683 597892 673684 597956
rect 673748 597892 673749 597956
rect 673683 597891 673749 597892
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 42014 592242 42074 597211
rect 42195 596460 42261 596461
rect 42195 596396 42196 596460
rect 42260 596396 42261 596460
rect 42195 596395 42261 596396
rect 41462 592182 42074 592242
rect 40539 589660 40605 589661
rect 40539 589596 40540 589660
rect 40604 589596 40605 589660
rect 40539 589595 40605 589596
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 581365 40418 584563
rect 40355 581364 40421 581365
rect 40355 581300 40356 581364
rect 40420 581300 40421 581364
rect 40355 581299 40421 581300
rect 40542 576877 40602 589595
rect 40723 589524 40789 589525
rect 40723 589460 40724 589524
rect 40788 589460 40789 589524
rect 40723 589459 40789 589460
rect 40726 578237 40786 589459
rect 40907 589292 40973 589293
rect 40907 589228 40908 589292
rect 40972 589228 40973 589292
rect 40907 589227 40973 589228
rect 40723 578236 40789 578237
rect 40723 578172 40724 578236
rect 40788 578172 40789 578236
rect 40723 578171 40789 578172
rect 40910 577557 40970 589227
rect 40907 577556 40973 577557
rect 40907 577492 40908 577556
rect 40972 577492 40973 577556
rect 40907 577491 40973 577492
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 573341 41522 592182
rect 42198 589290 42258 596395
rect 673686 592653 673746 597891
rect 673683 592652 673749 592653
rect 673683 592588 673684 592652
rect 673748 592588 673749 592652
rect 673683 592587 673749 592588
rect 43851 591564 43917 591565
rect 43851 591500 43852 591564
rect 43916 591500 43917 591564
rect 43851 591499 43917 591500
rect 41646 589230 42258 589290
rect 41459 573340 41525 573341
rect 41459 573276 41460 573340
rect 41524 573276 41525 573340
rect 41459 573275 41525 573276
rect 41646 572117 41706 589230
rect 42379 584900 42445 584901
rect 42379 584836 42380 584900
rect 42444 584836 42445 584900
rect 42379 584835 42445 584836
rect 41827 584628 41893 584629
rect 41827 584564 41828 584628
rect 41892 584564 41893 584628
rect 41827 584563 41893 584564
rect 41643 572116 41709 572117
rect 41643 572052 41644 572116
rect 41708 572052 41709 572116
rect 41643 572051 41709 572052
rect 41830 570213 41890 584563
rect 42195 584356 42261 584357
rect 42195 584292 42196 584356
rect 42260 584292 42261 584356
rect 42195 584291 42261 584292
rect 42198 580277 42258 584291
rect 42382 582045 42442 584835
rect 42379 582044 42445 582045
rect 42379 581980 42380 582044
rect 42444 581980 42445 582044
rect 42379 581979 42445 581980
rect 42195 580276 42261 580277
rect 42195 580212 42196 580276
rect 42260 580212 42261 580276
rect 42195 580211 42261 580212
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 535261 40602 545395
rect 40726 537029 40786 545667
rect 40723 537028 40789 537029
rect 40723 536964 40724 537028
rect 40788 536964 40789 537028
rect 40723 536963 40789 536964
rect 40539 535260 40605 535261
rect 40539 535196 40540 535260
rect 40604 535196 40605 535260
rect 40539 535195 40605 535196
rect 41462 529957 41522 553350
rect 41827 553212 41893 553213
rect 41827 553210 41828 553212
rect 41646 553150 41828 553210
rect 41459 529956 41525 529957
rect 41459 529892 41460 529956
rect 41524 529892 41525 529956
rect 41459 529891 41525 529892
rect 41646 529141 41706 553150
rect 41827 553148 41828 553150
rect 41892 553148 41893 553212
rect 41827 553147 41893 553148
rect 41827 551988 41893 551989
rect 41827 551924 41828 551988
rect 41892 551924 41893 551988
rect 41827 551923 41893 551924
rect 41830 529413 41890 551923
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 41643 529140 41709 529141
rect 41643 529076 41644 529140
rect 41708 529076 41709 529140
rect 41643 529075 41709 529076
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41462 424630 41890 424690
rect 40723 418844 40789 418845
rect 40723 418780 40724 418844
rect 40788 418780 40789 418844
rect 40723 418779 40789 418780
rect 40355 418572 40421 418573
rect 40355 418508 40356 418572
rect 40420 418508 40421 418572
rect 40355 418507 40421 418508
rect 40358 412650 40418 418507
rect 40358 412590 40602 412650
rect 40542 403885 40602 412590
rect 40726 409461 40786 418779
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 401845 41522 424630
rect 41827 421292 41893 421293
rect 41827 421290 41828 421292
rect 41646 421230 41828 421290
rect 41646 402990 41706 421230
rect 41827 421228 41828 421230
rect 41892 421228 41893 421292
rect 41827 421227 41893 421228
rect 42014 408510 42074 424763
rect 41830 408450 42074 408510
rect 41830 406333 41890 408450
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41459 401844 41525 401845
rect 41459 401780 41460 401844
rect 41524 401780 41525 401844
rect 41459 401779 41525 401780
rect 41830 398853 41890 402930
rect 41827 398852 41893 398853
rect 41827 398788 41828 398852
rect 41892 398788 41893 398852
rect 41827 398787 41893 398788
rect 41275 387564 41341 387565
rect 41275 387500 41276 387564
rect 41340 387500 41341 387564
rect 41275 387499 41341 387500
rect 41278 387290 41338 387499
rect 41827 387292 41893 387293
rect 41827 387290 41828 387292
rect 41278 387230 41828 387290
rect 41827 387228 41828 387230
rect 41892 387228 41893 387292
rect 41827 387227 41893 387228
rect 41643 381444 41709 381445
rect 41643 381380 41644 381444
rect 41708 381380 41709 381444
rect 41643 381379 41709 381380
rect 41646 379530 41706 381379
rect 41646 379470 41890 379530
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40355 375732 40421 375733
rect 40355 375668 40356 375732
rect 40420 375668 40421 375732
rect 40355 375667 40421 375668
rect 40358 368661 40418 375667
rect 40355 368660 40421 368661
rect 40355 368596 40356 368660
rect 40420 368596 40421 368660
rect 40355 368595 40421 368596
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363629 40786 378115
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364309 40970 377707
rect 41459 376956 41525 376957
rect 41459 376892 41460 376956
rect 41524 376892 41525 376956
rect 41459 376891 41525 376892
rect 40907 364308 40973 364309
rect 40907 364244 40908 364308
rect 40972 364244 40973 364308
rect 40907 364243 40973 364244
rect 40723 363628 40789 363629
rect 40723 363564 40724 363628
rect 40788 363564 40789 363628
rect 40723 363563 40789 363564
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 355741 41522 376891
rect 41830 362949 41890 379470
rect 42011 376548 42077 376549
rect 42011 376484 42012 376548
rect 42076 376484 42077 376548
rect 42011 376483 42077 376484
rect 41827 362948 41893 362949
rect 41827 362884 41828 362948
rect 41892 362884 41893 362948
rect 41827 362883 41893 362884
rect 42014 358733 42074 376483
rect 42011 358732 42077 358733
rect 42011 358668 42012 358732
rect 42076 358668 42077 358732
rect 42011 358667 42077 358668
rect 41459 355740 41525 355741
rect 41459 355676 41460 355740
rect 41524 355676 41525 355740
rect 41459 355675 41525 355676
rect 43854 354245 43914 591499
rect 674238 589933 674298 648891
rect 674419 642428 674485 642429
rect 674419 642364 674420 642428
rect 674484 642364 674485 642428
rect 674419 642363 674485 642364
rect 674422 637805 674482 642363
rect 674419 637804 674485 637805
rect 674419 637740 674420 637804
rect 674484 637740 674485 637804
rect 674419 637739 674485 637740
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674235 589932 674301 589933
rect 674235 589868 674236 589932
rect 674300 589868 674301 589932
rect 674235 589867 674301 589868
rect 673499 582588 673565 582589
rect 673499 582524 673500 582588
rect 673564 582524 673565 582588
rect 673499 582523 673565 582524
rect 673502 580413 673562 582523
rect 673499 580412 673565 580413
rect 673499 580348 673500 580412
rect 673564 580348 673565 580412
rect 673499 580347 673565 580348
rect 674422 533901 674482 602923
rect 674419 533900 674485 533901
rect 674419 533836 674420 533900
rect 674484 533836 674485 533900
rect 674419 533835 674485 533836
rect 674606 474877 674666 706283
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 687173 675402 696763
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 675339 687172 675405 687173
rect 675339 687108 675340 687172
rect 675404 687108 675405 687172
rect 675339 687107 675405 687108
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674971 645828 675037 645829
rect 674971 645764 674972 645828
rect 675036 645764 675037 645828
rect 674971 645763 675037 645764
rect 674974 637669 675034 645763
rect 675155 643244 675221 643245
rect 675155 643180 675156 643244
rect 675220 643180 675221 643244
rect 675155 643179 675221 643180
rect 675158 641341 675218 643179
rect 675155 641340 675221 641341
rect 675155 641276 675156 641340
rect 675220 641276 675221 641340
rect 675155 641275 675221 641276
rect 675342 637941 675402 652835
rect 675523 651540 675589 651541
rect 675523 651476 675524 651540
rect 675588 651476 675589 651540
rect 675523 651475 675589 651476
rect 675526 639437 675586 651475
rect 676811 644332 676877 644333
rect 676811 644268 676812 644332
rect 676876 644268 676877 644332
rect 676811 644267 676877 644268
rect 675523 639436 675589 639437
rect 675523 639372 675524 639436
rect 675588 639372 675589 639436
rect 675523 639371 675589 639372
rect 675339 637940 675405 637941
rect 675339 637876 675340 637940
rect 675404 637876 675405 637940
rect 675339 637875 675405 637876
rect 674971 637668 675037 637669
rect 674971 637604 674972 637668
rect 675036 637604 675037 637668
rect 674971 637603 675037 637604
rect 674971 636036 675037 636037
rect 674971 635972 674972 636036
rect 675036 635972 675037 636036
rect 674971 635971 675037 635972
rect 674974 629509 675034 635971
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 675155 629780 675221 629781
rect 675155 629716 675156 629780
rect 675220 629716 675221 629780
rect 675155 629715 675221 629716
rect 674971 629508 675037 629509
rect 674971 629444 674972 629508
rect 675036 629444 675037 629508
rect 674971 629443 675037 629444
rect 674971 599996 675037 599997
rect 674971 599932 674972 599996
rect 675036 599932 675037 599996
rect 674971 599931 675037 599932
rect 674974 597570 675034 599931
rect 674790 597510 675034 597570
rect 674790 596869 674850 597510
rect 674787 596868 674853 596869
rect 674787 596804 674788 596868
rect 674852 596804 674853 596868
rect 674787 596803 674853 596804
rect 675158 592925 675218 629715
rect 675523 607884 675589 607885
rect 675523 607820 675524 607884
rect 675588 607820 675589 607884
rect 675523 607819 675589 607820
rect 675526 593197 675586 607819
rect 676078 594693 676138 631347
rect 676075 594692 676141 594693
rect 676075 594628 676076 594692
rect 676140 594628 676141 594692
rect 676075 594627 676141 594628
rect 675523 593196 675589 593197
rect 675523 593132 675524 593196
rect 675588 593132 675589 593196
rect 675523 593131 675589 593132
rect 675155 592924 675221 592925
rect 675155 592860 675156 592924
rect 675220 592860 675221 592924
rect 675155 592859 675221 592860
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675523 562732 675589 562733
rect 675523 562730 675524 562732
rect 675342 562670 675524 562730
rect 675342 546005 675402 562670
rect 675523 562668 675524 562670
rect 675588 562668 675589 562732
rect 675523 562667 675589 562668
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 675339 546004 675405 546005
rect 675339 545940 675340 546004
rect 675404 545940 675405 546004
rect 675339 545939 675405 545940
rect 675526 545461 675586 561171
rect 675891 550628 675957 550629
rect 675891 550564 675892 550628
rect 675956 550564 675957 550628
rect 675891 550563 675957 550564
rect 675894 547637 675954 550563
rect 675891 547636 675957 547637
rect 675891 547572 675892 547636
rect 675956 547572 675957 547636
rect 675891 547571 675957 547572
rect 676078 546821 676138 586195
rect 676814 572797 676874 644267
rect 676998 619173 677058 694043
rect 676995 619172 677061 619173
rect 676995 619108 676996 619172
rect 677060 619108 677061 619172
rect 676995 619107 677061 619108
rect 676995 594692 677061 594693
rect 676995 594628 676996 594692
rect 677060 594628 677061 594692
rect 676995 594627 677061 594628
rect 676998 576061 677058 594627
rect 676995 576060 677061 576061
rect 676995 575996 676996 576060
rect 677060 575996 677061 576060
rect 676995 575995 677061 575996
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 676259 557564 676325 557565
rect 676259 557500 676260 557564
rect 676324 557500 676325 557564
rect 676259 557499 676325 557500
rect 676262 547637 676322 557499
rect 676811 553892 676877 553893
rect 676811 553828 676812 553892
rect 676876 553828 676877 553892
rect 676811 553827 676877 553828
rect 676259 547636 676325 547637
rect 676259 547572 676260 547636
rect 676324 547572 676325 547636
rect 676259 547571 676325 547572
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 675523 545460 675589 545461
rect 675523 545396 675524 545460
rect 675588 545396 675589 545460
rect 675523 545395 675589 545396
rect 676814 503437 676874 553827
rect 676995 550356 677061 550357
rect 676995 550292 676996 550356
rect 677060 550292 677061 550356
rect 676995 550291 677061 550292
rect 676998 503709 677058 550291
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 503436 676877 503437
rect 676811 503372 676812 503436
rect 676876 503372 676877 503436
rect 676811 503371 676877 503372
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 675894 488610 675954 488819
rect 675894 488550 676874 488610
rect 674603 474876 674669 474877
rect 674603 474812 674604 474876
rect 674668 474812 674669 474876
rect 674603 474811 674669 474812
rect 675339 453932 675405 453933
rect 675339 453868 675340 453932
rect 675404 453868 675405 453932
rect 675339 453867 675405 453868
rect 675342 410549 675402 453867
rect 675339 410548 675405 410549
rect 675339 410484 675340 410548
rect 675404 410484 675405 410548
rect 675339 410483 675405 410484
rect 676814 401301 676874 488550
rect 676811 401300 676877 401301
rect 676811 401236 676812 401300
rect 676876 401236 676877 401300
rect 676811 401235 676877 401236
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 389060 675957 389061
rect 675891 388996 675892 389060
rect 675956 388996 675957 389060
rect 675891 388995 675957 388996
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 377908 674853 377909
rect 674787 377844 674788 377908
rect 674852 377844 674853 377908
rect 674787 377843 674853 377844
rect 674790 372605 674850 377843
rect 675894 373013 675954 388995
rect 676078 378045 676138 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676075 378044 676141 378045
rect 676075 377980 676076 378044
rect 676140 377980 676141 378044
rect 676075 377979 676141 377980
rect 676262 377365 676322 395115
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676446 380629 676506 394707
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 675891 373012 675957 373013
rect 675891 372948 675892 373012
rect 675956 372948 675957 373012
rect 675891 372947 675957 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 43851 354244 43917 354245
rect 43851 354180 43852 354244
rect 43916 354180 43917 354244
rect 43851 354179 43917 354180
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 44219 353836 44285 353837
rect 44219 353772 44220 353836
rect 44284 353772 44285 353836
rect 44219 353771 44285 353772
rect 44222 342685 44282 353771
rect 675339 353020 675405 353021
rect 675339 352956 675340 353020
rect 675404 352956 675405 353020
rect 675339 352955 675405 352956
rect 673867 348532 673933 348533
rect 673867 348468 673868 348532
rect 673932 348468 673933 348532
rect 673867 348467 673933 348468
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 342684 44285 342685
rect 44219 342620 44220 342684
rect 44284 342620 44285 342684
rect 44219 342619 44285 342620
rect 44406 342410 44466 342891
rect 44222 342350 44466 342410
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 41459 338196 41525 338197
rect 41459 338132 41460 338196
rect 41524 338132 41525 338196
rect 41459 338131 41525 338132
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316709 40602 336907
rect 40723 335340 40789 335341
rect 40723 335276 40724 335340
rect 40788 335276 40789 335340
rect 40723 335275 40789 335276
rect 40726 317525 40786 335275
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40910 325413 40970 333643
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41462 319973 41522 338131
rect 41827 337788 41893 337789
rect 41827 337724 41828 337788
rect 41892 337724 41893 337788
rect 41827 337723 41893 337724
rect 41643 336564 41709 336565
rect 41643 336500 41644 336564
rect 41708 336500 41709 336564
rect 41643 336499 41709 336500
rect 41646 325710 41706 336499
rect 41830 326773 41890 337723
rect 42931 337380 42997 337381
rect 42931 337316 42932 337380
rect 42996 337316 42997 337380
rect 42931 337315 42997 337316
rect 42747 335748 42813 335749
rect 42747 335684 42748 335748
rect 42812 335684 42813 335748
rect 42747 335683 42813 335684
rect 42750 334389 42810 335683
rect 42747 334388 42813 334389
rect 42747 334324 42748 334388
rect 42812 334324 42813 334388
rect 42747 334323 42813 334324
rect 41827 326772 41893 326773
rect 41827 326708 41828 326772
rect 41892 326708 41893 326772
rect 41827 326707 41893 326708
rect 41646 325650 41890 325710
rect 41830 324869 41890 325650
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41459 319972 41525 319973
rect 41459 319908 41460 319972
rect 41524 319908 41525 319972
rect 41459 319907 41525 319908
rect 40723 317524 40789 317525
rect 40723 317460 40724 317524
rect 40788 317460 40789 317524
rect 40723 317459 40789 317460
rect 40539 316708 40605 316709
rect 40539 316644 40540 316708
rect 40604 316644 40605 316708
rect 40539 316643 40605 316644
rect 42934 312765 42994 337315
rect 43115 336972 43181 336973
rect 43115 336908 43116 336972
rect 43180 336908 43181 336972
rect 43115 336907 43181 336908
rect 43118 316029 43178 336907
rect 43115 316028 43181 316029
rect 43115 315964 43116 316028
rect 43180 315964 43181 316028
rect 43115 315963 43181 315964
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 43670 297669 43730 340443
rect 44222 311541 44282 342350
rect 44403 342140 44469 342141
rect 44403 342076 44404 342140
rect 44468 342076 44469 342140
rect 44403 342075 44469 342076
rect 44219 311540 44285 311541
rect 44219 311476 44220 311540
rect 44284 311476 44285 311540
rect 44219 311475 44285 311476
rect 44406 311269 44466 342075
rect 44403 311268 44469 311269
rect 44403 311204 44404 311268
rect 44468 311204 44469 311268
rect 44403 311203 44469 311204
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 294130 41890 295563
rect 40726 294070 41890 294130
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 40726 277677 40786 294070
rect 41827 292772 41893 292773
rect 41827 292770 41828 292772
rect 41784 292708 41828 292770
rect 41892 292708 41893 292772
rect 41784 292707 41893 292708
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 41784 292590 41844 292707
rect 40907 292527 40973 292528
rect 41462 292530 41844 292590
rect 40910 277949 40970 292527
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40723 277676 40789 277677
rect 40723 277612 40724 277676
rect 40788 277612 40789 277676
rect 40723 277611 40789 277612
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 292530
rect 41827 292364 41893 292365
rect 41827 292300 41828 292364
rect 41892 292300 41893 292364
rect 41827 292299 41893 292300
rect 41830 289830 41890 292299
rect 41646 289770 41890 289830
rect 41646 287070 41706 289770
rect 41646 287010 41890 287070
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 287010
rect 42014 281485 42074 296379
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 673870 278629 673930 348467
rect 675342 337245 675402 352955
rect 675526 340890 675586 354179
rect 675707 353836 675773 353837
rect 675707 353772 675708 353836
rect 675772 353772 675773 353836
rect 675707 353771 675773 353772
rect 675710 346490 675770 353771
rect 675894 351190 676506 351250
rect 675894 350981 675954 351190
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675894 350490 676322 350550
rect 675894 350301 675954 350490
rect 675891 350300 675957 350301
rect 675891 350236 675892 350300
rect 675956 350236 675957 350300
rect 675891 350235 675957 350236
rect 675710 346430 676092 346490
rect 676032 346410 676092 346430
rect 676032 346350 676138 346410
rect 675526 340830 675954 340890
rect 675894 339421 675954 340830
rect 675891 339420 675957 339421
rect 675891 339356 675892 339420
rect 675956 339356 675957 339420
rect 675891 339355 675957 339356
rect 675339 337244 675405 337245
rect 675339 337180 675340 337244
rect 675404 337180 675405 337244
rect 675339 337179 675405 337180
rect 674787 335884 674853 335885
rect 674787 335820 674788 335884
rect 674852 335820 674853 335884
rect 674787 335819 674853 335820
rect 674790 326909 674850 335819
rect 676078 328405 676138 346350
rect 676262 340373 676322 350490
rect 676259 340372 676325 340373
rect 676259 340308 676260 340372
rect 676324 340308 676325 340372
rect 676259 340307 676325 340308
rect 676446 336565 676506 351190
rect 676627 346628 676693 346629
rect 676627 346564 676628 346628
rect 676692 346564 676693 346628
rect 676627 346563 676693 346564
rect 676443 336564 676509 336565
rect 676443 336500 676444 336564
rect 676508 336500 676509 336564
rect 676443 336499 676509 336500
rect 676630 332349 676690 346563
rect 676627 332348 676693 332349
rect 676627 332284 676628 332348
rect 676692 332284 676693 332348
rect 676627 332283 676693 332284
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 674787 326908 674853 326909
rect 674787 326844 674788 326908
rect 674852 326844 674853 326908
rect 674787 326843 674853 326844
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 302250 675770 308755
rect 675891 306780 675957 306781
rect 675891 306716 675892 306780
rect 675956 306716 675957 306780
rect 675891 306715 675957 306716
rect 675894 306370 675954 306715
rect 675894 306310 676874 306370
rect 675891 305964 675957 305965
rect 675891 305900 675892 305964
rect 675956 305900 675957 305964
rect 675891 305899 675957 305900
rect 675894 305690 675954 305899
rect 675894 305630 676506 305690
rect 676029 305148 676095 305149
rect 676029 305084 676030 305148
rect 676094 305146 676095 305148
rect 676094 305084 676138 305146
rect 676029 305083 676138 305084
rect 676078 305010 676138 305083
rect 676078 304950 676322 305010
rect 675710 302190 676138 302250
rect 675707 299436 675773 299437
rect 675707 299372 675708 299436
rect 675772 299372 675773 299436
rect 675707 299371 675773 299372
rect 675339 296852 675405 296853
rect 675339 296788 675340 296852
rect 675404 296788 675405 296852
rect 675339 296787 675405 296788
rect 675342 289917 675402 296787
rect 675523 296580 675589 296581
rect 675523 296516 675524 296580
rect 675588 296516 675589 296580
rect 675523 296515 675589 296516
rect 675526 292093 675586 296515
rect 675523 292092 675589 292093
rect 675523 292028 675524 292092
rect 675588 292028 675589 292092
rect 675523 292027 675589 292028
rect 675339 289916 675405 289917
rect 675339 289852 675340 289916
rect 675404 289852 675405 289916
rect 675339 289851 675405 289852
rect 675710 282845 675770 299371
rect 675891 297396 675957 297397
rect 675891 297332 675892 297396
rect 675956 297332 675957 297396
rect 675891 297331 675957 297332
rect 675707 282844 675773 282845
rect 675707 282780 675708 282844
rect 675772 282780 675773 282844
rect 675707 282779 675773 282780
rect 675894 281213 675954 297331
rect 676078 283661 676138 302190
rect 676262 287061 676322 304950
rect 676446 291549 676506 305630
rect 676814 295221 676874 306310
rect 676811 295220 676877 295221
rect 676811 295156 676812 295220
rect 676876 295156 676877 295220
rect 676811 295155 676877 295156
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 281212 675957 281213
rect 675891 281148 675892 281212
rect 675956 281148 675957 281212
rect 675891 281147 675957 281148
rect 673867 278628 673933 278629
rect 673867 278564 673868 278628
rect 673932 278564 673933 278628
rect 673867 278563 673933 278564
rect 673867 277676 673933 277677
rect 673867 277612 673868 277676
rect 673932 277612 673933 277676
rect 673867 277611 673933 277612
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 40539 251428 40605 251429
rect 40539 251364 40540 251428
rect 40604 251364 40605 251428
rect 40539 251363 40605 251364
rect 40542 240141 40602 251363
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 40539 240140 40605 240141
rect 40539 240076 40540 240140
rect 40604 240076 40605 240140
rect 40539 240075 40605 240076
rect 40726 235925 40786 249731
rect 673870 249661 673930 277611
rect 674971 263668 675037 263669
rect 674971 263604 674972 263668
rect 675036 263604 675037 263668
rect 674971 263603 675037 263604
rect 674974 258090 675034 263603
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 674790 258030 675034 258090
rect 674790 249661 674850 258030
rect 676078 249661 676138 262379
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 673867 249660 673933 249661
rect 673867 249596 673868 249660
rect 673932 249596 673933 249660
rect 673867 249595 673933 249596
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 674603 246260 674669 246261
rect 674603 246196 674604 246260
rect 674668 246196 674669 246260
rect 674603 246195 674669 246196
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 673683 237420 673749 237421
rect 673683 237356 673684 237420
rect 673748 237356 673749 237420
rect 673683 237355 673749 237356
rect 40723 235924 40789 235925
rect 40723 235860 40724 235924
rect 40788 235860 40789 235924
rect 40723 235859 40789 235860
rect 42014 227357 42074 237355
rect 671291 234564 671357 234565
rect 671291 234500 671292 234564
rect 671356 234500 671357 234564
rect 671291 234499 671357 234500
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 670739 225452 670805 225453
rect 670739 225388 670740 225452
rect 670804 225388 670805 225452
rect 670739 225387 670805 225388
rect 670742 223957 670802 225387
rect 670739 223956 670805 223957
rect 670739 223892 670740 223956
rect 670804 223892 670805 223956
rect 670739 223891 670805 223892
rect 562366 219950 563530 220010
rect 518939 219740 519005 219741
rect 518939 219676 518940 219740
rect 519004 219676 519005 219740
rect 518939 219675 519005 219676
rect 528875 219740 528941 219741
rect 528875 219676 528876 219740
rect 528940 219676 528941 219740
rect 528875 219675 528941 219676
rect 499435 218924 499501 218925
rect 499435 218860 499436 218924
rect 499500 218860 499501 218924
rect 499435 218859 499501 218860
rect 496675 218652 496741 218653
rect 496675 218588 496676 218652
rect 496740 218650 496741 218652
rect 499438 218650 499498 218859
rect 496740 218590 499498 218650
rect 496740 218588 496741 218590
rect 496675 218587 496741 218588
rect 501091 217564 501157 217565
rect 501091 217500 501092 217564
rect 501156 217500 501157 217564
rect 501091 217499 501157 217500
rect 503299 217564 503365 217565
rect 503299 217500 503300 217564
rect 503364 217500 503365 217564
rect 503299 217499 503365 217500
rect 503667 217564 503733 217565
rect 503667 217500 503668 217564
rect 503732 217500 503733 217564
rect 503667 217499 503733 217500
rect 506059 217564 506125 217565
rect 506059 217500 506060 217564
rect 506124 217500 506125 217564
rect 506059 217499 506125 217500
rect 509187 217564 509253 217565
rect 509187 217500 509188 217564
rect 509252 217500 509253 217564
rect 509187 217499 509253 217500
rect 501094 215933 501154 217499
rect 503302 217021 503362 217499
rect 503299 217020 503365 217021
rect 503299 216956 503300 217020
rect 503364 216956 503365 217020
rect 503299 216955 503365 216956
rect 503670 216205 503730 217499
rect 503667 216204 503733 216205
rect 503667 216140 503668 216204
rect 503732 216140 503733 216204
rect 503667 216139 503733 216140
rect 501091 215932 501157 215933
rect 501091 215868 501092 215932
rect 501156 215868 501157 215932
rect 501091 215867 501157 215868
rect 506062 215389 506122 217499
rect 509190 215661 509250 217499
rect 518942 216477 519002 219675
rect 528878 216477 528938 219675
rect 562366 219469 562426 219950
rect 563470 219469 563530 219950
rect 571934 219950 572914 220010
rect 571934 219469 571994 219950
rect 562363 219468 562429 219469
rect 562363 219404 562364 219468
rect 562428 219404 562429 219468
rect 562363 219403 562429 219404
rect 563467 219468 563533 219469
rect 563467 219404 563468 219468
rect 563532 219404 563533 219468
rect 563467 219403 563533 219404
rect 571931 219468 571997 219469
rect 571931 219404 571932 219468
rect 571996 219404 571997 219468
rect 571931 219403 571997 219404
rect 572854 219197 572914 219950
rect 572851 219196 572917 219197
rect 572851 219132 572852 219196
rect 572916 219132 572917 219196
rect 572851 219131 572917 219132
rect 572483 218924 572549 218925
rect 572483 218860 572484 218924
rect 572548 218860 572549 218924
rect 572483 218859 572549 218860
rect 572486 217290 572546 218859
rect 666323 218652 666389 218653
rect 666323 218588 666324 218652
rect 666388 218588 666389 218652
rect 666323 218587 666389 218588
rect 573219 218108 573285 218109
rect 573219 218044 573220 218108
rect 573284 218044 573285 218108
rect 573219 218043 573285 218044
rect 573222 217290 573282 218043
rect 592171 217836 592237 217837
rect 592171 217772 592172 217836
rect 592236 217772 592237 217836
rect 592171 217771 592237 217772
rect 572486 217230 573282 217290
rect 591803 217292 591869 217293
rect 591803 217228 591804 217292
rect 591868 217290 591869 217292
rect 592174 217290 592234 217771
rect 591868 217230 592234 217290
rect 591868 217228 591869 217230
rect 591803 217227 591869 217228
rect 586651 217020 586717 217021
rect 586651 216956 586652 217020
rect 586716 216956 586717 217020
rect 586651 216955 586717 216956
rect 518939 216476 519005 216477
rect 518939 216412 518940 216476
rect 519004 216412 519005 216476
rect 518939 216411 519005 216412
rect 528691 216476 528757 216477
rect 528691 216412 528692 216476
rect 528756 216412 528757 216476
rect 528691 216411 528757 216412
rect 528875 216476 528941 216477
rect 528875 216412 528876 216476
rect 528940 216412 528941 216476
rect 528875 216411 528941 216412
rect 509187 215660 509253 215661
rect 509187 215596 509188 215660
rect 509252 215596 509253 215660
rect 509187 215595 509253 215596
rect 506059 215388 506125 215389
rect 506059 215324 506060 215388
rect 506124 215324 506125 215388
rect 506059 215323 506125 215324
rect 528694 215117 528754 216411
rect 586654 215117 586714 216955
rect 528691 215116 528757 215117
rect 528691 215052 528692 215116
rect 528756 215052 528757 215116
rect 528691 215051 528757 215052
rect 586651 215116 586717 215117
rect 586651 215052 586652 215116
rect 586716 215052 586717 215116
rect 586651 215051 586717 215052
rect 41459 208996 41525 208997
rect 41459 208932 41460 208996
rect 41524 208932 41525 208996
rect 41459 208931 41525 208932
rect 40539 208180 40605 208181
rect 40539 208116 40540 208180
rect 40604 208116 40605 208180
rect 40539 208115 40605 208116
rect 40542 197165 40602 208115
rect 40907 207364 40973 207365
rect 40907 207300 40908 207364
rect 40972 207300 40973 207364
rect 40907 207299 40973 207300
rect 40723 206956 40789 206957
rect 40723 206892 40724 206956
rect 40788 206892 40789 206956
rect 40723 206891 40789 206892
rect 40539 197164 40605 197165
rect 40539 197100 40540 197164
rect 40604 197100 40605 197164
rect 40539 197099 40605 197100
rect 40726 194170 40786 206891
rect 40910 195397 40970 207299
rect 41462 205650 41522 208931
rect 42011 205732 42077 205733
rect 42011 205668 42012 205732
rect 42076 205668 42077 205732
rect 42011 205667 42077 205668
rect 41462 205590 41706 205650
rect 40907 195396 40973 195397
rect 40907 195332 40908 195396
rect 40972 195332 40973 195396
rect 40907 195331 40973 195332
rect 41646 194850 41706 205590
rect 41827 202196 41893 202197
rect 41827 202132 41828 202196
rect 41892 202132 41893 202196
rect 41827 202131 41893 202132
rect 41830 195805 41890 202131
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 42014 195125 42074 205667
rect 666326 205650 666386 218587
rect 667979 215660 668045 215661
rect 667979 215596 667980 215660
rect 668044 215596 668045 215660
rect 667979 215595 668045 215596
rect 669451 215660 669517 215661
rect 669451 215596 669452 215660
rect 669516 215596 669517 215660
rect 669451 215595 669517 215596
rect 666326 205590 666570 205650
rect 42011 195124 42077 195125
rect 42011 195060 42012 195124
rect 42076 195060 42077 195124
rect 42011 195059 42077 195060
rect 41646 194790 42258 194850
rect 40726 194110 41522 194170
rect 41462 187237 41522 194110
rect 42011 193220 42077 193221
rect 42011 193156 42012 193220
rect 42076 193156 42077 193220
rect 42011 193155 42077 193156
rect 41459 187236 41525 187237
rect 41459 187172 41460 187236
rect 41524 187172 41525 187236
rect 41459 187171 41525 187172
rect 42014 186421 42074 193155
rect 42011 186420 42077 186421
rect 42011 186356 42012 186420
rect 42076 186356 42077 186420
rect 42011 186355 42077 186356
rect 42198 185877 42258 194790
rect 666510 189821 666570 205590
rect 666507 189820 666573 189821
rect 666507 189756 666508 189820
rect 666572 189756 666573 189820
rect 666507 189755 666573 189756
rect 42195 185876 42261 185877
rect 42195 185812 42196 185876
rect 42260 185812 42261 185876
rect 42195 185811 42261 185812
rect 667982 130661 668042 215595
rect 669454 214573 669514 215595
rect 669451 214572 669517 214573
rect 669451 214508 669452 214572
rect 669516 214508 669517 214572
rect 669451 214507 669517 214508
rect 669451 214028 669517 214029
rect 669451 213964 669452 214028
rect 669516 213964 669517 214028
rect 669451 213963 669517 213964
rect 669267 205732 669333 205733
rect 669267 205668 669268 205732
rect 669332 205668 669333 205732
rect 669267 205667 669333 205668
rect 669270 205461 669330 205667
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 669267 196076 669333 196077
rect 669267 196074 669268 196076
rect 669086 196014 669268 196074
rect 669086 186330 669146 196014
rect 669267 196012 669268 196014
rect 669332 196012 669333 196076
rect 669267 196011 669333 196012
rect 669454 186330 669514 213963
rect 669635 211172 669701 211173
rect 669635 211108 669636 211172
rect 669700 211108 669701 211172
rect 669635 211107 669701 211108
rect 669638 205733 669698 211107
rect 669635 205732 669701 205733
rect 669635 205668 669636 205732
rect 669700 205668 669701 205732
rect 669635 205667 669701 205668
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669638 196077 669698 205395
rect 669635 196076 669701 196077
rect 669635 196012 669636 196076
rect 669700 196012 669701 196076
rect 669635 196011 669701 196012
rect 669086 186270 669330 186330
rect 669454 186270 669698 186330
rect 669270 186010 669330 186270
rect 669270 185950 669514 186010
rect 669454 176670 669514 185950
rect 669270 176610 669514 176670
rect 669270 176490 669330 176610
rect 669270 176430 669514 176490
rect 669454 157350 669514 176430
rect 669638 167109 669698 186270
rect 669635 167108 669701 167109
rect 669635 167044 669636 167108
rect 669700 167044 669701 167108
rect 669635 167043 669701 167044
rect 669270 157290 669514 157350
rect 669270 138030 669330 157290
rect 671294 145349 671354 234499
rect 673686 232525 673746 237355
rect 673683 232524 673749 232525
rect 673683 232460 673684 232524
rect 673748 232460 673749 232524
rect 673683 232459 673749 232460
rect 673683 231844 673749 231845
rect 673683 231780 673684 231844
rect 673748 231780 673749 231844
rect 673683 231779 673749 231780
rect 673315 231572 673381 231573
rect 673315 231508 673316 231572
rect 673380 231508 673381 231572
rect 673315 231507 673381 231508
rect 671475 230076 671541 230077
rect 671475 230012 671476 230076
rect 671540 230012 671541 230076
rect 671475 230011 671541 230012
rect 671478 224090 671538 230011
rect 672947 226812 673013 226813
rect 672947 226748 672948 226812
rect 673012 226748 673013 226812
rect 672947 226747 673013 226748
rect 673131 226812 673197 226813
rect 673131 226748 673132 226812
rect 673196 226748 673197 226812
rect 673131 226747 673197 226748
rect 672950 225861 673010 226747
rect 671659 225860 671725 225861
rect 671659 225796 671660 225860
rect 671724 225796 671725 225860
rect 671659 225795 671725 225796
rect 672947 225860 673013 225861
rect 672947 225796 672948 225860
rect 673012 225796 673013 225860
rect 672947 225795 673013 225796
rect 671662 224365 671722 225795
rect 672763 225724 672829 225725
rect 672763 225660 672764 225724
rect 672828 225660 672829 225724
rect 672763 225659 672829 225660
rect 671659 224364 671725 224365
rect 671659 224300 671660 224364
rect 671724 224300 671725 224364
rect 671659 224299 671725 224300
rect 671659 224092 671725 224093
rect 671659 224090 671660 224092
rect 671478 224030 671660 224090
rect 671659 224028 671660 224030
rect 671724 224028 671725 224092
rect 671659 224027 671725 224028
rect 672766 223957 672826 225659
rect 673134 224093 673194 226747
rect 673131 224092 673197 224093
rect 673131 224028 673132 224092
rect 673196 224028 673197 224092
rect 673131 224027 673197 224028
rect 672763 223956 672829 223957
rect 672763 223892 672764 223956
rect 672828 223892 672829 223956
rect 672763 223891 672829 223892
rect 673318 222210 673378 231507
rect 673499 230076 673565 230077
rect 673499 230012 673500 230076
rect 673564 230012 673565 230076
rect 673499 230011 673565 230012
rect 672950 222150 673378 222210
rect 672395 221916 672461 221917
rect 672395 221852 672396 221916
rect 672460 221852 672461 221916
rect 672395 221851 672461 221852
rect 672398 220830 672458 221851
rect 672398 220770 672642 220830
rect 672582 214029 672642 220770
rect 672579 214028 672645 214029
rect 672579 213964 672580 214028
rect 672644 213964 672645 214028
rect 672579 213963 672645 213964
rect 672950 183565 673010 222150
rect 673131 220964 673197 220965
rect 673131 220900 673132 220964
rect 673196 220900 673197 220964
rect 673131 220899 673197 220900
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 671291 145348 671357 145349
rect 671291 145284 671292 145348
rect 671356 145284 671357 145348
rect 671291 145283 671357 145284
rect 669270 137970 669514 138030
rect 669454 137461 669514 137970
rect 669451 137460 669517 137461
rect 669451 137396 669452 137460
rect 669516 137396 669517 137460
rect 669451 137395 669517 137396
rect 673134 133925 673194 220899
rect 673131 133924 673197 133925
rect 673131 133860 673132 133924
rect 673196 133860 673197 133924
rect 673131 133859 673197 133860
rect 667979 130660 668045 130661
rect 667979 130596 667980 130660
rect 668044 130596 668045 130660
rect 667979 130595 668045 130596
rect 673502 128485 673562 230011
rect 673686 142221 673746 231779
rect 674235 229532 674301 229533
rect 674235 229468 674236 229532
rect 674300 229468 674301 229532
rect 674235 229467 674301 229468
rect 673867 225588 673933 225589
rect 673867 225524 673868 225588
rect 673932 225524 673933 225588
rect 673867 225523 673933 225524
rect 673870 222210 673930 225523
rect 674238 222869 674298 229467
rect 674606 223821 674666 246195
rect 676814 245581 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 245580 676877 245581
rect 676811 245516 676812 245580
rect 676876 245516 676877 245580
rect 676811 245515 676877 245516
rect 675339 245308 675405 245309
rect 675339 245244 675340 245308
rect 675404 245244 675405 245308
rect 675339 245243 675405 245244
rect 675155 245036 675221 245037
rect 675155 244972 675156 245036
rect 675220 244972 675221 245036
rect 675155 244971 675221 244972
rect 675158 237285 675218 244971
rect 675342 240277 675402 245243
rect 675339 240276 675405 240277
rect 675339 240212 675340 240276
rect 675404 240212 675405 240276
rect 675339 240211 675405 240212
rect 675155 237284 675221 237285
rect 675155 237220 675156 237284
rect 675220 237220 675221 237284
rect 675155 237219 675221 237220
rect 676811 235108 676877 235109
rect 676811 235044 676812 235108
rect 676876 235044 676877 235108
rect 676811 235043 676877 235044
rect 674971 228852 675037 228853
rect 674971 228788 674972 228852
rect 675036 228788 675037 228852
rect 674971 228787 675037 228788
rect 674787 228580 674853 228581
rect 674787 228516 674788 228580
rect 674852 228516 674853 228580
rect 674787 228515 674853 228516
rect 674603 223820 674669 223821
rect 674603 223756 674604 223820
rect 674668 223756 674669 223820
rect 674603 223755 674669 223756
rect 674235 222868 674301 222869
rect 674235 222804 674236 222868
rect 674300 222804 674301 222868
rect 674235 222803 674301 222804
rect 673870 222150 674114 222210
rect 674054 220149 674114 222150
rect 674790 220965 674850 228515
rect 674787 220964 674853 220965
rect 674787 220900 674788 220964
rect 674852 220900 674853 220964
rect 674787 220899 674853 220900
rect 674051 220148 674117 220149
rect 674051 220084 674052 220148
rect 674116 220084 674117 220148
rect 674051 220083 674117 220084
rect 674974 217970 675034 228787
rect 676814 224970 676874 235043
rect 676262 224910 676874 224970
rect 675891 222732 675957 222733
rect 675891 222668 675892 222732
rect 675956 222730 675957 222732
rect 676262 222730 676322 224910
rect 675956 222670 676322 222730
rect 675956 222668 675957 222670
rect 675891 222667 675957 222668
rect 675523 219060 675589 219061
rect 675523 218996 675524 219060
rect 675588 218996 675589 219060
rect 675523 218995 675589 218996
rect 674606 217910 675034 217970
rect 674606 217701 674666 217910
rect 674603 217700 674669 217701
rect 674603 217636 674604 217700
rect 674668 217636 674669 217700
rect 674603 217635 674669 217636
rect 674051 212124 674117 212125
rect 674051 212060 674052 212124
rect 674116 212060 674117 212124
rect 674051 212059 674117 212060
rect 673683 142220 673749 142221
rect 673683 142156 673684 142220
rect 673748 142156 673749 142220
rect 673683 142155 673749 142156
rect 673499 128484 673565 128485
rect 673499 128420 673500 128484
rect 673564 128420 673565 128484
rect 673499 128419 673565 128420
rect 674054 128213 674114 212059
rect 675526 204237 675586 218995
rect 676029 218244 676095 218245
rect 676029 218180 676030 218244
rect 676094 218180 676095 218244
rect 676029 218179 676095 218180
rect 676032 217970 676092 218179
rect 676032 217910 676506 217970
rect 675891 217020 675957 217021
rect 675891 216956 675892 217020
rect 675956 216956 675957 217020
rect 675891 216955 675957 216956
rect 675707 215388 675773 215389
rect 675707 215324 675708 215388
rect 675772 215324 675773 215388
rect 675707 215323 675773 215324
rect 675710 205650 675770 215323
rect 675894 210490 675954 216955
rect 676259 215150 676325 215151
rect 676259 215086 676260 215150
rect 676324 215086 676325 215150
rect 676259 215085 676325 215086
rect 675894 210430 676138 210490
rect 675710 205590 675954 205650
rect 675523 204236 675589 204237
rect 675523 204172 675524 204236
rect 675588 204172 675589 204236
rect 675523 204171 675589 204172
rect 675894 195261 675954 205590
rect 675891 195260 675957 195261
rect 675891 195196 675892 195260
rect 675956 195196 675957 195260
rect 675891 195195 675957 195196
rect 676078 191589 676138 210430
rect 676262 197165 676322 215085
rect 676446 205597 676506 217910
rect 676995 211172 677061 211173
rect 676995 211170 676996 211172
rect 676814 211110 676996 211170
rect 676443 205596 676509 205597
rect 676443 205532 676444 205596
rect 676508 205532 676509 205596
rect 676443 205531 676509 205532
rect 676814 200701 676874 211110
rect 676995 211108 676996 211110
rect 677060 211108 677061 211172
rect 676995 211107 677061 211108
rect 676811 200700 676877 200701
rect 676811 200636 676812 200700
rect 676876 200636 676877 200700
rect 676811 200635 676877 200636
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675710 171050 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675710 170990 676138 171050
rect 675707 170372 675773 170373
rect 675707 170308 675708 170372
rect 675772 170308 675773 170372
rect 675707 170307 675773 170308
rect 675710 150381 675770 170307
rect 675891 167516 675957 167517
rect 675891 167452 675892 167516
rect 675956 167452 675957 167516
rect 675891 167451 675957 167452
rect 675707 150380 675773 150381
rect 675707 150316 675708 150380
rect 675772 150316 675773 150380
rect 675707 150315 675773 150316
rect 675894 147661 675954 167451
rect 676078 148477 676138 170990
rect 676262 151605 676322 172350
rect 676446 159357 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159356 676509 159357
rect 676443 159292 676444 159356
rect 676508 159292 676509 159356
rect 676443 159291 676509 159292
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 151604 676325 151605
rect 676259 151540 676260 151604
rect 676324 151540 676325 151604
rect 676259 151539 676325 151540
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675891 147660 675957 147661
rect 675891 147596 675892 147660
rect 675956 147596 675957 147660
rect 675891 147595 675957 147596
rect 676627 128620 676693 128621
rect 676627 128556 676628 128620
rect 676692 128556 676693 128620
rect 676627 128555 676693 128556
rect 674051 128212 674117 128213
rect 674051 128148 674052 128212
rect 674116 128148 674117 128212
rect 674051 128147 674117 128148
rect 676443 126580 676509 126581
rect 676443 126516 676444 126580
rect 676508 126516 676509 126580
rect 676443 126515 676509 126516
rect 675891 124948 675957 124949
rect 675891 124884 675892 124948
rect 675956 124884 675957 124948
rect 675891 124883 675957 124884
rect 672947 122772 673013 122773
rect 672947 122708 672948 122772
rect 673012 122708 673013 122772
rect 672947 122707 673013 122708
rect 672950 122229 673010 122707
rect 672947 122228 673013 122229
rect 672947 122164 672948 122228
rect 673012 122164 673013 122228
rect 672947 122163 673013 122164
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 103189 675770 117267
rect 675894 108085 675954 124883
rect 676446 122850 676506 126515
rect 676262 122790 676506 122850
rect 676075 122092 676141 122093
rect 676075 122028 676076 122092
rect 676140 122028 676141 122092
rect 676075 122027 676141 122028
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 675707 103188 675773 103189
rect 675707 103124 675708 103188
rect 675772 103124 675773 103188
rect 675707 103123 675773 103124
rect 676078 102509 676138 122027
rect 676075 102508 676141 102509
rect 676075 102444 676076 102508
rect 676140 102444 676141 102508
rect 676075 102443 676141 102444
rect 676262 101421 676322 122790
rect 676443 118012 676509 118013
rect 676443 117948 676444 118012
rect 676508 117948 676509 118012
rect 676443 117947 676509 117948
rect 676446 109037 676506 117947
rect 676630 113117 676690 128555
rect 676811 124540 676877 124541
rect 676811 124476 676812 124540
rect 676876 124476 676877 124540
rect 676811 124475 676877 124476
rect 676814 118013 676874 124475
rect 676811 118012 676877 118013
rect 676811 117948 676812 118012
rect 676876 117948 676877 118012
rect 676811 117947 676877 117948
rect 676627 113116 676693 113117
rect 676627 113052 676628 113116
rect 676692 113052 676693 113116
rect 676627 113051 676693 113052
rect 676443 109036 676509 109037
rect 676443 108972 676444 109036
rect 676508 108972 676509 109036
rect 676443 108971 676509 108972
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 634675 96116 634741 96117
rect 634675 96052 634676 96116
rect 634740 96052 634741 96116
rect 634675 96051 634741 96052
rect 634678 77621 634738 96051
rect 637254 84210 637314 96867
rect 647187 96116 647253 96117
rect 647187 96052 647188 96116
rect 647252 96052 647253 96116
rect 647187 96051 647253 96052
rect 647190 94298 647250 96051
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 637070 77893 637130 84150
rect 637067 77892 637133 77893
rect 637067 77828 637068 77892
rect 637132 77828 637133 77892
rect 637067 77827 637133 77828
rect 634675 77620 634741 77621
rect 634675 77556 634676 77620
rect 634740 77556 634741 77620
rect 634675 77555 634741 77556
rect 462635 54772 462701 54773
rect 462635 54708 462636 54772
rect 462700 54708 462701 54772
rect 462635 54707 462701 54708
rect 462638 53685 462698 54707
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 194363 48924 194429 48925
rect 194363 48860 194364 48924
rect 194428 48860 194429 48924
rect 194363 48859 194429 48860
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40493 141802 43963
rect 194366 42125 194426 48859
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 463739 44436 463805 44437
rect 463739 44372 463740 44436
rect 463804 44372 463805 44436
rect 463739 44371 463805 44372
rect 440187 43892 440253 43893
rect 440187 43828 440188 43892
rect 440252 43890 440253 43892
rect 440923 43892 440989 43893
rect 440923 43890 440924 43892
rect 440252 43830 440924 43890
rect 440252 43828 440253 43830
rect 440187 43827 440253 43828
rect 440923 43828 440924 43830
rect 440988 43828 440989 43892
rect 440923 43827 440989 43828
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 463742 41938 463802 44371
rect 464107 44300 464173 44301
rect 464107 44236 464108 44300
rect 464172 44236 464173 44300
rect 464107 44235 464173 44236
rect 365483 41852 365549 41853
rect 365483 41788 365484 41852
rect 365548 41788 365549 41852
rect 403019 41852 403085 41853
rect 403019 41850 403020 41852
rect 365483 41787 365549 41788
rect 402286 41790 403020 41850
rect 365486 41258 365546 41787
rect 402286 41258 402346 41790
rect 403019 41788 403020 41790
rect 403084 41788 403085 41852
rect 403019 41787 403085 41788
rect 421971 41852 422037 41853
rect 421971 41788 421972 41852
rect 422036 41850 422037 41852
rect 422036 41790 422162 41850
rect 422036 41788 422037 41790
rect 421971 41787 422037 41788
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 464110 41853 464170 44235
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 464107 41852 464173 41853
rect 464107 41788 464108 41852
rect 464172 41788 464173 41852
rect 464107 41787 464173 41788
rect 425102 40578 425162 41702
rect 141739 40492 141805 40493
rect 141739 40428 141740 40492
rect 141804 40428 141805 40492
rect 141739 40427 141805 40428
<< via4 >>
rect 172566 997102 172802 997338
rect 245614 997252 245850 997338
rect 245614 997188 245700 997252
rect 245700 997188 245764 997252
rect 245764 997188 245850 997252
rect 245614 997102 245850 997188
rect 246350 997102 246586 997338
rect 278550 997102 278786 997338
rect 524006 997102 524242 997338
rect 532102 997102 532338 997338
rect 557126 997102 557362 997338
rect 634406 997102 634642 997338
rect 537990 993022 538226 993258
rect 572582 993022 572818 993258
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 361902 41852 362138 41938
rect 361902 41788 361988 41852
rect 361988 41788 362052 41852
rect 362052 41788 362138 41852
rect 361902 41702 362138 41788
rect 422162 41702 422398 41938
rect 425014 41702 425250 41938
rect 441390 41702 441626 41938
rect 463654 41702 463890 41938
rect 365398 41022 365634 41258
rect 402198 41022 402434 41258
rect 425014 40342 425250 40578
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 172524 997338 245892 997380
rect 172524 997102 172566 997338
rect 172802 997102 245614 997338
rect 245850 997102 245892 997338
rect 172524 997060 245892 997102
rect 246308 997338 278828 997380
rect 246308 997102 246350 997338
rect 246586 997102 278550 997338
rect 278786 997102 278828 997338
rect 246308 997060 278828 997102
rect 523964 997338 532380 997380
rect 523964 997102 524006 997338
rect 524242 997102 532102 997338
rect 532338 997102 532380 997338
rect 523964 997060 532380 997102
rect 557084 997338 634684 997380
rect 557084 997102 557126 997338
rect 557362 997102 634406 997338
rect 634642 997102 634684 997338
rect 557084 997060 634684 997102
rect 537948 993258 572860 993300
rect 537948 993022 537990 993258
rect 538226 993022 572582 993258
rect 572818 993022 572860 993258
rect 537948 992980 572860 993022
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 361860 41938 403120 41980
rect 361860 41702 361902 41938
rect 362138 41702 403120 41938
rect 361860 41660 403120 41702
rect 402800 41300 403120 41660
rect 403444 41660 412044 41980
rect 403444 41300 403764 41660
rect 365356 41258 402476 41300
rect 365356 41022 365398 41258
rect 365634 41022 402198 41258
rect 402434 41022 402476 41258
rect 365356 40980 402476 41022
rect 402800 40980 403764 41300
rect 411724 41300 412044 41660
rect 412460 41660 421796 41980
rect 422120 41938 423820 41980
rect 422120 41702 422162 41938
rect 422398 41702 423820 41938
rect 422120 41660 423820 41702
rect 424972 41938 441668 41980
rect 424972 41702 425014 41938
rect 425250 41702 441390 41938
rect 441626 41702 441668 41938
rect 424972 41660 441668 41702
rect 442084 41660 450684 41980
rect 412460 41300 412780 41660
rect 411724 40980 412780 41300
rect 421476 41300 421796 41660
rect 423500 41300 423820 41660
rect 442084 41300 442404 41660
rect 421476 40980 422440 41300
rect 423500 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41938 463932 41980
rect 451100 41702 463654 41938
rect 463890 41702 463932 41938
rect 451100 41660 463932 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 422120 40620 422440 40980
rect 422120 40578 425292 40620
rect 422120 40342 425014 40578
rect 425250 40342 425292 40578
rect 422120 40300 425292 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo ~/caravel_top_level/mag
timestamp 1638586901
transform 1 0 269370 0 1 5100
box -2520 0 15000 15560
use caravel_motto  caravel_motto ~/caravel_top_level/mag
timestamp 1637698310
transform 1 0 -54372 0 1 -4446
box 373080 14838 395618 19242
use caravel_power_routing  caravel_power_routing ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 0 0 1 0
box 6022 30806 711814 1031696
use caravel_clocking  clock_ctrl ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use copyright_block  copyright_block ~/caravel_top_level/mag
timestamp 1665519328
transform 1 0 149582 0 1 16298
box -262 -10348 35048 2764
use buff_flash_clkrst  flash_clkrst_buffers ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\] ~/caravel_top_level/mag
timestamp 1666360185
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666360185
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666360185
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666360185
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666360185
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666360185
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666360185
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666360185
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666360185
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666360185
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666360185
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1666360185
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1666360185
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1666360185
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1666360185
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1666360185
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666360185
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666360185
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666360185
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666360185
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666360185
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666360185
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666360185
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666360185
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666360185
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666360185
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666360185
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666360185
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666360185
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666360185
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666360185
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666360185
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1666360185
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1666360185
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1666360185
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1666360185
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1666360185
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1666360185
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0 ~/caravel_top_level/mag
timestamp 1666360185
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666360185
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666360185
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666360185
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666360185
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666360185
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666360185
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666360185
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666360185
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666360185
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666360185
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666360185
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666360185
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666360185
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1666360185
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1666360185
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1666360185
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1666360185
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1666360185
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1666360185
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1666360185
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1666360185
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1666360185
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1666360185
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1666360185
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666360185
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666360185
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666360185
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666360185
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666360185
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666360185
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666360185
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666360185
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666360185
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666360185
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666360185
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666360185
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666360185
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use mgmt_protect  mgmt_buffers ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use user_project_wrapper  mprj ~/caravel_top_level/mag
timestamp 1637147503
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use open_source  open_source ~/caravel_top_level/mag
timestamp 1666123577
transform 1 0 206098 0 1 2054
box 752 5164 29030 16242
use chip_io  padframe ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level ~/caravel_top_level/mag
timestamp 1666360185
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use gpio_signal_buffering  sigbuf ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
use mgmt_core_wrapper  soc ~/caravel_top_level/mag
timestamp 1665963385
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use spare_logic_block  spare_logic\[0\] ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666360185
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1666360185
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666360185
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock ~/caravel_top_level/mag
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use user_id_programming  user_id_value ~/caravel_top_level/mag
timestamp 1666360185
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal output
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal output
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal output
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal output
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19620 80934 0 FreeSans 16000 0 0 0 vccd
port 45 nsew power bidirectional
flabel metal5 s 697980 909666 711433 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew power bidirectional
flabel metal5 s 6167 914054 19620 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew power bidirectional
flabel metal5 s 624222 6811 636390 18976 0 FreeSans 16000 0 0 0 vdda
port 48 nsew power bidirectional
flabel metal5 s 698624 819822 710789 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew power bidirectional
flabel metal5 s 698624 505222 710789 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew power bidirectional
flabel metal5 s 6811 484410 18976 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew power bidirectional
flabel metal5 s 6811 111610 18976 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew power bidirectional
flabel metal5 s 6811 871210 18976 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew power bidirectional
flabel metal5 s 80222 6811 92390 18976 0 FreeSans 16000 0 0 0 vssa
port 54 nsew ground bidirectional
flabel metal5 s 577010 1018624 589178 1030789 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew ground bidirectional
flabel metal5 s 698624 417022 710789 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew ground bidirectional
flabel metal5 s 6811 829010 18976 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew ground bidirectional
flabel metal5 s 243266 6167 254146 19620 0 FreeSans 16000 0 0 0 vssd
port 58 nsew ground bidirectional
flabel metal5 s 697980 461866 711433 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew ground bidirectional
flabel metal5 s 6167 442854 19620 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew ground bidirectional
flabel metal5 s 570422 6811 582590 18976 0 FreeSans 16000 0 0 0 vssio
port 61 nsew ground bidirectional
flabel metal5 s 334810 1018624 346978 1030789 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
string LEFclass BLOCK
<< end >>
