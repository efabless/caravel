magic
tech sky130A
magscale 1 2
timestamp 1665259416
<< metal1 >>
rect 41866 995682 675734 995734
rect 41866 42225 41918 995682
rect 411070 42466 411076 42518
rect 411128 42506 411134 42518
rect 419718 42506 419724 42518
rect 411128 42478 419724 42506
rect 411128 42466 411134 42478
rect 419718 42466 419724 42478
rect 419776 42466 419782 42518
rect 465810 42476 465816 42528
rect 465868 42516 465874 42528
rect 474458 42516 474464 42528
rect 465868 42488 474464 42516
rect 465868 42476 465874 42488
rect 474458 42476 474464 42488
rect 474516 42476 474522 42528
rect 409230 42340 409236 42392
rect 409288 42380 409294 42392
rect 412266 42380 412272 42392
rect 409288 42352 412272 42380
rect 409288 42340 409294 42352
rect 412266 42340 412272 42352
rect 412324 42380 412330 42392
rect 415394 42380 415400 42392
rect 412324 42352 415400 42380
rect 412324 42340 412330 42352
rect 415394 42340 415400 42352
rect 415452 42340 415458 42392
rect 464004 42328 464010 42380
rect 464062 42368 464068 42380
rect 467040 42368 467046 42380
rect 464062 42340 467046 42368
rect 464062 42328 464068 42340
rect 467040 42328 467046 42340
rect 467098 42368 467104 42380
rect 470167 42368 470173 42380
rect 467098 42340 470173 42368
rect 467098 42328 467104 42340
rect 470167 42328 470173 42340
rect 470225 42328 470231 42380
rect 518802 42340 518808 42392
rect 518860 42380 518866 42392
rect 524966 42380 524972 42392
rect 518860 42352 524972 42380
rect 518860 42340 518866 42352
rect 524966 42340 524972 42352
rect 525024 42340 525030 42392
rect 675682 42225 675734 995682
rect 41866 42173 145035 42225
rect 145207 42173 195328 42225
rect 195380 42173 199653 42225
rect 199705 42173 303929 42225
rect 303981 42173 308066 42225
rect 308118 42173 358732 42225
rect 358784 42173 363053 42225
rect 363105 42173 413524 42225
rect 413576 42173 417858 42225
rect 417910 42173 468330 42225
rect 468382 42173 472656 42225
rect 472708 42173 523126 42225
rect 523178 42173 527457 42225
rect 527509 42173 675734 42225
rect 186548 42089 188522 42141
rect 188574 42089 192845 42141
rect 192897 42089 201494 42141
rect 201546 42089 202717 42141
rect 202769 42089 202775 42141
rect 295162 42089 297125 42141
rect 297177 42089 299607 42141
rect 299659 42089 305774 42141
rect 305826 42089 311317 42141
rect 311369 42089 311375 42141
rect 349962 42089 351925 42141
rect 351977 42089 354406 42141
rect 354458 42089 360570 42141
rect 360622 42089 366117 42141
rect 366169 42089 366175 42141
rect 404762 42089 406719 42141
rect 406771 42089 420917 42141
rect 420969 42089 420975 42141
rect 459562 42089 461524 42141
rect 461576 42089 475717 42141
rect 475769 42089 475775 42141
rect 514362 42089 516320 42141
rect 516372 42089 530517 42141
rect 530569 42089 530575 42141
rect 186548 42005 189163 42057
rect 189215 42005 191003 42057
rect 191055 42005 192202 42057
rect 192254 42005 193489 42057
rect 193541 42005 196528 42057
rect 196580 42005 197170 42057
rect 197222 42005 197813 42057
rect 197865 42005 198368 42057
rect 198420 42005 200206 42057
rect 200258 42005 200857 42057
rect 200909 42005 202563 42057
rect 202615 42005 202621 42057
rect 295162 42005 297768 42057
rect 297820 42005 300804 42057
rect 300856 42005 301451 42057
rect 301503 42005 302094 42057
rect 302146 42005 302643 42057
rect 302695 42005 305133 42057
rect 305185 42005 306418 42057
rect 306470 42005 308809 42057
rect 308861 42005 309452 42057
rect 309504 42005 311163 42057
rect 311215 42005 311221 42057
rect 349962 42005 352568 42057
rect 352620 42005 355600 42057
rect 355652 42005 356246 42057
rect 356298 42005 356889 42057
rect 356941 42005 357444 42057
rect 357496 42005 359928 42057
rect 359980 42005 361217 42057
rect 361269 42005 363607 42057
rect 363659 42005 364252 42057
rect 364304 42005 365963 42057
rect 366015 42005 366021 42057
rect 404762 42005 407367 42057
rect 407419 42005 410398 42057
rect 410450 42005 411691 42057
rect 411743 42005 414725 42057
rect 414777 42005 416013 42057
rect 416065 42005 418404 42057
rect 418456 42005 419045 42057
rect 419097 42005 420763 42057
rect 420815 42005 420821 42057
rect 459562 42005 462162 42057
rect 462214 42005 465201 42057
rect 465253 42005 466488 42057
rect 466540 42005 469522 42057
rect 469574 42005 470810 42057
rect 470862 42005 473201 42057
rect 473253 42005 473849 42057
rect 473901 42005 475563 42057
rect 475615 42005 475621 42057
rect 514362 42005 516969 42057
rect 517021 42005 520004 42057
rect 520056 42005 521293 42057
rect 521345 42005 524328 42057
rect 524380 42005 525615 42057
rect 525667 42005 528009 42057
rect 528061 42005 528652 42057
rect 528704 42005 530363 42057
rect 530415 42005 530421 42057
rect 186548 41921 187968 41973
rect 188020 41921 195973 41973
rect 196025 41921 202162 41973
rect 295162 41921 296576 41973
rect 296628 41921 304577 41973
rect 304629 41921 310827 41973
rect 349962 41921 351375 41973
rect 351427 41921 359374 41973
rect 359426 41921 365627 41973
rect 404762 41921 406170 41973
rect 406222 41921 414174 41973
rect 414226 41921 420427 41973
rect 459562 41921 460971 41973
rect 461023 41921 468967 41973
rect 469019 41921 475227 41973
rect 514362 41921 515772 41973
rect 515824 41921 523773 41973
rect 523825 41921 530027 41973
rect 186548 41837 186683 41889
rect 186735 41837 194688 41889
rect 194740 41837 199012 41889
rect 199064 41837 202162 41889
rect 295162 41837 295283 41889
rect 295335 41837 303290 41889
rect 303342 41837 307616 41889
rect 307668 41837 310827 41889
rect 349962 41837 350086 41889
rect 350138 41837 358090 41889
rect 358142 41837 362412 41889
rect 362464 41837 365627 41889
rect 404762 41837 404877 41889
rect 404929 41837 412888 41889
rect 412940 41837 417210 41889
rect 417262 41837 420427 41889
rect 459562 41837 459678 41889
rect 459730 41837 467684 41889
rect 467736 41837 472010 41889
rect 472062 41837 475227 41889
rect 514362 41837 514487 41889
rect 514539 41837 522486 41889
rect 522538 41837 526810 41889
rect 526862 41837 530027 41889
rect 140990 40073 140996 40125
rect 141048 40118 141054 40125
rect 141986 40118 141992 40125
rect 141048 40080 141992 40118
rect 141048 40073 141054 40080
rect 141986 40073 141992 40080
rect 142044 40118 142050 40125
rect 143062 40118 143068 40125
rect 142044 40080 143068 40118
rect 142044 40073 142050 40080
rect 143062 40073 143068 40080
rect 143120 40118 143126 40125
rect 143401 40118 143407 40125
rect 143120 40080 143407 40118
rect 143120 40073 143126 40080
rect 143401 40073 143407 40080
rect 143519 40118 143525 40125
rect 144597 40118 144603 40125
rect 143519 40080 144603 40118
rect 143519 40073 143525 40080
rect 144597 40073 144603 40080
rect 144655 40073 144661 40125
<< via1 >>
rect 411076 42466 411128 42518
rect 419724 42466 419776 42518
rect 465816 42476 465868 42528
rect 474464 42476 474516 42528
rect 409236 42340 409288 42392
rect 412272 42340 412324 42392
rect 415400 42340 415452 42392
rect 464010 42328 464062 42380
rect 467046 42328 467098 42380
rect 470173 42328 470225 42380
rect 518808 42340 518860 42392
rect 524972 42340 525024 42392
rect 145035 42173 145207 42225
rect 195328 42173 195380 42225
rect 199653 42173 199705 42225
rect 303929 42173 303981 42225
rect 308066 42173 308118 42225
rect 358732 42173 358784 42225
rect 363053 42173 363105 42225
rect 413524 42173 413576 42225
rect 417858 42173 417910 42225
rect 468330 42173 468382 42225
rect 472656 42173 472708 42225
rect 523126 42173 523178 42225
rect 527457 42173 527509 42225
rect 188522 42089 188574 42141
rect 192845 42089 192897 42141
rect 201494 42089 201546 42141
rect 202717 42089 202769 42141
rect 297125 42089 297177 42141
rect 299607 42089 299659 42141
rect 305774 42089 305826 42141
rect 311317 42089 311369 42141
rect 351925 42089 351977 42141
rect 354406 42089 354458 42141
rect 360570 42089 360622 42141
rect 366117 42089 366169 42141
rect 406719 42089 406771 42141
rect 420917 42089 420969 42141
rect 461524 42089 461576 42141
rect 475717 42089 475769 42141
rect 516320 42089 516372 42141
rect 530517 42089 530569 42141
rect 189163 42005 189215 42057
rect 191003 42005 191055 42057
rect 192202 42005 192254 42057
rect 193489 42005 193541 42057
rect 196528 42005 196580 42057
rect 197170 42005 197222 42057
rect 197813 42005 197865 42057
rect 198368 42005 198420 42057
rect 200206 42005 200258 42057
rect 200857 42005 200909 42057
rect 202563 42005 202615 42057
rect 297768 42005 297820 42057
rect 300804 42005 300856 42057
rect 301451 42005 301503 42057
rect 302094 42005 302146 42057
rect 302643 42005 302695 42057
rect 305133 42005 305185 42057
rect 306418 42005 306470 42057
rect 308809 42005 308861 42057
rect 309452 42005 309504 42057
rect 311163 42005 311215 42057
rect 352568 42005 352620 42057
rect 355600 42005 355652 42057
rect 356246 42005 356298 42057
rect 356889 42005 356941 42057
rect 357444 42005 357496 42057
rect 359928 42005 359980 42057
rect 361217 42005 361269 42057
rect 363607 42005 363659 42057
rect 364252 42005 364304 42057
rect 365963 42005 366015 42057
rect 407367 42005 407419 42057
rect 410398 42005 410450 42057
rect 411691 42005 411743 42057
rect 414725 42005 414777 42057
rect 416013 42005 416065 42057
rect 418404 42005 418456 42057
rect 419045 42005 419097 42057
rect 420763 42005 420815 42057
rect 462162 42005 462214 42057
rect 465201 42005 465253 42057
rect 466488 42005 466540 42057
rect 469522 42005 469574 42057
rect 470810 42005 470862 42057
rect 473201 42005 473253 42057
rect 473849 42005 473901 42057
rect 475563 42005 475615 42057
rect 516969 42005 517021 42057
rect 520004 42005 520056 42057
rect 521293 42005 521345 42057
rect 524328 42005 524380 42057
rect 525615 42005 525667 42057
rect 528009 42005 528061 42057
rect 528652 42005 528704 42057
rect 530363 42005 530415 42057
rect 187968 41921 188020 41973
rect 195973 41921 196025 41973
rect 296576 41921 296628 41973
rect 304577 41921 304629 41973
rect 351375 41921 351427 41973
rect 359374 41921 359426 41973
rect 406170 41921 406222 41973
rect 414174 41921 414226 41973
rect 460971 41921 461023 41973
rect 468967 41921 469019 41973
rect 515772 41921 515824 41973
rect 523773 41921 523825 41973
rect 186683 41837 186735 41889
rect 194688 41837 194740 41889
rect 199012 41837 199064 41889
rect 295283 41837 295335 41889
rect 303290 41837 303342 41889
rect 307616 41837 307668 41889
rect 350086 41837 350138 41889
rect 358090 41837 358142 41889
rect 362412 41837 362464 41889
rect 404877 41837 404929 41889
rect 412888 41837 412940 41889
rect 417210 41837 417262 41889
rect 459678 41837 459730 41889
rect 467684 41837 467736 41889
rect 472010 41837 472062 41889
rect 514487 41837 514539 41889
rect 522486 41837 522538 41889
rect 526810 41837 526862 41889
rect 140996 40073 141048 40125
rect 141992 40073 142044 40125
rect 143068 40073 143120 40125
rect 143407 40073 143519 40125
rect 144603 40073 144655 40125
<< metal2 >>
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 90021 995407 90077 995887
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 141421 995407 141477 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192821 995407 192877 995887
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244221 995407 244277 995887
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 295821 995407 295877 995887
rect 297017 995407 297073 995887
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 397621 995407 397677 995887
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 486621 995407 486677 995887
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 538021 995407 538077 995887
rect 539217 995407 539273 995887
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639821 995407 639877 995887
rect 641017 995407 641073 995887
rect 41713 969217 42193 969273
rect 41713 968021 42193 968077
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 41713 965537 42193 965593
rect 675407 965407 675887 965463
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 675407 963567 675887 963623
rect 41713 963053 42193 963109
rect 675407 963015 675887 963071
rect 41713 962501 42193 962557
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 675407 959243 675887 959299
rect 41713 958729 42193 958785
rect 675407 958691 675887 958747
rect 41713 958177 42193 958233
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 41713 956337 42193 956393
rect 675407 956207 675887 956263
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675407 953723 675887 953779
rect 675407 952527 675887 952583
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 864523 675887 864579
rect 675407 863327 675887 863383
rect 41713 799417 42193 799473
rect 41713 798221 42193 798277
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 775323 675887 775379
rect 675407 774127 675887 774183
rect 41713 756217 42193 756273
rect 41713 755021 42193 755077
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41713 743337 42193 743393
rect 675407 743295 675887 743351
rect 41713 742693 42193 742749
rect 675407 742651 675887 742707
rect 41713 742049 42193 742105
rect 675407 742007 675887 742063
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 730323 675887 730379
rect 675407 729127 675887 729183
rect 41713 713017 42193 713073
rect 41713 711821 42193 711877
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 685323 675887 685379
rect 675407 684127 675887 684183
rect 41713 669817 42193 669873
rect 41713 668621 42193 668677
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 640123 675887 640179
rect 675407 638927 675887 638983
rect 41713 626617 42193 626673
rect 41713 625421 42193 625477
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 595123 675887 595179
rect 675407 593927 675887 593983
rect 41713 583417 42193 583473
rect 41713 582221 42193 582277
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 549923 675887 549979
rect 675407 548727 675887 548783
rect 41713 540217 42193 540273
rect 41713 539021 42193 539077
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 412617 42193 412673
rect 41713 411421 42193 411477
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 372723 675887 372779
rect 675407 371527 675887 371583
rect 41713 369417 42193 369473
rect 41713 368221 42193 368277
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 327523 675887 327579
rect 675407 326327 675887 326383
rect 41713 326217 42193 326273
rect 41713 325021 42193 325077
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 41713 283017 42193 283073
rect 675407 282523 675887 282579
rect 41713 281821 42193 281877
rect 675407 281327 675887 281383
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 41713 239817 42193 239873
rect 41713 238621 42193 238677
rect 675407 238167 675887 238223
rect 41713 237977 42193 238033
rect 675407 237523 675887 237579
rect 675407 236327 675887 236383
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 41713 196617 42193 196673
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 41713 195421 42193 195477
rect 41713 194777 42193 194833
rect 675407 194807 675887 194863
rect 41713 192937 42193 192993
rect 675407 192967 675887 193023
rect 675407 192323 675887 192379
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 675407 191127 675887 191183
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 147323 675887 147379
rect 675407 146127 675887 146183
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 102123 675887 102179
rect 675407 100927 675887 100983
rect 465816 42528 465868 42534
rect 411076 42518 411128 42524
rect 411076 42460 411128 42466
rect 419724 42518 419776 42524
rect 465816 42470 465868 42476
rect 474464 42528 474516 42534
rect 474464 42470 474516 42476
rect 419724 42460 419776 42466
rect 409236 42392 409288 42398
rect 409236 42334 409288 42340
rect 195331 42231 195387 42242
rect 199655 42231 199711 42243
rect 303931 42231 303987 42240
rect 145035 42225 145207 42231
rect 195328 42225 195387 42231
rect 145035 42167 145207 42173
rect 140996 40125 141048 40131
rect 141992 40125 142044 40131
rect 140996 40067 141048 40073
rect 141986 40073 141992 40120
rect 143068 40125 143120 40131
rect 142044 40073 142050 40120
rect 141004 39990 141042 40067
rect 141667 39934 141813 40000
rect 141986 39998 142050 40073
rect 143407 40125 143519 40131
rect 144603 40125 144655 40131
rect 143068 40067 143120 40073
rect 143078 39996 143110 40067
rect 143398 40034 143407 40090
rect 143519 40034 143528 40090
rect 144603 40067 144655 40073
rect 144610 39990 144652 40067
rect 145106 39990 145136 42167
rect 186683 41889 186735 41895
rect 186683 41831 186735 41837
rect 187327 41713 187383 42193
rect 188522 42141 188574 42147
rect 188522 42083 188574 42089
rect 192845 42141 192897 42147
rect 192845 42083 192897 42089
rect 189163 42057 189215 42063
rect 189163 41999 189215 42005
rect 191003 42057 191055 42063
rect 191003 41999 191055 42005
rect 192202 42057 192254 42063
rect 192202 41999 192254 42005
rect 193489 42057 193541 42063
rect 193489 41999 193541 42005
rect 187968 41973 188020 41979
rect 187968 41915 188020 41921
rect 194043 41713 194099 42193
rect 195380 42173 195387 42225
rect 195328 42167 195387 42173
rect 199653 42225 199711 42231
rect 199705 42173 199711 42225
rect 199653 42167 199711 42173
rect 303929 42225 303987 42231
rect 303981 42173 303987 42225
rect 308065 42225 308121 42248
rect 303929 42167 303987 42173
rect 195331 42137 195387 42167
rect 199655 42137 199711 42167
rect 201494 42141 201546 42147
rect 201494 42083 201546 42089
rect 202717 42141 202769 42147
rect 196528 42057 196580 42063
rect 196528 41999 196580 42005
rect 197170 42057 197222 42063
rect 197170 41999 197222 42005
rect 197813 42057 197865 42063
rect 197813 41999 197865 42005
rect 198368 42057 198420 42063
rect 198368 41999 198420 42005
rect 200206 42057 200258 42063
rect 200206 41999 200258 42005
rect 200857 42057 200909 42063
rect 200857 41999 200909 42005
rect 202563 42057 202615 42063
rect 195973 41973 196025 41979
rect 195973 41915 196025 41921
rect 194688 41889 194740 41895
rect 194688 41831 194740 41837
rect 199012 41889 199064 41895
rect 199012 41831 199064 41837
rect 202563 40955 202615 42005
rect 202559 40946 202619 40955
rect 202559 40877 202619 40886
rect 202717 40782 202769 42089
rect 297125 42141 297177 42147
rect 297125 42083 297177 42089
rect 299607 42141 299659 42147
rect 303931 42137 303987 42167
rect 305774 42141 305826 42147
rect 299607 42083 299659 42089
rect 305774 42083 305826 42089
rect 297768 42057 297820 42063
rect 297768 41999 297820 42005
rect 300804 42057 300856 42063
rect 300804 41999 300856 42005
rect 301451 42057 301503 42063
rect 301451 41999 301503 42005
rect 302094 42057 302146 42063
rect 302094 41999 302146 42005
rect 302643 42057 302695 42063
rect 302643 41999 302695 42005
rect 305133 42057 305185 42063
rect 305133 41999 305185 42005
rect 306418 42057 306470 42063
rect 306418 41999 306470 42005
rect 296576 41973 296628 41979
rect 296576 41915 296628 41921
rect 304577 41973 304629 41979
rect 304577 41915 304629 41921
rect 295283 41889 295335 41895
rect 295283 41831 295335 41837
rect 303290 41889 303342 41895
rect 303290 41831 303342 41837
rect 306967 41713 307023 42193
rect 308065 42173 308066 42225
rect 308118 42173 308121 42225
rect 358731 42225 358787 42240
rect 363055 42231 363111 42240
rect 308065 42129 308121 42173
rect 308255 42129 308311 42193
rect 308065 42073 308311 42129
rect 307616 41889 307668 41895
rect 307616 41831 307668 41837
rect 308255 41713 308311 42073
rect 308809 42057 308861 42063
rect 308809 41999 308861 42005
rect 309452 42057 309504 42063
rect 309452 41999 309504 42005
rect 310095 41713 310151 42193
rect 358731 42173 358732 42225
rect 358784 42173 358787 42225
rect 363053 42225 363111 42231
rect 311317 42141 311369 42147
rect 311163 42057 311215 42063
rect 311163 40955 311215 42005
rect 311159 40946 311219 40955
rect 311159 40877 311219 40886
rect 311317 40782 311369 42089
rect 351925 42141 351977 42147
rect 351925 42083 351977 42089
rect 354406 42141 354458 42147
rect 358731 42137 358787 42173
rect 360570 42141 360622 42147
rect 354406 42083 354458 42089
rect 360570 42083 360622 42089
rect 352568 42057 352620 42063
rect 352568 41999 352620 42005
rect 355600 42057 355652 42063
rect 355600 41999 355652 42005
rect 356246 42057 356298 42063
rect 356246 41999 356298 42005
rect 356889 42057 356941 42063
rect 356889 41999 356941 42005
rect 357444 42057 357496 42063
rect 357444 41999 357496 42005
rect 359928 42057 359980 42063
rect 359928 41999 359980 42005
rect 361217 42057 361269 42063
rect 361217 41999 361269 42005
rect 351375 41973 351427 41979
rect 351375 41915 351427 41921
rect 359374 41973 359426 41979
rect 359374 41915 359426 41921
rect 350086 41889 350138 41895
rect 350086 41831 350138 41837
rect 358090 41889 358142 41895
rect 358090 41831 358142 41837
rect 361767 41713 361823 42193
rect 363105 42173 363111 42225
rect 363053 42167 363111 42173
rect 363055 42137 363111 42167
rect 363607 42057 363659 42063
rect 363607 41999 363659 42005
rect 364252 42057 364304 42063
rect 364252 41999 364304 42005
rect 362412 41889 362464 41895
rect 362412 41831 362464 41837
rect 364895 41713 364951 42193
rect 366117 42141 366169 42147
rect 365963 42057 366015 42063
rect 365963 40955 366015 42005
rect 365959 40946 366019 40955
rect 365959 40877 366019 40886
rect 366117 40782 366169 42089
rect 404877 41889 404929 41895
rect 404877 41831 404929 41837
rect 405527 41713 405583 42193
rect 406719 42141 406771 42147
rect 406719 42083 406771 42089
rect 407367 42057 407419 42063
rect 407367 41999 407419 42005
rect 406170 41973 406222 41979
rect 406170 41915 406222 41921
rect 409248 41820 409276 42334
rect 410398 42057 410450 42063
rect 410398 41999 410450 42005
rect 411088 41820 411116 42460
rect 412272 42392 412324 42398
rect 412272 42334 412324 42340
rect 415400 42392 415452 42398
rect 415400 42334 415452 42340
rect 412284 42193 412312 42334
rect 413531 42231 413587 42240
rect 411691 42057 411743 42063
rect 411691 41999 411743 42005
rect 412243 41820 412312 42193
rect 413524 42225 413587 42231
rect 413576 42173 413587 42225
rect 413524 42167 413587 42173
rect 413531 42135 413587 42167
rect 414725 42057 414777 42063
rect 414725 41999 414777 42005
rect 414174 41973 414226 41979
rect 414174 41915 414226 41921
rect 412888 41889 412940 41895
rect 412888 41831 412940 41837
rect 415412 41820 415440 42334
rect 417855 42225 417911 42236
rect 416013 42057 416065 42063
rect 416013 41999 416065 42005
rect 412243 41713 412299 41820
rect 416567 41713 416623 42193
rect 417855 42173 417858 42225
rect 417910 42173 417911 42225
rect 419736 42193 419764 42460
rect 464010 42380 464062 42386
rect 417855 42137 417911 42173
rect 418404 42057 418456 42063
rect 418404 41999 418456 42005
rect 419045 42057 419097 42063
rect 419045 41999 419097 42005
rect 417210 41889 417262 41895
rect 417210 41831 417262 41837
rect 419695 41820 419764 42193
rect 420917 42141 420969 42147
rect 420763 42057 420815 42063
rect 419695 41713 419751 41820
rect 420763 40955 420815 42005
rect 420759 40946 420819 40955
rect 420759 40877 420819 40886
rect 420917 40782 420969 42089
rect 459678 41889 459730 41895
rect 459678 41831 459730 41837
rect 460327 41713 460383 42193
rect 464010 42180 464062 42328
rect 461524 42141 461576 42147
rect 461524 42083 461576 42089
rect 462162 42057 462214 42063
rect 462162 41999 462214 42005
rect 465201 42057 465253 42063
rect 465201 41999 465253 42005
rect 460971 41973 461023 41979
rect 460971 41915 461023 41921
rect 465828 41834 465856 42470
rect 467046 42380 467098 42386
rect 467046 42193 467098 42328
rect 470173 42380 470225 42386
rect 468331 42231 468387 42245
rect 468330 42225 468387 42231
rect 466488 42057 466540 42063
rect 466488 41999 466540 42005
rect 465828 41806 465875 41834
rect 467043 41713 467099 42193
rect 468382 42173 468387 42225
rect 470173 42181 470225 42328
rect 472655 42225 472711 42235
rect 468330 42167 468387 42173
rect 468331 42135 468387 42167
rect 469522 42057 469574 42063
rect 469522 41999 469574 42005
rect 470810 42057 470862 42063
rect 470810 41999 470862 42005
rect 468967 41973 469019 41979
rect 468967 41915 469019 41921
rect 467684 41889 467736 41895
rect 467684 41831 467736 41837
rect 471367 41713 471423 42193
rect 472655 42173 472656 42225
rect 472708 42173 472711 42225
rect 472655 42132 472711 42173
rect 474476 42193 474504 42470
rect 518808 42392 518860 42398
rect 518808 42334 518860 42340
rect 524972 42392 525024 42398
rect 524972 42334 525024 42340
rect 473201 42057 473253 42063
rect 473201 41999 473253 42005
rect 473849 42057 473901 42063
rect 473849 41999 473901 42005
rect 472010 41889 472062 41895
rect 472010 41831 472062 41837
rect 474476 41806 474551 42193
rect 475717 42141 475769 42147
rect 474495 41713 474551 41806
rect 475563 42057 475615 42063
rect 475563 40955 475615 42005
rect 475559 40946 475619 40955
rect 475559 40877 475619 40886
rect 475717 40782 475769 42089
rect 514487 41889 514539 41895
rect 514487 41831 514539 41837
rect 515127 41713 515183 42193
rect 516320 42141 516372 42147
rect 516320 42083 516372 42089
rect 516969 42057 517021 42063
rect 516969 41999 517021 42005
rect 515772 41973 515824 41979
rect 515772 41915 515824 41921
rect 518820 41820 518848 42334
rect 523131 42231 523187 42251
rect 523126 42225 523187 42231
rect 520004 42057 520056 42063
rect 520004 41999 520056 42005
rect 520647 41713 520703 42193
rect 521293 42057 521345 42063
rect 521293 41999 521345 42005
rect 521843 41713 521899 42193
rect 523178 42173 523187 42225
rect 524984 42193 525012 42334
rect 527455 42225 527511 42249
rect 523126 42167 523187 42173
rect 523131 42128 523187 42167
rect 524328 42057 524380 42063
rect 524328 41999 524380 42005
rect 523773 41973 523825 41979
rect 523773 41915 523825 41921
rect 522486 41889 522538 41895
rect 522486 41831 522538 41837
rect 524971 41713 525027 42193
rect 525615 42057 525667 42063
rect 525615 41999 525667 42005
rect 526167 41713 526223 42193
rect 527455 42173 527457 42225
rect 527509 42173 527511 42225
rect 527455 42120 527511 42173
rect 528009 42057 528061 42063
rect 528009 41999 528061 42005
rect 528652 42057 528704 42063
rect 528652 41999 528704 42005
rect 526810 41889 526862 41895
rect 526810 41831 526862 41837
rect 529295 41713 529351 42193
rect 530517 42141 530569 42147
rect 530363 42057 530415 42063
rect 530363 40955 530415 42005
rect 530359 40946 530419 40955
rect 530359 40877 530419 40886
rect 530517 40782 530569 42089
rect 145830 40774 145888 40781
rect 145828 40772 145888 40774
rect 145828 40716 145830 40772
rect 145886 40716 145888 40772
rect 145828 40703 145888 40716
rect 202713 40773 202773 40782
rect 202713 40704 202773 40713
rect 311313 40773 311373 40782
rect 311313 40704 311373 40713
rect 366113 40773 366173 40782
rect 366113 40704 366173 40713
rect 420913 40773 420973 40782
rect 420913 40704 420973 40713
rect 475713 40773 475773 40782
rect 475713 40704 475773 40713
rect 530513 40773 530573 40782
rect 530513 40704 530573 40713
rect 145852 40134 145888 40703
rect 145828 40074 145837 40134
rect 145897 40074 145906 40134
<< via2 >>
rect 143407 40073 143519 40090
rect 143407 40034 143519 40073
rect 202559 40886 202619 40946
rect 311159 40886 311219 40946
rect 365959 40886 366019 40946
rect 420759 40886 420819 40946
rect 475559 40886 475619 40946
rect 530359 40886 530419 40946
rect 145830 40716 145886 40772
rect 202713 40713 202773 40773
rect 311313 40713 311373 40773
rect 366113 40713 366173 40773
rect 420913 40713 420973 40773
rect 475713 40713 475773 40773
rect 530513 40713 530573 40773
rect 145837 40074 145897 40134
<< metal3 >>
rect 40854 926876 46818 926940
rect 40854 922268 44294 926876
rect 46702 922268 46818 926876
rect 40854 922151 46818 922268
rect 670772 922374 676724 922500
rect 40854 921736 46818 921852
rect 40854 917280 41096 921736
rect 43504 917280 46818 921736
rect 670772 917822 674136 922374
rect 676496 917822 676724 922374
rect 670772 917700 676724 917822
rect 40854 917190 46818 917280
rect 670772 917268 676724 917410
rect 40854 916770 46818 916900
rect 40854 912162 44274 916770
rect 46682 912162 46818 916770
rect 670772 912862 670974 917268
rect 673314 912862 676724 917268
rect 670772 912748 676724 912862
rect 40854 912100 46818 912162
rect 670772 912322 676724 912449
rect 670772 907790 674170 912322
rect 676504 907790 676724 912322
rect 670772 907660 676724 907790
rect 670794 474564 676878 474700
rect 670794 470046 670926 474564
rect 673294 470046 676878 474564
rect 670794 469900 676878 470046
rect 670794 469480 676878 469600
rect 670794 465058 674144 469480
rect 676512 465058 676878 469480
rect 670794 464949 676878 465058
rect 670794 464548 676878 464649
rect 670794 460030 670932 464548
rect 673300 460030 676878 464548
rect 670794 459860 676878 460030
rect 41220 455654 46828 455740
rect 43508 451042 46828 455654
rect 41220 450951 46828 451042
rect 41220 450528 46828 450651
rect 41220 446104 44290 450528
rect 46690 446104 46828 450528
rect 41220 446000 46828 446104
rect 41220 445596 46828 445700
rect 43488 440984 46828 445596
rect 41220 440900 46828 440984
rect 202554 40946 202624 40951
rect 311154 40946 311224 40951
rect 365954 40946 366024 40951
rect 420754 40946 420824 40951
rect 475554 40946 475624 40951
rect 530354 40946 530424 40951
rect 202554 40886 202559 40946
rect 202619 40886 204878 40946
rect 202554 40881 202624 40886
rect 145825 40774 145891 40777
rect 145825 40772 148252 40774
rect 145825 40716 145830 40772
rect 145886 40716 148252 40772
rect 145825 40714 148252 40716
rect 202708 40773 202778 40778
rect 145825 40711 145891 40714
rect 202708 40713 202713 40773
rect 202773 40713 203064 40773
rect 204818 40713 204878 40886
rect 311154 40886 311159 40946
rect 311219 40886 314473 40946
rect 311154 40881 311224 40886
rect 311308 40773 311378 40778
rect 311308 40713 311313 40773
rect 311373 40713 312684 40773
rect 202708 40708 202778 40713
rect 311308 40708 311378 40713
rect 314413 40704 314473 40886
rect 365954 40886 365959 40946
rect 366019 40886 369270 40946
rect 365954 40881 366024 40886
rect 366108 40773 366178 40778
rect 366108 40713 366113 40773
rect 366173 40713 367484 40773
rect 369210 40716 369270 40886
rect 420754 40886 420759 40946
rect 420819 40886 424060 40946
rect 420754 40881 420824 40886
rect 420908 40773 420978 40778
rect 420908 40713 420913 40773
rect 420973 40713 422262 40773
rect 366108 40708 366178 40713
rect 420908 40708 420978 40713
rect 424000 40712 424060 40886
rect 475554 40886 475559 40946
rect 475619 40886 478875 40946
rect 475554 40881 475624 40886
rect 475708 40773 475778 40778
rect 475708 40713 475713 40773
rect 475773 40713 477055 40773
rect 475708 40708 475778 40713
rect 478815 40712 478875 40886
rect 530354 40886 530359 40946
rect 530419 40886 533657 40946
rect 530354 40881 530424 40886
rect 530508 40773 530578 40778
rect 530508 40713 530513 40773
rect 530573 40713 531856 40773
rect 530508 40708 530578 40713
rect 533597 40712 533657 40886
rect 148901 40316 149351 40338
rect 133094 40158 144010 40218
rect 133094 39984 133154 40158
rect 143407 40095 143519 40097
rect 143402 40090 143524 40095
rect 143402 40034 143407 40090
rect 143519 40034 143524 40090
rect 143402 39992 143524 40034
rect 143950 39984 144010 40158
rect 145832 40134 145902 40148
rect 145832 40074 145837 40134
rect 145897 40074 145902 40134
rect 145832 39982 145902 40074
rect 148901 40054 149134 40316
rect 149314 40054 149351 40316
rect 148901 31600 149351 40054
rect 149537 40321 149918 40342
rect 149537 39976 149634 40321
rect 149814 39976 149918 40321
rect 149537 38153 149918 39976
rect 149537 37372 149563 38153
rect 149891 37372 149918 38153
rect 149537 37340 149918 37372
rect 203701 40316 204151 40338
rect 203701 40054 203934 40316
rect 204114 40054 204151 40316
rect 148901 30843 148940 31600
rect 149305 30843 149351 31600
rect 148901 30806 149351 30843
rect 203701 31600 204151 40054
rect 204337 40321 204718 40342
rect 204337 39976 204434 40321
rect 204614 39976 204718 40321
rect 204337 38153 204718 39976
rect 204337 37372 204363 38153
rect 204691 37372 204718 38153
rect 204337 37340 204718 37372
rect 313301 40316 313751 40338
rect 313301 40054 313534 40316
rect 313714 40054 313751 40316
rect 203701 30843 203740 31600
rect 204105 30843 204151 31600
rect 203701 30806 204151 30843
rect 313301 31600 313751 40054
rect 313937 40321 314318 40342
rect 313937 39976 314034 40321
rect 314214 39976 314318 40321
rect 313937 38153 314318 39976
rect 313937 37372 313963 38153
rect 314291 37372 314318 38153
rect 313937 37340 314318 37372
rect 368101 40316 368551 40338
rect 368101 40054 368334 40316
rect 368514 40054 368551 40316
rect 313301 30843 313340 31600
rect 313705 30843 313751 31600
rect 313301 30806 313751 30843
rect 368101 31600 368551 40054
rect 368737 40321 369118 40342
rect 368737 39976 368834 40321
rect 369014 39976 369118 40321
rect 368737 38153 369118 39976
rect 368737 37372 368763 38153
rect 369091 37372 369118 38153
rect 368737 37340 369118 37372
rect 422901 40316 423351 40338
rect 422901 40054 423134 40316
rect 423314 40054 423351 40316
rect 368101 30843 368140 31600
rect 368505 30843 368551 31600
rect 368101 30806 368551 30843
rect 422901 31600 423351 40054
rect 423537 40321 423918 40342
rect 423537 39976 423634 40321
rect 423814 39976 423918 40321
rect 423537 38153 423918 39976
rect 423537 37372 423563 38153
rect 423891 37372 423918 38153
rect 423537 37340 423918 37372
rect 477701 40316 478151 40338
rect 477701 40054 477934 40316
rect 478114 40054 478151 40316
rect 422901 30843 422940 31600
rect 423305 30843 423351 31600
rect 422901 30806 423351 30843
rect 477701 31600 478151 40054
rect 478337 40321 478718 40342
rect 478337 39976 478434 40321
rect 478614 39976 478718 40321
rect 478337 38153 478718 39976
rect 478337 37372 478363 38153
rect 478691 37372 478718 38153
rect 478337 37340 478718 37372
rect 532501 40316 532951 40338
rect 532501 40054 532734 40316
rect 532914 40054 532951 40316
rect 477701 30843 477740 31600
rect 478105 30843 478151 31600
rect 477701 30806 478151 30843
rect 532501 31600 532951 40054
rect 533137 40321 533518 40342
rect 533137 39976 533234 40321
rect 533414 39976 533518 40321
rect 533137 38153 533518 39976
rect 533137 37372 533163 38153
rect 533491 37372 533518 38153
rect 533137 37340 533518 37372
rect 532501 30843 532540 31600
rect 532905 30843 532951 31600
rect 532501 30806 532951 30843
<< via3 >>
rect 44294 922268 46702 926876
rect 41096 917280 43504 921736
rect 674136 917822 676496 922374
rect 44274 912162 46682 916770
rect 670974 912862 673314 917268
rect 674170 907790 676504 912322
rect 670926 470046 673294 474564
rect 674144 465058 676512 469480
rect 670932 460030 673300 464548
rect 41142 451042 43508 455654
rect 44290 446104 46690 450528
rect 41122 440984 43488 445596
rect 149134 40054 149314 40316
rect 149634 39976 149814 40321
rect 149563 37372 149891 38153
rect 203934 40054 204114 40316
rect 148940 30843 149305 31600
rect 204434 39976 204614 40321
rect 204363 37372 204691 38153
rect 313534 40054 313714 40316
rect 203740 30843 204105 31600
rect 314034 39976 314214 40321
rect 313963 37372 314291 38153
rect 368334 40054 368514 40316
rect 313340 30843 313705 31600
rect 368834 39976 369014 40321
rect 368763 37372 369091 38153
rect 423134 40054 423314 40316
rect 368140 30843 368505 31600
rect 423634 39976 423814 40321
rect 423563 37372 423891 38153
rect 477934 40054 478114 40316
rect 422940 30843 423305 31600
rect 478434 39976 478614 40321
rect 478363 37372 478691 38153
rect 532734 40054 532914 40316
rect 477740 30843 478105 31600
rect 533234 39976 533414 40321
rect 533163 37372 533491 38153
rect 532540 30843 532905 31600
<< metal4 >>
rect 44198 926876 46800 926958
rect 44198 922268 44294 926876
rect 46702 922268 46800 926876
rect 44198 922154 46800 922268
rect 674010 922374 676616 922486
rect 40982 921736 43584 921844
rect 40982 917280 41096 921736
rect 43504 917280 43584 921736
rect 674010 917822 674136 922374
rect 676496 917822 676616 922374
rect 674010 917716 676616 917822
rect 40982 917186 43584 917280
rect 670826 917268 673434 917414
rect 44194 916770 46796 916898
rect 44194 912162 44274 916770
rect 46682 912162 46796 916770
rect 670826 912862 670974 917268
rect 673314 912862 673434 917268
rect 670826 912756 673434 912862
rect 44194 912094 46796 912162
rect 674016 912322 676622 912440
rect 674016 907790 674170 912322
rect 676504 907790 676622 912322
rect 674016 907670 676622 907790
rect 670824 474564 673424 474684
rect 670824 470046 670926 474564
rect 673294 470046 673424 474564
rect 670824 469900 673424 470046
rect 674024 469480 676618 469590
rect 674024 465058 674144 469480
rect 676512 465058 676618 469480
rect 674024 464954 676618 465058
rect 670826 464548 673426 464648
rect 670826 460030 670932 464548
rect 673300 460030 673426 464548
rect 670826 459864 673426 460030
rect 28653 440800 28719 455800
rect 36323 455607 37013 455799
rect 41008 455654 43618 455758
rect 41008 451042 41142 455654
rect 43508 451042 43618 455654
rect 41008 450950 43618 451042
rect 44202 450528 46812 450636
rect 44202 446104 44290 450528
rect 46690 446104 46812 450528
rect 44202 446016 46812 446104
rect 40994 445596 43604 445704
rect 40994 440984 41122 445596
rect 43488 440984 43604 445596
rect 40994 440896 43604 440984
rect 149632 40321 149816 40323
rect 149132 40316 149316 40318
rect 149132 40054 149134 40316
rect 149314 40054 149316 40316
rect 149132 40052 149316 40054
rect 149632 39976 149634 40321
rect 149814 39976 149816 40321
rect 204432 40321 204616 40323
rect 203932 40316 204116 40318
rect 203932 40054 203934 40316
rect 204114 40054 204116 40316
rect 203932 40052 204116 40054
rect 149632 39974 149816 39976
rect 204432 39976 204434 40321
rect 204614 39976 204616 40321
rect 314032 40321 314216 40323
rect 313532 40316 313716 40318
rect 313532 40054 313534 40316
rect 313714 40054 313716 40316
rect 313532 40052 313716 40054
rect 204432 39974 204616 39976
rect 314032 39976 314034 40321
rect 314214 39976 314216 40321
rect 368832 40321 369016 40323
rect 368332 40316 368516 40318
rect 368332 40054 368334 40316
rect 368514 40054 368516 40316
rect 368332 40052 368516 40054
rect 314032 39974 314216 39976
rect 368832 39976 368834 40321
rect 369014 39976 369016 40321
rect 423632 40321 423816 40323
rect 423132 40316 423316 40318
rect 423132 40054 423134 40316
rect 423314 40054 423316 40316
rect 423132 40052 423316 40054
rect 368832 39974 369016 39976
rect 423632 39976 423634 40321
rect 423814 39976 423816 40321
rect 478432 40321 478616 40323
rect 477932 40316 478116 40318
rect 477932 40054 477934 40316
rect 478114 40054 478116 40316
rect 477932 40052 478116 40054
rect 423632 39974 423816 39976
rect 478432 39976 478434 40321
rect 478614 39976 478616 40321
rect 533232 40321 533416 40323
rect 532732 40316 532916 40318
rect 532732 40054 532734 40316
rect 532914 40054 532916 40316
rect 532732 40052 532916 40054
rect 478432 39974 478616 39976
rect 533232 39976 533234 40321
rect 533414 39976 533416 40321
rect 533232 39974 533416 39976
rect 132600 36323 132792 37013
<< via4 >>
rect 44294 922268 46702 926876
rect 41096 917280 43504 921736
rect 674136 917822 676496 922374
rect 44274 912162 46682 916770
rect 670974 912862 673314 917268
rect 674170 907790 676504 912322
rect 670926 470046 673294 474564
rect 674144 465058 676512 469480
rect 670932 460030 673300 464548
rect 41142 451042 43508 455654
rect 44290 446104 46690 450528
rect 41122 440984 43488 445596
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 348400 1007147 348466 1008947
rect 348400 1004968 348466 1005617
rect 348400 1000607 348527 1001257
rect 6598 956440 19088 968960
rect 6167 914054 19619 924934
rect 40998 921736 43598 995004
rect 40998 917280 41096 921736
rect 43504 917280 43598 921736
rect 6811 871210 18975 883378
rect 6811 829010 18975 841178
rect 6598 786640 19088 799160
rect 6598 743440 19088 755960
rect 6598 700240 19088 712760
rect 6598 657040 19088 669560
rect 6598 613840 19088 626360
rect 6598 570640 19088 583160
rect 6598 527440 19088 539960
rect 6811 484410 18975 496578
rect 40998 455654 43598 917280
rect 6167 442854 19619 453734
rect 40998 451042 41142 455654
rect 43508 451042 43598 455654
rect 40998 445596 43598 451042
rect 40998 440984 41122 445596
rect 43488 440984 43598 445596
rect 6598 399840 19088 412360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 6598 227040 19088 239560
rect 6598 183840 19088 196360
rect 40998 179300 43598 440984
rect 44198 926876 46798 995004
rect 44198 922268 44294 926876
rect 46702 922268 46798 926876
rect 44198 916770 46798 922268
rect 44198 912162 44274 916770
rect 46682 912162 46798 916770
rect 44198 450528 46798 912162
rect 44198 446104 44290 450528
rect 46690 446104 46798 450528
rect 44198 179300 46798 446104
rect 670820 917268 673420 992714
rect 670820 912862 670974 917268
rect 673314 912862 673420 917268
rect 670820 474564 673420 912862
rect 670820 470046 670926 474564
rect 673294 470046 673420 474564
rect 670820 464548 673420 470046
rect 670820 460030 670932 464548
rect 673300 460030 673420 464548
rect 6811 111610 18975 123778
rect 670820 95156 673420 460030
rect 674020 922374 676620 992714
rect 698512 952840 711002 965360
rect 674020 917822 674136 922374
rect 676496 917822 676620 922374
rect 674020 912322 676620 917822
rect 674020 907790 674170 912322
rect 676504 907790 676620 912322
rect 697980 909666 711432 920546
rect 674020 469480 676620 907790
rect 698512 863640 711002 876160
rect 698624 819822 710788 831990
rect 698512 774440 711002 786960
rect 698512 729440 711002 741960
rect 698512 684440 711002 696960
rect 698512 639240 711002 651760
rect 698512 594240 711002 606760
rect 698512 549040 711002 561560
rect 698624 505222 710788 517390
rect 674020 465058 674144 469480
rect 676512 465058 676620 469480
rect 674020 95156 676620 465058
rect 697980 461866 711432 472746
rect 698624 417022 710788 429190
rect 698512 371840 711002 384360
rect 698512 326640 711002 339160
rect 698512 281640 711002 294160
rect 698512 236640 711002 249160
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__com_bus_slice_20um  FILLER_5 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1663859327
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1663859327
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1663859327
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1663859327
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1663859327
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1663859327
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1663859327
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1663859327
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1663859327
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1663859327
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1663859327
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1663859327
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1663859327
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1663859327
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1663859327
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1663859327
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1663859327
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1663859327
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1663859327
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1663859327
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1663859327
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1663859327
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1663859327
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1663859327
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1663859327
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1663859327
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1663859327
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1663859327
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1663859327
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1663859327
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1663859327
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1663859327
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1663859327
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1663859327
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1663859327
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1663859327
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1663859327
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1663859327
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1663859327
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1663859327
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1663859327
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1663859327
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1663859327
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1663859327
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1663859327
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1663859327
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1663859327
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1663859327
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1663859327
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1663859327
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1663859327
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1663859327
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1663859327
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1663859327
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1663859327
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1663859327
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1663859327
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1663859327
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1663859327
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1663859327
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1663859327
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1663859327
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1663859327
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1663859327
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1663859327
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1663859327
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1663859327
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1663859327
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1663859327
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1663859327
transform 1 0 350400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1663859327
transform 1 0 354400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1663859327
transform 1 0 358400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1663859327
transform 1 0 362400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1663859327
transform 1 0 366400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1663859327
transform 1 0 370400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1663859327
transform 1 0 374400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1663859327
transform 1 0 378400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_94
timestamp 1663859327
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1663859327
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1663859327
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1663859327
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1663859327
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1663859327
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1663859327
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1663859327
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1663859327
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1663859327
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1663859327
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1663859327
transform 1 0 431800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1663859327
transform 1 0 435800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1663859327
transform 1 0 439800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1663859327
transform 1 0 443800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1663859327
transform 1 0 447800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1663859327
transform 1 0 451800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1663859327
transform 1 0 455800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1663859327
transform 1 0 459800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1663859327
transform 1 0 463800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1663859327
transform 1 0 467800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_116
timestamp 1663859327
transform 1 0 471800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1663859327
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1663859327
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1663859327
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1663859327
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1663859327
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1663859327
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1663859327
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1663859327
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_126
timestamp 1663859327
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_127
timestamp 1663859327
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_128
timestamp 1663859327
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_129
timestamp 1663859327
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1663859327
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1663859327
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1663859327
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1663859327
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1663859327
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1663859327
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1663859327
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1663859327
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_139
timestamp 1663859327
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_140
timestamp 1663859327
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1663859327
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_142
timestamp 1663859327
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1663859327
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1663859327
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1663859327
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1663859327
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1663859327
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_149
timestamp 1663859327
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1663859327
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1663859327
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_152
timestamp 1663859327
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_153
timestamp 1663859327
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1663859327
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1663859327
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1663859327
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1663859327
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1663859327
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_160
timestamp 1663859327
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1663859327
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1663859327
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1663859327
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1663859327
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_165
timestamp 1663859327
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_166
timestamp 1663859327
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1663859327
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1663859327
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1663859327
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1663859327
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_171
timestamp 1663859327
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_172
timestamp 1663859327
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1663859327
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1663859327
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_181
timestamp 1663859327
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_182
timestamp 1663859327
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_183
timestamp 1663859327
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1663859327
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1663859327
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1663859327
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_188
timestamp 1663859327
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_189
timestamp 1663859327
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1663859327
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1663859327
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1663859327
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_199
timestamp 1663859327
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_200
timestamp 1663859327
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1663859327
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1663859327
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1663859327
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_205
timestamp 1663859327
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_206
timestamp 1663859327
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1663859327
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1663859327
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1663859327
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_216
timestamp 1663859327
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_217
timestamp 1663859327
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1663859327
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1663859327
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1663859327
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_222
timestamp 1663859327
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_223
timestamp 1663859327
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1663859327
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1663859327
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1663859327
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_233
timestamp 1663859327
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_234
timestamp 1663859327
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1663859327
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1663859327
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1663859327
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1663859327
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_240
timestamp 1663859327
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1663859327
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1663859327
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1663859327
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_250
timestamp 1663859327
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_251
timestamp 1663859327
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1663859327
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1663859327
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_255
timestamp 1663859327
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_256
timestamp 1663859327
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_257
timestamp 1663859327
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1663859327
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1663859327
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1663859327
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_267
timestamp 1663859327
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_268
timestamp 1663859327
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1663859327
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1663859327
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1663859327
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_273
timestamp 1663859327
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_274
timestamp 1663859327
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1663859327
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1663859327
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1663859327
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1663859327
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_285
timestamp 1663859327
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1663859327
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1663859327
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_289
timestamp 1663859327
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_290
timestamp 1663859327
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_291
timestamp 1663859327
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1663859327
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1663859327
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_300
timestamp 1663859327
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_301
timestamp 1663859327
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_302
timestamp 1663859327
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1663859327
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1663859327
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1663859327
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_307
timestamp 1663859327
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_308
timestamp 1663859327
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1663859327
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1663859327
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1663859327
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_318
timestamp 1663859327
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_319
timestamp 1663859327
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1663859327
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1663859327
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1663859327
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_324
timestamp 1663859327
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_325
timestamp 1663859327
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1663859327
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1663859327
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1663859327
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_335
timestamp 1663859327
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_336
timestamp 1663859327
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1663859327
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1663859327
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1663859327
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_341
timestamp 1663859327
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_342
timestamp 1663859327
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1663859327
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1663859327
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1663859327
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_352
timestamp 1663859327
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_353
timestamp 1663859327
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1663859327
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1663859327
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1663859327
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1663859327
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1663859327
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1663859327
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1663859327
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1663859327
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_369
timestamp 1663859327
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_370
timestamp 1663859327
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1663859327
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1663859327
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1663859327
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1663859327
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1663859327
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1663859327
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1663859327
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1663859327
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1663859327
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_380
timestamp 1663859327
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_381
timestamp 1663859327
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_382
timestamp 1663859327
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1663859327
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1663859327
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1663859327
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_387
timestamp 1663859327
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1663859327
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1663859327
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_390
timestamp 1663859327
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_391
timestamp 1663859327
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_392
timestamp 1663859327
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1663859327
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1663859327
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1663859327
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_397
timestamp 1663859327
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_398
timestamp 1663859327
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1663859327
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_400
timestamp 1663859327
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_401
timestamp 1663859327
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_402
timestamp 1663859327
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1663859327
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1663859327
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_407
timestamp 1663859327
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_408
timestamp 1663859327
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_409
timestamp 1663859327
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1663859327
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_411
timestamp 1663859327
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_412
timestamp 1663859327
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_413
timestamp 1663859327
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1663859327
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1663859327
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1663859327
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_418
timestamp 1663859327
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_419
timestamp 1663859327
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1663859327
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_421
timestamp 1663859327
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_422
timestamp 1663859327
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_423
timestamp 1663859327
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1663859327
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1663859327
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1663859327
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_428
timestamp 1663859327
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_429
timestamp 1663859327
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_430
timestamp 1663859327
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_431
timestamp 1663859327
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_432
timestamp 1663859327
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_433
timestamp 1663859327
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1663859327
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1663859327
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1663859327
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_438
timestamp 1663859327
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_439
timestamp 1663859327
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1663859327
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_441
timestamp 1663859327
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_442
timestamp 1663859327
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1663859327
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1663859327
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1663859327
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1663859327
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1663859327
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_449
timestamp 1663859327
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1663859327
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_451
timestamp 1663859327
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_452
timestamp 1663859327
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_453
timestamp 1663859327
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1663859327
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1663859327
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1663859327
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1663859327
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_459
timestamp 1663859327
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1663859327
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_461
timestamp 1663859327
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_462
timestamp 1663859327
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_463
timestamp 1663859327
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1663859327
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1663859327
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1663859327
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_468
timestamp 1663859327
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1663859327
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1663859327
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_471
timestamp 1663859327
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_472
timestamp 1663859327
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_473
timestamp 1663859327
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1663859327
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1663859327
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1663859327
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_478
timestamp 1663859327
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_479
timestamp 1663859327
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_480
timestamp 1663859327
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_481
timestamp 1663859327
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_482
timestamp 1663859327
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_483
timestamp 1663859327
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1663859327
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1663859327
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1663859327
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_488
timestamp 1663859327
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_489
timestamp 1663859327
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_490
timestamp 1663859327
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_491
timestamp 1663859327
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_492
timestamp 1663859327
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1663859327
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1663859327
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1663859327
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1663859327
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1663859327
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1663859327
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_500
timestamp 1663859327
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_501
timestamp 1663859327
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_502
timestamp 1663859327
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1663859327
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1663859327
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1663859327
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1663859327
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1663859327
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1663859327
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1663859327
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_511
timestamp 1663859327
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_512
timestamp 1663859327
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1663859327
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1663859327
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1663859327
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1663859327
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1663859327
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1663859327
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1663859327
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_521
timestamp 1663859327
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_522
timestamp 1663859327
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1663859327
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1663859327
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1663859327
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1663859327
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_528
timestamp 1663859327
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_529
timestamp 1663859327
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1663859327
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_531
timestamp 1663859327
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_532
timestamp 1663859327
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_533
timestamp 1663859327
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1663859327
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1663859327
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1663859327
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_538
timestamp 1663859327
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_539
timestamp 1663859327
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_540
timestamp 1663859327
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_541
timestamp 1663859327
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_542
timestamp 1663859327
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_543
timestamp 1663859327
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1663859327
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1663859327
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1663859327
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1663859327
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1663859327
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_550
timestamp 1663859327
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_551
timestamp 1663859327
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_552
timestamp 1663859327
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1663859327
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1663859327
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1663859327
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1663859327
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_558
timestamp 1663859327
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1663859327
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1663859327
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_561
timestamp 1663859327
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_562
timestamp 1663859327
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_563
timestamp 1663859327
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1663859327
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1663859327
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1663859327
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_568
timestamp 1663859327
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_569
timestamp 1663859327
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1663859327
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_571
timestamp 1663859327
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_572
timestamp 1663859327
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_573
timestamp 1663859327
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1663859327
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1663859327
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1663859327
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_578
timestamp 1663859327
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_579
timestamp 1663859327
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1663859327
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_581
timestamp 1663859327
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_582
timestamp 1663859327
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_583
timestamp 1663859327
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1663859327
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1663859327
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1663859327
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1663859327
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_589
timestamp 1663859327
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1663859327
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_591
timestamp 1663859327
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_592
timestamp 1663859327
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1663859327
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1663859327
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1663859327
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1663859327
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1663859327
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1663859327
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1663859327
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_601
timestamp 1663859327
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_602
timestamp 1663859327
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_603
timestamp 1663859327
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_604
timestamp 1663859327
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1663859327
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1663859327
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1663859327
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1663859327
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1663859327
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1663859327
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1663859327
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_612
timestamp 1663859327
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1663859327
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1663859327
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1663859327
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1663859327
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1663859327
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1663859327
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1663859327
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_622
timestamp 1663859327
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1663859327
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1663859327
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1663859327
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1663859327
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1663859327
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1663859327
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1663859327
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_631
timestamp 1663859327
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1663859327
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1663859327
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1663859327
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1663859327
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1663859327
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1663859327
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1663859327
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1663859327
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_641
timestamp 1663859327
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1663859327
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1663859327
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1663859327
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1663859327
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1663859327
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1663859327
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1663859327
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_650
timestamp 1663859327
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_651
timestamp 1663859327
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1663859327
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1663859327
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1663859327
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1663859327
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1663859327
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1663859327
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1663859327
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_660
timestamp 1663859327
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1663859327
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1663859327
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1663859327
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1663859327
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1663859327
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1663859327
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1663859327
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_669
timestamp 1663859327
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1663859327
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1663859327
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1663859327
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1663859327
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1663859327
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1663859327
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1663859327
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_678
timestamp 1663859327
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_679
timestamp 1663859327
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1663859327
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1663859327
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1663859327
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1663859327
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1663859327
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1663859327
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1663859327
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_688
timestamp 1663859327
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1663859327
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1663859327
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1663859327
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1663859327
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1663859327
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1663859327
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1663859327
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_697
timestamp 1663859327
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1663859327
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1663859327
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1663859327
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1663859327
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1663859327
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1663859327
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1663859327
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1663859327
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_707
timestamp 1663859327
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1663859327
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1663859327
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1663859327
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1663859327
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1663859327
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1663859327
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1663859327
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_716
timestamp 1663859327
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1663859327
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1663859327
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1663859327
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1663859327
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1663859327
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1663859327
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1663859327
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_725
timestamp 1663859327
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_726
timestamp 1663859327
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1663859327
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1663859327
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1663859327
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1663859327
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1663859327
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1663859327
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1663859327
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_735
timestamp 1663859327
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1663859327
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1663859327
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1663859327
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1663859327
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1663859327
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1663859327
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1663859327
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_744
timestamp 1663859327
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_745
timestamp 1663859327
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1663859327
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1663859327
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1663859327
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1663859327
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1663859327
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1663859327
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1663859327
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_754
timestamp 1663859327
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1663859327
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1663859327
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1663859327
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1663859327
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1663859327
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1663859327
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1663859327
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_763
timestamp 1663859327
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1663859327
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1663859327
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1663859327
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1663859327
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1663859327
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1663859327
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1663859327
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_772
timestamp 1663859327
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_773
timestamp 1663859327
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1663859327
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1663859327
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1663859327
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1663859327
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1663859327
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1663859327
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1663859327
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_782
timestamp 1663859327
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1663859327
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1663859327
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1663859327
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1663859327
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1663859327
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_789
timestamp 1663859327
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_790
timestamp 1663859327
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_791
timestamp 1663859327
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_792
timestamp 1663859327
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1663859327
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1663859327
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1663859327
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1663859327
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_798
timestamp 1663859327
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_799
timestamp 1663859327
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_800
timestamp 1663859327
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_801
timestamp 1663859327
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1663859327
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1663859327
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1663859327
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1663859327
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1663859327
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_808
timestamp 1663859327
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_809
timestamp 1663859327
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_810
timestamp 1663859327
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_811
timestamp 1663859327
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB1
timestamp 1663859327
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB2
timestamp 1663859327
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB3
timestamp 1663859327
transform 1 0 349400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1663859327
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1663859327
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1663859327
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1663859327
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1663859327
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1663859327
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1663859327
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1663859327
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1663859327
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1663859327
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1663859327
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1663859327
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1663859327
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1663859327
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1663859327
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1663859327
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1663859327
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1663859327
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1663859327
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1663859327
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1663859327
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1663859327
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1663859327
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1663859327
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1663859327
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1663859327
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1663859327
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1663859327
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1663859327
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1663859327
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1663859327
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1663859327
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1663859327
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1663859327
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1663859327
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1663859327
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1663859327
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1663859327
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1663859327
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1663859327
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1663859327
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1663859327
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1663859327
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1663859327
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1663859327
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1663859327
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1663859327
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1663859327
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1663859327
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1663859327
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1663859327
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1663859327
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1663859327
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1663859327
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1663859327
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1663859327
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1663859327
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1663859327
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1663859327
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1663859327
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1663859327
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1663859327
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1663859327
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1663859327
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1663859327
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1663859327
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1663859327
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1663859327
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1663859327
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1663859327
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1663859327
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use chip_io_gpio_connects  chip_io_gpio_connects_0
timestamp 1665248140
transform 1 0 0 0 1 0
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_1
timestamp 1665248140
transform 1 0 0 0 1 45200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_2
timestamp 1665248140
transform 1 0 0 0 1 90200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_3
timestamp 1665248140
transform 1 0 0 0 1 135400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_4
timestamp 1665248140
transform 1 0 0 0 1 180400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_5
timestamp 1665248140
transform 1 0 0 0 1 225400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_6
timestamp 1665248140
transform 1 0 0 0 1 270600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_7
timestamp 1665248140
transform 1 0 0 0 1 447800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_8
timestamp 1665248140
transform 1 0 0 0 1 493000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_9
timestamp 1665248140
transform 1 0 0 0 1 538000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_10
timestamp 1665248140
transform 1 0 0 0 1 583200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_11
timestamp 1665248140
transform 1 0 0 0 1 628200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_12
timestamp 1665248140
transform 1 0 0 0 1 673200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_13
timestamp 1665248140
transform 1 0 0 0 1 762400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_14
timestamp 1665248140
transform 1 0 0 0 1 851600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_15
timestamp 1665248140
transform -1 0 717600 0 -1 297600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_16
timestamp 1665248140
transform 0 -1 742000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_17
timestamp 1665248140
transform 0 -1 640200 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_18
timestamp 1665248140
transform 0 -1 588800 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_19
timestamp 1665248140
transform 0 -1 499800 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_21
timestamp 1665248140
transform 0 -1 398000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_22
timestamp 1665248140
transform 0 -1 346400 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_23
timestamp 1665248140
transform 0 -1 295000 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_24
timestamp 1665248140
transform 0 -1 243600 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_25
timestamp 1665248140
transform 0 -1 192200 1 0 320000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_26
timestamp 1665248140
transform -1 0 717600 0 -1 1070200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_27
timestamp 1665248140
transform -1 0 717600 0 -1 900400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_28
timestamp 1665248140
transform -1 0 717600 0 -1 857200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_29
timestamp 1665248140
transform -1 0 717600 0 -1 814000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_30
timestamp 1665248140
transform -1 0 717600 0 -1 770800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_31
timestamp 1665248140
transform -1 0 717600 0 -1 727600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_32
timestamp 1665248140
transform -1 0 717600 0 -1 684400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_33
timestamp 1665248140
transform -1 0 717600 0 -1 641200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_34
timestamp 1665248140
transform -1 0 717600 0 -1 513600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_35
timestamp 1665248140
transform -1 0 717600 0 -1 470400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_36
timestamp 1665248140
transform -1 0 717600 0 -1 427200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_37
timestamp 1665248140
transform -1 0 717600 0 -1 384000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_38
timestamp 1665248140
transform -1 0 717600 0 -1 340800
box 675407 99896 675887 115709
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 202400 0 -1 42193
box -32 0 16032 42193
use constant_block  constant_block_0
timestamp 1665259416
transform -1 0 151016 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_1
timestamp 1665259416
transform -1 0 205816 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_2
timestamp 1665259416
transform -1 0 315416 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_3
timestamp 1665259416
transform -1 0 370216 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_4
timestamp 1665259416
transform -1 0 425016 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_5
timestamp 1665259416
transform -1 0 479816 0 1 39452
box 0 496 2800 2224
use constant_block  constant_block_6
timestamp 1665259416
transform -1 0 534616 0 1 39452
box 0 496 2800 2224
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 348400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1663859327
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1663859327
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1663859327
transform -1 0 365800 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1663859327
transform -1 0 311000 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1663859327
transform -1 0 420600 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1663859327
transform -1 0 475400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1663859327
transform -1 0 530200 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1663859327
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1663859327
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1663859327
transform 0 1 675407 -1 0 116000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1663859327
transform 0 1 675407 -1 0 161200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1663859327
transform 0 1 675407 -1 0 206200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1663859327
transform 0 1 675407 -1 0 251400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1663859327
transform 0 1 675407 -1 0 296400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1663859327
transform 0 1 675407 -1 0 341400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1663859327
transform 0 1 675407 -1 0 386600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1663859327
transform 0 1 675407 -1 0 563800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1663859327
transform 0 1 675407 -1 0 609000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1663859327
transform 0 1 675407 -1 0 654000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1663859327
transform 0 1 675407 -1 0 699200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1663859327
transform 0 1 675407 -1 0 744200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1663859327
transform 0 1 675407 -1 0 789200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1663859327
transform 0 1 675407 -1 0 878400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1663859327
transform 0 1 675407 -1 0 967600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1663859327
transform 1 0 626000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1663859327
transform 1 0 524200 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1663859327
transform 1 0 472800 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[18\]
timestamp 1663859327
transform 1 0 383800 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1663859327
transform 1 0 282000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1663859327
transform 1 0 230400 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1663859327
transform 1 0 179000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1663859327
transform 1 0 127600 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1663859327
transform 1 0 76200 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1663859327
transform 0 -1 42193 1 0 954200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1663859327
transform 0 -1 42193 1 0 784400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1663859327
transform 0 -1 42193 1 0 741200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1663859327
transform 0 -1 42193 1 0 698000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1663859327
transform 0 -1 42193 1 0 654800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1663859327
transform 0 -1 42193 1 0 611600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1663859327
transform 0 -1 42193 1 0 568400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1663859327
transform 0 -1 42193 1 0 525200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1663859327
transform 0 -1 42193 1 0 397600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1663859327
transform 0 -1 42193 1 0 354400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1663859327
transform 0 -1 42193 1 0 311200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1663859327
transform 0 -1 42193 1 0 268000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1663859327
transform 0 -1 42193 1 0 224800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1663859327
transform 0 -1 42193 1 0 181600
box -32 0 16032 42193
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__corner_pad  user1_corner
timestamp 1663859327
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user1_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 1 678007 -1 0 922600
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1663859327
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1663859327
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user1_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 1 678007 -1 0 474800
box 0 -2177 17187 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1663859327
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user2_vccd_lvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 912000
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user2_vssd_lvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 440800
box 0 -2177 17187 39593
<< labels >>
flabel metal5 s 187640 6598 200180 19088 6 FreeSans 320 0 0 0 clock
port 0 nsew signal input
flabel metal2 s 187327 41713 187383 42193 0 FreeSans 320 90 0 0 clock_core
port 1 nsew signal tristate
flabel metal2 s 194043 41713 194099 42193 0 FreeSans 320 90 0 0 por
port 2 nsew signal input
flabel metal5 s 351040 6598 363580 19088 6 FreeSans 320 0 0 0 flash_clk
port 3 nsew signal tristate
flabel metal2 s 361767 41713 361823 42193 0 FreeSans 320 90 0 0 flash_clk_core
port 4 nsew signal input
flabel metal2 s 364895 41713 364951 42193 0 FreeSans 320 90 0 0 flash_clk_oeb_core
port 6 nsew signal input
flabel metal5 s 296240 6598 308780 19088 6 FreeSans 320 0 0 0 flash_csb
port 7 nsew signal tristate
flabel metal2 s 306967 41713 307023 42193 0 FreeSans 320 90 0 0 flash_csb_core
port 8 nsew signal input
flabel metal2 s 310095 41713 310151 42193 0 FreeSans 320 90 0 0 flash_csb_oeb_core
port 10 nsew signal input
flabel metal5 s 405840 6598 418380 19088 6 FreeSans 320 0 0 0 flash_io0
port 11 nsew signal bidirectional
flabel metal2 s 405527 41713 405583 42193 0 FreeSans 320 90 0 0 flash_io0_di_core
port 12 nsew signal tristate
flabel metal2 s 416567 41713 416623 42193 0 FreeSans 320 90 0 0 flash_io0_do_core
port 13 nsew signal input
flabel metal2 s 412243 41713 412299 42193 0 FreeSans 320 90 0 0 flash_io0_ieb_core
port 14 nsew signal input
flabel metal2 s 419695 41713 419751 42193 0 FreeSans 320 90 0 0 flash_io0_oeb_core
port 15 nsew signal input
flabel metal5 s 460640 6598 473180 19088 6 FreeSans 320 0 0 0 flash_io1
port 16 nsew signal bidirectional
flabel metal2 s 460327 41713 460383 42193 0 FreeSans 320 90 0 0 flash_io1_di_core
port 17 nsew signal tristate
flabel metal2 s 471367 41713 471423 42193 0 FreeSans 320 90 0 0 flash_io1_do_core
port 18 nsew signal input
flabel metal2 s 474495 41713 474551 42193 0 FreeSans 320 90 0 0 flash_io1_oeb_core
port 20 nsew signal input
flabel metal5 s 515440 6598 527980 19088 6 FreeSans 320 0 0 0 gpio
port 21 nsew signal bidirectional
flabel metal2 s 515127 41713 515183 42193 0 FreeSans 320 90 0 0 gpio_in_core
port 22 nsew signal tristate
flabel metal2 s 521843 41713 521899 42193 0 FreeSans 320 90 0 0 gpio_inenb_core
port 23 nsew signal input
flabel metal2 s 520647 41713 520703 42193 0 FreeSans 320 90 0 0 gpio_mode0_core
port 24 nsew signal input
flabel metal2 s 524971 41713 525027 42193 0 FreeSans 320 90 0 0 gpio_mode1_core
port 25 nsew signal input
flabel metal2 s 526167 41713 526223 42193 0 FreeSans 320 90 0 0 gpio_out_core
port 26 nsew signal input
flabel metal2 s 529295 41713 529351 42193 0 FreeSans 320 90 0 0 gpio_outenb_core
port 27 nsew signal input
flabel metal5 s 6167 70054 19619 80934 6 FreeSans 320 0 0 0 vccd_pad
port 28 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 6 FreeSans 320 0 0 0 vdda_pad
port 29 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 6 FreeSans 320 0 0 0 vddio_pad
port 30 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 6 FreeSans 320 0 0 0 vddio_pad2
port 31 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 6 FreeSans 320 0 0 0 vssa_pad
port 32 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 6 FreeSans 320 0 0 0 vssd_pad
port 33 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 6 FreeSans 320 0 0 0 vssio_pad
port 34 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 6 FreeSans 320 0 0 0 vssio_pad2
port 35 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 6 FreeSans 320 0 0 0 mprj_io[0]
port 36 nsew signal bidirectional
flabel metal2 s 675407 105803 675887 105859 0 FreeSans 320 0 0 0 mprj_io_analog_en[0]
port 37 nsew signal input
flabel metal2 s 675407 107091 675887 107147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[0]
port 38 nsew signal input
flabel metal2 s 675407 110127 675887 110183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[0]
port 39 nsew signal input
flabel metal2 s 675407 106447 675887 106503 0 FreeSans 320 0 0 0 mprj_io_dm[0]
port 40 nsew signal input
flabel metal2 s 675407 104607 675887 104663 0 FreeSans 320 0 0 0 mprj_io_dm[1]
port 41 nsew signal input
flabel metal2 s 675407 110771 675887 110827 0 FreeSans 320 0 0 0 mprj_io_dm[2]
port 42 nsew signal input
flabel metal2 s 675407 111415 675887 111471 0 FreeSans 320 0 0 0 mprj_io_holdover[0]
port 43 nsew signal input
flabel metal2 s 675407 114451 675887 114507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
flabel metal2 s 675407 107643 675887 107699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[0]
port 45 nsew signal input
flabel metal2 s 675407 115095 675887 115151 0 FreeSans 320 0 0 0 mprj_io_oeb[0]
port 46 nsew signal input
flabel metal2 s 675407 111967 675887 112023 0 FreeSans 320 0 0 0 mprj_io_out[0]
port 47 nsew signal input
flabel metal2 s 675407 102767 675887 102823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[0]
port 48 nsew signal input
flabel metal2 s 675407 113807 675887 113863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[0]
port 49 nsew signal input
flabel metal2 s 675407 100927 675887 100983 0 FreeSans 320 0 0 0 mprj_io_in[0]
port 50 nsew signal tristate
flabel metal2 s 675407 686611 675887 686667 0 FreeSans 320 0 0 0 mprj_analog_io[3]
port 51 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 6 FreeSans 320 0 0 0 mprj_io[10]
port 52 nsew signal bidirectional
flabel metal2 s 675407 689003 675887 689059 0 FreeSans 320 0 0 0 mprj_io_analog_en[10]
port 53 nsew signal input
flabel metal2 s 675407 690291 675887 690347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[10]
port 54 nsew signal input
flabel metal2 s 675407 693327 675887 693383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[10]
port 55 nsew signal input
flabel metal2 s 675407 689647 675887 689703 0 FreeSans 320 0 0 0 mprj_io_dm[30]
port 56 nsew signal input
flabel metal2 s 675407 687807 675887 687863 0 FreeSans 320 0 0 0 mprj_io_dm[31]
port 57 nsew signal input
flabel metal2 s 675407 693971 675887 694027 0 FreeSans 320 0 0 0 mprj_io_dm[32]
port 58 nsew signal input
flabel metal2 s 675407 694615 675887 694671 0 FreeSans 320 0 0 0 mprj_io_holdover[10]
port 59 nsew signal input
flabel metal2 s 675407 697651 675887 697707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[10]
port 60 nsew signal input
flabel metal2 s 675407 690843 675887 690899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[10]
port 61 nsew signal input
flabel metal2 s 675407 698295 675887 698351 0 FreeSans 320 0 0 0 mprj_io_oeb[10]
port 62 nsew signal input
flabel metal2 s 675407 695167 675887 695223 0 FreeSans 320 0 0 0 mprj_io_out[10]
port 63 nsew signal input
flabel metal2 s 675407 685967 675887 686023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[10]
port 64 nsew signal input
flabel metal2 s 675407 697007 675887 697063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[10]
port 65 nsew signal input
flabel metal2 s 675407 684127 675887 684183 0 FreeSans 320 0 0 0 mprj_io_in[10]
port 66 nsew signal tristate
flabel metal2 s 675407 731611 675887 731667 0 FreeSans 320 0 0 0 mprj_analog_io[4]
port 67 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 6 FreeSans 320 0 0 0 mprj_io[11]
port 68 nsew signal bidirectional
flabel metal2 s 675407 734003 675887 734059 0 FreeSans 320 0 0 0 mprj_io_analog_en[11]
port 69 nsew signal input
flabel metal2 s 675407 735291 675887 735347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[11]
port 70 nsew signal input
flabel metal2 s 675407 738327 675887 738383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[11]
port 71 nsew signal input
flabel metal2 s 675407 734647 675887 734703 0 FreeSans 320 0 0 0 mprj_io_dm[33]
port 72 nsew signal input
flabel metal2 s 675407 732807 675887 732863 0 FreeSans 320 0 0 0 mprj_io_dm[34]
port 73 nsew signal input
flabel metal2 s 675407 738971 675887 739027 0 FreeSans 320 0 0 0 mprj_io_dm[35]
port 74 nsew signal input
flabel metal2 s 675407 739615 675887 739671 0 FreeSans 320 0 0 0 mprj_io_holdover[11]
port 75 nsew signal input
flabel metal2 s 675407 742651 675887 742707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[11]
port 76 nsew signal input
flabel metal2 s 675407 735843 675887 735899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[11]
port 77 nsew signal input
flabel metal2 s 675407 743295 675887 743351 0 FreeSans 320 0 0 0 mprj_io_oeb[11]
port 78 nsew signal input
flabel metal2 s 675407 740167 675887 740223 0 FreeSans 320 0 0 0 mprj_io_out[11]
port 79 nsew signal input
flabel metal2 s 675407 730967 675887 731023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[11]
port 80 nsew signal input
flabel metal2 s 675407 742007 675887 742063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[11]
port 81 nsew signal input
flabel metal2 s 675407 729127 675887 729183 0 FreeSans 320 0 0 0 mprj_io_in[11]
port 82 nsew signal tristate
flabel metal2 s 675407 776611 675887 776667 0 FreeSans 320 0 0 0 mprj_analog_io[5]
port 83 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 6 FreeSans 320 0 0 0 mprj_io[12]
port 84 nsew signal bidirectional
flabel metal2 s 675407 779003 675887 779059 0 FreeSans 320 0 0 0 mprj_io_analog_en[12]
port 85 nsew signal input
flabel metal2 s 675407 780291 675887 780347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[12]
port 86 nsew signal input
flabel metal2 s 675407 783327 675887 783383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[12]
port 87 nsew signal input
flabel metal2 s 675407 779647 675887 779703 0 FreeSans 320 0 0 0 mprj_io_dm[36]
port 88 nsew signal input
flabel metal2 s 675407 777807 675887 777863 0 FreeSans 320 0 0 0 mprj_io_dm[37]
port 89 nsew signal input
flabel metal2 s 675407 783971 675887 784027 0 FreeSans 320 0 0 0 mprj_io_dm[38]
port 90 nsew signal input
flabel metal2 s 675407 784615 675887 784671 0 FreeSans 320 0 0 0 mprj_io_holdover[12]
port 91 nsew signal input
flabel metal2 s 675407 787651 675887 787707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[12]
port 92 nsew signal input
flabel metal2 s 675407 780843 675887 780899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[12]
port 93 nsew signal input
flabel metal2 s 675407 788295 675887 788351 0 FreeSans 320 0 0 0 mprj_io_oeb[12]
port 94 nsew signal input
flabel metal2 s 675407 785167 675887 785223 0 FreeSans 320 0 0 0 mprj_io_out[12]
port 95 nsew signal input
flabel metal2 s 675407 775967 675887 776023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[12]
port 96 nsew signal input
flabel metal2 s 675407 787007 675887 787063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[12]
port 97 nsew signal input
flabel metal2 s 675407 774127 675887 774183 0 FreeSans 320 0 0 0 mprj_io_in[12]
port 98 nsew signal tristate
flabel metal2 s 675407 865811 675887 865867 0 FreeSans 320 0 0 0 mprj_analog_io[6]
port 99 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 6 FreeSans 320 0 0 0 mprj_io[13]
port 100 nsew signal bidirectional
flabel metal2 s 675407 868203 675887 868259 0 FreeSans 320 0 0 0 mprj_io_analog_en[13]
port 101 nsew signal input
flabel metal2 s 675407 869491 675887 869547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[13]
port 102 nsew signal input
flabel metal2 s 675407 872527 675887 872583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[13]
port 103 nsew signal input
flabel metal2 s 675407 868847 675887 868903 0 FreeSans 320 0 0 0 mprj_io_dm[39]
port 104 nsew signal input
flabel metal2 s 675407 867007 675887 867063 0 FreeSans 320 0 0 0 mprj_io_dm[40]
port 105 nsew signal input
flabel metal2 s 675407 873171 675887 873227 0 FreeSans 320 0 0 0 mprj_io_dm[41]
port 106 nsew signal input
flabel metal2 s 675407 873815 675887 873871 0 FreeSans 320 0 0 0 mprj_io_holdover[13]
port 107 nsew signal input
flabel metal2 s 675407 876851 675887 876907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[13]
port 108 nsew signal input
flabel metal2 s 675407 870043 675887 870099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[13]
port 109 nsew signal input
flabel metal2 s 675407 877495 675887 877551 0 FreeSans 320 0 0 0 mprj_io_oeb[13]
port 110 nsew signal input
flabel metal2 s 675407 874367 675887 874423 0 FreeSans 320 0 0 0 mprj_io_out[13]
port 111 nsew signal input
flabel metal2 s 675407 865167 675887 865223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[13]
port 112 nsew signal input
flabel metal2 s 675407 876207 675887 876263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[13]
port 113 nsew signal input
flabel metal2 s 675407 863327 675887 863383 0 FreeSans 320 0 0 0 mprj_io_in[13]
port 114 nsew signal tristate
flabel metal2 s 675407 955011 675887 955067 0 FreeSans 320 0 0 0 mprj_analog_io[7]
port 115 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965380 6 FreeSans 320 0 0 0 mprj_io[14]
port 116 nsew signal bidirectional
flabel metal2 s 675407 957403 675887 957459 0 FreeSans 320 0 0 0 mprj_io_analog_en[14]
port 117 nsew signal input
flabel metal2 s 675407 958691 675887 958747 0 FreeSans 320 0 0 0 mprj_io_analog_pol[14]
port 118 nsew signal input
flabel metal2 s 675407 961727 675887 961783 0 FreeSans 320 0 0 0 mprj_io_analog_sel[14]
port 119 nsew signal input
flabel metal2 s 675407 958047 675887 958103 0 FreeSans 320 0 0 0 mprj_io_dm[42]
port 120 nsew signal input
flabel metal2 s 675407 956207 675887 956263 0 FreeSans 320 0 0 0 mprj_io_dm[43]
port 121 nsew signal input
flabel metal2 s 675407 962371 675887 962427 0 FreeSans 320 0 0 0 mprj_io_dm[44]
port 122 nsew signal input
flabel metal2 s 675407 963015 675887 963071 0 FreeSans 320 0 0 0 mprj_io_holdover[14]
port 123 nsew signal input
flabel metal2 s 675407 966051 675887 966107 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[14]
port 124 nsew signal input
flabel metal2 s 675407 959243 675887 959299 0 FreeSans 320 0 0 0 mprj_io_inp_dis[14]
port 125 nsew signal input
flabel metal2 s 675407 966695 675887 966751 0 FreeSans 320 0 0 0 mprj_io_oeb[14]
port 126 nsew signal input
flabel metal2 s 675407 963567 675887 963623 0 FreeSans 320 0 0 0 mprj_io_out[14]
port 127 nsew signal input
flabel metal2 s 675407 954367 675887 954423 0 FreeSans 320 0 0 0 mprj_io_slow_sel[14]
port 128 nsew signal input
flabel metal2 s 675407 965407 675887 965463 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[14]
port 129 nsew signal input
flabel metal2 s 675407 952527 675887 952583 0 FreeSans 320 0 0 0 mprj_io_in[14]
port 130 nsew signal tristate
flabel metal2 s 638533 995407 638589 995887 0 FreeSans 320 90 0 0 mprj_analog_io[8]
port 131 nsew signal bidirectional
flabel metal5 s 628220 1018512 640760 1031002 6 FreeSans 320 0 0 0 mprj_io[15]
port 132 nsew signal bidirectional
flabel metal2 s 636141 995407 636197 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[15]
port 133 nsew signal input
flabel metal2 s 634853 995407 634909 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[15]
port 134 nsew signal input
flabel metal2 s 631817 995407 631873 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[15]
port 135 nsew signal input
flabel metal2 s 635497 995407 635553 995887 0 FreeSans 320 90 0 0 mprj_io_dm[45]
port 136 nsew signal input
flabel metal2 s 637337 995407 637393 995887 0 FreeSans 320 90 0 0 mprj_io_dm[46]
port 137 nsew signal input
flabel metal2 s 631173 995407 631229 995887 0 FreeSans 320 90 0 0 mprj_io_dm[47]
port 138 nsew signal input
flabel metal2 s 630529 995407 630585 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[15]
port 139 nsew signal input
flabel metal2 s 627493 995407 627549 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[15]
port 140 nsew signal input
flabel metal2 s 634301 995407 634357 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[15]
port 141 nsew signal input
flabel metal2 s 626849 995407 626905 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[15]
port 142 nsew signal input
flabel metal2 s 629977 995407 630033 995887 0 FreeSans 320 90 0 0 mprj_io_out[15]
port 143 nsew signal input
flabel metal2 s 639177 995407 639233 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[15]
port 144 nsew signal input
flabel metal2 s 628137 995407 628193 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[15]
port 145 nsew signal input
flabel metal2 s 641017 995407 641073 995887 0 FreeSans 320 90 0 0 mprj_io_in[15]
port 146 nsew signal tristate
flabel metal2 s 536733 995407 536789 995887 0 FreeSans 320 90 0 0 mprj_analog_io[9]
port 147 nsew signal bidirectional
flabel metal5 s 526420 1018512 538960 1031002 6 FreeSans 320 0 0 0 mprj_io[16]
port 148 nsew signal bidirectional
flabel metal2 s 534341 995407 534397 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[16]
port 149 nsew signal input
flabel metal2 s 533053 995407 533109 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[16]
port 150 nsew signal input
flabel metal2 s 530017 995407 530073 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[16]
port 151 nsew signal input
flabel metal2 s 533697 995407 533753 995887 0 FreeSans 320 90 0 0 mprj_io_dm[48]
port 152 nsew signal input
flabel metal2 s 535537 995407 535593 995887 0 FreeSans 320 90 0 0 mprj_io_dm[49]
port 153 nsew signal input
flabel metal2 s 529373 995407 529429 995887 0 FreeSans 320 90 0 0 mprj_io_dm[50]
port 154 nsew signal input
flabel metal2 s 528729 995407 528785 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[16]
port 155 nsew signal input
flabel metal2 s 525693 995407 525749 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[16]
port 156 nsew signal input
flabel metal2 s 532501 995407 532557 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[16]
port 157 nsew signal input
flabel metal2 s 525049 995407 525105 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[16]
port 158 nsew signal input
flabel metal2 s 528177 995407 528233 995887 0 FreeSans 320 90 0 0 mprj_io_out[16]
port 159 nsew signal input
flabel metal2 s 537377 995407 537433 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[16]
port 160 nsew signal input
flabel metal2 s 526337 995407 526393 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[16]
port 161 nsew signal input
flabel metal2 s 539217 995407 539273 995887 0 FreeSans 320 90 0 0 mprj_io_in[16]
port 162 nsew signal tristate
flabel metal2 s 485333 995407 485389 995887 0 FreeSans 320 90 0 0 mprj_analog_io[10]
port 163 nsew signal bidirectional
flabel metal5 s 475020 1018512 487560 1031002 6 FreeSans 320 0 0 0 mprj_io[17]
port 164 nsew signal bidirectional
flabel metal2 s 482941 995407 482997 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[17]
port 165 nsew signal input
flabel metal2 s 481653 995407 481709 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[17]
port 166 nsew signal input
flabel metal2 s 478617 995407 478673 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[17]
port 167 nsew signal input
flabel metal2 s 482297 995407 482353 995887 0 FreeSans 320 90 0 0 mprj_io_dm[51]
port 168 nsew signal input
flabel metal2 s 484137 995407 484193 995887 0 FreeSans 320 90 0 0 mprj_io_dm[52]
port 169 nsew signal input
flabel metal2 s 477973 995407 478029 995887 0 FreeSans 320 90 0 0 mprj_io_dm[53]
port 170 nsew signal input
flabel metal2 s 477329 995407 477385 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[17]
port 171 nsew signal input
flabel metal2 s 474293 995407 474349 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[17]
port 172 nsew signal input
flabel metal2 s 481101 995407 481157 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[17]
port 173 nsew signal input
flabel metal2 s 473649 995407 473705 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[17]
port 174 nsew signal input
flabel metal2 s 476777 995407 476833 995887 0 FreeSans 320 90 0 0 mprj_io_out[17]
port 175 nsew signal input
flabel metal2 s 485977 995407 486033 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[17]
port 176 nsew signal input
flabel metal2 s 474937 995407 474993 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[17]
port 177 nsew signal input
flabel metal2 s 487817 995407 487873 995887 0 FreeSans 320 90 0 0 mprj_io_in[17]
port 178 nsew signal tristate
flabel metal2 s 396333 995407 396389 995887 0 FreeSans 320 90 0 0 mprj_analog_io[11]
port 179 nsew signal bidirectional
flabel metal5 s 386020 1018512 398560 1031002 6 FreeSans 320 0 0 0 mprj_io[18]
port 180 nsew signal bidirectional
flabel metal2 s 393941 995407 393997 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[18]
port 181 nsew signal input
flabel metal2 s 392653 995407 392709 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[18]
port 182 nsew signal input
flabel metal2 s 389617 995407 389673 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[18]
port 183 nsew signal input
flabel metal2 s 393297 995407 393353 995887 0 FreeSans 320 90 0 0 mprj_io_dm[54]
port 184 nsew signal input
flabel metal2 s 395137 995407 395193 995887 0 FreeSans 320 90 0 0 mprj_io_dm[55]
port 185 nsew signal input
flabel metal2 s 388973 995407 389029 995887 0 FreeSans 320 90 0 0 mprj_io_dm[56]
port 186 nsew signal input
flabel metal2 s 388329 995407 388385 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[18]
port 187 nsew signal input
flabel metal2 s 385293 995407 385349 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[18]
port 188 nsew signal input
flabel metal2 s 392101 995407 392157 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[18]
port 189 nsew signal input
flabel metal2 s 384649 995407 384705 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[18]
port 190 nsew signal input
flabel metal2 s 387777 995407 387833 995887 0 FreeSans 320 90 0 0 mprj_io_out[18]
port 191 nsew signal input
flabel metal2 s 396977 995407 397033 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[18]
port 192 nsew signal input
flabel metal2 s 385937 995407 385993 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[18]
port 193 nsew signal input
flabel metal2 s 398817 995407 398873 995887 0 FreeSans 320 90 0 0 mprj_io_in[18]
port 194 nsew signal tristate
flabel metal5 s 698512 146440 711002 158980 6 FreeSans 320 0 0 0 mprj_io[1]
port 195 nsew signal bidirectional
flabel metal2 s 675407 151003 675887 151059 0 FreeSans 320 0 0 0 mprj_io_analog_en[1]
port 196 nsew signal input
flabel metal2 s 675407 152291 675887 152347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[1]
port 197 nsew signal input
flabel metal2 s 675407 155327 675887 155383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[1]
port 198 nsew signal input
flabel metal2 s 675407 151647 675887 151703 0 FreeSans 320 0 0 0 mprj_io_dm[3]
port 199 nsew signal input
flabel metal2 s 675407 149807 675887 149863 0 FreeSans 320 0 0 0 mprj_io_dm[4]
port 200 nsew signal input
flabel metal2 s 675407 155971 675887 156027 0 FreeSans 320 0 0 0 mprj_io_dm[5]
port 201 nsew signal input
flabel metal2 s 675407 156615 675887 156671 0 FreeSans 320 0 0 0 mprj_io_holdover[1]
port 202 nsew signal input
flabel metal2 s 675407 159651 675887 159707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[1]
port 203 nsew signal input
flabel metal2 s 675407 152843 675887 152899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[1]
port 204 nsew signal input
flabel metal2 s 675407 160295 675887 160351 0 FreeSans 320 0 0 0 mprj_io_oeb[1]
port 205 nsew signal input
flabel metal2 s 675407 157167 675887 157223 0 FreeSans 320 0 0 0 mprj_io_out[1]
port 206 nsew signal input
flabel metal2 s 675407 147967 675887 148023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[1]
port 207 nsew signal input
flabel metal2 s 675407 159007 675887 159063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[1]
port 208 nsew signal input
flabel metal2 s 675407 146127 675887 146183 0 FreeSans 320 0 0 0 mprj_io_in[1]
port 209 nsew signal tristate
flabel metal5 s 698512 191440 711002 203980 6 FreeSans 320 0 0 0 mprj_io[2]
port 210 nsew signal bidirectional
flabel metal2 s 675407 196003 675887 196059 0 FreeSans 320 0 0 0 mprj_io_analog_en[2]
port 211 nsew signal input
flabel metal2 s 675407 197291 675887 197347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[2]
port 212 nsew signal input
flabel metal2 s 675407 200327 675887 200383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[2]
port 213 nsew signal input
flabel metal2 s 675407 196647 675887 196703 0 FreeSans 320 0 0 0 mprj_io_dm[6]
port 214 nsew signal input
flabel metal2 s 675407 194807 675887 194863 0 FreeSans 320 0 0 0 mprj_io_dm[7]
port 215 nsew signal input
flabel metal2 s 675407 200971 675887 201027 0 FreeSans 320 0 0 0 mprj_io_dm[8]
port 216 nsew signal input
flabel metal2 s 675407 201615 675887 201671 0 FreeSans 320 0 0 0 mprj_io_holdover[2]
port 217 nsew signal input
flabel metal2 s 675407 204651 675887 204707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[2]
port 218 nsew signal input
flabel metal2 s 675407 197843 675887 197899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[2]
port 219 nsew signal input
flabel metal2 s 675407 205295 675887 205351 0 FreeSans 320 0 0 0 mprj_io_oeb[2]
port 220 nsew signal input
flabel metal2 s 675407 202167 675887 202223 0 FreeSans 320 0 0 0 mprj_io_out[2]
port 221 nsew signal input
flabel metal2 s 675407 192967 675887 193023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[2]
port 222 nsew signal input
flabel metal2 s 675407 204007 675887 204063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[2]
port 223 nsew signal input
flabel metal2 s 675407 191127 675887 191183 0 FreeSans 320 0 0 0 mprj_io_in[2]
port 224 nsew signal tristate
flabel metal5 s 698512 236640 711002 249180 6 FreeSans 320 0 0 0 mprj_io[3]
port 225 nsew signal bidirectional
flabel metal2 s 675407 241203 675887 241259 0 FreeSans 320 0 0 0 mprj_io_analog_en[3]
port 226 nsew signal input
flabel metal2 s 675407 242491 675887 242547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[3]
port 227 nsew signal input
flabel metal2 s 675407 245527 675887 245583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[3]
port 228 nsew signal input
flabel metal2 s 675407 240007 675887 240063 0 FreeSans 320 0 0 0 mprj_io_dm[10]
port 229 nsew signal input
flabel metal2 s 675407 246171 675887 246227 0 FreeSans 320 0 0 0 mprj_io_dm[11]
port 230 nsew signal input
flabel metal2 s 675407 241847 675887 241903 0 FreeSans 320 0 0 0 mprj_io_dm[9]
port 231 nsew signal input
flabel metal2 s 675407 246815 675887 246871 0 FreeSans 320 0 0 0 mprj_io_holdover[3]
port 232 nsew signal input
flabel metal2 s 675407 249851 675887 249907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[3]
port 233 nsew signal input
flabel metal2 s 675407 243043 675887 243099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[3]
port 234 nsew signal input
flabel metal2 s 675407 250495 675887 250551 0 FreeSans 320 0 0 0 mprj_io_oeb[3]
port 235 nsew signal input
flabel metal2 s 675407 247367 675887 247423 0 FreeSans 320 0 0 0 mprj_io_out[3]
port 236 nsew signal input
flabel metal2 s 675407 238167 675887 238223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[3]
port 237 nsew signal input
flabel metal2 s 675407 249207 675887 249263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[3]
port 238 nsew signal input
flabel metal2 s 675407 236327 675887 236383 0 FreeSans 320 0 0 0 mprj_io_in[3]
port 239 nsew signal tristate
flabel metal5 s 698512 281640 711002 294180 6 FreeSans 320 0 0 0 mprj_io[4]
port 240 nsew signal bidirectional
flabel metal2 s 675407 286203 675887 286259 0 FreeSans 320 0 0 0 mprj_io_analog_en[4]
port 241 nsew signal input
flabel metal2 s 675407 287491 675887 287547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[4]
port 242 nsew signal input
flabel metal2 s 675407 290527 675887 290583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[4]
port 243 nsew signal input
flabel metal2 s 675407 286847 675887 286903 0 FreeSans 320 0 0 0 mprj_io_dm[12]
port 244 nsew signal input
flabel metal2 s 675407 285007 675887 285063 0 FreeSans 320 0 0 0 mprj_io_dm[13]
port 245 nsew signal input
flabel metal2 s 675407 291171 675887 291227 0 FreeSans 320 0 0 0 mprj_io_dm[14]
port 246 nsew signal input
flabel metal2 s 675407 291815 675887 291871 0 FreeSans 320 0 0 0 mprj_io_holdover[4]
port 247 nsew signal input
flabel metal2 s 675407 294851 675887 294907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[4]
port 248 nsew signal input
flabel metal2 s 675407 288043 675887 288099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[4]
port 249 nsew signal input
flabel metal2 s 675407 295495 675887 295551 0 FreeSans 320 0 0 0 mprj_io_oeb[4]
port 250 nsew signal input
flabel metal2 s 675407 292367 675887 292423 0 FreeSans 320 0 0 0 mprj_io_out[4]
port 251 nsew signal input
flabel metal2 s 675407 283167 675887 283223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[4]
port 252 nsew signal input
flabel metal2 s 675407 294207 675887 294263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[4]
port 253 nsew signal input
flabel metal2 s 675407 281327 675887 281383 0 FreeSans 320 0 0 0 mprj_io_in[4]
port 254 nsew signal tristate
flabel metal5 s 698512 326640 711002 339180 6 FreeSans 320 0 0 0 mprj_io[5]
port 255 nsew signal bidirectional
flabel metal2 s 675407 331203 675887 331259 0 FreeSans 320 0 0 0 mprj_io_analog_en[5]
port 256 nsew signal input
flabel metal2 s 675407 332491 675887 332547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[5]
port 257 nsew signal input
flabel metal2 s 675407 335527 675887 335583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[5]
port 258 nsew signal input
flabel metal2 s 675407 331847 675887 331903 0 FreeSans 320 0 0 0 mprj_io_dm[15]
port 259 nsew signal input
flabel metal2 s 675407 330007 675887 330063 0 FreeSans 320 0 0 0 mprj_io_dm[16]
port 260 nsew signal input
flabel metal2 s 675407 336171 675887 336227 0 FreeSans 320 0 0 0 mprj_io_dm[17]
port 261 nsew signal input
flabel metal2 s 675407 336815 675887 336871 0 FreeSans 320 0 0 0 mprj_io_holdover[5]
port 262 nsew signal input
flabel metal2 s 675407 339851 675887 339907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[5]
port 263 nsew signal input
flabel metal2 s 675407 333043 675887 333099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[5]
port 264 nsew signal input
flabel metal2 s 675407 340495 675887 340551 0 FreeSans 320 0 0 0 mprj_io_oeb[5]
port 265 nsew signal input
flabel metal2 s 675407 337367 675887 337423 0 FreeSans 320 0 0 0 mprj_io_out[5]
port 266 nsew signal input
flabel metal2 s 675407 328167 675887 328223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[5]
port 267 nsew signal input
flabel metal2 s 675407 339207 675887 339263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[5]
port 268 nsew signal input
flabel metal2 s 675407 326327 675887 326383 0 FreeSans 320 0 0 0 mprj_io_in[5]
port 269 nsew signal tristate
flabel metal5 s 698512 371840 711002 384380 6 FreeSans 320 0 0 0 mprj_io[6]
port 270 nsew signal bidirectional
flabel metal2 s 675407 376403 675887 376459 0 FreeSans 320 0 0 0 mprj_io_analog_en[6]
port 271 nsew signal input
flabel metal2 s 675407 377691 675887 377747 0 FreeSans 320 0 0 0 mprj_io_analog_pol[6]
port 272 nsew signal input
flabel metal2 s 675407 380727 675887 380783 0 FreeSans 320 0 0 0 mprj_io_analog_sel[6]
port 273 nsew signal input
flabel metal2 s 675407 377047 675887 377103 0 FreeSans 320 0 0 0 mprj_io_dm[18]
port 274 nsew signal input
flabel metal2 s 675407 375207 675887 375263 0 FreeSans 320 0 0 0 mprj_io_dm[19]
port 275 nsew signal input
flabel metal2 s 675407 381371 675887 381427 0 FreeSans 320 0 0 0 mprj_io_dm[20]
port 276 nsew signal input
flabel metal2 s 675407 382015 675887 382071 0 FreeSans 320 0 0 0 mprj_io_holdover[6]
port 277 nsew signal input
flabel metal2 s 675407 385051 675887 385107 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[6]
port 278 nsew signal input
flabel metal2 s 675407 378243 675887 378299 0 FreeSans 320 0 0 0 mprj_io_inp_dis[6]
port 279 nsew signal input
flabel metal2 s 675407 385695 675887 385751 0 FreeSans 320 0 0 0 mprj_io_oeb[6]
port 280 nsew signal input
flabel metal2 s 675407 382567 675887 382623 0 FreeSans 320 0 0 0 mprj_io_out[6]
port 281 nsew signal input
flabel metal2 s 675407 373367 675887 373423 0 FreeSans 320 0 0 0 mprj_io_slow_sel[6]
port 282 nsew signal input
flabel metal2 s 675407 384407 675887 384463 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[6]
port 283 nsew signal input
flabel metal2 s 675407 371527 675887 371583 0 FreeSans 320 0 0 0 mprj_io_in[6]
port 284 nsew signal tristate
flabel metal2 s 675407 551211 675887 551267 0 FreeSans 320 0 0 0 mprj_analog_io[0]
port 285 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 6 FreeSans 320 0 0 0 mprj_io[7]
port 286 nsew signal bidirectional
flabel metal2 s 675407 553603 675887 553659 0 FreeSans 320 0 0 0 mprj_io_analog_en[7]
port 287 nsew signal input
flabel metal2 s 675407 554891 675887 554947 0 FreeSans 320 0 0 0 mprj_io_analog_pol[7]
port 288 nsew signal input
flabel metal2 s 675407 557927 675887 557983 0 FreeSans 320 0 0 0 mprj_io_analog_sel[7]
port 289 nsew signal input
flabel metal2 s 675407 554247 675887 554303 0 FreeSans 320 0 0 0 mprj_io_dm[21]
port 290 nsew signal input
flabel metal2 s 675407 552407 675887 552463 0 FreeSans 320 0 0 0 mprj_io_dm[22]
port 291 nsew signal input
flabel metal2 s 675407 558571 675887 558627 0 FreeSans 320 0 0 0 mprj_io_dm[23]
port 292 nsew signal input
flabel metal2 s 675407 559215 675887 559271 0 FreeSans 320 0 0 0 mprj_io_holdover[7]
port 293 nsew signal input
flabel metal2 s 675407 562251 675887 562307 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[7]
port 294 nsew signal input
flabel metal2 s 675407 555443 675887 555499 0 FreeSans 320 0 0 0 mprj_io_inp_dis[7]
port 295 nsew signal input
flabel metal2 s 675407 562895 675887 562951 0 FreeSans 320 0 0 0 mprj_io_oeb[7]
port 296 nsew signal input
flabel metal2 s 675407 559767 675887 559823 0 FreeSans 320 0 0 0 mprj_io_out[7]
port 297 nsew signal input
flabel metal2 s 675407 550567 675887 550623 0 FreeSans 320 0 0 0 mprj_io_slow_sel[7]
port 298 nsew signal input
flabel metal2 s 675407 561607 675887 561663 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[7]
port 299 nsew signal input
flabel metal2 s 675407 548727 675887 548783 0 FreeSans 320 0 0 0 mprj_io_in[7]
port 300 nsew signal tristate
flabel metal2 s 675407 596411 675887 596467 0 FreeSans 320 0 0 0 mprj_analog_io[1]
port 301 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 6 FreeSans 320 0 0 0 mprj_io[8]
port 302 nsew signal bidirectional
flabel metal2 s 675407 598803 675887 598859 0 FreeSans 320 0 0 0 mprj_io_analog_en[8]
port 303 nsew signal input
flabel metal2 s 675407 600091 675887 600147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[8]
port 304 nsew signal input
flabel metal2 s 675407 603127 675887 603183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[8]
port 305 nsew signal input
flabel metal2 s 675407 599447 675887 599503 0 FreeSans 320 0 0 0 mprj_io_dm[24]
port 306 nsew signal input
flabel metal2 s 675407 597607 675887 597663 0 FreeSans 320 0 0 0 mprj_io_dm[25]
port 307 nsew signal input
flabel metal2 s 675407 603771 675887 603827 0 FreeSans 320 0 0 0 mprj_io_dm[26]
port 308 nsew signal input
flabel metal2 s 675407 604415 675887 604471 0 FreeSans 320 0 0 0 mprj_io_holdover[8]
port 309 nsew signal input
flabel metal2 s 675407 607451 675887 607507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[8]
port 310 nsew signal input
flabel metal2 s 675407 600643 675887 600699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[8]
port 311 nsew signal input
flabel metal2 s 675407 608095 675887 608151 0 FreeSans 320 0 0 0 mprj_io_oeb[8]
port 312 nsew signal input
flabel metal2 s 675407 604967 675887 605023 0 FreeSans 320 0 0 0 mprj_io_out[8]
port 313 nsew signal input
flabel metal2 s 675407 595767 675887 595823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[8]
port 314 nsew signal input
flabel metal2 s 675407 606807 675887 606863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[8]
port 315 nsew signal input
flabel metal2 s 675407 593927 675887 593983 0 FreeSans 320 0 0 0 mprj_io_in[8]
port 316 nsew signal tristate
flabel metal2 s 675407 641411 675887 641467 0 FreeSans 320 0 0 0 mprj_analog_io[2]
port 317 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 6 FreeSans 320 0 0 0 mprj_io[9]
port 318 nsew signal bidirectional
flabel metal2 s 675407 643803 675887 643859 0 FreeSans 320 0 0 0 mprj_io_analog_en[9]
port 319 nsew signal input
flabel metal2 s 675407 645091 675887 645147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[9]
port 320 nsew signal input
flabel metal2 s 675407 648127 675887 648183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[9]
port 321 nsew signal input
flabel metal2 s 675407 644447 675887 644503 0 FreeSans 320 0 0 0 mprj_io_dm[27]
port 322 nsew signal input
flabel metal2 s 675407 642607 675887 642663 0 FreeSans 320 0 0 0 mprj_io_dm[28]
port 323 nsew signal input
flabel metal2 s 675407 648771 675887 648827 0 FreeSans 320 0 0 0 mprj_io_dm[29]
port 324 nsew signal input
flabel metal2 s 675407 649415 675887 649471 0 FreeSans 320 0 0 0 mprj_io_holdover[9]
port 325 nsew signal input
flabel metal2 s 675407 652451 675887 652507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[9]
port 326 nsew signal input
flabel metal2 s 675407 645643 675887 645699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[9]
port 327 nsew signal input
flabel metal2 s 675407 653095 675887 653151 0 FreeSans 320 0 0 0 mprj_io_oeb[9]
port 328 nsew signal input
flabel metal2 s 675407 649967 675887 650023 0 FreeSans 320 0 0 0 mprj_io_out[9]
port 329 nsew signal input
flabel metal2 s 675407 640767 675887 640823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[9]
port 330 nsew signal input
flabel metal2 s 675407 651807 675887 651863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[9]
port 331 nsew signal input
flabel metal2 s 675407 638927 675887 638983 0 FreeSans 320 0 0 0 mprj_io_in[9]
port 332 nsew signal tristate
flabel metal2 s 294533 995407 294589 995887 0 FreeSans 320 90 0 0 mprj_analog_io[12]
port 333 nsew signal bidirectional
flabel metal5 s 284220 1018512 296760 1031002 6 FreeSans 320 0 0 0 mprj_io[19]
port 334 nsew signal bidirectional
flabel metal2 s 292141 995407 292197 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[19]
port 335 nsew signal input
flabel metal2 s 290853 995407 290909 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[19]
port 336 nsew signal input
flabel metal2 s 287817 995407 287873 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[19]
port 337 nsew signal input
flabel metal2 s 291497 995407 291553 995887 0 FreeSans 320 90 0 0 mprj_io_dm[57]
port 338 nsew signal input
flabel metal2 s 293337 995407 293393 995887 0 FreeSans 320 90 0 0 mprj_io_dm[58]
port 339 nsew signal input
flabel metal2 s 287173 995407 287229 995887 0 FreeSans 320 90 0 0 mprj_io_dm[59]
port 340 nsew signal input
flabel metal2 s 286529 995407 286585 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[19]
port 341 nsew signal input
flabel metal2 s 283493 995407 283549 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[19]
port 342 nsew signal input
flabel metal2 s 290301 995407 290357 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[19]
port 343 nsew signal input
flabel metal2 s 282849 995407 282905 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[19]
port 344 nsew signal input
flabel metal2 s 285977 995407 286033 995887 0 FreeSans 320 90 0 0 mprj_io_out[19]
port 345 nsew signal input
flabel metal2 s 295177 995407 295233 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[19]
port 346 nsew signal input
flabel metal2 s 284137 995407 284193 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[19]
port 347 nsew signal input
flabel metal2 s 297017 995407 297073 995887 0 FreeSans 320 90 0 0 mprj_io_in[19]
port 348 nsew signal tristate
flabel metal2 s 41713 624133 42193 624189 0 FreeSans 320 0 0 0 mprj_analog_io[22]
port 349 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 6 FreeSans 320 0 0 0 mprj_io[29]
port 350 nsew signal bidirectional
flabel metal2 s 41713 621741 42193 621797 0 FreeSans 320 0 0 0 mprj_io_analog_en[29]
port 351 nsew signal input
flabel metal2 s 41713 620453 42193 620509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[29]
port 352 nsew signal input
flabel metal2 s 41713 617417 42193 617473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[29]
port 353 nsew signal input
flabel metal2 s 41713 621097 42193 621153 0 FreeSans 320 0 0 0 mprj_io_dm[87]
port 354 nsew signal input
flabel metal2 s 41713 622937 42193 622993 0 FreeSans 320 0 0 0 mprj_io_dm[88]
port 355 nsew signal input
flabel metal2 s 41713 616773 42193 616829 0 FreeSans 320 0 0 0 mprj_io_dm[89]
port 356 nsew signal input
flabel metal2 s 41713 616129 42193 616185 0 FreeSans 320 0 0 0 mprj_io_holdover[29]
port 357 nsew signal input
flabel metal2 s 41713 613093 42193 613149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[29]
port 358 nsew signal input
flabel metal2 s 41713 619901 42193 619957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[29]
port 359 nsew signal input
flabel metal2 s 41713 612449 42193 612505 0 FreeSans 320 0 0 0 mprj_io_oeb[29]
port 360 nsew signal input
flabel metal2 s 41713 615577 42193 615633 0 FreeSans 320 0 0 0 mprj_io_out[29]
port 361 nsew signal input
flabel metal2 s 41713 624777 42193 624833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[29]
port 362 nsew signal input
flabel metal2 s 41713 613737 42193 613793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[29]
port 363 nsew signal input
flabel metal2 s 41713 626617 42193 626673 0 FreeSans 320 0 0 0 mprj_io_in[29]
port 364 nsew signal tristate
flabel metal2 s 41713 580933 42193 580989 0 FreeSans 320 0 0 0 mprj_analog_io[23]
port 365 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 6 FreeSans 320 0 0 0 mprj_io[30]
port 366 nsew signal bidirectional
flabel metal2 s 41713 578541 42193 578597 0 FreeSans 320 0 0 0 mprj_io_analog_en[30]
port 367 nsew signal input
flabel metal2 s 41713 577253 42193 577309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[30]
port 368 nsew signal input
flabel metal2 s 41713 574217 42193 574273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[30]
port 369 nsew signal input
flabel metal2 s 41713 577897 42193 577953 0 FreeSans 320 0 0 0 mprj_io_dm[90]
port 370 nsew signal input
flabel metal2 s 41713 579737 42193 579793 0 FreeSans 320 0 0 0 mprj_io_dm[91]
port 371 nsew signal input
flabel metal2 s 41713 573573 42193 573629 0 FreeSans 320 0 0 0 mprj_io_dm[92]
port 372 nsew signal input
flabel metal2 s 41713 572929 42193 572985 0 FreeSans 320 0 0 0 mprj_io_holdover[30]
port 373 nsew signal input
flabel metal2 s 41713 569893 42193 569949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[30]
port 374 nsew signal input
flabel metal2 s 41713 576701 42193 576757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[30]
port 375 nsew signal input
flabel metal2 s 41713 569249 42193 569305 0 FreeSans 320 0 0 0 mprj_io_oeb[30]
port 376 nsew signal input
flabel metal2 s 41713 572377 42193 572433 0 FreeSans 320 0 0 0 mprj_io_out[30]
port 377 nsew signal input
flabel metal2 s 41713 581577 42193 581633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[30]
port 378 nsew signal input
flabel metal2 s 41713 570537 42193 570593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[30]
port 379 nsew signal input
flabel metal2 s 41713 583417 42193 583473 0 FreeSans 320 0 0 0 mprj_io_in[30]
port 380 nsew signal tristate
flabel metal2 s 41713 537733 42193 537789 0 FreeSans 320 0 0 0 mprj_analog_io[24]
port 381 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 6 FreeSans 320 0 0 0 mprj_io[31]
port 382 nsew signal bidirectional
flabel metal2 s 41713 535341 42193 535397 0 FreeSans 320 0 0 0 mprj_io_analog_en[31]
port 383 nsew signal input
flabel metal2 s 41713 534053 42193 534109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[31]
port 384 nsew signal input
flabel metal2 s 41713 531017 42193 531073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[31]
port 385 nsew signal input
flabel metal2 s 41713 534697 42193 534753 0 FreeSans 320 0 0 0 mprj_io_dm[93]
port 386 nsew signal input
flabel metal2 s 41713 536537 42193 536593 0 FreeSans 320 0 0 0 mprj_io_dm[94]
port 387 nsew signal input
flabel metal2 s 41713 530373 42193 530429 0 FreeSans 320 0 0 0 mprj_io_dm[95]
port 388 nsew signal input
flabel metal2 s 41713 529729 42193 529785 0 FreeSans 320 0 0 0 mprj_io_holdover[31]
port 389 nsew signal input
flabel metal2 s 41713 526693 42193 526749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[31]
port 390 nsew signal input
flabel metal2 s 41713 533501 42193 533557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[31]
port 391 nsew signal input
flabel metal2 s 41713 526049 42193 526105 0 FreeSans 320 0 0 0 mprj_io_oeb[31]
port 392 nsew signal input
flabel metal2 s 41713 529177 42193 529233 0 FreeSans 320 0 0 0 mprj_io_out[31]
port 393 nsew signal input
flabel metal2 s 41713 538377 42193 538433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[31]
port 394 nsew signal input
flabel metal2 s 41713 527337 42193 527393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[31]
port 395 nsew signal input
flabel metal2 s 41713 540217 42193 540273 0 FreeSans 320 0 0 0 mprj_io_in[31]
port 396 nsew signal tristate
flabel metal2 s 41713 410133 42193 410189 0 FreeSans 320 0 0 0 mprj_analog_io[25]
port 397 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 6 FreeSans 320 0 0 0 mprj_io[32]
port 398 nsew signal bidirectional
flabel metal2 s 41713 407741 42193 407797 0 FreeSans 320 0 0 0 mprj_io_analog_en[32]
port 399 nsew signal input
flabel metal2 s 41713 406453 42193 406509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[32]
port 400 nsew signal input
flabel metal2 s 41713 403417 42193 403473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[32]
port 401 nsew signal input
flabel metal2 s 41713 407097 42193 407153 0 FreeSans 320 0 0 0 mprj_io_dm[96]
port 402 nsew signal input
flabel metal2 s 41713 408937 42193 408993 0 FreeSans 320 0 0 0 mprj_io_dm[97]
port 403 nsew signal input
flabel metal2 s 41713 402773 42193 402829 0 FreeSans 320 0 0 0 mprj_io_dm[98]
port 404 nsew signal input
flabel metal2 s 41713 402129 42193 402185 0 FreeSans 320 0 0 0 mprj_io_holdover[32]
port 405 nsew signal input
flabel metal2 s 41713 399093 42193 399149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[32]
port 406 nsew signal input
flabel metal2 s 41713 405901 42193 405957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[32]
port 407 nsew signal input
flabel metal2 s 41713 398449 42193 398505 0 FreeSans 320 0 0 0 mprj_io_oeb[32]
port 408 nsew signal input
flabel metal2 s 41713 401577 42193 401633 0 FreeSans 320 0 0 0 mprj_io_out[32]
port 409 nsew signal input
flabel metal2 s 41713 410777 42193 410833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[32]
port 410 nsew signal input
flabel metal2 s 41713 399737 42193 399793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[32]
port 411 nsew signal input
flabel metal2 s 41713 412617 42193 412673 0 FreeSans 320 0 0 0 mprj_io_in[32]
port 412 nsew signal tristate
flabel metal2 s 41713 366933 42193 366989 0 FreeSans 320 0 0 0 mprj_analog_io[26]
port 413 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 6 FreeSans 320 0 0 0 mprj_io[33]
port 414 nsew signal bidirectional
flabel metal2 s 41713 364541 42193 364597 0 FreeSans 320 0 0 0 mprj_io_analog_en[33]
port 415 nsew signal input
flabel metal2 s 41713 363253 42193 363309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[33]
port 416 nsew signal input
flabel metal2 s 41713 360217 42193 360273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[33]
port 417 nsew signal input
flabel metal2 s 41713 365737 42193 365793 0 FreeSans 320 0 0 0 mprj_io_dm[100]
port 418 nsew signal input
flabel metal2 s 41713 359573 42193 359629 0 FreeSans 320 0 0 0 mprj_io_dm[101]
port 419 nsew signal input
flabel metal2 s 41713 363897 42193 363953 0 FreeSans 320 0 0 0 mprj_io_dm[99]
port 420 nsew signal input
flabel metal2 s 41713 358929 42193 358985 0 FreeSans 320 0 0 0 mprj_io_holdover[33]
port 421 nsew signal input
flabel metal2 s 41713 355893 42193 355949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[33]
port 422 nsew signal input
flabel metal2 s 41713 362701 42193 362757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[33]
port 423 nsew signal input
flabel metal2 s 41713 355249 42193 355305 0 FreeSans 320 0 0 0 mprj_io_oeb[33]
port 424 nsew signal input
flabel metal2 s 41713 358377 42193 358433 0 FreeSans 320 0 0 0 mprj_io_out[33]
port 425 nsew signal input
flabel metal2 s 41713 367577 42193 367633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[33]
port 426 nsew signal input
flabel metal2 s 41713 356537 42193 356593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[33]
port 427 nsew signal input
flabel metal2 s 41713 369417 42193 369473 0 FreeSans 320 0 0 0 mprj_io_in[33]
port 428 nsew signal tristate
flabel metal2 s 41713 323733 42193 323789 0 FreeSans 320 0 0 0 mprj_analog_io[27]
port 429 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 6 FreeSans 320 0 0 0 mprj_io[34]
port 430 nsew signal bidirectional
flabel metal2 s 41713 321341 42193 321397 0 FreeSans 320 0 0 0 mprj_io_analog_en[34]
port 431 nsew signal input
flabel metal2 s 41713 320053 42193 320109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[34]
port 432 nsew signal input
flabel metal2 s 41713 317017 42193 317073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[34]
port 433 nsew signal input
flabel metal2 s 41713 320697 42193 320753 0 FreeSans 320 0 0 0 mprj_io_dm[102]
port 434 nsew signal input
flabel metal2 s 41713 322537 42193 322593 0 FreeSans 320 0 0 0 mprj_io_dm[103]
port 435 nsew signal input
flabel metal2 s 41713 316373 42193 316429 0 FreeSans 320 0 0 0 mprj_io_dm[104]
port 436 nsew signal input
flabel metal2 s 41713 315729 42193 315785 0 FreeSans 320 0 0 0 mprj_io_holdover[34]
port 437 nsew signal input
flabel metal2 s 41713 312693 42193 312749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[34]
port 438 nsew signal input
flabel metal2 s 41713 319501 42193 319557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[34]
port 439 nsew signal input
flabel metal2 s 41713 312049 42193 312105 0 FreeSans 320 0 0 0 mprj_io_oeb[34]
port 440 nsew signal input
flabel metal2 s 41713 315177 42193 315233 0 FreeSans 320 0 0 0 mprj_io_out[34]
port 441 nsew signal input
flabel metal2 s 41713 324377 42193 324433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[34]
port 442 nsew signal input
flabel metal2 s 41713 313337 42193 313393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[34]
port 443 nsew signal input
flabel metal2 s 41713 326217 42193 326273 0 FreeSans 320 0 0 0 mprj_io_in[34]
port 444 nsew signal tristate
flabel metal2 s 41713 280533 42193 280589 0 FreeSans 320 0 0 0 mprj_analog_io[28]
port 445 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 6 FreeSans 320 0 0 0 mprj_io[35]
port 446 nsew signal bidirectional
flabel metal2 s 41713 278141 42193 278197 0 FreeSans 320 0 0 0 mprj_io_analog_en[35]
port 447 nsew signal input
flabel metal2 s 41713 276853 42193 276909 0 FreeSans 320 0 0 0 mprj_io_analog_pol[35]
port 448 nsew signal input
flabel metal2 s 41713 273817 42193 273873 0 FreeSans 320 0 0 0 mprj_io_analog_sel[35]
port 449 nsew signal input
flabel metal2 s 41713 277497 42193 277553 0 FreeSans 320 0 0 0 mprj_io_dm[105]
port 450 nsew signal input
flabel metal2 s 41713 279337 42193 279393 0 FreeSans 320 0 0 0 mprj_io_dm[106]
port 451 nsew signal input
flabel metal2 s 41713 273173 42193 273229 0 FreeSans 320 0 0 0 mprj_io_dm[107]
port 452 nsew signal input
flabel metal2 s 41713 272529 42193 272585 0 FreeSans 320 0 0 0 mprj_io_holdover[35]
port 453 nsew signal input
flabel metal2 s 41713 269493 42193 269549 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[35]
port 454 nsew signal input
flabel metal2 s 41713 276301 42193 276357 0 FreeSans 320 0 0 0 mprj_io_inp_dis[35]
port 455 nsew signal input
flabel metal2 s 41713 268849 42193 268905 0 FreeSans 320 0 0 0 mprj_io_oeb[35]
port 456 nsew signal input
flabel metal2 s 41713 271977 42193 272033 0 FreeSans 320 0 0 0 mprj_io_out[35]
port 457 nsew signal input
flabel metal2 s 41713 281177 42193 281233 0 FreeSans 320 0 0 0 mprj_io_slow_sel[35]
port 458 nsew signal input
flabel metal2 s 41713 270137 42193 270193 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[35]
port 459 nsew signal input
flabel metal2 s 41713 283017 42193 283073 0 FreeSans 320 0 0 0 mprj_io_in[35]
port 460 nsew signal tristate
flabel metal5 s 6598 227020 19088 239560 6 FreeSans 320 0 0 0 mprj_io[36]
port 461 nsew signal bidirectional
flabel metal2 s 41713 234941 42193 234997 0 FreeSans 320 0 0 0 mprj_io_analog_en[36]
port 462 nsew signal input
flabel metal2 s 41713 233653 42193 233709 0 FreeSans 320 0 0 0 mprj_io_analog_pol[36]
port 463 nsew signal input
flabel metal2 s 41713 230617 42193 230673 0 FreeSans 320 0 0 0 mprj_io_analog_sel[36]
port 464 nsew signal input
flabel metal2 s 41713 234297 42193 234353 0 FreeSans 320 0 0 0 mprj_io_dm[108]
port 465 nsew signal input
flabel metal2 s 41713 236137 42193 236193 0 FreeSans 320 0 0 0 mprj_io_dm[109]
port 466 nsew signal input
flabel metal2 s 41713 229973 42193 230029 0 FreeSans 320 0 0 0 mprj_io_dm[110]
port 467 nsew signal input
flabel metal2 s 41713 229329 42193 229385 0 FreeSans 320 0 0 0 mprj_io_holdover[36]
port 468 nsew signal input
flabel metal2 s 41713 226293 42193 226349 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[36]
port 469 nsew signal input
flabel metal2 s 41713 233101 42193 233157 0 FreeSans 320 0 0 0 mprj_io_inp_dis[36]
port 470 nsew signal input
flabel metal2 s 41713 225649 42193 225705 0 FreeSans 320 0 0 0 mprj_io_oeb[36]
port 471 nsew signal input
flabel metal2 s 41713 228777 42193 228833 0 FreeSans 320 0 0 0 mprj_io_out[36]
port 472 nsew signal input
flabel metal2 s 41713 237977 42193 238033 0 FreeSans 320 0 0 0 mprj_io_slow_sel[36]
port 473 nsew signal input
flabel metal2 s 41713 226937 42193 226993 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[36]
port 474 nsew signal input
flabel metal2 s 41713 239817 42193 239873 0 FreeSans 320 0 0 0 mprj_io_in[36]
port 475 nsew signal tristate
flabel metal5 s 6598 183820 19088 196360 6 FreeSans 320 0 0 0 mprj_io[37]
port 476 nsew signal bidirectional
flabel metal2 s 41713 191741 42193 191797 0 FreeSans 320 0 0 0 mprj_io_analog_en[37]
port 477 nsew signal input
flabel metal2 s 41713 190453 42193 190509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[37]
port 478 nsew signal input
flabel metal2 s 41713 187417 42193 187473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[37]
port 479 nsew signal input
flabel metal2 s 41713 191097 42193 191153 0 FreeSans 320 0 0 0 mprj_io_dm[111]
port 480 nsew signal input
flabel metal2 s 41713 192937 42193 192993 0 FreeSans 320 0 0 0 mprj_io_dm[112]
port 481 nsew signal input
flabel metal2 s 41713 186773 42193 186829 0 FreeSans 320 0 0 0 mprj_io_dm[113]
port 482 nsew signal input
flabel metal2 s 41713 186129 42193 186185 0 FreeSans 320 0 0 0 mprj_io_holdover[37]
port 483 nsew signal input
flabel metal2 s 41713 183093 42193 183149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[37]
port 484 nsew signal input
flabel metal2 s 41713 189901 42193 189957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[37]
port 485 nsew signal input
flabel metal2 s 41713 182449 42193 182505 0 FreeSans 320 0 0 0 mprj_io_oeb[37]
port 486 nsew signal input
flabel metal2 s 41713 185577 42193 185633 0 FreeSans 320 0 0 0 mprj_io_out[37]
port 487 nsew signal input
flabel metal2 s 41713 194777 42193 194833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[37]
port 488 nsew signal input
flabel metal2 s 41713 183737 42193 183793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[37]
port 489 nsew signal input
flabel metal2 s 41713 196617 42193 196673 0 FreeSans 320 0 0 0 mprj_io_in[37]
port 490 nsew signal tristate
flabel metal2 s 242933 995407 242989 995887 0 FreeSans 320 90 0 0 mprj_analog_io[13]
port 491 nsew signal bidirectional
flabel metal5 s 232620 1018512 245160 1031002 6 FreeSans 320 0 0 0 mprj_io[20]
port 492 nsew signal bidirectional
flabel metal2 s 240541 995407 240597 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[20]
port 493 nsew signal input
flabel metal2 s 239253 995407 239309 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[20]
port 494 nsew signal input
flabel metal2 s 236217 995407 236273 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[20]
port 495 nsew signal input
flabel metal2 s 239897 995407 239953 995887 0 FreeSans 320 90 0 0 mprj_io_dm[60]
port 496 nsew signal input
flabel metal2 s 241737 995407 241793 995887 0 FreeSans 320 90 0 0 mprj_io_dm[61]
port 497 nsew signal input
flabel metal2 s 235573 995407 235629 995887 0 FreeSans 320 90 0 0 mprj_io_dm[62]
port 498 nsew signal input
flabel metal2 s 234929 995407 234985 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[20]
port 499 nsew signal input
flabel metal2 s 231893 995407 231949 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[20]
port 500 nsew signal input
flabel metal2 s 238701 995407 238757 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[20]
port 501 nsew signal input
flabel metal2 s 231249 995407 231305 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[20]
port 502 nsew signal input
flabel metal2 s 234377 995407 234433 995887 0 FreeSans 320 90 0 0 mprj_io_out[20]
port 503 nsew signal input
flabel metal2 s 243577 995407 243633 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[20]
port 504 nsew signal input
flabel metal2 s 232537 995407 232593 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[20]
port 505 nsew signal input
flabel metal2 s 245417 995407 245473 995887 0 FreeSans 320 90 0 0 mprj_io_in[20]
port 506 nsew signal tristate
flabel metal2 s 191533 995407 191589 995887 0 FreeSans 320 90 0 0 mprj_analog_io[14]
port 507 nsew signal bidirectional
flabel metal5 s 181220 1018512 193760 1031002 6 FreeSans 320 0 0 0 mprj_io[21]
port 508 nsew signal bidirectional
flabel metal2 s 189141 995407 189197 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[21]
port 509 nsew signal input
flabel metal2 s 187853 995407 187909 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[21]
port 510 nsew signal input
flabel metal2 s 184817 995407 184873 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[21]
port 511 nsew signal input
flabel metal2 s 188497 995407 188553 995887 0 FreeSans 320 90 0 0 mprj_io_dm[63]
port 512 nsew signal input
flabel metal2 s 190337 995407 190393 995887 0 FreeSans 320 90 0 0 mprj_io_dm[64]
port 513 nsew signal input
flabel metal2 s 184173 995407 184229 995887 0 FreeSans 320 90 0 0 mprj_io_dm[65]
port 514 nsew signal input
flabel metal2 s 183529 995407 183585 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[21]
port 515 nsew signal input
flabel metal2 s 180493 995407 180549 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[21]
port 516 nsew signal input
flabel metal2 s 187301 995407 187357 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[21]
port 517 nsew signal input
flabel metal2 s 179849 995407 179905 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[21]
port 518 nsew signal input
flabel metal2 s 182977 995407 183033 995887 0 FreeSans 320 90 0 0 mprj_io_out[21]
port 519 nsew signal input
flabel metal2 s 192177 995407 192233 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[21]
port 520 nsew signal input
flabel metal2 s 181137 995407 181193 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[21]
port 521 nsew signal input
flabel metal2 s 194017 995407 194073 995887 0 FreeSans 320 90 0 0 mprj_io_in[21]
port 522 nsew signal tristate
flabel metal2 s 140133 995407 140189 995887 0 FreeSans 320 90 0 0 mprj_analog_io[15]
port 523 nsew signal bidirectional
flabel metal5 s 129820 1018512 142360 1031002 6 FreeSans 320 0 0 0 mprj_io[22]
port 524 nsew signal bidirectional
flabel metal2 s 137741 995407 137797 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[22]
port 525 nsew signal input
flabel metal2 s 136453 995407 136509 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[22]
port 526 nsew signal input
flabel metal2 s 133417 995407 133473 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[22]
port 527 nsew signal input
flabel metal2 s 137097 995407 137153 995887 0 FreeSans 320 90 0 0 mprj_io_dm[66]
port 528 nsew signal input
flabel metal2 s 138937 995407 138993 995887 0 FreeSans 320 90 0 0 mprj_io_dm[67]
port 529 nsew signal input
flabel metal2 s 132773 995407 132829 995887 0 FreeSans 320 90 0 0 mprj_io_dm[68]
port 530 nsew signal input
flabel metal2 s 132129 995407 132185 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[22]
port 531 nsew signal input
flabel metal2 s 129093 995407 129149 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[22]
port 532 nsew signal input
flabel metal2 s 135901 995407 135957 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[22]
port 533 nsew signal input
flabel metal2 s 128449 995407 128505 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[22]
port 534 nsew signal input
flabel metal2 s 131577 995407 131633 995887 0 FreeSans 320 90 0 0 mprj_io_out[22]
port 535 nsew signal input
flabel metal2 s 140777 995407 140833 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[22]
port 536 nsew signal input
flabel metal2 s 129737 995407 129793 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[22]
port 537 nsew signal input
flabel metal2 s 142617 995407 142673 995887 0 FreeSans 320 90 0 0 mprj_io_in[22]
port 538 nsew signal tristate
flabel metal2 s 88733 995407 88789 995887 0 FreeSans 320 90 0 0 mprj_analog_io[16]
port 539 nsew signal bidirectional
flabel metal5 s 78420 1018512 90960 1031002 6 FreeSans 320 0 0 0 mprj_io[23]
port 540 nsew signal bidirectional
flabel metal2 s 86341 995407 86397 995887 0 FreeSans 320 90 0 0 mprj_io_analog_en[23]
port 541 nsew signal input
flabel metal2 s 85053 995407 85109 995887 0 FreeSans 320 90 0 0 mprj_io_analog_pol[23]
port 542 nsew signal input
flabel metal2 s 82017 995407 82073 995887 0 FreeSans 320 90 0 0 mprj_io_analog_sel[23]
port 543 nsew signal input
flabel metal2 s 85697 995407 85753 995887 0 FreeSans 320 90 0 0 mprj_io_dm[69]
port 544 nsew signal input
flabel metal2 s 87537 995407 87593 995887 0 FreeSans 320 90 0 0 mprj_io_dm[70]
port 545 nsew signal input
flabel metal2 s 81373 995407 81429 995887 0 FreeSans 320 90 0 0 mprj_io_dm[71]
port 546 nsew signal input
flabel metal2 s 80729 995407 80785 995887 0 FreeSans 320 90 0 0 mprj_io_holdover[23]
port 547 nsew signal input
flabel metal2 s 77693 995407 77749 995887 0 FreeSans 320 90 0 0 mprj_io_ib_mode_sel[23]
port 548 nsew signal input
flabel metal2 s 84501 995407 84557 995887 0 FreeSans 320 90 0 0 mprj_io_inp_dis[23]
port 549 nsew signal input
flabel metal2 s 77049 995407 77105 995887 0 FreeSans 320 90 0 0 mprj_io_oeb[23]
port 550 nsew signal input
flabel metal2 s 80177 995407 80233 995887 0 FreeSans 320 90 0 0 mprj_io_out[23]
port 551 nsew signal input
flabel metal2 s 89377 995407 89433 995887 0 FreeSans 320 90 0 0 mprj_io_slow_sel[23]
port 552 nsew signal input
flabel metal2 s 78337 995407 78393 995887 0 FreeSans 320 90 0 0 mprj_io_vtrip_sel[23]
port 553 nsew signal input
flabel metal2 s 91217 995407 91273 995887 0 FreeSans 320 90 0 0 mprj_io_in[23]
port 554 nsew signal tristate
flabel metal2 s 41713 966733 42193 966789 0 FreeSans 320 0 0 0 mprj_analog_io[17]
port 555 nsew signal bidirectional
flabel metal5 s 6598 956420 19088 968960 6 FreeSans 320 0 0 0 mprj_io[24]
port 556 nsew signal bidirectional
flabel metal2 s 41713 964341 42193 964397 0 FreeSans 320 0 0 0 mprj_io_analog_en[24]
port 557 nsew signal input
flabel metal2 s 41713 963053 42193 963109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[24]
port 558 nsew signal input
flabel metal2 s 41713 960017 42193 960073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[24]
port 559 nsew signal input
flabel metal2 s 41713 963697 42193 963753 0 FreeSans 320 0 0 0 mprj_io_dm[72]
port 560 nsew signal input
flabel metal2 s 41713 965537 42193 965593 0 FreeSans 320 0 0 0 mprj_io_dm[73]
port 561 nsew signal input
flabel metal2 s 41713 959373 42193 959429 0 FreeSans 320 0 0 0 mprj_io_dm[74]
port 562 nsew signal input
flabel metal2 s 41713 958729 42193 958785 0 FreeSans 320 0 0 0 mprj_io_holdover[24]
port 563 nsew signal input
flabel metal2 s 41713 955693 42193 955749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[24]
port 564 nsew signal input
flabel metal2 s 41713 962501 42193 962557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[24]
port 565 nsew signal input
flabel metal2 s 41713 955049 42193 955105 0 FreeSans 320 0 0 0 mprj_io_oeb[24]
port 566 nsew signal input
flabel metal2 s 41713 958177 42193 958233 0 FreeSans 320 0 0 0 mprj_io_out[24]
port 567 nsew signal input
flabel metal2 s 41713 967377 42193 967433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[24]
port 568 nsew signal input
flabel metal2 s 41713 956337 42193 956393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[24]
port 569 nsew signal input
flabel metal2 s 41713 969217 42193 969273 0 FreeSans 320 0 0 0 mprj_io_in[24]
port 570 nsew signal tristate
flabel metal2 s 41713 796933 42193 796989 0 FreeSans 320 0 0 0 mprj_analog_io[18]
port 571 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 6 FreeSans 320 0 0 0 mprj_io[25]
port 572 nsew signal bidirectional
flabel metal2 s 41713 794541 42193 794597 0 FreeSans 320 0 0 0 mprj_io_analog_en[25]
port 573 nsew signal input
flabel metal2 s 41713 793253 42193 793309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[25]
port 574 nsew signal input
flabel metal2 s 41713 790217 42193 790273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[25]
port 575 nsew signal input
flabel metal2 s 41713 793897 42193 793953 0 FreeSans 320 0 0 0 mprj_io_dm[75]
port 576 nsew signal input
flabel metal2 s 41713 795737 42193 795793 0 FreeSans 320 0 0 0 mprj_io_dm[76]
port 577 nsew signal input
flabel metal2 s 41713 789573 42193 789629 0 FreeSans 320 0 0 0 mprj_io_dm[77]
port 578 nsew signal input
flabel metal2 s 41713 788929 42193 788985 0 FreeSans 320 0 0 0 mprj_io_holdover[25]
port 579 nsew signal input
flabel metal2 s 41713 785893 42193 785949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[25]
port 580 nsew signal input
flabel metal2 s 41713 792701 42193 792757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[25]
port 581 nsew signal input
flabel metal2 s 41713 785249 42193 785305 0 FreeSans 320 0 0 0 mprj_io_oeb[25]
port 582 nsew signal input
flabel metal2 s 41713 788377 42193 788433 0 FreeSans 320 0 0 0 mprj_io_out[25]
port 583 nsew signal input
flabel metal2 s 41713 797577 42193 797633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[25]
port 584 nsew signal input
flabel metal2 s 41713 786537 42193 786593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[25]
port 585 nsew signal input
flabel metal2 s 41713 799417 42193 799473 0 FreeSans 320 0 0 0 mprj_io_in[25]
port 586 nsew signal tristate
flabel metal2 s 41713 753733 42193 753789 0 FreeSans 320 0 0 0 mprj_analog_io[19]
port 587 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 6 FreeSans 320 0 0 0 mprj_io[26]
port 588 nsew signal bidirectional
flabel metal2 s 41713 751341 42193 751397 0 FreeSans 320 0 0 0 mprj_io_analog_en[26]
port 589 nsew signal input
flabel metal2 s 41713 750053 42193 750109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[26]
port 590 nsew signal input
flabel metal2 s 41713 747017 42193 747073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[26]
port 591 nsew signal input
flabel metal2 s 41713 750697 42193 750753 0 FreeSans 320 0 0 0 mprj_io_dm[78]
port 592 nsew signal input
flabel metal2 s 41713 752537 42193 752593 0 FreeSans 320 0 0 0 mprj_io_dm[79]
port 593 nsew signal input
flabel metal2 s 41713 746373 42193 746429 0 FreeSans 320 0 0 0 mprj_io_dm[80]
port 594 nsew signal input
flabel metal2 s 41713 745729 42193 745785 0 FreeSans 320 0 0 0 mprj_io_holdover[26]
port 595 nsew signal input
flabel metal2 s 41713 742693 42193 742749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[26]
port 596 nsew signal input
flabel metal2 s 41713 749501 42193 749557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[26]
port 597 nsew signal input
flabel metal2 s 41713 742049 42193 742105 0 FreeSans 320 0 0 0 mprj_io_oeb[26]
port 598 nsew signal input
flabel metal2 s 41713 745177 42193 745233 0 FreeSans 320 0 0 0 mprj_io_out[26]
port 599 nsew signal input
flabel metal2 s 41713 754377 42193 754433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[26]
port 600 nsew signal input
flabel metal2 s 41713 743337 42193 743393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[26]
port 601 nsew signal input
flabel metal2 s 41713 756217 42193 756273 0 FreeSans 320 0 0 0 mprj_io_in[26]
port 602 nsew signal tristate
flabel metal2 s 41713 710533 42193 710589 0 FreeSans 320 0 0 0 mprj_analog_io[20]
port 603 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 6 FreeSans 320 0 0 0 mprj_io[27]
port 604 nsew signal bidirectional
flabel metal2 s 41713 708141 42193 708197 0 FreeSans 320 0 0 0 mprj_io_analog_en[27]
port 605 nsew signal input
flabel metal2 s 41713 706853 42193 706909 0 FreeSans 320 0 0 0 mprj_io_analog_pol[27]
port 606 nsew signal input
flabel metal2 s 41713 703817 42193 703873 0 FreeSans 320 0 0 0 mprj_io_analog_sel[27]
port 607 nsew signal input
flabel metal2 s 41713 707497 42193 707553 0 FreeSans 320 0 0 0 mprj_io_dm[81]
port 608 nsew signal input
flabel metal2 s 41713 709337 42193 709393 0 FreeSans 320 0 0 0 mprj_io_dm[82]
port 609 nsew signal input
flabel metal2 s 41713 703173 42193 703229 0 FreeSans 320 0 0 0 mprj_io_dm[83]
port 610 nsew signal input
flabel metal2 s 41713 702529 42193 702585 0 FreeSans 320 0 0 0 mprj_io_holdover[27]
port 611 nsew signal input
flabel metal2 s 41713 699493 42193 699549 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[27]
port 612 nsew signal input
flabel metal2 s 41713 706301 42193 706357 0 FreeSans 320 0 0 0 mprj_io_inp_dis[27]
port 613 nsew signal input
flabel metal2 s 41713 698849 42193 698905 0 FreeSans 320 0 0 0 mprj_io_oeb[27]
port 614 nsew signal input
flabel metal2 s 41713 701977 42193 702033 0 FreeSans 320 0 0 0 mprj_io_out[27]
port 615 nsew signal input
flabel metal2 s 41713 711177 42193 711233 0 FreeSans 320 0 0 0 mprj_io_slow_sel[27]
port 616 nsew signal input
flabel metal2 s 41713 700137 42193 700193 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[27]
port 617 nsew signal input
flabel metal2 s 41713 713017 42193 713073 0 FreeSans 320 0 0 0 mprj_io_in[27]
port 618 nsew signal tristate
flabel metal2 s 41713 667333 42193 667389 0 FreeSans 320 0 0 0 mprj_analog_io[21]
port 619 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 6 FreeSans 320 0 0 0 mprj_io[28]
port 620 nsew signal bidirectional
flabel metal2 s 41713 664941 42193 664997 0 FreeSans 320 0 0 0 mprj_io_analog_en[28]
port 621 nsew signal input
flabel metal2 s 41713 663653 42193 663709 0 FreeSans 320 0 0 0 mprj_io_analog_pol[28]
port 622 nsew signal input
flabel metal2 s 41713 660617 42193 660673 0 FreeSans 320 0 0 0 mprj_io_analog_sel[28]
port 623 nsew signal input
flabel metal2 s 41713 664297 42193 664353 0 FreeSans 320 0 0 0 mprj_io_dm[84]
port 624 nsew signal input
flabel metal2 s 41713 666137 42193 666193 0 FreeSans 320 0 0 0 mprj_io_dm[85]
port 625 nsew signal input
flabel metal2 s 41713 659973 42193 660029 0 FreeSans 320 0 0 0 mprj_io_dm[86]
port 626 nsew signal input
flabel metal2 s 41713 659329 42193 659385 0 FreeSans 320 0 0 0 mprj_io_holdover[28]
port 627 nsew signal input
flabel metal2 s 41713 656293 42193 656349 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[28]
port 628 nsew signal input
flabel metal2 s 41713 663101 42193 663157 0 FreeSans 320 0 0 0 mprj_io_inp_dis[28]
port 629 nsew signal input
flabel metal2 s 41713 655649 42193 655705 0 FreeSans 320 0 0 0 mprj_io_oeb[28]
port 630 nsew signal input
flabel metal2 s 41713 658777 42193 658833 0 FreeSans 320 0 0 0 mprj_io_out[28]
port 631 nsew signal input
flabel metal2 s 41713 667977 42193 668033 0 FreeSans 320 0 0 0 mprj_io_slow_sel[28]
port 632 nsew signal input
flabel metal2 s 41713 656937 42193 656993 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[28]
port 633 nsew signal input
flabel metal2 s 41713 669817 42193 669873 0 FreeSans 320 0 0 0 mprj_io_in[28]
port 634 nsew signal tristate
flabel metal5 s 136713 7143 144149 18309 6 FreeSans 320 0 0 0 resetb
port 636 nsew signal input
flabel metal4 s 132600 36323 132792 37013 6 FreeSans 320 0 0 0 vdda
port 638 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 6 FreeSans 320 0 0 0 vccd1_pad
port 641 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 6 FreeSans 320 0 0 0 vdda1_pad
port 642 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 6 FreeSans 320 0 0 0 vdda1_pad2
port 643 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 6 FreeSans 320 0 0 0 vssa1_pad
port 644 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 6 FreeSans 320 0 0 0 vssa1_pad2
port 645 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 6 FreeSans 320 0 0 0 vssd1_pad
port 650 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 6 FreeSans 320 0 0 0 vccd2_pad
port 651 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 6 FreeSans 320 0 0 0 vdda2_pad
port 652 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 6 FreeSans 320 0 0 0 vssa2_pad
port 653 nsew signal bidirectional
flabel metal4 s 36323 455607 37013 455799 6 FreeSans 320 0 0 0 vdda2
port 656 nsew signal bidirectional
flabel metal4 s 28653 440800 28719 455800 6 FreeSans 320 0 0 0 vssa2
port 658 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 6 FreeSans 320 0 0 0 vssd2_pad
port 660 nsew signal bidirectional
flabel metal2 141667 39934 141813 40000 0 FreeSans 320 0 0 0 resetb_core_h
port 637 nsew signal tristate
flabel metal5 41130 179416 43498 180132 0 FreeSans 3200 0 0 0 vssd2
port 659 nsew signal bidirectional
flabel metal5 44242 179326 46748 180098 0 FreeSans 3200 0 0 0 vccd2
port 655 nsew signal bidirectional
flabel metal5 670926 95262 673290 96090 0 FreeSans 3200 180 0 0 vssd1
port 649 nsew signal bidirectional
flabel metal5 674122 95266 676502 96062 0 FreeSans 3200 180 0 0 vccd1
port 646 nsew signal bidirectional
flabel metal2 675407 102123 675887 102179 0 FreeSans 320 0 0 0 mprj_io_one[0]
port 661 nsew
flabel metal2 675407 147323 675887 147379 0 FreeSans 320 0 0 0 mprj_io_one[1]
port 662 nsew
flabel metal2 675407 192323 675887 192379 0 FreeSans 320 0 0 0 mprj_io_one[2]
port 663 nsew
flabel metal2 675407 237523 675887 237579 0 FreeSans 320 0 0 0 mprj_io_one[3]
port 664 nsew
flabel metal2 675407 282523 675887 282579 0 FreeSans 320 0 0 0 mprj_io_one[4]
port 665 nsew
flabel metal2 675407 327523 675887 327579 0 FreeSans 320 0 0 0 mprj_io_one[5]
port 666 nsew
flabel metal2 675407 372723 675887 372779 0 FreeSans 320 0 0 0 mprj_io_one[6]
port 667 nsew
flabel metal2 675407 549923 675887 549979 0 FreeSans 320 0 0 0 mprj_io_one[7]
port 668 nsew
flabel metal2 675407 595123 675887 595179 0 FreeSans 320 0 0 0 mprj_io_one[8]
port 669 nsew
flabel metal2 675407 640123 675887 640179 0 FreeSans 320 0 0 0 mprj_io_one[9]
port 670 nsew
flabel metal2 675407 685323 675887 685379 0 FreeSans 320 0 0 0 mprj_io_one[10]
port 671 nsew
flabel metal2 675407 730323 675887 730379 0 FreeSans 320 0 0 0 mprj_io_one[11]
port 672 nsew
flabel metal2 675407 775323 675887 775379 0 FreeSans 320 0 0 0 mprj_io_one[12]
port 673 nsew
flabel metal2 675407 864523 675887 864579 0 FreeSans 320 0 0 0 mprj_io_one[13]
port 674 nsew
flabel metal2 675407 953723 675887 953779 0 FreeSans 320 0 0 0 mprj_io_one[14]
port 675 nsew
flabel metal2 639821 995407 639877 995887 0 FreeSans 320 90 0 0 mprj_io_one[15]
port 676 nsew
flabel metal2 538021 995407 538077 995887 0 FreeSans 320 90 0 0 mprj_io_one[16]
port 677 nsew
flabel metal2 486621 995407 486677 995887 0 FreeSans 320 90 0 0 mprj_io_one[17]
port 678 nsew
flabel metal2 397621 995407 397677 995887 0 FreeSans 320 90 0 0 mprj_io_one[18]
port 679 nsew
flabel metal2 295821 995407 295877 995887 0 FreeSans 320 90 0 0 mprj_io_one[19]
port 680 nsew
flabel metal2 244221 995407 244277 995887 0 FreeSans 320 90 0 0 mprj_io_one[20]
port 681 nsew
flabel metal2 192821 995407 192877 995887 0 FreeSans 320 90 0 0 mprj_io_one[21]
port 682 nsew
flabel metal2 141421 995407 141477 995887 0 FreeSans 320 90 0 0 mprj_io_one[22]
port 683 nsew
flabel metal2 90021 995407 90077 995887 0 FreeSans 320 90 0 0 mprj_io_one[23]
port 684 nsew
flabel metal2 41713 968021 42193 968077 0 FreeSans 320 0 0 0 mprj_io_one[24]
port 686 nsew
flabel metal2 41713 798221 42193 798277 0 FreeSans 320 0 0 0 mprj_io_one[25]
port 687 nsew
flabel metal2 41713 755021 42193 755077 0 FreeSans 320 0 0 0 mprj_io_one[26]
port 688 nsew
flabel metal2 41713 711821 42193 711877 0 FreeSans 320 0 0 0 mprj_io_one[27]
port 689 nsew
flabel metal2 41713 668621 42193 668677 0 FreeSans 320 0 0 0 mprj_io_one[28]
port 690 nsew
flabel metal2 41713 625421 42193 625477 0 FreeSans 320 0 0 0 mprj_io_one[29]
port 691 nsew
flabel metal2 41713 582221 42193 582277 0 FreeSans 320 0 0 0 mprj_io_one[30]
port 692 nsew
flabel metal2 41713 539021 42193 539077 0 FreeSans 320 0 0 0 mprj_io_one[31]
port 693 nsew
flabel metal2 41713 411421 42193 411477 0 FreeSans 320 0 0 0 mprj_io_one[32]
port 694 nsew
flabel metal2 41713 368221 42193 368277 0 FreeSans 320 0 0 0 mprj_io_one[33]
port 695 nsew
flabel metal2 41713 325021 42193 325077 0 FreeSans 320 0 0 0 mprj_io_one[34]
port 696 nsew
flabel metal2 41713 281821 42193 281877 0 FreeSans 320 0 0 0 mprj_io_one[35]
port 697 nsew
flabel metal2 41713 238621 42193 238677 0 FreeSans 320 0 0 0 mprj_io_one[36]
port 698 nsew
flabel metal2 41713 195421 42193 195477 0 FreeSans 320 0 0 0 mprj_io_one[37]
port 699 nsew
flabel metal2 s 467043 41713 467099 42193 0 FreeSans 320 90 0 0 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal3 140494 40183 140494 40183 1 xresloop
rlabel metal1 142538 40100 142538 40100 1 xres_vss_loop
flabel metal2 308255 41713 308311 42193 0 FreeSans 320 90 0 0 porb_h
port 700 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
