VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping_alt
  CLASS BLOCK ;
  FOREIGN housekeeping_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 410.230 BY 550.950 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 366.640 10.640 368.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 289.840 10.640 291.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.040 10.640 214.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.240 10.640 137.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.440 10.640 61.040 538.800 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
  END VPWR
  PIN debug_in
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END debug_in
  PIN debug_mode
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END debug_mode
  PIN debug_oeb
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END debug_oeb
  PIN debug_out
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END debug_out
  PIN irq[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END irq[0]
  PIN irq[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END irq[1]
  PIN irq[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 54.440 410.230 55.040 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 299.240 410.230 299.840 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 323.720 410.230 324.320 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 348.200 410.230 348.800 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 372.680 410.230 373.280 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 397.160 410.230 397.760 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 421.640 410.230 422.240 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 446.120 410.230 446.720 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 470.600 410.230 471.200 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 495.080 410.230 495.680 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 519.560 410.230 520.160 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 78.920 410.230 79.520 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 233.770 546.950 234.050 550.950 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 242.050 546.950 242.330 550.950 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 250.330 546.950 250.610 550.950 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 258.610 546.950 258.890 550.950 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 266.890 546.950 267.170 550.950 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 275.170 546.950 275.450 550.950 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 546.950 283.730 550.950 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 291.730 546.950 292.010 550.950 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 300.010 546.950 300.290 550.950 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 308.290 546.950 308.570 550.950 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 103.400 410.230 104.000 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 316.570 546.950 316.850 550.950 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 324.850 546.950 325.130 550.950 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.130 546.950 333.410 550.950 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 546.950 341.690 550.950 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.690 546.950 349.970 550.950 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 357.970 546.950 358.250 550.950 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 366.250 546.950 366.530 550.950 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 374.530 546.950 374.810 550.950 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 127.880 410.230 128.480 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 152.360 410.230 152.960 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 176.840 410.230 177.440 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 201.320 410.230 201.920 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 225.800 410.230 226.400 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 250.280 410.230 250.880 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 406.230 274.760 410.230 275.360 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 62.600 410.230 63.200 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 307.400 410.230 308.000 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 331.880 410.230 332.480 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 356.360 410.230 356.960 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 380.840 410.230 381.440 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 405.320 410.230 405.920 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 429.800 410.230 430.400 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 454.280 410.230 454.880 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 478.760 410.230 479.360 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 503.240 410.230 503.840 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 527.720 410.230 528.320 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 87.080 410.230 87.680 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.530 546.950 236.810 550.950 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 546.950 245.090 550.950 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 253.090 546.950 253.370 550.950 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 546.950 261.650 550.950 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 546.950 269.930 550.950 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 546.950 278.210 550.950 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 286.210 546.950 286.490 550.950 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 294.490 546.950 294.770 550.950 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 546.950 303.050 550.950 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 311.050 546.950 311.330 550.950 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 111.560 410.230 112.160 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 319.330 546.950 319.610 550.950 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 327.610 546.950 327.890 550.950 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 546.950 336.170 550.950 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 344.170 546.950 344.450 550.950 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 546.950 352.730 550.950 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 546.950 361.010 550.950 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 369.010 546.950 369.290 550.950 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 377.290 546.950 377.570 550.950 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 136.040 410.230 136.640 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 160.520 410.230 161.120 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 185.000 410.230 185.600 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 209.480 410.230 210.080 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 233.960 410.230 234.560 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 258.440 410.230 259.040 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 282.920 410.230 283.520 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 70.760 410.230 71.360 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 315.560 410.230 316.160 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 340.040 410.230 340.640 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 364.520 410.230 365.120 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 389.000 410.230 389.600 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 406.230 413.480 410.230 414.080 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 406.230 437.960 410.230 438.560 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 462.440 410.230 463.040 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 486.920 410.230 487.520 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 511.400 410.230 512.000 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 535.880 410.230 536.480 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 95.240 410.230 95.840 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 239.290 546.950 239.570 550.950 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 546.950 247.850 550.950 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 255.850 546.950 256.130 550.950 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 264.130 546.950 264.410 550.950 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 272.410 546.950 272.690 550.950 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 280.690 546.950 280.970 550.950 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 288.970 546.950 289.250 550.950 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 297.250 546.950 297.530 550.950 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 305.530 546.950 305.810 550.950 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 546.950 314.090 550.950 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 119.720 410.230 120.320 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 322.090 546.950 322.370 550.950 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 330.370 546.950 330.650 550.950 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 546.950 338.930 550.950 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 346.930 546.950 347.210 550.950 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 355.210 546.950 355.490 550.950 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 363.490 546.950 363.770 550.950 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 371.770 546.950 372.050 550.950 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 546.950 380.330 550.950 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 144.200 410.230 144.800 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 168.680 410.230 169.280 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 193.160 410.230 193.760 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 217.640 410.230 218.240 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 242.120 410.230 242.720 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 266.600 410.230 267.200 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 406.230 291.080 410.230 291.680 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oeb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END pad_flash_clk_oeb
  PIN pad_flash_csb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oeb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END pad_flash_csb_oeb
  PIN pad_flash_io0_di
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ieb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END pad_flash_io0_ieb
  PIN pad_flash_io0_oeb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END pad_flash_io0_oeb
  PIN pad_flash_io1_di
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ieb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END pad_flash_io1_ieb
  PIN pad_flash_io1_oeb
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END pad_flash_io1_oeb
  PIN pll90_sel[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END pwr_ctrl_out[0]
  PIN pwr_ctrl_out[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END pwr_ctrl_out[1]
  PIN pwr_ctrl_out[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END pwr_ctrl_out[2]
  PIN pwr_ctrl_out[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END pwr_ctrl_out[3]
  PIN qspi_enabled
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END qspi_enabled
  PIN reset
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END reset
  PIN ser_rx
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END ser_rx
  PIN ser_tx
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END ser_tx
  PIN serial_clock
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 13.640 410.230 14.240 ;
    END
  END serial_clock
  PIN serial_data_1
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 38.120 410.230 38.720 ;
    END
  END serial_data_1
  PIN serial_data_2
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 46.280 410.230 46.880 ;
    END
  END serial_data_2
  PIN serial_load
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 29.960 410.230 30.560 ;
    END
  END serial_load
  PIN serial_resetn
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 406.230 21.800 410.230 22.400 ;
    END
  END serial_resetn
  PIN spi_csb
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END spi_csb
  PIN spi_enabled
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END spi_enabled
  PIN spi_sck
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END spi_sck
  PIN spi_sdi
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END spi_sdi
  PIN spi_sdo
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END trap
  PIN uart_enabled
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END uart_enabled
  PIN user_clock
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END user_clock
  PIN usr1_vcc_pwrgood
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 222.730 546.950 223.010 550.950 ;
    END
  END usr1_vcc_pwrgood
  PIN usr1_vdd_pwrgood
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 228.250 546.950 228.530 550.950 ;
    END
  END usr1_vdd_pwrgood
  PIN usr2_vcc_pwrgood
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 225.490 546.950 225.770 550.950 ;
    END
  END usr2_vcc_pwrgood
  PIN usr2_vdd_pwrgood
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 231.010 546.950 231.290 550.950 ;
    END
  END usr2_vdd_pwrgood
  PIN wb_ack_o
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.530 546.950 29.810 550.950 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 57.130 546.950 57.410 550.950 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.890 546.950 60.170 550.950 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.650 546.950 62.930 550.950 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 65.410 546.950 65.690 550.950 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 68.170 546.950 68.450 550.950 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.930 546.950 71.210 550.950 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.690 546.950 73.970 550.950 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 76.450 546.950 76.730 550.950 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.210 546.950 79.490 550.950 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.970 546.950 82.250 550.950 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 546.950 32.570 550.950 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.730 546.950 85.010 550.950 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.490 546.950 87.770 550.950 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 546.950 90.530 550.950 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.010 546.950 93.290 550.950 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.770 546.950 96.050 550.950 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.530 546.950 98.810 550.950 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 101.290 546.950 101.570 550.950 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 104.050 546.950 104.330 550.950 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.810 546.950 107.090 550.950 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 546.950 109.850 550.950 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.050 546.950 35.330 550.950 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.330 546.950 112.610 550.950 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 115.090 546.950 115.370 550.950 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.810 546.950 38.090 550.950 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.570 546.950 40.850 550.950 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 43.330 546.950 43.610 550.950 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 46.090 546.950 46.370 550.950 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.850 546.950 49.130 550.950 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 546.950 51.890 550.950 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.370 546.950 54.650 550.950 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 219.970 546.950 220.250 550.950 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 117.850 546.950 118.130 550.950 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 145.450 546.950 145.730 550.950 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 148.210 546.950 148.490 550.950 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 150.970 546.950 151.250 550.950 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 153.730 546.950 154.010 550.950 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 156.490 546.950 156.770 550.950 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 159.250 546.950 159.530 550.950 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.010 546.950 162.290 550.950 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.770 546.950 165.050 550.950 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 167.530 546.950 167.810 550.950 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.290 546.950 170.570 550.950 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 120.610 546.950 120.890 550.950 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.050 546.950 173.330 550.950 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.810 546.950 176.090 550.950 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 178.570 546.950 178.850 550.950 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 181.330 546.950 181.610 550.950 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 184.090 546.950 184.370 550.950 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 546.950 187.130 550.950 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 189.610 546.950 189.890 550.950 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 192.370 546.950 192.650 550.950 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.130 546.950 195.410 550.950 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 197.890 546.950 198.170 550.950 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 123.370 546.950 123.650 550.950 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 200.650 546.950 200.930 550.950 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 203.410 546.950 203.690 550.950 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 126.130 546.950 126.410 550.950 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 546.950 129.170 550.950 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.650 546.950 131.930 550.950 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 134.410 546.950 134.690 550.950 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 137.170 546.950 137.450 550.950 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 139.930 546.950 140.210 550.950 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 142.690 546.950 142.970 550.950 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 546.950 206.450 550.950 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.930 546.950 209.210 550.950 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 211.690 546.950 211.970 550.950 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 214.450 546.950 214.730 550.950 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END wb_stb_i
  PIN wb_we_i
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.210 546.950 217.490 550.950 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 404.340 538.645 ;
      LAYER met1 ;
        RECT 4.670 6.840 409.790 538.800 ;
      LAYER met2 ;
        RECT 4.690 546.670 29.250 547.130 ;
        RECT 30.090 546.670 32.010 547.130 ;
        RECT 32.850 546.670 34.770 547.130 ;
        RECT 35.610 546.670 37.530 547.130 ;
        RECT 38.370 546.670 40.290 547.130 ;
        RECT 41.130 546.670 43.050 547.130 ;
        RECT 43.890 546.670 45.810 547.130 ;
        RECT 46.650 546.670 48.570 547.130 ;
        RECT 49.410 546.670 51.330 547.130 ;
        RECT 52.170 546.670 54.090 547.130 ;
        RECT 54.930 546.670 56.850 547.130 ;
        RECT 57.690 546.670 59.610 547.130 ;
        RECT 60.450 546.670 62.370 547.130 ;
        RECT 63.210 546.670 65.130 547.130 ;
        RECT 65.970 546.670 67.890 547.130 ;
        RECT 68.730 546.670 70.650 547.130 ;
        RECT 71.490 546.670 73.410 547.130 ;
        RECT 74.250 546.670 76.170 547.130 ;
        RECT 77.010 546.670 78.930 547.130 ;
        RECT 79.770 546.670 81.690 547.130 ;
        RECT 82.530 546.670 84.450 547.130 ;
        RECT 85.290 546.670 87.210 547.130 ;
        RECT 88.050 546.670 89.970 547.130 ;
        RECT 90.810 546.670 92.730 547.130 ;
        RECT 93.570 546.670 95.490 547.130 ;
        RECT 96.330 546.670 98.250 547.130 ;
        RECT 99.090 546.670 101.010 547.130 ;
        RECT 101.850 546.670 103.770 547.130 ;
        RECT 104.610 546.670 106.530 547.130 ;
        RECT 107.370 546.670 109.290 547.130 ;
        RECT 110.130 546.670 112.050 547.130 ;
        RECT 112.890 546.670 114.810 547.130 ;
        RECT 115.650 546.670 117.570 547.130 ;
        RECT 118.410 546.670 120.330 547.130 ;
        RECT 121.170 546.670 123.090 547.130 ;
        RECT 123.930 546.670 125.850 547.130 ;
        RECT 126.690 546.670 128.610 547.130 ;
        RECT 129.450 546.670 131.370 547.130 ;
        RECT 132.210 546.670 134.130 547.130 ;
        RECT 134.970 546.670 136.890 547.130 ;
        RECT 137.730 546.670 139.650 547.130 ;
        RECT 140.490 546.670 142.410 547.130 ;
        RECT 143.250 546.670 145.170 547.130 ;
        RECT 146.010 546.670 147.930 547.130 ;
        RECT 148.770 546.670 150.690 547.130 ;
        RECT 151.530 546.670 153.450 547.130 ;
        RECT 154.290 546.670 156.210 547.130 ;
        RECT 157.050 546.670 158.970 547.130 ;
        RECT 159.810 546.670 161.730 547.130 ;
        RECT 162.570 546.670 164.490 547.130 ;
        RECT 165.330 546.670 167.250 547.130 ;
        RECT 168.090 546.670 170.010 547.130 ;
        RECT 170.850 546.670 172.770 547.130 ;
        RECT 173.610 546.670 175.530 547.130 ;
        RECT 176.370 546.670 178.290 547.130 ;
        RECT 179.130 546.670 181.050 547.130 ;
        RECT 181.890 546.670 183.810 547.130 ;
        RECT 184.650 546.670 186.570 547.130 ;
        RECT 187.410 546.670 189.330 547.130 ;
        RECT 190.170 546.670 192.090 547.130 ;
        RECT 192.930 546.670 194.850 547.130 ;
        RECT 195.690 546.670 197.610 547.130 ;
        RECT 198.450 546.670 200.370 547.130 ;
        RECT 201.210 546.670 203.130 547.130 ;
        RECT 203.970 546.670 205.890 547.130 ;
        RECT 206.730 546.670 208.650 547.130 ;
        RECT 209.490 546.670 211.410 547.130 ;
        RECT 212.250 546.670 214.170 547.130 ;
        RECT 215.010 546.670 216.930 547.130 ;
        RECT 217.770 546.670 219.690 547.130 ;
        RECT 220.530 546.670 222.450 547.130 ;
        RECT 223.290 546.670 225.210 547.130 ;
        RECT 226.050 546.670 227.970 547.130 ;
        RECT 228.810 546.670 230.730 547.130 ;
        RECT 231.570 546.670 233.490 547.130 ;
        RECT 234.330 546.670 236.250 547.130 ;
        RECT 237.090 546.670 239.010 547.130 ;
        RECT 239.850 546.670 241.770 547.130 ;
        RECT 242.610 546.670 244.530 547.130 ;
        RECT 245.370 546.670 247.290 547.130 ;
        RECT 248.130 546.670 250.050 547.130 ;
        RECT 250.890 546.670 252.810 547.130 ;
        RECT 253.650 546.670 255.570 547.130 ;
        RECT 256.410 546.670 258.330 547.130 ;
        RECT 259.170 546.670 261.090 547.130 ;
        RECT 261.930 546.670 263.850 547.130 ;
        RECT 264.690 546.670 266.610 547.130 ;
        RECT 267.450 546.670 269.370 547.130 ;
        RECT 270.210 546.670 272.130 547.130 ;
        RECT 272.970 546.670 274.890 547.130 ;
        RECT 275.730 546.670 277.650 547.130 ;
        RECT 278.490 546.670 280.410 547.130 ;
        RECT 281.250 546.670 283.170 547.130 ;
        RECT 284.010 546.670 285.930 547.130 ;
        RECT 286.770 546.670 288.690 547.130 ;
        RECT 289.530 546.670 291.450 547.130 ;
        RECT 292.290 546.670 294.210 547.130 ;
        RECT 295.050 546.670 296.970 547.130 ;
        RECT 297.810 546.670 299.730 547.130 ;
        RECT 300.570 546.670 302.490 547.130 ;
        RECT 303.330 546.670 305.250 547.130 ;
        RECT 306.090 546.670 308.010 547.130 ;
        RECT 308.850 546.670 310.770 547.130 ;
        RECT 311.610 546.670 313.530 547.130 ;
        RECT 314.370 546.670 316.290 547.130 ;
        RECT 317.130 546.670 319.050 547.130 ;
        RECT 319.890 546.670 321.810 547.130 ;
        RECT 322.650 546.670 324.570 547.130 ;
        RECT 325.410 546.670 327.330 547.130 ;
        RECT 328.170 546.670 330.090 547.130 ;
        RECT 330.930 546.670 332.850 547.130 ;
        RECT 333.690 546.670 335.610 547.130 ;
        RECT 336.450 546.670 338.370 547.130 ;
        RECT 339.210 546.670 341.130 547.130 ;
        RECT 341.970 546.670 343.890 547.130 ;
        RECT 344.730 546.670 346.650 547.130 ;
        RECT 347.490 546.670 349.410 547.130 ;
        RECT 350.250 546.670 352.170 547.130 ;
        RECT 353.010 546.670 354.930 547.130 ;
        RECT 355.770 546.670 357.690 547.130 ;
        RECT 358.530 546.670 360.450 547.130 ;
        RECT 361.290 546.670 363.210 547.130 ;
        RECT 364.050 546.670 365.970 547.130 ;
        RECT 366.810 546.670 368.730 547.130 ;
        RECT 369.570 546.670 371.490 547.130 ;
        RECT 372.330 546.670 374.250 547.130 ;
        RECT 375.090 546.670 377.010 547.130 ;
        RECT 377.850 546.670 379.770 547.130 ;
        RECT 380.610 546.670 410.160 547.130 ;
        RECT 4.690 4.280 410.160 546.670 ;
        RECT 4.690 3.670 14.070 4.280 ;
        RECT 14.910 3.670 18.210 4.280 ;
        RECT 19.050 3.670 22.350 4.280 ;
        RECT 23.190 3.670 26.490 4.280 ;
        RECT 27.330 3.670 30.630 4.280 ;
        RECT 31.470 3.670 34.770 4.280 ;
        RECT 35.610 3.670 38.910 4.280 ;
        RECT 39.750 3.670 43.050 4.280 ;
        RECT 43.890 3.670 47.190 4.280 ;
        RECT 48.030 3.670 51.330 4.280 ;
        RECT 52.170 3.670 55.470 4.280 ;
        RECT 56.310 3.670 59.610 4.280 ;
        RECT 60.450 3.670 63.750 4.280 ;
        RECT 64.590 3.670 67.890 4.280 ;
        RECT 68.730 3.670 72.030 4.280 ;
        RECT 72.870 3.670 76.170 4.280 ;
        RECT 77.010 3.670 80.310 4.280 ;
        RECT 81.150 3.670 84.450 4.280 ;
        RECT 85.290 3.670 88.590 4.280 ;
        RECT 89.430 3.670 92.730 4.280 ;
        RECT 93.570 3.670 96.870 4.280 ;
        RECT 97.710 3.670 101.010 4.280 ;
        RECT 101.850 3.670 105.150 4.280 ;
        RECT 105.990 3.670 109.290 4.280 ;
        RECT 110.130 3.670 113.430 4.280 ;
        RECT 114.270 3.670 117.570 4.280 ;
        RECT 118.410 3.670 121.710 4.280 ;
        RECT 122.550 3.670 125.850 4.280 ;
        RECT 126.690 3.670 129.990 4.280 ;
        RECT 130.830 3.670 134.130 4.280 ;
        RECT 134.970 3.670 138.270 4.280 ;
        RECT 139.110 3.670 142.410 4.280 ;
        RECT 143.250 3.670 146.550 4.280 ;
        RECT 147.390 3.670 150.690 4.280 ;
        RECT 151.530 3.670 154.830 4.280 ;
        RECT 155.670 3.670 158.970 4.280 ;
        RECT 159.810 3.670 163.110 4.280 ;
        RECT 163.950 3.670 167.250 4.280 ;
        RECT 168.090 3.670 171.390 4.280 ;
        RECT 172.230 3.670 175.530 4.280 ;
        RECT 176.370 3.670 179.670 4.280 ;
        RECT 180.510 3.670 183.810 4.280 ;
        RECT 184.650 3.670 187.950 4.280 ;
        RECT 188.790 3.670 192.090 4.280 ;
        RECT 192.930 3.670 196.230 4.280 ;
        RECT 197.070 3.670 200.370 4.280 ;
        RECT 201.210 3.670 204.510 4.280 ;
        RECT 205.350 3.670 208.650 4.280 ;
        RECT 209.490 3.670 212.790 4.280 ;
        RECT 213.630 3.670 216.930 4.280 ;
        RECT 217.770 3.670 221.070 4.280 ;
        RECT 221.910 3.670 225.210 4.280 ;
        RECT 226.050 3.670 229.350 4.280 ;
        RECT 230.190 3.670 233.490 4.280 ;
        RECT 234.330 3.670 237.630 4.280 ;
        RECT 238.470 3.670 241.770 4.280 ;
        RECT 242.610 3.670 245.910 4.280 ;
        RECT 246.750 3.670 250.050 4.280 ;
        RECT 250.890 3.670 254.190 4.280 ;
        RECT 255.030 3.670 258.330 4.280 ;
        RECT 259.170 3.670 262.470 4.280 ;
        RECT 263.310 3.670 266.610 4.280 ;
        RECT 267.450 3.670 270.750 4.280 ;
        RECT 271.590 3.670 274.890 4.280 ;
        RECT 275.730 3.670 279.030 4.280 ;
        RECT 279.870 3.670 283.170 4.280 ;
        RECT 284.010 3.670 287.310 4.280 ;
        RECT 288.150 3.670 291.450 4.280 ;
        RECT 292.290 3.670 295.590 4.280 ;
        RECT 296.430 3.670 299.730 4.280 ;
        RECT 300.570 3.670 303.870 4.280 ;
        RECT 304.710 3.670 308.010 4.280 ;
        RECT 308.850 3.670 312.150 4.280 ;
        RECT 312.990 3.670 316.290 4.280 ;
        RECT 317.130 3.670 320.430 4.280 ;
        RECT 321.270 3.670 324.570 4.280 ;
        RECT 325.410 3.670 328.710 4.280 ;
        RECT 329.550 3.670 332.850 4.280 ;
        RECT 333.690 3.670 336.990 4.280 ;
        RECT 337.830 3.670 341.130 4.280 ;
        RECT 341.970 3.670 345.270 4.280 ;
        RECT 346.110 3.670 349.410 4.280 ;
        RECT 350.250 3.670 353.550 4.280 ;
        RECT 354.390 3.670 357.690 4.280 ;
        RECT 358.530 3.670 361.830 4.280 ;
        RECT 362.670 3.670 365.970 4.280 ;
        RECT 366.810 3.670 370.110 4.280 ;
        RECT 370.950 3.670 374.250 4.280 ;
        RECT 375.090 3.670 378.390 4.280 ;
        RECT 379.230 3.670 382.530 4.280 ;
        RECT 383.370 3.670 386.670 4.280 ;
        RECT 387.510 3.670 390.810 4.280 ;
        RECT 391.650 3.670 394.950 4.280 ;
        RECT 395.790 3.670 410.160 4.280 ;
      LAYER met3 ;
        RECT 4.400 539.560 409.795 540.425 ;
        RECT 4.000 536.880 409.795 539.560 ;
        RECT 4.000 535.480 405.830 536.880 ;
        RECT 4.000 532.800 409.795 535.480 ;
        RECT 4.400 531.400 409.795 532.800 ;
        RECT 4.000 528.720 409.795 531.400 ;
        RECT 4.000 527.320 405.830 528.720 ;
        RECT 4.000 524.640 409.795 527.320 ;
        RECT 4.400 523.240 409.795 524.640 ;
        RECT 4.000 520.560 409.795 523.240 ;
        RECT 4.000 519.160 405.830 520.560 ;
        RECT 4.000 516.480 409.795 519.160 ;
        RECT 4.400 515.080 409.795 516.480 ;
        RECT 4.000 512.400 409.795 515.080 ;
        RECT 4.000 511.000 405.830 512.400 ;
        RECT 4.000 508.320 409.795 511.000 ;
        RECT 4.400 506.920 409.795 508.320 ;
        RECT 4.000 504.240 409.795 506.920 ;
        RECT 4.000 502.840 405.830 504.240 ;
        RECT 4.000 500.160 409.795 502.840 ;
        RECT 4.400 498.760 409.795 500.160 ;
        RECT 4.000 496.080 409.795 498.760 ;
        RECT 4.000 494.680 405.830 496.080 ;
        RECT 4.000 492.000 409.795 494.680 ;
        RECT 4.400 490.600 409.795 492.000 ;
        RECT 4.000 487.920 409.795 490.600 ;
        RECT 4.000 486.520 405.830 487.920 ;
        RECT 4.000 483.840 409.795 486.520 ;
        RECT 4.400 482.440 409.795 483.840 ;
        RECT 4.000 479.760 409.795 482.440 ;
        RECT 4.000 478.360 405.830 479.760 ;
        RECT 4.000 475.680 409.795 478.360 ;
        RECT 4.400 474.280 409.795 475.680 ;
        RECT 4.000 471.600 409.795 474.280 ;
        RECT 4.000 470.200 405.830 471.600 ;
        RECT 4.000 467.520 409.795 470.200 ;
        RECT 4.400 466.120 409.795 467.520 ;
        RECT 4.000 463.440 409.795 466.120 ;
        RECT 4.000 462.040 405.830 463.440 ;
        RECT 4.000 459.360 409.795 462.040 ;
        RECT 4.400 457.960 409.795 459.360 ;
        RECT 4.000 455.280 409.795 457.960 ;
        RECT 4.000 453.880 405.830 455.280 ;
        RECT 4.000 451.200 409.795 453.880 ;
        RECT 4.400 449.800 409.795 451.200 ;
        RECT 4.000 447.120 409.795 449.800 ;
        RECT 4.000 445.720 405.830 447.120 ;
        RECT 4.000 443.040 409.795 445.720 ;
        RECT 4.400 441.640 409.795 443.040 ;
        RECT 4.000 438.960 409.795 441.640 ;
        RECT 4.000 437.560 405.830 438.960 ;
        RECT 4.000 434.880 409.795 437.560 ;
        RECT 4.400 433.480 409.795 434.880 ;
        RECT 4.000 430.800 409.795 433.480 ;
        RECT 4.000 429.400 405.830 430.800 ;
        RECT 4.000 426.720 409.795 429.400 ;
        RECT 4.400 425.320 409.795 426.720 ;
        RECT 4.000 422.640 409.795 425.320 ;
        RECT 4.000 421.240 405.830 422.640 ;
        RECT 4.000 418.560 409.795 421.240 ;
        RECT 4.400 417.160 409.795 418.560 ;
        RECT 4.000 414.480 409.795 417.160 ;
        RECT 4.000 413.080 405.830 414.480 ;
        RECT 4.000 410.400 409.795 413.080 ;
        RECT 4.400 409.000 409.795 410.400 ;
        RECT 4.000 406.320 409.795 409.000 ;
        RECT 4.000 404.920 405.830 406.320 ;
        RECT 4.000 402.240 409.795 404.920 ;
        RECT 4.400 400.840 409.795 402.240 ;
        RECT 4.000 398.160 409.795 400.840 ;
        RECT 4.000 396.760 405.830 398.160 ;
        RECT 4.000 394.080 409.795 396.760 ;
        RECT 4.400 392.680 409.795 394.080 ;
        RECT 4.000 390.000 409.795 392.680 ;
        RECT 4.000 388.600 405.830 390.000 ;
        RECT 4.000 385.920 409.795 388.600 ;
        RECT 4.400 384.520 409.795 385.920 ;
        RECT 4.000 381.840 409.795 384.520 ;
        RECT 4.000 380.440 405.830 381.840 ;
        RECT 4.000 377.760 409.795 380.440 ;
        RECT 4.400 376.360 409.795 377.760 ;
        RECT 4.000 373.680 409.795 376.360 ;
        RECT 4.000 372.280 405.830 373.680 ;
        RECT 4.000 369.600 409.795 372.280 ;
        RECT 4.400 368.200 409.795 369.600 ;
        RECT 4.000 365.520 409.795 368.200 ;
        RECT 4.000 364.120 405.830 365.520 ;
        RECT 4.000 361.440 409.795 364.120 ;
        RECT 4.400 360.040 409.795 361.440 ;
        RECT 4.000 357.360 409.795 360.040 ;
        RECT 4.000 355.960 405.830 357.360 ;
        RECT 4.000 353.280 409.795 355.960 ;
        RECT 4.400 351.880 409.795 353.280 ;
        RECT 4.000 349.200 409.795 351.880 ;
        RECT 4.000 347.800 405.830 349.200 ;
        RECT 4.000 345.120 409.795 347.800 ;
        RECT 4.400 343.720 409.795 345.120 ;
        RECT 4.000 341.040 409.795 343.720 ;
        RECT 4.000 339.640 405.830 341.040 ;
        RECT 4.000 336.960 409.795 339.640 ;
        RECT 4.400 335.560 409.795 336.960 ;
        RECT 4.000 332.880 409.795 335.560 ;
        RECT 4.000 331.480 405.830 332.880 ;
        RECT 4.000 328.800 409.795 331.480 ;
        RECT 4.400 327.400 409.795 328.800 ;
        RECT 4.000 324.720 409.795 327.400 ;
        RECT 4.000 323.320 405.830 324.720 ;
        RECT 4.000 320.640 409.795 323.320 ;
        RECT 4.400 319.240 409.795 320.640 ;
        RECT 4.000 316.560 409.795 319.240 ;
        RECT 4.000 315.160 405.830 316.560 ;
        RECT 4.000 312.480 409.795 315.160 ;
        RECT 4.400 311.080 409.795 312.480 ;
        RECT 4.000 308.400 409.795 311.080 ;
        RECT 4.000 307.000 405.830 308.400 ;
        RECT 4.000 304.320 409.795 307.000 ;
        RECT 4.400 302.920 409.795 304.320 ;
        RECT 4.000 300.240 409.795 302.920 ;
        RECT 4.000 298.840 405.830 300.240 ;
        RECT 4.000 296.160 409.795 298.840 ;
        RECT 4.400 294.760 409.795 296.160 ;
        RECT 4.000 292.080 409.795 294.760 ;
        RECT 4.000 290.680 405.830 292.080 ;
        RECT 4.000 288.000 409.795 290.680 ;
        RECT 4.400 286.600 409.795 288.000 ;
        RECT 4.000 283.920 409.795 286.600 ;
        RECT 4.000 282.520 405.830 283.920 ;
        RECT 4.000 279.840 409.795 282.520 ;
        RECT 4.400 278.440 409.795 279.840 ;
        RECT 4.000 275.760 409.795 278.440 ;
        RECT 4.000 274.360 405.830 275.760 ;
        RECT 4.000 271.680 409.795 274.360 ;
        RECT 4.400 270.280 409.795 271.680 ;
        RECT 4.000 267.600 409.795 270.280 ;
        RECT 4.000 266.200 405.830 267.600 ;
        RECT 4.000 263.520 409.795 266.200 ;
        RECT 4.400 262.120 409.795 263.520 ;
        RECT 4.000 259.440 409.795 262.120 ;
        RECT 4.000 258.040 405.830 259.440 ;
        RECT 4.000 255.360 409.795 258.040 ;
        RECT 4.400 253.960 409.795 255.360 ;
        RECT 4.000 251.280 409.795 253.960 ;
        RECT 4.000 249.880 405.830 251.280 ;
        RECT 4.000 247.200 409.795 249.880 ;
        RECT 4.400 245.800 409.795 247.200 ;
        RECT 4.000 243.120 409.795 245.800 ;
        RECT 4.000 241.720 405.830 243.120 ;
        RECT 4.000 239.040 409.795 241.720 ;
        RECT 4.400 237.640 409.795 239.040 ;
        RECT 4.000 234.960 409.795 237.640 ;
        RECT 4.000 233.560 405.830 234.960 ;
        RECT 4.000 230.880 409.795 233.560 ;
        RECT 4.400 229.480 409.795 230.880 ;
        RECT 4.000 226.800 409.795 229.480 ;
        RECT 4.000 225.400 405.830 226.800 ;
        RECT 4.000 222.720 409.795 225.400 ;
        RECT 4.400 221.320 409.795 222.720 ;
        RECT 4.000 218.640 409.795 221.320 ;
        RECT 4.000 217.240 405.830 218.640 ;
        RECT 4.000 214.560 409.795 217.240 ;
        RECT 4.400 213.160 409.795 214.560 ;
        RECT 4.000 210.480 409.795 213.160 ;
        RECT 4.000 209.080 405.830 210.480 ;
        RECT 4.000 206.400 409.795 209.080 ;
        RECT 4.400 205.000 409.795 206.400 ;
        RECT 4.000 202.320 409.795 205.000 ;
        RECT 4.000 200.920 405.830 202.320 ;
        RECT 4.000 198.240 409.795 200.920 ;
        RECT 4.400 196.840 409.795 198.240 ;
        RECT 4.000 194.160 409.795 196.840 ;
        RECT 4.000 192.760 405.830 194.160 ;
        RECT 4.000 190.080 409.795 192.760 ;
        RECT 4.400 188.680 409.795 190.080 ;
        RECT 4.000 186.000 409.795 188.680 ;
        RECT 4.000 184.600 405.830 186.000 ;
        RECT 4.000 181.920 409.795 184.600 ;
        RECT 4.400 180.520 409.795 181.920 ;
        RECT 4.000 177.840 409.795 180.520 ;
        RECT 4.000 176.440 405.830 177.840 ;
        RECT 4.000 173.760 409.795 176.440 ;
        RECT 4.400 172.360 409.795 173.760 ;
        RECT 4.000 169.680 409.795 172.360 ;
        RECT 4.000 168.280 405.830 169.680 ;
        RECT 4.000 165.600 409.795 168.280 ;
        RECT 4.400 164.200 409.795 165.600 ;
        RECT 4.000 161.520 409.795 164.200 ;
        RECT 4.000 160.120 405.830 161.520 ;
        RECT 4.000 157.440 409.795 160.120 ;
        RECT 4.400 156.040 409.795 157.440 ;
        RECT 4.000 153.360 409.795 156.040 ;
        RECT 4.000 151.960 405.830 153.360 ;
        RECT 4.000 149.280 409.795 151.960 ;
        RECT 4.400 147.880 409.795 149.280 ;
        RECT 4.000 145.200 409.795 147.880 ;
        RECT 4.000 143.800 405.830 145.200 ;
        RECT 4.000 141.120 409.795 143.800 ;
        RECT 4.400 139.720 409.795 141.120 ;
        RECT 4.000 137.040 409.795 139.720 ;
        RECT 4.000 135.640 405.830 137.040 ;
        RECT 4.000 132.960 409.795 135.640 ;
        RECT 4.400 131.560 409.795 132.960 ;
        RECT 4.000 128.880 409.795 131.560 ;
        RECT 4.000 127.480 405.830 128.880 ;
        RECT 4.000 124.800 409.795 127.480 ;
        RECT 4.400 123.400 409.795 124.800 ;
        RECT 4.000 120.720 409.795 123.400 ;
        RECT 4.000 119.320 405.830 120.720 ;
        RECT 4.000 116.640 409.795 119.320 ;
        RECT 4.400 115.240 409.795 116.640 ;
        RECT 4.000 112.560 409.795 115.240 ;
        RECT 4.000 111.160 405.830 112.560 ;
        RECT 4.000 108.480 409.795 111.160 ;
        RECT 4.400 107.080 409.795 108.480 ;
        RECT 4.000 104.400 409.795 107.080 ;
        RECT 4.000 103.000 405.830 104.400 ;
        RECT 4.000 100.320 409.795 103.000 ;
        RECT 4.400 98.920 409.795 100.320 ;
        RECT 4.000 96.240 409.795 98.920 ;
        RECT 4.000 94.840 405.830 96.240 ;
        RECT 4.000 92.160 409.795 94.840 ;
        RECT 4.400 90.760 409.795 92.160 ;
        RECT 4.000 88.080 409.795 90.760 ;
        RECT 4.000 86.680 405.830 88.080 ;
        RECT 4.000 84.000 409.795 86.680 ;
        RECT 4.400 82.600 409.795 84.000 ;
        RECT 4.000 79.920 409.795 82.600 ;
        RECT 4.000 78.520 405.830 79.920 ;
        RECT 4.000 75.840 409.795 78.520 ;
        RECT 4.400 74.440 409.795 75.840 ;
        RECT 4.000 71.760 409.795 74.440 ;
        RECT 4.000 70.360 405.830 71.760 ;
        RECT 4.000 67.680 409.795 70.360 ;
        RECT 4.400 66.280 409.795 67.680 ;
        RECT 4.000 63.600 409.795 66.280 ;
        RECT 4.000 62.200 405.830 63.600 ;
        RECT 4.000 59.520 409.795 62.200 ;
        RECT 4.400 58.120 409.795 59.520 ;
        RECT 4.000 55.440 409.795 58.120 ;
        RECT 4.000 54.040 405.830 55.440 ;
        RECT 4.000 51.360 409.795 54.040 ;
        RECT 4.400 49.960 409.795 51.360 ;
        RECT 4.000 47.280 409.795 49.960 ;
        RECT 4.000 45.880 405.830 47.280 ;
        RECT 4.000 43.200 409.795 45.880 ;
        RECT 4.400 41.800 409.795 43.200 ;
        RECT 4.000 39.120 409.795 41.800 ;
        RECT 4.000 37.720 405.830 39.120 ;
        RECT 4.000 35.040 409.795 37.720 ;
        RECT 4.400 33.640 409.795 35.040 ;
        RECT 4.000 30.960 409.795 33.640 ;
        RECT 4.000 29.560 405.830 30.960 ;
        RECT 4.000 26.880 409.795 29.560 ;
        RECT 4.400 25.480 409.795 26.880 ;
        RECT 4.000 22.800 409.795 25.480 ;
        RECT 4.000 21.400 405.830 22.800 ;
        RECT 4.000 18.720 409.795 21.400 ;
        RECT 4.400 17.320 409.795 18.720 ;
        RECT 4.000 14.640 409.795 17.320 ;
        RECT 4.000 13.240 405.830 14.640 ;
        RECT 4.000 10.560 409.795 13.240 ;
        RECT 4.400 9.160 409.795 10.560 ;
        RECT 4.000 7.655 409.795 9.160 ;
      LAYER met4 ;
        RECT 8.575 13.095 20.640 534.985 ;
        RECT 23.040 13.095 59.040 534.985 ;
        RECT 61.440 13.095 97.440 534.985 ;
        RECT 99.840 13.095 135.840 534.985 ;
        RECT 138.240 13.095 174.240 534.985 ;
        RECT 176.640 13.095 212.640 534.985 ;
        RECT 215.040 13.095 251.040 534.985 ;
        RECT 253.440 13.095 289.440 534.985 ;
        RECT 291.840 13.095 327.840 534.985 ;
        RECT 330.240 13.095 366.240 534.985 ;
        RECT 368.640 13.095 401.745 534.985 ;
  END
END housekeeping_alt
END LIBRARY

