VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3165.000 BY 4767.000 ;
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 725.135 -2.000 725.415 4.000 ;
    END
  END clock_core
  PIN flash_clk_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1597.335 -2.000 1597.615 4.000 ;
    END
  END flash_clk_frame
  PIN flash_clk_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1612.975 -2.000 1613.255 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb_frame
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1323.335 -2.000 1323.615 4.000 ;
    END
  END flash_csb_frame
  PIN flash_csb_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1338.975 -2.000 1339.255 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1816.135 -2.000 1816.415 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1871.335 -2.000 1871.615 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1849.715 -2.000 1849.995 4.000 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1886.975 -2.000 1887.255 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2090.135 -2.000 2090.415 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2145.335 -2.000 2145.615 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2123.715 -2.000 2123.995 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2160.975 -2.000 2161.255 4.000 ;
    END
  END flash_io1_oeb
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2364.135 -2.000 2364.415 4.000 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2397.715 -2.000 2397.995 4.000 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2391.735 -2.000 2392.015 4.000 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2413.355 -2.000 2413.635 4.000 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2419.335 -2.000 2419.615 4.000 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2434.975 -2.000 2435.255 4.000 ;
    END
  END gpio_outenb_core
  PIN mprj_analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2545.395 3167.185 2545.995 ;
    END
  END mprj_analog_io[0]
  PIN mprj_analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2215.165 4763.000 2215.445 4768.935 ;
    END
  END mprj_analog_io[10]
  PIN mprj_analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1770.165 4763.000 1770.445 4768.935 ;
    END
  END mprj_analog_io[11]
  PIN mprj_analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1261.165 4763.000 1261.445 4768.935 ;
    END
  END mprj_analog_io[12]
  PIN mprj_analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1003.165 4763.000 1003.445 4768.935 ;
    END
  END mprj_analog_io[13]
  PIN mprj_analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 746.165 4763.000 746.445 4768.935 ;
    END
  END mprj_analog_io[14]
  PIN mprj_analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 489.165 4763.000 489.445 4768.935 ;
    END
  END mprj_analog_io[15]
  PIN mprj_analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 232.165 4763.000 232.445 4768.935 ;
    END
  END mprj_analog_io[16]
  PIN mprj_analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4623.005 4.000 4623.605 ;
    END
  END mprj_analog_io[17]
  PIN mprj_analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3774.005 4.000 3774.605 ;
    END
  END mprj_analog_io[18]
  PIN mprj_analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3558.005 4.000 3558.605 ;
    END
  END mprj_analog_io[19]
  PIN mprj_analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2771.395 3167.185 2771.995 ;
    END
  END mprj_analog_io[1]
  PIN mprj_analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3342.005 4.000 3342.605 ;
    END
  END mprj_analog_io[20]
  PIN mprj_analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3126.005 4.000 3126.605 ;
    END
  END mprj_analog_io[21]
  PIN mprj_analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2910.005 4.000 2910.605 ;
    END
  END mprj_analog_io[22]
  PIN mprj_analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2694.005 4.000 2694.605 ;
    END
  END mprj_analog_io[23]
  PIN mprj_analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2478.005 4.000 2478.605 ;
    END
  END mprj_analog_io[24]
  PIN mprj_analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1840.005 4.000 1840.605 ;
    END
  END mprj_analog_io[25]
  PIN mprj_analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1624.005 4.000 1624.605 ;
    END
  END mprj_analog_io[26]
  PIN mprj_analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1408.005 4.000 1408.605 ;
    END
  END mprj_analog_io[27]
  PIN mprj_analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1192.005 4.000 1192.605 ;
    END
  END mprj_analog_io[28]
  PIN mprj_analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2996.395 3167.185 2996.995 ;
    END
  END mprj_analog_io[2]
  PIN mprj_analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3222.395 3167.185 3222.995 ;
    END
  END mprj_analog_io[3]
  PIN mprj_analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3447.395 3167.185 3447.995 ;
    END
  END mprj_analog_io[4]
  PIN mprj_analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3672.395 3167.185 3672.995 ;
    END
  END mprj_analog_io[5]
  PIN mprj_analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4118.395 3167.185 4118.995 ;
    END
  END mprj_analog_io[6]
  PIN mprj_analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4564.395 3167.185 4564.995 ;
    END
  END mprj_analog_io[7]
  PIN mprj_analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2981.165 4763.000 2981.445 4768.935 ;
    END
  END mprj_analog_io[8]
  PIN mprj_analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2472.165 4763.000 2472.445 4768.935 ;
    END
  END mprj_analog_io[9]
  PIN mprj_io_analog_en[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 318.355 3167.185 318.955 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_en[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3234.355 3167.185 3234.955 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_en[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3459.355 3167.185 3459.955 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_en[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3684.355 3167.185 3684.955 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_en[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4130.355 3167.185 4130.955 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_en[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4576.355 3167.185 4576.955 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_en[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2969.205 4763.000 2969.485 4768.935 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_en[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2460.205 4763.000 2460.485 4768.935 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_en[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2203.205 4763.000 2203.485 4768.935 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_en[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1758.205 4763.000 1758.485 4768.935 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_en[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1249.205 4763.000 1249.485 4768.935 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_en[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 544.355 3167.185 544.955 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_en[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 991.205 4763.000 991.485 4768.935 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_en[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 734.205 4763.000 734.485 4768.935 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_en[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 477.205 4763.000 477.485 4768.935 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_en[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 220.205 4763.000 220.485 4768.935 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_en[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4611.045 4.000 4611.645 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_en[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3762.045 4.000 3762.645 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_en[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3546.045 4.000 3546.645 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_en[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3330.045 4.000 3330.645 ;
    END
  END mprj_io_analog_en[27]
  PIN mprj_io_analog_en[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3114.045 4.000 3114.645 ;
    END
  END mprj_io_analog_en[28]
  PIN mprj_io_analog_en[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2898.045 4.000 2898.645 ;
    END
  END mprj_io_analog_en[29]
  PIN mprj_io_analog_en[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 769.355 3167.185 769.955 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_en[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2682.045 4.000 2682.645 ;
    END
  END mprj_io_analog_en[30]
  PIN mprj_io_analog_en[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2466.045 4.000 2466.645 ;
    END
  END mprj_io_analog_en[31]
  PIN mprj_io_analog_en[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1828.045 4.000 1828.645 ;
    END
  END mprj_io_analog_en[32]
  PIN mprj_io_analog_en[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1612.045 4.000 1612.645 ;
    END
  END mprj_io_analog_en[33]
  PIN mprj_io_analog_en[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1396.045 4.000 1396.645 ;
    END
  END mprj_io_analog_en[34]
  PIN mprj_io_analog_en[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1180.045 4.000 1180.645 ;
    END
  END mprj_io_analog_en[35]
  PIN mprj_io_analog_en[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 964.045 4.000 964.645 ;
    END
  END mprj_io_analog_en[36]
  PIN mprj_io_analog_en[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 748.045 4.000 748.645 ;
    END
  END mprj_io_analog_en[37]
  PIN mprj_io_analog_en[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 995.355 3167.185 995.955 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_en[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1220.355 3167.185 1220.955 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_en[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1445.355 3167.185 1445.955 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_en[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1671.355 3167.185 1671.955 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_en[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2557.355 3167.185 2557.955 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_en[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2783.355 3167.185 2783.955 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_en[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3008.355 3167.185 3008.955 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 324.795 3167.185 325.395 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_pol[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3240.795 3167.185 3241.395 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_pol[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3465.795 3167.185 3466.395 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_pol[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3690.795 3167.185 3691.395 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_pol[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4136.795 3167.185 4137.395 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_pol[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4582.795 3167.185 4583.395 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_pol[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2962.765 4763.000 2963.045 4768.935 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_pol[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2453.765 4763.000 2454.045 4768.935 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_pol[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2196.765 4763.000 2197.045 4768.935 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_pol[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1751.765 4763.000 1752.045 4768.935 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_pol[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1242.765 4763.000 1243.045 4768.935 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_pol[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 550.795 3167.185 551.395 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_pol[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 984.765 4763.000 985.045 4768.935 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_pol[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 727.765 4763.000 728.045 4768.935 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_pol[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 470.765 4763.000 471.045 4768.935 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_pol[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 213.765 4763.000 214.045 4768.935 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_pol[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4604.605 4.000 4605.205 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_pol[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3755.605 4.000 3756.205 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_pol[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3539.605 4.000 3540.205 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_pol[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3323.605 4.290 3324.205 ;
    END
  END mprj_io_analog_pol[27]
  PIN mprj_io_analog_pol[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3107.605 4.000 3108.205 ;
    END
  END mprj_io_analog_pol[28]
  PIN mprj_io_analog_pol[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2891.605 4.000 2892.205 ;
    END
  END mprj_io_analog_pol[29]
  PIN mprj_io_analog_pol[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 775.795 3167.185 776.395 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_pol[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2675.605 4.000 2676.205 ;
    END
  END mprj_io_analog_pol[30]
  PIN mprj_io_analog_pol[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2459.605 4.000 2460.205 ;
    END
  END mprj_io_analog_pol[31]
  PIN mprj_io_analog_pol[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1821.605 4.000 1822.205 ;
    END
  END mprj_io_analog_pol[32]
  PIN mprj_io_analog_pol[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1605.605 4.000 1606.205 ;
    END
  END mprj_io_analog_pol[33]
  PIN mprj_io_analog_pol[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1389.605 4.000 1390.205 ;
    END
  END mprj_io_analog_pol[34]
  PIN mprj_io_analog_pol[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1173.605 4.000 1174.205 ;
    END
  END mprj_io_analog_pol[35]
  PIN mprj_io_analog_pol[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 957.605 4.000 958.205 ;
    END
  END mprj_io_analog_pol[36]
  PIN mprj_io_analog_pol[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 741.605 4.000 742.205 ;
    END
  END mprj_io_analog_pol[37]
  PIN mprj_io_analog_pol[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1001.795 3167.185 1002.395 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_pol[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1226.795 3167.185 1227.395 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_pol[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1451.795 3167.185 1452.395 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_pol[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1677.795 3167.185 1678.395 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_pol[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2563.795 3167.185 2564.395 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_pol[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2789.795 3167.185 2790.395 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_pol[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3014.795 3167.185 3015.395 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 339.975 3167.185 340.575 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_analog_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3255.975 3167.185 3256.575 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_analog_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3480.975 3167.185 3481.575 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_analog_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3705.975 3167.185 3706.575 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_analog_sel[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4151.975 3167.185 4152.575 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_analog_sel[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4597.975 3167.185 4598.575 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_analog_sel[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2947.585 4763.000 2947.865 4768.935 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_analog_sel[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2438.585 4763.000 2438.865 4768.935 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_analog_sel[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2181.585 4763.000 2181.865 4768.935 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_analog_sel[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1736.585 4763.000 1736.865 4768.935 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_analog_sel[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1227.585 4763.000 1227.865 4768.935 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_analog_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 565.975 3167.185 566.575 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_analog_sel[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 969.585 4763.000 969.865 4768.935 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_analog_sel[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 712.585 4763.000 712.865 4768.935 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_analog_sel[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 455.585 4763.000 455.865 4768.935 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_analog_sel[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 198.585 4763.000 198.865 4768.935 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_analog_sel[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4589.425 4.000 4590.025 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_analog_sel[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3740.425 4.000 3741.025 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_analog_sel[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3524.425 4.000 3525.025 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_analog_sel[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3308.425 4.000 3309.025 ;
    END
  END mprj_io_analog_sel[27]
  PIN mprj_io_analog_sel[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3092.425 4.000 3093.025 ;
    END
  END mprj_io_analog_sel[28]
  PIN mprj_io_analog_sel[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2876.425 4.000 2877.025 ;
    END
  END mprj_io_analog_sel[29]
  PIN mprj_io_analog_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 790.975 3167.185 791.575 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_analog_sel[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2660.425 4.000 2661.025 ;
    END
  END mprj_io_analog_sel[30]
  PIN mprj_io_analog_sel[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2444.425 4.000 2445.025 ;
    END
  END mprj_io_analog_sel[31]
  PIN mprj_io_analog_sel[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1806.425 4.000 1807.025 ;
    END
  END mprj_io_analog_sel[32]
  PIN mprj_io_analog_sel[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1590.425 4.000 1591.025 ;
    END
  END mprj_io_analog_sel[33]
  PIN mprj_io_analog_sel[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1374.425 4.000 1375.025 ;
    END
  END mprj_io_analog_sel[34]
  PIN mprj_io_analog_sel[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1158.425 4.000 1159.025 ;
    END
  END mprj_io_analog_sel[35]
  PIN mprj_io_analog_sel[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 942.425 4.000 943.025 ;
    END
  END mprj_io_analog_sel[36]
  PIN mprj_io_analog_sel[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 726.425 4.000 727.025 ;
    END
  END mprj_io_analog_sel[37]
  PIN mprj_io_analog_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1016.975 3167.185 1017.575 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_analog_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1241.975 3167.185 1242.575 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_analog_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1466.975 3167.185 1467.575 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_analog_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1692.975 3167.185 1693.575 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_analog_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2578.975 3167.185 2579.575 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_analog_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2804.975 3167.185 2805.575 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_analog_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3029.975 3167.185 3030.575 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 321.575 3167.185 322.175 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1618.025 4.000 1618.625 ;
    END
  END mprj_io_dm[100]
  PIN mprj_io_dm[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1587.205 4.000 1587.805 ;
    END
  END mprj_io_dm[101]
  PIN mprj_io_dm[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1392.825 4.000 1393.425 ;
    END
  END mprj_io_dm[102]
  PIN mprj_io_dm[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1402.025 4.000 1402.625 ;
    END
  END mprj_io_dm[103]
  PIN mprj_io_dm[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1371.205 4.000 1371.805 ;
    END
  END mprj_io_dm[104]
  PIN mprj_io_dm[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1176.825 4.000 1177.425 ;
    END
  END mprj_io_dm[105]
  PIN mprj_io_dm[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1186.025 4.000 1186.625 ;
    END
  END mprj_io_dm[106]
  PIN mprj_io_dm[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1155.205 4.000 1155.805 ;
    END
  END mprj_io_dm[107]
  PIN mprj_io_dm[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 960.825 4.000 961.425 ;
    END
  END mprj_io_dm[108]
  PIN mprj_io_dm[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 970.025 4.000 970.625 ;
    END
  END mprj_io_dm[109]
  PIN mprj_io_dm[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 989.375 3167.185 989.975 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 939.205 4.000 939.805 ;
    END
  END mprj_io_dm[110]
  PIN mprj_io_dm[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 744.825 4.000 745.425 ;
    END
  END mprj_io_dm[111]
  PIN mprj_io_dm[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 754.025 4.000 754.625 ;
    END
  END mprj_io_dm[112]
  PIN mprj_io_dm[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 723.205 4.000 723.805 ;
    END
  END mprj_io_dm[113]
  PIN mprj_io_dm[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1020.195 3167.185 1020.795 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1223.575 3167.185 1224.175 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1214.375 3167.185 1214.975 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1245.195 3167.185 1245.795 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_dm[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1448.575 3167.185 1449.175 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1439.375 3167.185 1439.975 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1470.195 3167.185 1470.795 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_dm[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1674.575 3167.185 1675.175 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1665.375 3167.185 1665.975 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 312.375 3167.185 312.975 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1696.195 3167.185 1696.795 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_dm[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2560.575 3167.185 2561.175 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2551.375 3167.185 2551.975 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2582.195 3167.185 2582.795 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_dm[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2786.575 3167.185 2787.175 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2777.375 3167.185 2777.975 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2808.195 3167.185 2808.795 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_dm[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3011.575 3167.185 3012.175 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3002.375 3167.185 3002.975 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3033.195 3167.185 3033.795 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_dm[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 343.195 3167.185 343.795 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_dm[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3237.575 3167.185 3238.175 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3228.375 3167.185 3228.975 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3259.195 3167.185 3259.795 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_dm[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3462.575 3167.185 3463.175 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3453.375 3167.185 3453.975 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3484.195 3167.185 3484.795 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_dm[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3687.575 3167.185 3688.175 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3678.375 3167.185 3678.975 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3709.195 3167.185 3709.795 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_dm[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4133.575 3167.185 4134.175 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 547.575 3167.185 548.175 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4124.375 3167.185 4124.975 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4155.195 3167.185 4155.795 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_dm[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4579.575 3167.185 4580.175 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4570.375 3167.185 4570.975 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4601.195 3167.185 4601.795 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_dm[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2965.985 4763.000 2966.265 4768.935 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2975.185 4763.000 2975.465 4768.935 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2944.365 4763.000 2944.645 4768.935 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_dm[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2456.985 4763.000 2457.265 4768.935 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2466.185 4763.000 2466.465 4768.935 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 538.375 3167.185 538.975 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2435.365 4763.000 2435.645 4768.935 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_dm[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2199.985 4763.000 2200.265 4768.935 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2209.185 4763.000 2209.465 4768.935 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2178.365 4763.000 2178.645 4768.935 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_dm[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1754.985 4763.000 1755.265 4768.935 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1764.185 4763.000 1764.465 4768.935 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1733.365 4763.000 1733.645 4768.935 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_dm[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1245.985 4763.000 1246.265 4768.935 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1255.185 4763.000 1255.465 4768.935 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1224.365 4763.000 1224.645 4768.935 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_dm[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 569.195 3167.185 569.795 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_dm[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 987.985 4763.000 988.265 4768.935 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 997.185 4763.000 997.465 4768.935 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 966.365 4763.000 966.645 4768.935 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_dm[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 730.985 4763.000 731.265 4768.935 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 740.185 4763.000 740.465 4768.935 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 709.365 4763.000 709.645 4768.935 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_dm[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 473.985 4763.000 474.265 4768.935 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 483.185 4763.000 483.465 4768.935 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 452.365 4763.000 452.645 4768.935 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_dm[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 216.985 4763.000 217.265 4768.935 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 772.575 3167.185 773.175 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 226.185 4763.000 226.465 4768.935 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 195.365 4763.000 195.645 4768.935 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_dm[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4607.825 4.000 4608.425 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4617.025 4.000 4617.625 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4586.205 4.000 4586.805 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_dm[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3758.825 4.000 3759.425 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3768.025 4.000 3768.625 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3737.205 4.000 3737.805 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_dm[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3542.825 4.000 3543.425 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3552.025 4.000 3552.625 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 763.375 3167.185 763.975 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3521.205 4.000 3521.805 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_dm[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3326.825 4.000 3327.425 ;
    END
  END mprj_io_dm[81]
  PIN mprj_io_dm[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3336.025 4.000 3336.625 ;
    END
  END mprj_io_dm[82]
  PIN mprj_io_dm[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3305.205 4.000 3305.805 ;
    END
  END mprj_io_dm[83]
  PIN mprj_io_dm[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3110.825 4.000 3111.425 ;
    END
  END mprj_io_dm[84]
  PIN mprj_io_dm[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3120.025 4.000 3120.625 ;
    END
  END mprj_io_dm[85]
  PIN mprj_io_dm[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3089.205 4.000 3089.805 ;
    END
  END mprj_io_dm[86]
  PIN mprj_io_dm[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2894.825 4.000 2895.425 ;
    END
  END mprj_io_dm[87]
  PIN mprj_io_dm[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2904.025 4.000 2904.625 ;
    END
  END mprj_io_dm[88]
  PIN mprj_io_dm[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2873.205 4.000 2873.805 ;
    END
  END mprj_io_dm[89]
  PIN mprj_io_dm[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 794.195 3167.185 794.795 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_dm[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2678.825 4.000 2679.425 ;
    END
  END mprj_io_dm[90]
  PIN mprj_io_dm[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2688.025 4.000 2688.625 ;
    END
  END mprj_io_dm[91]
  PIN mprj_io_dm[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2657.205 4.000 2657.805 ;
    END
  END mprj_io_dm[92]
  PIN mprj_io_dm[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2462.825 4.000 2463.425 ;
    END
  END mprj_io_dm[93]
  PIN mprj_io_dm[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2472.025 4.000 2472.625 ;
    END
  END mprj_io_dm[94]
  PIN mprj_io_dm[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2441.205 4.000 2441.805 ;
    END
  END mprj_io_dm[95]
  PIN mprj_io_dm[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1824.825 4.000 1825.425 ;
    END
  END mprj_io_dm[96]
  PIN mprj_io_dm[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1834.025 4.000 1834.625 ;
    END
  END mprj_io_dm[97]
  PIN mprj_io_dm[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1803.205 4.000 1803.805 ;
    END
  END mprj_io_dm[98]
  PIN mprj_io_dm[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1608.825 4.000 1609.425 ;
    END
  END mprj_io_dm[99]
  PIN mprj_io_dm[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 998.575 3167.185 999.175 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 346.415 3167.185 347.015 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_holdover[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3262.415 3167.185 3263.015 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_holdover[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3487.415 3167.185 3488.015 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_holdover[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3712.415 3167.185 3713.015 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_holdover[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4158.415 3167.185 4159.015 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_holdover[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4604.415 3167.185 4605.015 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_holdover[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2941.145 4763.000 2941.425 4768.935 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_holdover[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2432.145 4763.000 2432.425 4768.935 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_holdover[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2175.145 4763.000 2175.425 4768.935 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_holdover[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1730.145 4763.000 1730.425 4768.935 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_holdover[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1221.145 4763.000 1221.425 4768.935 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_holdover[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 572.415 3167.185 573.015 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_holdover[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 963.145 4763.000 963.425 4768.935 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_holdover[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 706.145 4763.000 706.425 4768.935 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_holdover[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 449.145 4763.000 449.425 4768.935 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_holdover[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 192.145 4763.000 192.425 4768.935 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_holdover[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4582.985 4.000 4583.585 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_holdover[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3733.985 4.000 3734.585 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_holdover[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3517.985 4.000 3518.585 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_holdover[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3301.985 4.000 3302.585 ;
    END
  END mprj_io_holdover[27]
  PIN mprj_io_holdover[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3085.985 4.000 3086.585 ;
    END
  END mprj_io_holdover[28]
  PIN mprj_io_holdover[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2869.985 4.000 2870.585 ;
    END
  END mprj_io_holdover[29]
  PIN mprj_io_holdover[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 797.415 3167.185 798.015 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_holdover[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2653.985 4.000 2654.585 ;
    END
  END mprj_io_holdover[30]
  PIN mprj_io_holdover[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2437.985 4.000 2438.585 ;
    END
  END mprj_io_holdover[31]
  PIN mprj_io_holdover[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1799.985 4.000 1800.585 ;
    END
  END mprj_io_holdover[32]
  PIN mprj_io_holdover[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1583.985 4.000 1584.585 ;
    END
  END mprj_io_holdover[33]
  PIN mprj_io_holdover[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1367.985 4.000 1368.585 ;
    END
  END mprj_io_holdover[34]
  PIN mprj_io_holdover[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1151.985 4.000 1152.585 ;
    END
  END mprj_io_holdover[35]
  PIN mprj_io_holdover[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 935.985 4.000 936.585 ;
    END
  END mprj_io_holdover[36]
  PIN mprj_io_holdover[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 719.985 4.000 720.585 ;
    END
  END mprj_io_holdover[37]
  PIN mprj_io_holdover[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1023.415 3167.185 1024.015 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_holdover[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1248.415 3167.185 1249.015 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_holdover[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1473.415 3167.185 1474.015 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_holdover[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1699.415 3167.185 1700.015 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_holdover[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2585.415 3167.185 2586.015 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_holdover[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2811.415 3167.185 2812.015 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_holdover[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3036.415 3167.185 3037.015 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 361.595 3167.185 362.195 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3277.595 3167.185 3278.195 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3502.595 3167.185 3503.195 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3727.595 3167.185 3728.195 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4173.595 3167.185 4174.195 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4619.595 3167.185 4620.195 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2925.965 4763.000 2926.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2416.965 4763.000 2417.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2159.965 4763.000 2160.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1714.965 4763.000 1715.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1205.965 4763.000 1206.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 587.595 3167.185 588.195 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 947.965 4763.000 948.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 690.965 4763.000 691.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 433.965 4763.000 434.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 176.965 4763.000 177.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4567.805 4.000 4568.405 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3718.805 4.000 3719.405 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3502.805 4.000 3503.405 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_ib_mode_sel[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3286.805 4.000 3287.405 ;
    END
  END mprj_io_ib_mode_sel[27]
  PIN mprj_io_ib_mode_sel[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3070.805 4.000 3071.405 ;
    END
  END mprj_io_ib_mode_sel[28]
  PIN mprj_io_ib_mode_sel[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2854.805 4.000 2855.405 ;
    END
  END mprj_io_ib_mode_sel[29]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 812.595 3167.185 813.195 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_ib_mode_sel[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2638.805 4.000 2639.405 ;
    END
  END mprj_io_ib_mode_sel[30]
  PIN mprj_io_ib_mode_sel[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2422.805 4.000 2423.405 ;
    END
  END mprj_io_ib_mode_sel[31]
  PIN mprj_io_ib_mode_sel[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1784.805 4.000 1785.405 ;
    END
  END mprj_io_ib_mode_sel[32]
  PIN mprj_io_ib_mode_sel[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1568.805 4.000 1569.405 ;
    END
  END mprj_io_ib_mode_sel[33]
  PIN mprj_io_ib_mode_sel[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1352.805 4.000 1353.405 ;
    END
  END mprj_io_ib_mode_sel[34]
  PIN mprj_io_ib_mode_sel[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1136.805 4.000 1137.405 ;
    END
  END mprj_io_ib_mode_sel[35]
  PIN mprj_io_ib_mode_sel[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 920.805 4.000 921.405 ;
    END
  END mprj_io_ib_mode_sel[36]
  PIN mprj_io_ib_mode_sel[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 704.805 4.290 705.405 ;
    END
  END mprj_io_ib_mode_sel[37]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1038.595 3167.185 1039.195 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1263.595 3167.185 1264.195 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1488.595 3167.185 1489.195 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1714.595 3167.185 1715.195 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2600.595 3167.185 2601.195 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2826.595 3167.185 2827.195 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3051.595 3167.185 3052.195 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 293.975 3167.185 294.575 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3209.975 3167.185 3210.575 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3434.975 3167.185 3435.575 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3659.975 3167.185 3660.575 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4105.975 3167.185 4106.575 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4551.975 3167.185 4552.575 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2993.585 4763.000 2993.865 4768.935 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2484.585 4763.000 2484.865 4768.935 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2227.585 4763.000 2227.865 4768.935 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1782.585 4763.000 1782.865 4768.935 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1273.585 4763.000 1273.865 4768.935 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 519.975 3167.185 520.575 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1015.585 4763.000 1015.865 4768.935 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 758.585 4763.000 758.865 4768.935 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 501.585 4763.000 501.865 4768.935 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 244.585 4763.000 244.865 4768.935 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4635.425 4.000 4636.025 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3786.425 4.000 3787.025 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3570.425 4.000 3571.025 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3354.425 4.000 3355.025 ;
    END
  END mprj_io_in[27]
  PIN mprj_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3138.425 4.000 3139.025 ;
    END
  END mprj_io_in[28]
  PIN mprj_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2922.425 4.000 2923.025 ;
    END
  END mprj_io_in[29]
  PIN mprj_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 744.975 3167.185 745.575 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2706.425 4.000 2707.025 ;
    END
  END mprj_io_in[30]
  PIN mprj_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2490.425 4.000 2491.025 ;
    END
  END mprj_io_in[31]
  PIN mprj_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1852.425 4.000 1853.025 ;
    END
  END mprj_io_in[32]
  PIN mprj_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1636.425 4.000 1637.025 ;
    END
  END mprj_io_in[33]
  PIN mprj_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1420.425 4.000 1421.025 ;
    END
  END mprj_io_in[34]
  PIN mprj_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1204.425 4.000 1205.025 ;
    END
  END mprj_io_in[35]
  PIN mprj_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 988.425 4.000 989.025 ;
    END
  END mprj_io_in[36]
  PIN mprj_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT -2.185 772.425 4.000 773.025 ;
    END
  END mprj_io_in[37]
  PIN mprj_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 970.975 3167.185 971.575 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1195.975 3167.185 1196.575 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1420.975 3167.185 1421.575 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1646.975 3167.185 1647.575 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2532.975 3167.185 2533.575 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2758.975 3167.185 2759.575 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2983.975 3167.185 2984.575 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_inp_dis[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 327.555 3167.185 328.155 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_inp_dis[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3243.555 3167.185 3244.155 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_inp_dis[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3468.555 3167.185 3469.155 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_inp_dis[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3693.555 3167.185 3694.155 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_inp_dis[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4139.555 3167.185 4140.155 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_inp_dis[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4585.555 3167.185 4586.155 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_inp_dis[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2960.005 4763.000 2960.285 4768.935 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_inp_dis[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2451.005 4763.000 2451.285 4768.935 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_inp_dis[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2194.005 4763.000 2194.285 4768.935 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_inp_dis[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1749.005 4763.000 1749.285 4768.935 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_inp_dis[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1240.005 4763.000 1240.285 4768.935 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_inp_dis[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 553.555 3167.185 554.155 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_inp_dis[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 982.005 4763.000 982.285 4768.935 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_inp_dis[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 725.005 4763.000 725.285 4768.935 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_inp_dis[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 468.005 4763.000 468.285 4768.935 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_inp_dis[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 211.005 4763.000 211.285 4768.935 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_inp_dis[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4601.845 4.000 4602.445 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_inp_dis[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3752.845 4.000 3753.445 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_inp_dis[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3536.845 4.000 3537.445 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_inp_dis[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3320.845 4.000 3321.445 ;
    END
  END mprj_io_inp_dis[27]
  PIN mprj_io_inp_dis[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3104.845 4.000 3105.445 ;
    END
  END mprj_io_inp_dis[28]
  PIN mprj_io_inp_dis[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2888.845 4.000 2889.445 ;
    END
  END mprj_io_inp_dis[29]
  PIN mprj_io_inp_dis[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 778.555 3167.185 779.155 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_inp_dis[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2672.845 4.000 2673.445 ;
    END
  END mprj_io_inp_dis[30]
  PIN mprj_io_inp_dis[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2456.845 4.000 2457.445 ;
    END
  END mprj_io_inp_dis[31]
  PIN mprj_io_inp_dis[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1818.845 4.000 1819.445 ;
    END
  END mprj_io_inp_dis[32]
  PIN mprj_io_inp_dis[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1602.845 4.000 1603.445 ;
    END
  END mprj_io_inp_dis[33]
  PIN mprj_io_inp_dis[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1386.845 4.000 1387.445 ;
    END
  END mprj_io_inp_dis[34]
  PIN mprj_io_inp_dis[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1170.845 4.000 1171.445 ;
    END
  END mprj_io_inp_dis[35]
  PIN mprj_io_inp_dis[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 954.845 4.000 955.445 ;
    END
  END mprj_io_inp_dis[36]
  PIN mprj_io_inp_dis[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 738.845 4.000 739.445 ;
    END
  END mprj_io_inp_dis[37]
  PIN mprj_io_inp_dis[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1004.555 3167.185 1005.155 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_inp_dis[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1229.555 3167.185 1230.155 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_inp_dis[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1454.555 3167.185 1455.155 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_inp_dis[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1680.555 3167.185 1681.155 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_inp_dis[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2566.555 3167.185 2567.155 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_inp_dis[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2792.555 3167.185 2793.155 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_inp_dis[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3017.555 3167.185 3018.155 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 364.815 3167.185 365.415 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3280.815 3167.185 3281.415 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3505.815 3167.185 3506.415 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3730.815 3167.185 3731.415 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4176.815 3167.185 4177.415 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4622.815 3167.185 4623.415 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2922.745 4763.000 2923.025 4768.935 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2413.745 4763.000 2414.025 4768.935 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2156.745 4763.000 2157.025 4768.935 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1711.745 4763.000 1712.025 4768.935 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1202.745 4763.000 1203.025 4768.935 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 590.815 3167.185 591.415 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 944.745 4763.000 945.025 4768.935 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 687.745 4763.000 688.025 4768.935 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 430.745 4763.000 431.025 4768.935 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 173.745 4763.000 174.025 4768.935 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4564.585 4.000 4565.185 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3715.585 4.000 3716.185 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3499.585 4.000 3500.185 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3283.585 4.000 3284.185 ;
    END
  END mprj_io_oeb[27]
  PIN mprj_io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3067.585 4.000 3068.185 ;
    END
  END mprj_io_oeb[28]
  PIN mprj_io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2851.585 4.000 2852.185 ;
    END
  END mprj_io_oeb[29]
  PIN mprj_io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 815.815 3167.185 816.415 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2635.585 4.000 2636.185 ;
    END
  END mprj_io_oeb[30]
  PIN mprj_io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2419.585 4.000 2420.185 ;
    END
  END mprj_io_oeb[31]
  PIN mprj_io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1781.585 4.000 1782.185 ;
    END
  END mprj_io_oeb[32]
  PIN mprj_io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1565.585 4.000 1566.185 ;
    END
  END mprj_io_oeb[33]
  PIN mprj_io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1349.585 4.000 1350.185 ;
    END
  END mprj_io_oeb[34]
  PIN mprj_io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1133.585 4.000 1134.185 ;
    END
  END mprj_io_oeb[35]
  PIN mprj_io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 917.585 4.000 918.185 ;
    END
  END mprj_io_oeb[36]
  PIN mprj_io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 701.585 4.000 702.185 ;
    END
  END mprj_io_oeb[37]
  PIN mprj_io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1041.815 3167.185 1042.415 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1266.815 3167.185 1267.415 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1491.815 3167.185 1492.415 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1717.815 3167.185 1718.415 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2603.815 3167.185 2604.415 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2829.815 3167.185 2830.415 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3054.815 3167.185 3055.415 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_one[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 299.955 3167.185 300.555 ;
    END
  END mprj_io_one[0]
  PIN mprj_io_one[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3215.955 3167.185 3216.555 ;
    END
  END mprj_io_one[10]
  PIN mprj_io_one[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3440.955 3167.185 3441.555 ;
    END
  END mprj_io_one[11]
  PIN mprj_io_one[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3665.955 3167.185 3666.555 ;
    END
  END mprj_io_one[12]
  PIN mprj_io_one[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4111.955 3167.185 4112.555 ;
    END
  END mprj_io_one[13]
  PIN mprj_io_one[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4557.955 3167.185 4558.555 ;
    END
  END mprj_io_one[14]
  PIN mprj_io_one[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2987.605 4763.000 2987.885 4768.935 ;
    END
  END mprj_io_one[15]
  PIN mprj_io_one[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2478.605 4763.000 2478.885 4768.935 ;
    END
  END mprj_io_one[16]
  PIN mprj_io_one[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2221.605 4763.000 2221.885 4768.935 ;
    END
  END mprj_io_one[17]
  PIN mprj_io_one[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1776.605 4763.000 1776.885 4768.935 ;
    END
  END mprj_io_one[18]
  PIN mprj_io_one[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1267.605 4763.000 1267.885 4768.935 ;
    END
  END mprj_io_one[19]
  PIN mprj_io_one[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 525.955 3167.185 526.555 ;
    END
  END mprj_io_one[1]
  PIN mprj_io_one[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1009.605 4763.000 1009.885 4768.935 ;
    END
  END mprj_io_one[20]
  PIN mprj_io_one[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 752.605 4763.000 752.885 4768.935 ;
    END
  END mprj_io_one[21]
  PIN mprj_io_one[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 495.605 4763.000 495.885 4768.935 ;
    END
  END mprj_io_one[22]
  PIN mprj_io_one[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.605 4763.000 238.885 4768.935 ;
    END
  END mprj_io_one[23]
  PIN mprj_io_one[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4629.445 4.000 4630.045 ;
    END
  END mprj_io_one[24]
  PIN mprj_io_one[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3780.445 4.000 3781.045 ;
    END
  END mprj_io_one[25]
  PIN mprj_io_one[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3564.445 4.000 3565.045 ;
    END
  END mprj_io_one[26]
  PIN mprj_io_one[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3348.445 4.000 3349.045 ;
    END
  END mprj_io_one[27]
  PIN mprj_io_one[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3132.445 4.000 3133.045 ;
    END
  END mprj_io_one[28]
  PIN mprj_io_one[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2916.445 4.000 2917.045 ;
    END
  END mprj_io_one[29]
  PIN mprj_io_one[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 750.955 3167.185 751.555 ;
    END
  END mprj_io_one[2]
  PIN mprj_io_one[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2700.445 4.000 2701.045 ;
    END
  END mprj_io_one[30]
  PIN mprj_io_one[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2484.445 4.000 2485.045 ;
    END
  END mprj_io_one[31]
  PIN mprj_io_one[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1846.445 4.000 1847.045 ;
    END
  END mprj_io_one[32]
  PIN mprj_io_one[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1630.445 4.000 1631.045 ;
    END
  END mprj_io_one[33]
  PIN mprj_io_one[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1414.445 4.000 1415.045 ;
    END
  END mprj_io_one[34]
  PIN mprj_io_one[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1198.445 4.000 1199.045 ;
    END
  END mprj_io_one[35]
  PIN mprj_io_one[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 982.445 4.000 983.045 ;
    END
  END mprj_io_one[36]
  PIN mprj_io_one[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT -2.185 766.445 4.000 767.045 ;
    END
  END mprj_io_one[37]
  PIN mprj_io_one[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 976.955 3167.185 977.555 ;
    END
  END mprj_io_one[3]
  PIN mprj_io_one[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1201.955 3167.185 1202.555 ;
    END
  END mprj_io_one[4]
  PIN mprj_io_one[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1426.955 3167.185 1427.555 ;
    END
  END mprj_io_one[5]
  PIN mprj_io_one[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1652.955 3167.185 1653.555 ;
    END
  END mprj_io_one[6]
  PIN mprj_io_one[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2538.955 3167.185 2539.555 ;
    END
  END mprj_io_one[7]
  PIN mprj_io_one[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2764.955 3167.185 2765.555 ;
    END
  END mprj_io_one[8]
  PIN mprj_io_one[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2989.955 3167.185 2990.555 ;
    END
  END mprj_io_one[9]
  PIN mprj_io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 349.175 3167.185 349.775 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3265.175 3167.185 3265.775 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3490.175 3167.185 3490.775 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3715.175 3167.185 3715.775 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4161.175 3167.185 4161.775 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4607.175 3167.185 4607.775 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2938.385 4763.000 2938.665 4768.935 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2429.385 4763.000 2429.665 4768.935 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2172.385 4763.000 2172.665 4768.935 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1727.385 4763.000 1727.665 4768.935 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1218.385 4763.000 1218.665 4768.935 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 575.175 3167.185 575.775 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 960.385 4763.000 960.665 4768.935 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 703.385 4763.000 703.665 4768.935 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 446.385 4763.000 446.665 4768.935 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 189.385 4763.000 189.665 4768.935 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4580.225 4.000 4580.825 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3731.225 4.000 3731.825 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3515.225 4.000 3515.825 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3299.225 4.000 3299.825 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3083.225 4.000 3083.825 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2867.225 4.000 2867.825 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 800.175 3167.185 800.775 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2651.225 4.000 2651.825 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2435.225 4.000 2435.825 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1797.225 4.000 1797.825 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1581.225 4.000 1581.825 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1365.225 4.000 1365.825 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1149.225 4.000 1149.825 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 933.225 4.000 933.825 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 717.225 4.000 717.825 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1026.175 3167.185 1026.775 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1251.175 3167.185 1251.775 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1476.175 3167.185 1476.775 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1702.175 3167.185 1702.775 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2588.175 3167.185 2588.775 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2814.175 3167.185 2814.775 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3039.175 3167.185 3039.775 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 303.175 3167.185 303.775 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_slow_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3219.175 3167.185 3219.775 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_slow_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3444.175 3167.185 3444.775 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_slow_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3669.175 3167.185 3669.775 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_slow_sel[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4115.175 3167.185 4115.775 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_slow_sel[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4561.175 3167.185 4561.775 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_slow_sel[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2984.385 4763.000 2984.665 4768.935 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_slow_sel[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2475.385 4763.000 2475.665 4768.935 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_slow_sel[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2218.385 4763.000 2218.665 4768.935 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_slow_sel[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1773.385 4763.000 1773.665 4768.935 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_slow_sel[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1264.385 4763.000 1264.665 4768.935 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_slow_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 529.175 3167.185 529.775 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_slow_sel[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1006.385 4763.000 1006.665 4768.935 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_slow_sel[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 749.385 4763.000 749.665 4768.935 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_slow_sel[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 492.385 4763.000 492.665 4768.935 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_slow_sel[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 235.385 4763.000 235.665 4768.935 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_slow_sel[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4626.225 4.000 4626.825 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_slow_sel[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3777.225 4.000 3777.825 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_slow_sel[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3561.225 4.000 3561.825 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_slow_sel[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3345.225 4.000 3345.825 ;
    END
  END mprj_io_slow_sel[27]
  PIN mprj_io_slow_sel[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3129.225 4.000 3129.825 ;
    END
  END mprj_io_slow_sel[28]
  PIN mprj_io_slow_sel[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2913.225 4.000 2913.825 ;
    END
  END mprj_io_slow_sel[29]
  PIN mprj_io_slow_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 754.175 3167.185 754.775 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_slow_sel[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2697.225 4.000 2697.825 ;
    END
  END mprj_io_slow_sel[30]
  PIN mprj_io_slow_sel[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2481.225 4.000 2481.825 ;
    END
  END mprj_io_slow_sel[31]
  PIN mprj_io_slow_sel[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1843.225 4.000 1843.825 ;
    END
  END mprj_io_slow_sel[32]
  PIN mprj_io_slow_sel[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1627.225 4.000 1627.825 ;
    END
  END mprj_io_slow_sel[33]
  PIN mprj_io_slow_sel[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1411.225 4.000 1411.825 ;
    END
  END mprj_io_slow_sel[34]
  PIN mprj_io_slow_sel[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1195.225 4.000 1195.825 ;
    END
  END mprj_io_slow_sel[35]
  PIN mprj_io_slow_sel[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 979.225 4.000 979.825 ;
    END
  END mprj_io_slow_sel[36]
  PIN mprj_io_slow_sel[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 763.225 4.000 763.825 ;
    END
  END mprj_io_slow_sel[37]
  PIN mprj_io_slow_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 980.175 3167.185 980.775 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_slow_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1205.175 3167.185 1205.775 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_slow_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1430.175 3167.185 1430.775 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_slow_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1656.175 3167.185 1656.775 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_slow_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2542.175 3167.185 2542.775 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_slow_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2768.175 3167.185 2768.775 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_slow_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2993.175 3167.185 2993.775 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 358.375 3167.185 358.975 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3274.375 3167.185 3274.975 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3499.375 3167.185 3499.975 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3724.375 3167.185 3724.975 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4170.375 3167.185 4170.975 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4616.375 3167.185 4616.975 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2929.185 4763.000 2929.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2420.185 4763.000 2420.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2163.185 4763.000 2163.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1718.185 4763.000 1718.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1209.185 4763.000 1209.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 584.375 3167.185 584.975 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 951.185 4763.000 951.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 694.185 4763.000 694.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 437.185 4763.000 437.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 180.185 4763.000 180.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 4571.025 4.000 4571.625 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3722.025 4.000 3722.625 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3506.025 4.000 3506.625 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_vtrip_sel[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3290.025 4.000 3290.625 ;
    END
  END mprj_io_vtrip_sel[27]
  PIN mprj_io_vtrip_sel[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 3074.025 4.000 3074.625 ;
    END
  END mprj_io_vtrip_sel[28]
  PIN mprj_io_vtrip_sel[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2858.025 4.000 2858.625 ;
    END
  END mprj_io_vtrip_sel[29]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 809.375 3167.185 809.975 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_vtrip_sel[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2642.025 4.000 2642.625 ;
    END
  END mprj_io_vtrip_sel[30]
  PIN mprj_io_vtrip_sel[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 2426.025 4.000 2426.625 ;
    END
  END mprj_io_vtrip_sel[31]
  PIN mprj_io_vtrip_sel[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1788.025 4.000 1788.625 ;
    END
  END mprj_io_vtrip_sel[32]
  PIN mprj_io_vtrip_sel[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1572.025 4.000 1572.625 ;
    END
  END mprj_io_vtrip_sel[33]
  PIN mprj_io_vtrip_sel[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1356.025 4.000 1356.625 ;
    END
  END mprj_io_vtrip_sel[34]
  PIN mprj_io_vtrip_sel[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 1140.025 4.000 1140.625 ;
    END
  END mprj_io_vtrip_sel[35]
  PIN mprj_io_vtrip_sel[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 924.025 4.000 924.625 ;
    END
  END mprj_io_vtrip_sel[36]
  PIN mprj_io_vtrip_sel[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT -2.185 708.025 4.000 708.625 ;
    END
  END mprj_io_vtrip_sel[37]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1035.375 3167.185 1035.975 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1260.375 3167.185 1260.975 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1485.375 3167.185 1485.975 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1711.375 3167.185 1711.975 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2597.375 3167.185 2597.975 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2823.375 3167.185 2823.975 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3048.375 3167.185 3048.975 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN por_l
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 758.715 -2.000 758.995 4.000 ;
    END
  END por_l
  PIN porb_h
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met2 ;
        RECT 1329.775 -2.000 1330.055 4.000 ;
    END
  END porb_h
  PIN rstb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 1.041900 ;
    PORT
      LAYER met2 ;
        RECT 496.835 -10.525 497.115 4.000 ;
    END
  END rstb_h
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.920 10.640 15.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3147.180 10.640 3152.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 11.880 3154.920 19.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4739.560 3154.920 4749.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.920 10.640 72.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3087.180 10.640 3089.180 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 10.640 130.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 835.505 130.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 4631.350 130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 10.640 230.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 835.505 230.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.920 4631.350 230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 10.640 330.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 835.505 330.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.920 4631.350 330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 10.640 430.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 835.505 430.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.920 4631.350 430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.920 10.640 530.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.920 835.505 530.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.920 4631.350 530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 10.640 630.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 835.505 630.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.920 4631.350 630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 10.640 730.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 835.505 730.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.920 4631.350 730.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 10.640 830.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 835.505 830.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 823.920 4631.350 830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.920 10.640 930.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.920 835.505 930.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.920 4631.350 930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.920 835.505 1030.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.920 4631.350 1030.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.920 10.640 1130.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.920 835.505 1130.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1123.920 4631.350 1130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.920 10.640 1230.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.920 835.505 1230.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.920 4631.350 1230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.920 10.640 1330.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.920 835.505 1330.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.920 4631.350 1330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.920 10.640 1430.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.920 835.505 1430.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.920 4631.350 1430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.920 10.640 1530.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.920 835.505 1530.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.920 4631.350 1530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 10.640 1630.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 835.505 1630.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1623.920 4631.350 1630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.920 10.640 1730.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.920 835.505 1730.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1723.920 4631.350 1730.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 10.640 1830.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 835.505 1830.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.920 4631.350 1830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 10.640 1930.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 835.505 1930.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1923.920 4631.350 1930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 10.640 2030.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 835.505 2030.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.920 4631.350 2030.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.920 10.640 2130.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.920 835.505 2130.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.920 4631.350 2130.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.920 10.640 2230.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.920 835.505 2230.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.920 4631.350 2230.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.920 10.640 2330.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.920 835.505 2330.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2323.920 4631.350 2330.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.920 10.640 2430.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.920 835.505 2430.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.920 4631.350 2430.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.920 10.640 2530.320 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.920 835.505 2530.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.920 4631.350 2530.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.920 10.640 2630.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2623.920 4631.350 2630.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 10.640 2730.320 266.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 797.820 2730.320 903.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2723.920 939.820 2730.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 103.620 2830.320 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 793.705 2830.320 903.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 939.820 2830.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.920 4631.350 2830.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 10.640 2930.320 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 793.705 2930.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2923.920 4631.350 2930.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 10.640 3030.320 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 793.705 3030.320 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 3023.920 4631.350 3030.320 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 212.680 555.260 219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 312.680 555.260 319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 412.680 555.260 419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 512.680 555.260 519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 612.680 555.260 619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 712.680 555.260 719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 812.680 555.260 819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 912.680 3154.920 919.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1012.680 3154.920 1019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1112.680 75.920 1119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1212.680 75.920 1219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1312.680 75.920 1319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1412.680 75.920 1419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1512.680 75.920 1519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1612.680 75.920 1619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1712.680 75.920 1719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1812.680 75.920 1819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1912.680 75.920 1919.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2112.680 75.920 2119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2312.680 75.920 2319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2412.680 75.920 2419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2512.680 75.920 2519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2612.680 75.920 2619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2712.680 75.920 2719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2812.680 75.920 2819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2912.680 75.920 2919.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3012.680 75.920 3019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3112.680 75.920 3119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3212.680 75.920 3219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3312.680 75.920 3319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3412.680 75.920 3419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3512.680 75.920 3519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3612.680 75.920 3619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3712.680 75.920 3719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3812.680 75.920 3819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4012.680 75.920 4019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4112.680 75.920 4119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4212.680 75.920 4219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4312.680 75.920 4319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4512.680 75.920 4519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4612.680 75.920 4619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 212.680 3154.920 219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 312.680 3154.920 319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 412.680 3154.920 419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 512.680 3154.920 519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 612.680 3154.920 619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 712.680 3154.920 719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 812.680 3154.920 819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1112.680 3154.920 1119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1212.680 3154.920 1219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1312.680 3154.920 1319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1412.680 3154.920 1419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1512.680 3154.920 1519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1612.680 3154.920 1619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1712.680 3154.920 1719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 1812.680 3154.920 1819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2012.680 3154.920 2019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2212.680 3154.920 2219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2412.680 3154.920 2419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2512.680 3154.920 2519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2612.680 3154.920 2619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2712.680 3154.920 2719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2812.680 3154.920 2819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 2912.680 3154.920 2919.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3012.680 3154.920 3019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3112.680 3154.920 3119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3212.680 3154.920 3219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3312.680 3154.920 3319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3412.680 3154.920 3419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3512.680 3154.920 3519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3612.680 3154.920 3619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3712.680 3154.920 3719.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 3812.680 3154.920 3819.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4012.680 3154.920 4019.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4112.680 3154.920 4119.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4212.680 3154.920 4219.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4312.680 3154.920 4319.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4412.680 3154.920 4419.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4512.680 3154.920 4519.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.180 4612.680 3154.920 4619.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 953.000 3154.920 967.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2968.375 10.640 2969.975 269.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 2968.375 793.605 2969.975 1032.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2968.375 4631.250 2969.975 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.280 886.480 2782.280 960.400 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.920 10.640 27.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3135.180 10.640 3140.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 31.080 3154.920 39.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4716.360 3154.920 4726.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 852.780 3154.920 857.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.720 10.640 1280.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.720 835.505 1280.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.720 4631.350 1280.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.720 10.640 1380.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.720 835.505 1380.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.720 4631.350 1380.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 10.640 1480.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 835.505 1480.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 4631.350 1480.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.640 10.640 270.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.640 850.960 270.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.640 4631.350 270.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.640 10.640 570.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.640 850.960 570.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.640 4631.350 570.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.640 10.640 1170.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.640 850.960 1170.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.640 4631.350 1170.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.640 10.640 1470.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.640 850.960 1470.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.640 4631.350 1470.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.640 10.640 1770.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.640 850.960 1770.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.640 4631.350 1770.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.640 10.640 2070.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.640 850.960 2070.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.640 4631.350 2070.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.640 10.640 2370.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.640 850.960 2370.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.640 4631.350 2370.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.640 10.640 2770.040 266.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.640 797.820 2770.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.640 4631.350 2770.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.640 10.640 970.040 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.640 850.960 970.040 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.640 4631.350 970.040 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1209.680 120.440 1212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1309.680 120.440 1312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1409.680 120.440 1412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1509.680 120.440 1512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1609.680 120.440 1612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1709.680 120.440 1712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1809.680 120.440 1812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1909.680 120.440 1912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2009.680 120.440 2012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2109.680 120.440 2112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2209.680 115.340 2212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2309.680 120.440 2312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2409.680 120.440 2412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2509.680 120.440 2512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2609.680 120.440 2612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2709.680 120.440 2712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2809.680 120.440 2812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2909.680 120.440 2912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3009.680 120.440 3012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3109.680 120.440 3112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3209.680 120.440 3212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3309.680 120.440 3312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3409.680 120.440 3412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3509.680 120.440 3512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3609.680 120.440 3612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3709.680 115.340 3712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3809.680 120.440 3812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3909.680 120.440 3912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4009.680 120.440 4012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4109.680 120.440 4112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4209.680 120.440 4212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4309.680 120.440 4312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4409.680 120.440 4412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4509.680 120.440 4512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1209.680 3154.920 1212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1309.680 3154.920 1312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1409.680 3154.920 1412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1509.680 3154.920 1512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1609.680 3154.920 1612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1709.680 3154.920 1712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1809.680 3154.920 1812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1909.680 3154.920 1912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2009.680 3154.920 2012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2109.680 3154.920 2112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2209.680 3154.920 2212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2309.680 3154.920 2312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2409.680 3154.920 2412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2509.680 3154.920 2512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2609.680 3154.920 2612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2709.680 3154.920 2712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2809.680 3154.920 2812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2909.680 3154.920 2912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3009.680 3154.920 3012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3109.680 3154.920 3112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3209.680 3154.920 3212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3309.680 3154.920 3312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3409.680 3154.920 3412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3509.680 3154.920 3512.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3609.680 3154.920 3612.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3709.680 3154.920 3712.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3809.680 3154.920 3812.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3909.680 3154.920 3912.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4009.680 3154.920 4012.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4109.680 3154.920 4112.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4209.680 3154.920 4212.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4309.680 3154.920 4312.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4409.680 3154.920 4412.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4509.680 3154.920 4512.080 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 64.920 10.640 69.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3093.180 10.640 3098.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 98.280 3154.920 106.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4635.160 3154.920 4645.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 866.380 3154.920 871.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.720 10.640 855.520 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.720 850.960 855.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.720 4631.350 855.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.720 10.640 905.520 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.720 850.960 905.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.720 4631.350 905.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1218.480 120.440 1220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1318.480 120.440 1320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1418.480 120.440 1420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1518.480 120.440 1520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1618.480 120.440 1620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1718.480 120.440 1720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1818.480 115.340 1820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1918.480 120.440 1920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2018.480 120.440 2020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2118.480 120.440 2120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2218.480 120.440 2220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2318.480 120.440 2320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2418.480 120.440 2420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2518.480 120.440 2520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2618.480 120.440 2620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2718.480 120.440 2720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2818.480 120.440 2820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2918.480 120.440 2920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3018.480 120.440 3020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3118.480 120.440 3120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3218.480 120.440 3220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3318.480 115.340 3320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3418.480 120.440 3420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3518.480 120.440 3520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3618.480 120.440 3620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3718.480 120.440 3720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3818.480 120.440 3820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3918.480 120.440 3920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4018.480 120.440 4020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4118.480 120.440 4120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4218.480 120.440 4220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4318.480 120.440 4320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4418.480 120.440 4420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4518.480 120.440 4520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1218.480 3154.920 1220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1318.480 3154.920 1320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1418.480 3154.920 1420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1518.480 3154.920 1520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1618.480 3154.920 1620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1718.480 3154.920 1720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1818.480 3154.920 1820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1918.480 3154.920 1920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2018.480 3154.920 2020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2118.480 3154.920 2120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2218.480 3154.920 2220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2318.480 3154.920 2320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2418.480 3154.920 2420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2518.480 3154.920 2520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2618.480 3154.920 2620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2718.480 3154.920 2720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2818.480 3154.920 2820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2918.480 3154.920 2920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3018.480 3154.920 3020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3118.480 3154.920 3120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3218.480 3154.920 3220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3318.480 3154.920 3320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3418.480 3154.920 3420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3518.480 3154.920 3520.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3618.480 3154.920 3620.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3718.480 3154.920 3720.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3818.480 3154.920 3820.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3918.480 3154.920 3920.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4018.480 3154.920 4020.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4118.480 3154.920 4120.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4218.480 3154.920 4220.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4318.480 3154.920 4320.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4418.480 3154.920 4420.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4518.480 3154.920 4520.880 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 52.920 10.640 57.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3105.180 10.640 3110.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 79.080 3154.920 87.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4658.360 3154.920 4668.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 879.980 3154.920 884.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1843.720 10.640 1848.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1843.720 835.505 1848.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1843.720 4631.350 1848.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.720 10.640 1888.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.720 835.505 1888.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.720 4631.350 1888.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1231.680 115.340 1234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1331.680 120.440 1334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1431.680 120.440 1434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1531.680 120.440 1534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1631.680 120.440 1634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1731.680 120.440 1734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1831.680 120.440 1834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1931.680 120.440 1934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2031.680 120.440 2034.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2131.680 120.440 2134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2231.680 120.440 2234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2331.680 120.440 2334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2431.680 120.440 2434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2531.680 120.440 2534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2631.680 120.440 2634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2731.680 115.340 2734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2831.680 120.440 2834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2931.680 120.440 2934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3031.680 120.440 3034.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3131.680 120.440 3134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3231.680 120.440 3234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3331.680 120.440 3334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3431.680 120.440 3434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3531.680 120.440 3534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3631.680 120.440 3634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3731.680 120.440 3734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3831.680 120.440 3834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3931.680 120.440 3934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4031.680 120.440 4034.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4131.680 120.440 4134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4231.680 115.340 4234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4331.680 120.440 4334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4431.680 120.440 4434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4531.680 120.440 4534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1231.680 3154.920 1234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1331.680 3154.920 1334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1431.680 3154.920 1434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1531.680 3154.920 1534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1631.680 3154.920 1634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1731.680 3154.920 1734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1831.680 3154.920 1834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1931.680 3154.920 1934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2131.680 3154.920 2134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2331.680 3154.920 2334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2531.680 3154.920 2534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2731.680 3154.920 2734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2931.680 3154.920 2934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3131.680 3154.920 3134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3231.680 3154.920 3234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3331.680 3154.920 3334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3431.680 3154.920 3434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3531.680 3154.920 3534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3631.680 3154.920 3634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3731.680 3154.920 3734.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3831.680 3154.920 3834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3931.680 3154.920 3934.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4031.680 3154.920 4034.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4131.680 3154.920 4134.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4231.680 3154.920 4234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4331.680 3154.920 4334.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4431.680 3154.920 4434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4531.680 3154.920 4534.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 2031.680 3154.920 2034.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 2231.680 3154.920 2234.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 2431.680 3154.920 2434.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 2631.680 3154.920 2634.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 2831.680 3154.920 2834.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3031.680 3154.920 3034.080 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.920 10.640 45.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3117.180 10.640 3122.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 59.880 3154.920 67.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4681.560 3154.920 4691.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 893.580 3154.920 898.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1859.720 10.640 1864.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1859.720 835.505 1864.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1859.720 4631.350 1864.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.720 10.640 1904.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.720 835.505 1904.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.720 4631.350 1904.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1236.080 120.440 1238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1336.080 120.440 1338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1436.080 120.440 1438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1536.080 120.440 1538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1636.080 120.440 1638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1736.080 120.440 1738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1836.080 120.440 1838.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1936.080 120.440 1938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2036.080 120.440 2038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2136.080 120.440 2138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2236.080 120.440 2238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2336.080 120.440 2338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2436.080 120.440 2438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2536.080 115.340 2538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2636.080 120.440 2638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2736.080 120.440 2738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2836.080 120.440 2838.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2936.080 120.440 2938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3036.080 120.440 3038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3136.080 120.440 3138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3236.080 120.440 3238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3336.080 120.440 3338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3436.080 120.440 3438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3536.080 120.440 3538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3636.080 120.440 3638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3736.080 120.440 3738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3836.080 120.440 3838.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3936.080 120.440 3938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4036.080 115.340 4038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4136.080 120.440 4138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4236.080 120.440 4238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4336.080 120.440 4338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4436.080 120.440 4438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4536.080 120.440 4538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1336.080 3154.920 1338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1536.080 3154.920 1538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1736.080 3154.920 1738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1936.080 3154.920 1938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2036.080 3154.920 2038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2136.080 3154.920 2138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2236.080 3154.920 2238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2336.080 3154.920 2338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2436.080 3154.920 2438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2536.080 3154.920 2538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2636.080 3154.920 2638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2736.080 3154.920 2738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2836.080 3154.920 2838.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2936.080 3154.920 2938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3036.080 3154.920 3038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3136.080 3154.920 3138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3236.080 3154.920 3238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3336.080 3154.920 3338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3436.080 3154.920 3438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3536.080 3154.920 3538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3636.080 3154.920 3638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3736.080 3154.920 3738.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3836.080 3154.920 3838.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3936.080 3154.920 3938.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4036.080 3154.920 4038.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4136.080 3154.920 4138.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4236.080 3154.920 4238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4336.080 3154.920 4338.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4436.080 3154.920 4438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4536.080 3154.920 4538.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 1236.080 3154.920 1238.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 1436.080 3154.920 1438.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 1636.080 3154.920 1638.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 1836.080 3154.920 1838.480 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 121.600 118.380 2681.365 124.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 2614.460 152.380 2681.365 158.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 2648.720 10.640 2653.520 1032.330 ;
    END
  END vddio
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.920 10.640 51.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3111.180 10.640 3116.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 69.480 3154.920 77.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4669.960 3154.920 4679.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 886.780 3154.920 891.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.720 10.640 1856.520 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.720 850.960 1856.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.720 4631.350 1856.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.720 10.640 1896.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.720 835.505 1896.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1891.720 4631.350 1896.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1227.280 120.440 1229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1327.280 120.440 1329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1427.280 115.340 1429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1527.280 120.440 1529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1627.280 120.440 1629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1727.280 120.440 1729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1827.280 120.440 1829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1927.280 120.440 1929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2027.280 120.440 2029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2127.280 120.440 2129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2227.280 120.440 2229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2327.280 120.440 2329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2427.280 120.440 2429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2527.280 120.440 2529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2627.280 120.440 2629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2727.280 120.440 2729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2827.280 120.440 2829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2927.280 115.340 2929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3027.280 120.440 3029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3127.280 120.440 3129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3227.280 120.440 3229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3327.280 120.440 3329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3427.280 120.440 3429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3527.280 120.440 3529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3627.280 120.440 3629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3727.280 120.440 3729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3827.280 120.440 3829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3927.280 120.440 3929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4027.280 120.440 4029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4127.280 120.440 4129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4227.280 120.440 4229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4327.280 120.440 4329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4427.280 115.340 4429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4527.280 120.440 4529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1227.280 3154.920 1229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1327.280 3154.920 1329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1427.280 3154.920 1429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1527.280 3154.920 1529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1627.280 3154.920 1629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1727.280 3154.920 1729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1827.280 3154.920 1829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1927.280 3154.920 1929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2027.280 3154.920 2029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2127.280 3154.920 2129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2227.280 3154.920 2229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2327.280 3154.920 2329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2427.280 3154.920 2429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2527.280 3154.920 2529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2627.280 3154.920 2629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2727.280 3154.920 2729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2827.280 3154.920 2829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2927.280 3154.920 2929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3127.280 3154.920 3129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3327.280 3154.920 3329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3527.280 3154.920 3529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3727.280 3154.920 3729.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3927.280 3154.920 3929.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4127.280 3154.920 4129.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4327.280 3154.920 4329.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4427.280 3154.920 4429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4527.280 3154.920 4529.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3027.280 3154.920 3029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3227.280 3154.920 3229.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3427.280 3154.920 3429.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3627.280 3154.920 3629.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 3827.280 3154.920 3829.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 4027.280 3154.920 4029.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 4227.280 3154.920 4229.680 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.920 10.640 39.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3123.180 10.640 3128.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 50.280 3154.920 58.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4693.160 3154.920 4703.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 900.380 3154.920 905.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.720 10.640 1872.520 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.720 850.960 1872.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1867.720 4631.350 1872.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.720 10.640 1912.520 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.720 850.960 1912.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1907.720 4631.350 1912.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1240.480 120.440 1242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1340.480 120.440 1342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1440.480 120.440 1442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1540.480 120.440 1542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1640.480 120.440 1642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1740.480 120.440 1742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1840.480 120.440 1842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1940.480 120.440 1942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2040.480 120.440 2042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2140.480 120.440 2142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2240.480 120.440 2242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2340.480 115.340 2342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2440.480 120.440 2442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2540.480 120.440 2542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2640.480 120.440 2642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2740.480 120.440 2742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2840.480 120.440 2842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2940.480 120.440 2942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3040.480 120.440 3042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3140.480 120.440 3142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3240.480 120.440 3242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3340.480 120.440 3342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3440.480 120.440 3442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3540.480 120.440 3542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3640.480 120.440 3642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3740.480 120.440 3742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3840.480 115.340 3842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3940.480 120.440 3942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4040.480 120.440 4042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4140.480 120.440 4142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4240.480 120.440 4242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4340.480 120.440 4342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4440.480 120.440 4442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4540.480 120.440 4542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1240.480 3154.920 1242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1340.480 3154.920 1342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1440.480 3154.920 1442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1540.480 3154.920 1542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1640.480 3154.920 1642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1740.480 3154.920 1742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1840.480 3154.920 1842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1940.480 3154.920 1942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2040.480 3154.920 2042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2140.480 3154.920 2142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2240.480 3154.920 2242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2340.480 3154.920 2342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2440.480 3154.920 2442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2540.480 3154.920 2542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2640.480 3154.920 2642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2740.480 3154.920 2742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2840.480 3154.920 2842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2940.480 3154.920 2942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3040.480 3154.920 3042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3140.480 3154.920 3142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3240.480 3154.920 3242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3340.480 3154.920 3342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3440.480 3154.920 3442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3540.480 3154.920 3542.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3640.480 3154.920 3642.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3740.480 3154.920 3742.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3840.480 3154.920 3842.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3940.480 3154.920 3942.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4040.480 3154.920 4042.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4140.480 3154.920 4142.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4240.480 3154.920 4242.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4340.480 3154.920 4342.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4440.480 3154.920 4442.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4540.480 3154.920 4542.880 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.920 10.640 21.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3141.180 10.640 3146.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 21.480 3154.920 29.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4727.960 3154.920 4737.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.920 10.640 75.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3090.180 10.640 3092.180 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.520 10.640 137.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.520 835.505 137.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.520 4631.350 137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 10.640 237.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 835.505 237.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.520 4631.350 237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 10.640 337.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 835.505 337.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.520 4631.350 337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 10.640 437.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 835.505 437.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 431.520 4631.350 437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.520 10.640 537.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.520 835.505 537.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.520 4631.350 537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 10.640 637.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 835.505 637.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 631.520 4631.350 637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 10.640 737.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 835.505 737.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.520 4631.350 737.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 10.640 837.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 835.505 837.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.520 4631.350 837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 10.640 937.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 835.505 937.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 4631.350 937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.520 835.505 1037.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.520 4631.350 1037.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.520 10.640 1137.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.520 835.505 1137.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.520 4631.350 1137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.520 10.640 1237.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.520 835.505 1237.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.520 4631.350 1237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1331.520 10.640 1337.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1331.520 835.505 1337.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1331.520 4631.350 1337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.520 10.640 1437.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.520 835.505 1437.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.520 4631.350 1437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.520 10.640 1537.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.520 835.505 1537.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.520 4631.350 1537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 10.640 1637.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 835.505 1637.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1631.520 4631.350 1637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.520 10.640 1737.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.520 835.505 1737.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.520 4631.350 1737.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 10.640 1837.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 835.505 1837.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.520 4631.350 1837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 10.640 1937.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 835.505 1937.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.520 4631.350 1937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 10.640 2037.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 835.505 2037.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2031.520 4631.350 2037.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.520 10.640 2137.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.520 835.505 2137.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.520 4631.350 2137.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.520 10.640 2237.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.520 835.505 2237.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.520 4631.350 2237.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.520 10.640 2337.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.520 835.505 2337.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2331.520 4631.350 2337.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2431.520 10.640 2437.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2431.520 835.505 2437.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2431.520 4631.350 2437.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2531.520 10.640 2537.920 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2531.520 835.505 2537.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2531.520 4631.350 2537.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.520 10.640 2637.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.520 4631.350 2637.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 10.640 2737.920 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 793.705 2737.920 903.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.520 939.820 2737.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 103.620 2837.920 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 793.705 2837.920 903.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 939.820 2837.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.520 4631.350 2837.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 10.640 2937.920 269.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 793.705 2937.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.520 4631.350 2937.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 10.640 3037.920 266.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 797.820 3037.920 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 3031.520 4631.350 3037.920 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 221.480 555.260 227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 321.480 555.260 327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 421.480 555.260 427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 521.480 555.260 527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 621.480 555.260 627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 721.480 555.260 727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 821.480 3154.920 827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 921.480 3154.920 927.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1021.480 3154.920 1027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1121.480 75.920 1127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1221.480 75.920 1227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1321.480 75.920 1327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1421.480 75.920 1427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1521.480 75.920 1527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1621.480 75.920 1627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1721.480 75.920 1727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1821.480 75.920 1827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1921.480 75.920 1927.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2121.480 75.920 2127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2321.480 75.920 2327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2421.480 75.920 2427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2521.480 75.920 2527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2621.480 75.920 2627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2721.480 75.920 2727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2821.480 75.920 2827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2921.480 75.920 2927.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3021.480 75.920 3027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3121.480 75.920 3127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3221.480 75.920 3227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3321.480 75.920 3327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3421.480 75.920 3427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3521.480 75.920 3527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3621.480 75.920 3627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3721.480 75.920 3727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3821.480 75.920 3827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4021.480 75.920 4027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4121.480 75.920 4127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4221.480 75.920 4227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4321.480 75.920 4327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4521.480 75.920 4527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4621.480 73.910 4627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 221.480 3154.920 227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 321.480 3154.920 327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 421.480 3154.920 427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 521.480 3154.920 527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 621.480 3154.920 627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 721.480 3154.920 727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1121.480 3154.920 1127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1221.480 3154.920 1227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1321.480 3154.920 1327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1421.480 3154.920 1427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1521.480 3154.920 1527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1621.480 3154.920 1627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1721.480 3154.920 1727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 1821.480 3154.920 1827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2021.480 3154.920 2027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2221.480 3154.920 2227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2421.480 3154.920 2427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2521.480 3154.920 2527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2621.480 3154.920 2627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2721.480 3154.920 2727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2821.480 3154.920 2827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 2921.480 3154.920 2927.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3021.480 3154.920 3027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3121.480 3154.920 3127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3221.480 3154.920 3227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3321.480 3154.920 3327.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3421.480 3154.920 3427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3521.480 3154.920 3527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3621.480 3154.920 3627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3721.480 3154.920 3727.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 3821.480 3154.920 3827.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 4021.480 3154.920 4027.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 4121.480 3154.920 4127.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 4221.480 3154.920 4227.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 4421.480 3154.920 4427.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3088.180 4521.480 3154.920 4527.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 3089.190 4621.480 3154.920 4627.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 969.800 3154.920 984.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2990.755 10.640 2992.355 269.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 2990.755 793.605 2992.355 1032.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2990.755 4631.250 2992.355 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2783.720 886.480 2788.720 960.400 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.920 10.640 33.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3129.180 10.640 3134.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 40.680 3154.920 48.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4704.760 3154.920 4714.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 859.580 3154.920 864.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.720 10.640 1288.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.720 835.505 1288.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.720 4631.350 1288.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1383.720 10.640 1388.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1383.720 835.505 1388.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1383.720 4631.350 1388.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1483.720 10.640 1488.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 1483.720 835.505 1488.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1483.720 4631.350 1488.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 10.640 262.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 850.960 262.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 4631.350 262.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.040 10.640 562.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.040 850.960 562.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.040 4631.350 562.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.040 10.640 1162.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.040 850.960 1162.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.040 4631.350 1162.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1456.040 10.640 1462.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1456.040 850.960 1462.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1456.040 4631.350 1462.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.040 10.640 1762.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.040 850.960 1762.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.040 4631.350 1762.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.040 10.640 2062.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.040 850.960 2062.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.040 4631.350 2062.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.040 10.640 2362.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.040 850.960 2362.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2356.040 4631.350 2362.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2756.040 10.640 2762.440 266.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2756.040 797.820 2762.440 903.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2756.040 939.820 2762.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2756.040 4631.350 2762.440 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.040 10.640 962.440 108.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.040 850.960 962.440 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.040 4631.350 962.440 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1214.080 120.440 1216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1314.080 120.440 1316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1414.080 120.440 1416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1514.080 120.440 1516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1614.080 120.440 1616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1714.080 120.440 1716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1814.080 120.440 1816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1914.080 120.440 1916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2014.080 115.340 2016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2114.080 120.440 2116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2214.080 120.440 2216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2314.080 120.440 2316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2414.080 120.440 2416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2514.080 120.440 2516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2614.080 120.440 2616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2714.080 120.440 2716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2814.080 120.440 2816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2914.080 120.440 2916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3014.080 120.440 3016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3114.080 120.440 3116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3214.080 120.440 3216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3314.080 120.440 3316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3414.080 120.440 3416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3514.080 115.340 3516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3614.080 120.440 3616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3714.080 120.440 3716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3814.080 120.440 3816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3914.080 120.440 3916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4014.080 120.440 4016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4114.080 120.440 4116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4214.080 120.440 4216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4314.080 120.440 4316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4414.080 120.440 4416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4514.080 120.440 4516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1214.080 3154.920 1216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1314.080 3154.920 1316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1414.080 3154.920 1416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1514.080 3154.920 1516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1614.080 3154.920 1616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1714.080 3154.920 1716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1814.080 3154.920 1816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1914.080 3154.920 1916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2014.080 3154.920 2016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2114.080 3154.920 2116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2214.080 3154.920 2216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2314.080 3154.920 2316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2414.080 3154.920 2416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2514.080 3154.920 2516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2614.080 3154.920 2616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2714.080 3154.920 2716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2814.080 3154.920 2816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2914.080 3154.920 2916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3014.080 3154.920 3016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3114.080 3154.920 3116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3214.080 3154.920 3216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3314.080 3154.920 3316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3414.080 3154.920 3416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3514.080 3154.920 3516.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3614.080 3154.920 3616.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3714.080 3154.920 3716.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3814.080 3154.920 3816.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3914.080 3154.920 3916.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4014.080 3154.920 4016.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4114.080 3154.920 4116.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4214.080 3154.920 4216.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4314.080 3154.920 4316.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4414.080 3154.920 4416.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4514.080 3154.920 4516.480 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 58.920 10.640 63.920 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3099.180 10.640 3104.180 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 88.680 3154.920 96.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4646.760 3154.920 4656.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 873.180 3154.920 877.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 10.640 863.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 835.505 863.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 4631.350 863.520 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 10.640 913.520 114.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 835.505 913.520 1032.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 4631.350 913.520 4754.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1222.880 120.440 1225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1322.880 120.440 1325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1422.880 120.440 1425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1522.880 120.440 1525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1622.880 115.340 1625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1722.880 120.440 1725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1822.880 120.440 1825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 1922.880 120.440 1925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2022.880 120.440 2025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2122.880 120.440 2125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2222.880 120.440 2225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2322.880 120.440 2325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2422.880 120.440 2425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2522.880 120.440 2525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2622.880 120.440 2625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2722.880 120.440 2725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2822.880 120.440 2825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 2922.880 120.440 2925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3022.880 120.440 3025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3122.880 115.340 3125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3222.880 120.440 3225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3322.880 120.440 3325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3422.880 120.440 3425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3522.880 120.440 3525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3622.880 120.440 3625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3722.880 120.440 3725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3822.880 120.440 3825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 3922.880 120.440 3925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4022.880 120.440 4025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4122.880 120.440 4125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4222.880 120.440 4225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4322.880 120.440 4325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4422.880 120.440 4425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.880 4522.880 120.440 4525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1222.880 3154.920 1225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1322.880 3154.920 1325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1422.880 3154.920 1425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1522.880 3154.920 1525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1622.880 3154.920 1625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1722.880 3154.920 1725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1822.880 3154.920 1825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 1922.880 3154.920 1925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2022.880 3154.920 2025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2122.880 3154.920 2125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2222.880 3154.920 2225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2322.880 3154.920 2325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2422.880 3154.920 2425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2522.880 3154.920 2525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2622.880 3154.920 2625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2722.880 3154.920 2725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2822.880 3154.920 2825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 2922.880 3154.920 2925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3022.880 3154.920 3025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3122.880 3154.920 3125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3222.880 3154.920 3225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3322.880 3154.920 3325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3422.880 3154.920 3425.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3522.880 3154.920 3525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3622.880 3154.920 3625.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3722.880 3154.920 3725.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3822.880 3154.920 3825.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 3922.880 3154.920 3925.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4022.880 3154.920 4025.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4122.880 3154.920 4125.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4322.880 3154.920 4325.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3043.040 4522.880 3154.920 4525.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 4222.880 3154.920 4225.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3048.140 4422.880 3154.920 4425.280 ;
    END
  END vssd2
  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 121.600 126.380 2681.365 132.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 2602.900 160.380 2720.455 166.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.520 10.640 2660.320 1032.330 ;
    END
  END vssio
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 3154.680 4754.645 ;
      LAYER met1 ;
        RECT 6.510 10.640 3161.970 4755.540 ;
      LAYER met2 ;
        RECT 6.530 4762.720 173.465 4763.810 ;
        RECT 174.305 4762.720 176.685 4763.810 ;
        RECT 177.525 4762.720 179.905 4763.810 ;
        RECT 180.745 4762.720 189.105 4763.810 ;
        RECT 189.945 4762.720 191.865 4763.810 ;
        RECT 192.705 4762.720 195.085 4763.810 ;
        RECT 195.925 4762.720 198.305 4763.810 ;
        RECT 199.145 4762.720 210.725 4763.810 ;
        RECT 211.565 4762.720 213.485 4763.810 ;
        RECT 214.325 4762.720 216.705 4763.810 ;
        RECT 217.545 4762.720 219.925 4763.810 ;
        RECT 220.765 4762.720 225.905 4763.810 ;
        RECT 226.745 4762.720 231.885 4763.810 ;
        RECT 232.725 4762.720 235.105 4763.810 ;
        RECT 235.945 4762.720 238.325 4763.810 ;
        RECT 239.165 4762.720 244.305 4763.810 ;
        RECT 245.145 4762.720 430.465 4763.810 ;
        RECT 431.305 4762.720 433.685 4763.810 ;
        RECT 434.525 4762.720 436.905 4763.810 ;
        RECT 437.745 4762.720 446.105 4763.810 ;
        RECT 446.945 4762.720 448.865 4763.810 ;
        RECT 449.705 4762.720 452.085 4763.810 ;
        RECT 452.925 4762.720 455.305 4763.810 ;
        RECT 456.145 4762.720 467.725 4763.810 ;
        RECT 468.565 4762.720 470.485 4763.810 ;
        RECT 471.325 4762.720 473.705 4763.810 ;
        RECT 474.545 4762.720 476.925 4763.810 ;
        RECT 477.765 4762.720 482.905 4763.810 ;
        RECT 483.745 4762.720 488.885 4763.810 ;
        RECT 489.725 4762.720 492.105 4763.810 ;
        RECT 492.945 4762.720 495.325 4763.810 ;
        RECT 496.165 4762.720 501.305 4763.810 ;
        RECT 502.145 4762.720 687.465 4763.810 ;
        RECT 688.305 4762.720 690.685 4763.810 ;
        RECT 691.525 4762.720 693.905 4763.810 ;
        RECT 694.745 4762.720 703.105 4763.810 ;
        RECT 703.945 4762.720 705.865 4763.810 ;
        RECT 706.705 4762.720 709.085 4763.810 ;
        RECT 709.925 4762.720 712.305 4763.810 ;
        RECT 713.145 4762.720 724.725 4763.810 ;
        RECT 725.565 4762.720 727.485 4763.810 ;
        RECT 728.325 4762.720 730.705 4763.810 ;
        RECT 731.545 4762.720 733.925 4763.810 ;
        RECT 734.765 4762.720 739.905 4763.810 ;
        RECT 740.745 4762.720 745.885 4763.810 ;
        RECT 746.725 4762.720 749.105 4763.810 ;
        RECT 749.945 4762.720 752.325 4763.810 ;
        RECT 753.165 4762.720 758.305 4763.810 ;
        RECT 759.145 4762.720 944.465 4763.810 ;
        RECT 945.305 4762.720 947.685 4763.810 ;
        RECT 948.525 4762.720 950.905 4763.810 ;
        RECT 951.745 4762.720 960.105 4763.810 ;
        RECT 960.945 4762.720 962.865 4763.810 ;
        RECT 963.705 4762.720 966.085 4763.810 ;
        RECT 966.925 4762.720 969.305 4763.810 ;
        RECT 970.145 4762.720 981.725 4763.810 ;
        RECT 982.565 4762.720 984.485 4763.810 ;
        RECT 985.325 4762.720 987.705 4763.810 ;
        RECT 988.545 4762.720 990.925 4763.810 ;
        RECT 991.765 4762.720 996.905 4763.810 ;
        RECT 997.745 4762.720 1002.885 4763.810 ;
        RECT 1003.725 4762.720 1006.105 4763.810 ;
        RECT 1006.945 4762.720 1009.325 4763.810 ;
        RECT 1010.165 4762.720 1015.305 4763.810 ;
        RECT 1016.145 4762.720 1202.465 4763.810 ;
        RECT 1203.305 4762.720 1205.685 4763.810 ;
        RECT 1206.525 4762.720 1208.905 4763.810 ;
        RECT 1209.745 4762.720 1218.105 4763.810 ;
        RECT 1218.945 4762.720 1220.865 4763.810 ;
        RECT 1221.705 4762.720 1224.085 4763.810 ;
        RECT 1224.925 4762.720 1227.305 4763.810 ;
        RECT 1228.145 4762.720 1239.725 4763.810 ;
        RECT 1240.565 4762.720 1242.485 4763.810 ;
        RECT 1243.325 4762.720 1245.705 4763.810 ;
        RECT 1246.545 4762.720 1248.925 4763.810 ;
        RECT 1249.765 4762.720 1254.905 4763.810 ;
        RECT 1255.745 4762.720 1260.885 4763.810 ;
        RECT 1261.725 4762.720 1264.105 4763.810 ;
        RECT 1264.945 4762.720 1267.325 4763.810 ;
        RECT 1268.165 4762.720 1273.305 4763.810 ;
        RECT 1274.145 4762.720 1711.465 4763.810 ;
        RECT 1712.305 4762.720 1714.685 4763.810 ;
        RECT 1715.525 4762.720 1717.905 4763.810 ;
        RECT 1718.745 4762.720 1727.105 4763.810 ;
        RECT 1727.945 4762.720 1729.865 4763.810 ;
        RECT 1730.705 4762.720 1733.085 4763.810 ;
        RECT 1733.925 4762.720 1736.305 4763.810 ;
        RECT 1737.145 4762.720 1748.725 4763.810 ;
        RECT 1749.565 4762.720 1751.485 4763.810 ;
        RECT 1752.325 4762.720 1754.705 4763.810 ;
        RECT 1755.545 4762.720 1757.925 4763.810 ;
        RECT 1758.765 4762.720 1763.905 4763.810 ;
        RECT 1764.745 4762.720 1769.885 4763.810 ;
        RECT 1770.725 4762.720 1773.105 4763.810 ;
        RECT 1773.945 4762.720 1776.325 4763.810 ;
        RECT 1777.165 4762.720 1782.305 4763.810 ;
        RECT 1783.145 4762.720 2156.465 4763.810 ;
        RECT 2157.305 4762.720 2159.685 4763.810 ;
        RECT 2160.525 4762.720 2162.905 4763.810 ;
        RECT 2163.745 4762.720 2172.105 4763.810 ;
        RECT 2172.945 4762.720 2174.865 4763.810 ;
        RECT 2175.705 4762.720 2178.085 4763.810 ;
        RECT 2178.925 4762.720 2181.305 4763.810 ;
        RECT 2182.145 4762.720 2193.725 4763.810 ;
        RECT 2194.565 4762.720 2196.485 4763.810 ;
        RECT 2197.325 4762.720 2199.705 4763.810 ;
        RECT 2200.545 4762.720 2202.925 4763.810 ;
        RECT 2203.765 4762.720 2208.905 4763.810 ;
        RECT 2209.745 4762.720 2214.885 4763.810 ;
        RECT 2215.725 4762.720 2218.105 4763.810 ;
        RECT 2218.945 4762.720 2221.325 4763.810 ;
        RECT 2222.165 4762.720 2227.305 4763.810 ;
        RECT 2228.145 4762.720 2413.465 4763.810 ;
        RECT 2414.305 4762.720 2416.685 4763.810 ;
        RECT 2417.525 4762.720 2419.905 4763.810 ;
        RECT 2420.745 4762.720 2429.105 4763.810 ;
        RECT 2429.945 4762.720 2431.865 4763.810 ;
        RECT 2432.705 4762.720 2435.085 4763.810 ;
        RECT 2435.925 4762.720 2438.305 4763.810 ;
        RECT 2439.145 4762.720 2450.725 4763.810 ;
        RECT 2451.565 4762.720 2453.485 4763.810 ;
        RECT 2454.325 4762.720 2456.705 4763.810 ;
        RECT 2457.545 4762.720 2459.925 4763.810 ;
        RECT 2460.765 4762.720 2465.905 4763.810 ;
        RECT 2466.745 4762.720 2471.885 4763.810 ;
        RECT 2472.725 4762.720 2475.105 4763.810 ;
        RECT 2475.945 4762.720 2478.325 4763.810 ;
        RECT 2479.165 4762.720 2484.305 4763.810 ;
        RECT 2485.145 4762.720 2922.465 4763.810 ;
        RECT 2923.305 4762.720 2925.685 4763.810 ;
        RECT 2926.525 4762.720 2928.905 4763.810 ;
        RECT 2929.745 4762.720 2938.105 4763.810 ;
        RECT 2938.945 4762.720 2940.865 4763.810 ;
        RECT 2941.705 4762.720 2944.085 4763.810 ;
        RECT 2944.925 4762.720 2947.305 4763.810 ;
        RECT 2948.145 4762.720 2959.725 4763.810 ;
        RECT 2960.565 4762.720 2962.485 4763.810 ;
        RECT 2963.325 4762.720 2965.705 4763.810 ;
        RECT 2966.545 4762.720 2968.925 4763.810 ;
        RECT 2969.765 4762.720 2974.905 4763.810 ;
        RECT 2975.745 4762.720 2980.885 4763.810 ;
        RECT 2981.725 4762.720 2984.105 4763.810 ;
        RECT 2984.945 4762.720 2987.325 4763.810 ;
        RECT 2988.165 4762.720 2993.305 4763.810 ;
        RECT 2994.145 4762.720 3161.950 4763.810 ;
        RECT 6.530 4.280 3161.950 4762.720 ;
        RECT 6.530 3.670 496.555 4.280 ;
        RECT 497.395 3.670 724.855 4.280 ;
        RECT 725.695 3.670 758.435 4.280 ;
        RECT 759.275 3.670 1323.055 4.280 ;
        RECT 1323.895 3.670 1329.495 4.280 ;
        RECT 1330.335 3.670 1338.695 4.280 ;
        RECT 1339.535 3.670 1597.055 4.280 ;
        RECT 1597.895 3.670 1612.695 4.280 ;
        RECT 1613.535 3.670 1815.855 4.280 ;
        RECT 1816.695 3.670 1849.435 4.280 ;
        RECT 1850.275 3.670 1871.055 4.280 ;
        RECT 1871.895 3.670 1886.695 4.280 ;
        RECT 1887.535 3.670 2089.855 4.280 ;
        RECT 2090.695 3.670 2123.435 4.280 ;
        RECT 2124.275 3.670 2145.055 4.280 ;
        RECT 2145.895 3.670 2160.695 4.280 ;
        RECT 2161.535 3.670 2363.855 4.280 ;
        RECT 2364.695 3.670 2391.455 4.280 ;
        RECT 2392.295 3.670 2397.435 4.280 ;
        RECT 2398.275 3.670 2413.075 4.280 ;
        RECT 2413.915 3.670 2419.055 4.280 ;
        RECT 2419.895 3.670 2434.695 4.280 ;
        RECT 2435.535 3.670 3161.950 4.280 ;
      LAYER met3 ;
        RECT 2666.935 4767.000 2690.965 4777.980 ;
        RECT 2716.840 4767.000 2740.870 4777.980 ;
        RECT 0.000 4636.425 3165.000 4767.000 ;
        RECT 4.400 4635.025 3165.000 4636.425 ;
        RECT 0.000 4630.445 3165.000 4635.025 ;
        RECT 4.400 4629.045 3165.000 4630.445 ;
        RECT 0.000 4627.225 3165.000 4629.045 ;
        RECT 4.400 4625.825 3165.000 4627.225 ;
        RECT 0.000 4624.005 3165.000 4625.825 ;
        RECT 4.400 4623.815 3165.000 4624.005 ;
        RECT 4.400 4622.605 3160.600 4623.815 ;
        RECT 0.000 4622.415 3160.600 4622.605 ;
        RECT 0.000 4620.595 3165.000 4622.415 ;
        RECT 0.000 4619.195 3160.600 4620.595 ;
        RECT 0.000 4618.025 3165.000 4619.195 ;
        RECT 4.400 4617.375 3165.000 4618.025 ;
        RECT 4.400 4616.625 3160.600 4617.375 ;
        RECT 0.000 4615.975 3160.600 4616.625 ;
        RECT 0.000 4612.045 3165.000 4615.975 ;
        RECT 4.400 4610.645 3165.000 4612.045 ;
        RECT 0.000 4608.825 3165.000 4610.645 ;
        RECT 4.400 4608.175 3165.000 4608.825 ;
        RECT 4.400 4607.425 3160.600 4608.175 ;
        RECT 0.000 4606.775 3160.600 4607.425 ;
        RECT 0.000 4605.605 3165.000 4606.775 ;
        RECT 4.400 4605.415 3165.000 4605.605 ;
        RECT 4.400 4604.205 3160.600 4605.415 ;
        RECT 0.000 4604.015 3160.600 4604.205 ;
        RECT 0.000 4602.845 3165.000 4604.015 ;
        RECT 4.400 4602.195 3165.000 4602.845 ;
        RECT 4.400 4601.445 3160.600 4602.195 ;
        RECT 0.000 4600.795 3160.600 4601.445 ;
        RECT 0.000 4598.975 3165.000 4600.795 ;
        RECT 0.000 4597.575 3160.600 4598.975 ;
        RECT 0.000 4590.425 3165.000 4597.575 ;
        RECT 4.400 4589.025 3165.000 4590.425 ;
        RECT 0.000 4587.205 3165.000 4589.025 ;
        RECT 4.400 4586.555 3165.000 4587.205 ;
        RECT 4.400 4585.805 3160.600 4586.555 ;
        RECT 0.000 4585.155 3160.600 4585.805 ;
        RECT 0.000 4583.985 3165.000 4585.155 ;
        RECT 4.400 4583.795 3165.000 4583.985 ;
        RECT 4.400 4582.585 3160.600 4583.795 ;
        RECT 0.000 4582.395 3160.600 4582.585 ;
        RECT 0.000 4581.225 3165.000 4582.395 ;
        RECT 4.400 4580.575 3165.000 4581.225 ;
        RECT 4.400 4579.825 3160.600 4580.575 ;
        RECT 0.000 4579.175 3160.600 4579.825 ;
        RECT 0.000 4577.355 3165.000 4579.175 ;
        RECT 0.000 4575.955 3160.600 4577.355 ;
        RECT 0.000 4572.025 3165.000 4575.955 ;
        RECT 4.400 4571.375 3165.000 4572.025 ;
        RECT 4.400 4570.625 3160.600 4571.375 ;
        RECT 0.000 4569.975 3160.600 4570.625 ;
        RECT 0.000 4568.805 3165.000 4569.975 ;
        RECT 4.400 4567.405 3165.000 4568.805 ;
        RECT 0.000 4565.585 3165.000 4567.405 ;
        RECT 4.400 4565.395 3165.000 4565.585 ;
        RECT 4.400 4564.185 3160.600 4565.395 ;
        RECT 0.000 4563.995 3160.600 4564.185 ;
        RECT 0.000 4562.175 3165.000 4563.995 ;
        RECT 0.000 4560.775 3160.600 4562.175 ;
        RECT 0.000 4558.955 3165.000 4560.775 ;
        RECT 0.000 4557.555 3160.600 4558.955 ;
        RECT 0.000 4552.975 3165.000 4557.555 ;
        RECT 0.000 4551.575 3160.600 4552.975 ;
        RECT 0.000 4543.280 3165.000 4551.575 ;
        RECT 0.000 4540.080 9.480 4543.280 ;
        RECT 120.840 4540.080 3042.640 4543.280 ;
        RECT 3155.320 4540.080 3165.000 4543.280 ;
        RECT 0.000 4538.880 3165.000 4540.080 ;
        RECT 0.000 4535.680 9.480 4538.880 ;
        RECT 120.840 4535.680 3042.640 4538.880 ;
        RECT 3155.320 4535.680 3165.000 4538.880 ;
        RECT 0.000 4534.480 3165.000 4535.680 ;
        RECT 0.000 4531.280 9.480 4534.480 ;
        RECT 120.840 4531.280 3042.640 4534.480 ;
        RECT 3155.320 4531.280 3165.000 4534.480 ;
        RECT 0.000 4530.080 3165.000 4531.280 ;
        RECT 0.000 4526.880 9.480 4530.080 ;
        RECT 120.840 4526.880 3042.640 4530.080 ;
        RECT 3155.320 4526.880 3165.000 4530.080 ;
        RECT 0.000 4525.680 3165.000 4526.880 ;
        RECT 0.000 4522.480 9.480 4525.680 ;
        RECT 120.840 4522.480 3042.640 4525.680 ;
        RECT 3155.320 4522.480 3165.000 4525.680 ;
        RECT 0.000 4521.280 3165.000 4522.480 ;
        RECT 0.000 4518.080 9.480 4521.280 ;
        RECT 120.840 4518.080 3042.640 4521.280 ;
        RECT 3155.320 4518.080 3165.000 4521.280 ;
        RECT 0.000 4516.880 3165.000 4518.080 ;
        RECT 0.000 4513.680 9.480 4516.880 ;
        RECT 120.840 4513.680 3042.640 4516.880 ;
        RECT 3155.320 4513.680 3165.000 4516.880 ;
        RECT 0.000 4512.480 3165.000 4513.680 ;
        RECT 0.000 4509.280 9.480 4512.480 ;
        RECT 120.840 4509.280 3042.640 4512.480 ;
        RECT 3155.320 4509.280 3165.000 4512.480 ;
        RECT 0.000 4443.280 3165.000 4509.280 ;
        RECT 0.000 4440.080 9.480 4443.280 ;
        RECT 120.840 4440.080 3042.640 4443.280 ;
        RECT 3155.320 4440.080 3165.000 4443.280 ;
        RECT 0.000 4438.880 3165.000 4440.080 ;
        RECT 0.000 4435.680 9.480 4438.880 ;
        RECT 120.840 4435.680 3042.640 4438.880 ;
        RECT 3155.320 4435.680 3165.000 4438.880 ;
        RECT 0.000 4434.480 3165.000 4435.680 ;
        RECT 0.000 4431.280 9.480 4434.480 ;
        RECT 120.840 4431.280 3042.640 4434.480 ;
        RECT 3155.320 4431.280 3165.000 4434.480 ;
        RECT 0.000 4430.080 3165.000 4431.280 ;
        RECT 0.000 4426.880 9.480 4430.080 ;
        RECT 115.740 4426.880 3042.640 4430.080 ;
        RECT 3155.320 4426.880 3165.000 4430.080 ;
        RECT 0.000 4425.680 3165.000 4426.880 ;
        RECT 0.000 4424.200 9.480 4425.680 ;
        RECT -16.080 4422.480 9.480 4424.200 ;
        RECT 120.840 4422.480 3047.740 4425.680 ;
        RECT 3155.320 4422.480 3165.000 4425.680 ;
        RECT -16.080 4421.280 3165.000 4422.480 ;
        RECT -16.080 4418.080 9.480 4421.280 ;
        RECT 120.840 4418.080 3042.640 4421.280 ;
        RECT 3155.320 4418.080 3165.000 4421.280 ;
        RECT -16.080 4416.880 3165.000 4418.080 ;
        RECT -16.080 4413.680 9.480 4416.880 ;
        RECT 120.840 4413.680 3042.640 4416.880 ;
        RECT 3155.320 4413.680 3165.000 4416.880 ;
        RECT -16.080 4412.480 3165.000 4413.680 ;
        RECT -16.080 4409.280 9.480 4412.480 ;
        RECT 120.840 4409.280 3042.640 4412.480 ;
        RECT 3155.320 4409.280 3165.000 4412.480 ;
        RECT -16.080 4402.000 3165.000 4409.280 ;
        RECT -16.080 4400.255 3178.020 4402.000 ;
        RECT 0.000 4398.650 3178.020 4400.255 ;
        RECT -11.000 4378.055 3178.020 4398.650 ;
        RECT -11.000 4376.450 3165.000 4378.055 ;
        RECT -11.000 4375.600 3176.020 4376.450 ;
        RECT 0.000 4374.000 3176.020 4375.600 ;
        RECT -16.080 4353.345 3176.020 4374.000 ;
        RECT -16.080 4351.745 3165.000 4353.345 ;
        RECT -16.080 4350.055 3178.020 4351.745 ;
        RECT 0.000 4343.280 3178.020 4350.055 ;
        RECT 0.000 4340.080 9.480 4343.280 ;
        RECT 120.840 4340.080 3042.640 4343.280 ;
        RECT 3155.320 4340.080 3178.020 4343.280 ;
        RECT 0.000 4338.880 3178.020 4340.080 ;
        RECT 0.000 4335.680 9.480 4338.880 ;
        RECT 120.840 4335.680 3042.640 4338.880 ;
        RECT 3155.320 4335.680 3178.020 4338.880 ;
        RECT 0.000 4334.480 3178.020 4335.680 ;
        RECT 0.000 4331.280 9.480 4334.480 ;
        RECT 120.840 4331.280 3042.640 4334.480 ;
        RECT 3155.320 4331.280 3178.020 4334.480 ;
        RECT 0.000 4330.080 3178.020 4331.280 ;
        RECT 0.000 4326.880 9.480 4330.080 ;
        RECT 120.840 4326.880 3042.640 4330.080 ;
        RECT 3155.320 4327.800 3178.020 4330.080 ;
        RECT 3155.320 4326.880 3165.000 4327.800 ;
        RECT 0.000 4325.680 3165.000 4326.880 ;
        RECT 0.000 4322.480 9.480 4325.680 ;
        RECT 120.840 4322.480 3042.640 4325.680 ;
        RECT 3155.320 4322.480 3165.000 4325.680 ;
        RECT 0.000 4321.280 3165.000 4322.480 ;
        RECT 0.000 4318.080 9.480 4321.280 ;
        RECT 120.840 4318.080 3042.640 4321.280 ;
        RECT 3155.320 4318.080 3165.000 4321.280 ;
        RECT 0.000 4316.880 3165.000 4318.080 ;
        RECT 0.000 4313.680 9.480 4316.880 ;
        RECT 120.840 4313.680 3042.640 4316.880 ;
        RECT 3155.320 4313.680 3165.000 4316.880 ;
        RECT 0.000 4312.480 3165.000 4313.680 ;
        RECT 0.000 4309.280 9.480 4312.480 ;
        RECT 120.840 4309.280 3042.640 4312.480 ;
        RECT 3155.320 4309.280 3165.000 4312.480 ;
        RECT 0.000 4243.280 3165.000 4309.280 ;
        RECT 0.000 4240.080 9.480 4243.280 ;
        RECT 120.840 4240.080 3042.640 4243.280 ;
        RECT 3155.320 4240.080 3165.000 4243.280 ;
        RECT 0.000 4238.880 3165.000 4240.080 ;
        RECT 0.000 4235.680 9.480 4238.880 ;
        RECT 120.840 4235.680 3042.640 4238.880 ;
        RECT 3155.320 4235.680 3165.000 4238.880 ;
        RECT 0.000 4234.480 3165.000 4235.680 ;
        RECT 0.000 4231.280 9.480 4234.480 ;
        RECT 115.740 4231.280 3042.640 4234.480 ;
        RECT 3155.320 4231.280 3165.000 4234.480 ;
        RECT 0.000 4230.080 3165.000 4231.280 ;
        RECT 0.000 4226.880 9.480 4230.080 ;
        RECT 120.840 4226.880 3047.740 4230.080 ;
        RECT 3155.320 4226.880 3165.000 4230.080 ;
        RECT 0.000 4225.680 3165.000 4226.880 ;
        RECT 0.000 4222.480 9.480 4225.680 ;
        RECT 120.840 4222.480 3047.740 4225.680 ;
        RECT 3155.320 4222.480 3165.000 4225.680 ;
        RECT 0.000 4221.280 3165.000 4222.480 ;
        RECT 0.000 4218.080 9.480 4221.280 ;
        RECT 120.840 4218.080 3042.640 4221.280 ;
        RECT 3155.320 4218.080 3165.000 4221.280 ;
        RECT 0.000 4216.880 3165.000 4218.080 ;
        RECT 0.000 4213.680 9.480 4216.880 ;
        RECT 120.840 4213.680 3042.640 4216.880 ;
        RECT 3155.320 4213.680 3165.000 4216.880 ;
        RECT 0.000 4212.480 3165.000 4213.680 ;
        RECT 0.000 4209.280 9.480 4212.480 ;
        RECT 120.840 4209.280 3042.640 4212.480 ;
        RECT 3155.320 4209.280 3165.000 4212.480 ;
        RECT 0.000 4177.815 3165.000 4209.280 ;
        RECT 0.000 4176.415 3160.600 4177.815 ;
        RECT 0.000 4174.595 3165.000 4176.415 ;
        RECT 0.000 4173.195 3160.600 4174.595 ;
        RECT 0.000 4171.375 3165.000 4173.195 ;
        RECT 0.000 4169.975 3160.600 4171.375 ;
        RECT 0.000 4162.175 3165.000 4169.975 ;
        RECT 0.000 4160.775 3160.600 4162.175 ;
        RECT 0.000 4159.415 3165.000 4160.775 ;
        RECT 0.000 4158.015 3160.600 4159.415 ;
        RECT 0.000 4156.195 3165.000 4158.015 ;
        RECT 0.000 4154.795 3160.600 4156.195 ;
        RECT 0.000 4152.975 3165.000 4154.795 ;
        RECT 0.000 4151.575 3160.600 4152.975 ;
        RECT 0.000 4143.280 3165.000 4151.575 ;
        RECT 0.000 4140.080 9.480 4143.280 ;
        RECT 120.840 4140.080 3042.640 4143.280 ;
        RECT 3155.320 4140.555 3165.000 4143.280 ;
        RECT 3155.320 4140.080 3160.600 4140.555 ;
        RECT 0.000 4139.155 3160.600 4140.080 ;
        RECT 0.000 4138.880 3165.000 4139.155 ;
        RECT 0.000 4135.680 9.480 4138.880 ;
        RECT 120.840 4135.680 3042.640 4138.880 ;
        RECT 3155.320 4137.795 3165.000 4138.880 ;
        RECT 3155.320 4136.395 3160.600 4137.795 ;
        RECT 3155.320 4135.680 3165.000 4136.395 ;
        RECT 0.000 4134.575 3165.000 4135.680 ;
        RECT 0.000 4134.480 3160.600 4134.575 ;
        RECT 0.000 4131.280 9.480 4134.480 ;
        RECT 120.840 4131.280 3042.640 4134.480 ;
        RECT 3155.320 4133.175 3160.600 4134.480 ;
        RECT 3155.320 4131.355 3165.000 4133.175 ;
        RECT 3155.320 4131.280 3160.600 4131.355 ;
        RECT 0.000 4130.080 3160.600 4131.280 ;
        RECT 0.000 4126.880 9.480 4130.080 ;
        RECT 120.840 4126.880 3042.640 4130.080 ;
        RECT 3155.320 4129.955 3160.600 4130.080 ;
        RECT 3155.320 4126.880 3165.000 4129.955 ;
        RECT 0.000 4125.680 3165.000 4126.880 ;
        RECT 0.000 4122.480 9.480 4125.680 ;
        RECT 120.840 4122.480 3042.640 4125.680 ;
        RECT 3155.320 4125.375 3165.000 4125.680 ;
        RECT 3155.320 4123.975 3160.600 4125.375 ;
        RECT 3155.320 4122.480 3165.000 4123.975 ;
        RECT 0.000 4121.280 3165.000 4122.480 ;
        RECT 0.000 4118.080 9.480 4121.280 ;
        RECT 120.840 4118.080 3042.640 4121.280 ;
        RECT 3155.320 4119.395 3165.000 4121.280 ;
        RECT 3155.320 4118.080 3160.600 4119.395 ;
        RECT 0.000 4117.995 3160.600 4118.080 ;
        RECT 0.000 4116.880 3165.000 4117.995 ;
        RECT 0.000 4113.680 9.480 4116.880 ;
        RECT 120.840 4113.680 3042.640 4116.880 ;
        RECT 3155.320 4116.175 3165.000 4116.880 ;
        RECT 3155.320 4114.775 3160.600 4116.175 ;
        RECT 3155.320 4113.680 3165.000 4114.775 ;
        RECT 0.000 4112.955 3165.000 4113.680 ;
        RECT 0.000 4112.480 3160.600 4112.955 ;
        RECT 0.000 4109.280 9.480 4112.480 ;
        RECT 120.840 4109.280 3042.640 4112.480 ;
        RECT 3155.320 4111.555 3160.600 4112.480 ;
        RECT 3155.320 4109.280 3165.000 4111.555 ;
        RECT 0.000 4106.975 3165.000 4109.280 ;
        RECT 0.000 4105.575 3160.600 4106.975 ;
        RECT 0.000 4043.280 3165.000 4105.575 ;
        RECT 0.000 4040.080 9.480 4043.280 ;
        RECT 120.840 4040.080 3042.640 4043.280 ;
        RECT 3155.320 4040.080 3165.000 4043.280 ;
        RECT 0.000 4038.880 3165.000 4040.080 ;
        RECT 0.000 4035.680 9.480 4038.880 ;
        RECT 115.740 4035.680 3042.640 4038.880 ;
        RECT 3155.320 4035.680 3165.000 4038.880 ;
        RECT 0.000 4034.480 3165.000 4035.680 ;
        RECT 0.000 4031.280 9.480 4034.480 ;
        RECT 120.840 4031.280 3042.640 4034.480 ;
        RECT 3155.320 4031.280 3165.000 4034.480 ;
        RECT 0.000 4030.080 3165.000 4031.280 ;
        RECT 0.000 4026.880 9.480 4030.080 ;
        RECT 120.840 4026.880 3047.740 4030.080 ;
        RECT 3155.320 4026.880 3165.000 4030.080 ;
        RECT 0.000 4025.680 3165.000 4026.880 ;
        RECT 0.000 4022.480 9.480 4025.680 ;
        RECT 120.840 4022.480 3042.640 4025.680 ;
        RECT 3155.320 4022.480 3165.000 4025.680 ;
        RECT 0.000 4021.280 3165.000 4022.480 ;
        RECT 0.000 4018.080 9.480 4021.280 ;
        RECT 120.840 4018.080 3042.640 4021.280 ;
        RECT 3155.320 4018.080 3165.000 4021.280 ;
        RECT 0.000 4016.880 3165.000 4018.080 ;
        RECT 0.000 4013.680 9.480 4016.880 ;
        RECT 120.840 4013.680 3042.640 4016.880 ;
        RECT 3155.320 4013.680 3165.000 4016.880 ;
        RECT 0.000 4012.480 3165.000 4013.680 ;
        RECT 0.000 4009.280 9.480 4012.480 ;
        RECT 120.840 4009.280 3042.640 4012.480 ;
        RECT 3155.320 4009.280 3165.000 4012.480 ;
        RECT 0.000 4001.790 3165.000 4009.280 ;
        RECT -16.080 3977.845 3165.000 4001.790 ;
        RECT 0.000 3956.005 3165.000 3977.845 ;
        RECT 0.000 3951.895 3178.020 3956.005 ;
        RECT -16.080 3943.280 3178.020 3951.895 ;
        RECT -16.080 3940.080 9.480 3943.280 ;
        RECT 120.840 3940.080 3042.640 3943.280 ;
        RECT 3155.320 3940.080 3178.020 3943.280 ;
        RECT -16.080 3938.880 3178.020 3940.080 ;
        RECT -16.080 3935.680 9.480 3938.880 ;
        RECT 120.840 3935.680 3042.640 3938.880 ;
        RECT 3155.320 3935.680 3178.020 3938.880 ;
        RECT -16.080 3934.480 3178.020 3935.680 ;
        RECT -16.080 3931.280 9.480 3934.480 ;
        RECT 120.840 3931.280 3042.640 3934.480 ;
        RECT 3155.320 3932.060 3178.020 3934.480 ;
        RECT 3155.320 3931.280 3165.000 3932.060 ;
        RECT -16.080 3930.080 3165.000 3931.280 ;
        RECT -16.080 3927.950 9.480 3930.080 ;
        RECT 0.000 3926.880 9.480 3927.950 ;
        RECT 120.840 3926.880 3042.640 3930.080 ;
        RECT 3155.320 3926.880 3165.000 3930.080 ;
        RECT 0.000 3925.680 3165.000 3926.880 ;
        RECT 0.000 3922.480 9.480 3925.680 ;
        RECT 120.840 3922.480 3042.640 3925.680 ;
        RECT 3155.320 3922.480 3165.000 3925.680 ;
        RECT 0.000 3921.280 3165.000 3922.480 ;
        RECT 0.000 3918.080 9.480 3921.280 ;
        RECT 120.840 3918.080 3042.640 3921.280 ;
        RECT 3155.320 3918.080 3165.000 3921.280 ;
        RECT 0.000 3916.880 3165.000 3918.080 ;
        RECT 0.000 3913.680 9.480 3916.880 ;
        RECT 120.840 3913.680 3042.640 3916.880 ;
        RECT 3155.320 3913.680 3165.000 3916.880 ;
        RECT 0.000 3912.480 3165.000 3913.680 ;
        RECT 0.000 3909.280 9.480 3912.480 ;
        RECT 120.840 3909.280 3042.640 3912.480 ;
        RECT 3155.320 3909.280 3165.000 3912.480 ;
        RECT 0.000 3906.090 3165.000 3909.280 ;
        RECT 0.000 3882.145 3178.020 3906.090 ;
        RECT 0.000 3843.280 3165.000 3882.145 ;
        RECT 0.000 3840.080 9.480 3843.280 ;
        RECT 115.740 3840.080 3042.640 3843.280 ;
        RECT 3155.320 3840.080 3165.000 3843.280 ;
        RECT 0.000 3838.880 3165.000 3840.080 ;
        RECT 0.000 3835.680 9.480 3838.880 ;
        RECT 120.840 3835.680 3042.640 3838.880 ;
        RECT 3155.320 3835.680 3165.000 3838.880 ;
        RECT 0.000 3834.480 3165.000 3835.680 ;
        RECT 0.000 3831.280 9.480 3834.480 ;
        RECT 120.840 3831.280 3042.640 3834.480 ;
        RECT 3155.320 3831.280 3165.000 3834.480 ;
        RECT 0.000 3830.080 3165.000 3831.280 ;
        RECT 0.000 3826.880 9.480 3830.080 ;
        RECT 120.840 3826.880 3047.740 3830.080 ;
        RECT 3155.320 3826.880 3165.000 3830.080 ;
        RECT 0.000 3825.680 3165.000 3826.880 ;
        RECT 0.000 3822.480 9.480 3825.680 ;
        RECT 120.840 3822.480 3042.640 3825.680 ;
        RECT 3155.320 3822.480 3165.000 3825.680 ;
        RECT 0.000 3821.280 3165.000 3822.480 ;
        RECT 0.000 3818.080 9.480 3821.280 ;
        RECT 120.840 3818.080 3042.640 3821.280 ;
        RECT 3155.320 3818.080 3165.000 3821.280 ;
        RECT 0.000 3816.880 3165.000 3818.080 ;
        RECT 0.000 3813.680 9.480 3816.880 ;
        RECT 120.840 3813.680 3042.640 3816.880 ;
        RECT 3155.320 3813.680 3165.000 3816.880 ;
        RECT 0.000 3812.480 3165.000 3813.680 ;
        RECT 0.000 3809.280 9.480 3812.480 ;
        RECT 120.840 3809.280 3042.640 3812.480 ;
        RECT 3155.320 3809.280 3165.000 3812.480 ;
        RECT 0.000 3787.425 3165.000 3809.280 ;
        RECT 4.400 3786.025 3165.000 3787.425 ;
        RECT 0.000 3781.445 3165.000 3786.025 ;
        RECT 4.400 3780.045 3165.000 3781.445 ;
        RECT 0.000 3778.225 3165.000 3780.045 ;
        RECT 4.400 3776.825 3165.000 3778.225 ;
        RECT 0.000 3775.005 3165.000 3776.825 ;
        RECT 4.400 3773.605 3165.000 3775.005 ;
        RECT 0.000 3769.025 3165.000 3773.605 ;
        RECT 4.400 3767.625 3165.000 3769.025 ;
        RECT 0.000 3763.045 3165.000 3767.625 ;
        RECT 4.400 3761.645 3165.000 3763.045 ;
        RECT 0.000 3759.825 3165.000 3761.645 ;
        RECT 4.400 3758.425 3165.000 3759.825 ;
        RECT 0.000 3756.605 3165.000 3758.425 ;
        RECT 4.400 3755.205 3165.000 3756.605 ;
        RECT 0.000 3753.845 3165.000 3755.205 ;
        RECT 4.400 3752.445 3165.000 3753.845 ;
        RECT 0.000 3743.280 3165.000 3752.445 ;
        RECT 0.000 3741.425 9.480 3743.280 ;
        RECT 4.400 3740.080 9.480 3741.425 ;
        RECT 120.840 3740.080 3042.640 3743.280 ;
        RECT 3155.320 3740.080 3165.000 3743.280 ;
        RECT 4.400 3740.025 3165.000 3740.080 ;
        RECT 0.000 3738.880 3165.000 3740.025 ;
        RECT 0.000 3738.205 9.480 3738.880 ;
        RECT 4.400 3736.805 9.480 3738.205 ;
        RECT 0.000 3735.680 9.480 3736.805 ;
        RECT 120.840 3735.680 3042.640 3738.880 ;
        RECT 3155.320 3735.680 3165.000 3738.880 ;
        RECT 0.000 3734.985 3165.000 3735.680 ;
        RECT 4.400 3734.480 3165.000 3734.985 ;
        RECT 4.400 3733.585 9.480 3734.480 ;
        RECT 0.000 3732.225 9.480 3733.585 ;
        RECT 4.400 3731.280 9.480 3732.225 ;
        RECT 120.840 3731.280 3042.640 3734.480 ;
        RECT 3155.320 3731.815 3165.000 3734.480 ;
        RECT 3155.320 3731.280 3160.600 3731.815 ;
        RECT 4.400 3730.825 3160.600 3731.280 ;
        RECT 0.000 3730.415 3160.600 3730.825 ;
        RECT 0.000 3730.080 3165.000 3730.415 ;
        RECT 0.000 3726.880 9.480 3730.080 ;
        RECT 120.840 3726.880 3042.640 3730.080 ;
        RECT 3155.320 3728.595 3165.000 3730.080 ;
        RECT 3155.320 3727.195 3160.600 3728.595 ;
        RECT 3155.320 3726.880 3165.000 3727.195 ;
        RECT 0.000 3725.680 3165.000 3726.880 ;
        RECT 0.000 3723.025 9.480 3725.680 ;
        RECT 4.400 3722.480 9.480 3723.025 ;
        RECT 120.840 3722.480 3042.640 3725.680 ;
        RECT 3155.320 3725.375 3165.000 3725.680 ;
        RECT 3155.320 3723.975 3160.600 3725.375 ;
        RECT 3155.320 3722.480 3165.000 3723.975 ;
        RECT 4.400 3721.625 3165.000 3722.480 ;
        RECT 0.000 3721.280 3165.000 3721.625 ;
        RECT 0.000 3719.805 9.480 3721.280 ;
        RECT 4.400 3718.405 9.480 3719.805 ;
        RECT 0.000 3718.080 9.480 3718.405 ;
        RECT 120.840 3718.080 3042.640 3721.280 ;
        RECT 3155.320 3718.080 3165.000 3721.280 ;
        RECT 0.000 3716.880 3165.000 3718.080 ;
        RECT 0.000 3716.585 9.480 3716.880 ;
        RECT 4.400 3715.185 9.480 3716.585 ;
        RECT 0.000 3713.680 9.480 3715.185 ;
        RECT 120.840 3713.680 3042.640 3716.880 ;
        RECT 3155.320 3716.175 3165.000 3716.880 ;
        RECT 3155.320 3714.775 3160.600 3716.175 ;
        RECT 3155.320 3713.680 3165.000 3714.775 ;
        RECT 0.000 3713.415 3165.000 3713.680 ;
        RECT 0.000 3712.480 3160.600 3713.415 ;
        RECT 0.000 3709.280 9.480 3712.480 ;
        RECT 115.740 3709.280 3042.640 3712.480 ;
        RECT 3155.320 3712.015 3160.600 3712.480 ;
        RECT 3155.320 3710.195 3165.000 3712.015 ;
        RECT 3155.320 3709.280 3160.600 3710.195 ;
        RECT 0.000 3708.795 3160.600 3709.280 ;
        RECT 0.000 3706.975 3165.000 3708.795 ;
        RECT 0.000 3705.575 3160.600 3706.975 ;
        RECT 0.000 3694.555 3165.000 3705.575 ;
        RECT 0.000 3693.155 3160.600 3694.555 ;
        RECT 0.000 3691.795 3165.000 3693.155 ;
        RECT 0.000 3690.395 3160.600 3691.795 ;
        RECT 0.000 3688.575 3165.000 3690.395 ;
        RECT 0.000 3687.175 3160.600 3688.575 ;
        RECT 0.000 3685.355 3165.000 3687.175 ;
        RECT 0.000 3683.955 3160.600 3685.355 ;
        RECT 0.000 3679.375 3165.000 3683.955 ;
        RECT 0.000 3677.975 3160.600 3679.375 ;
        RECT 0.000 3673.395 3165.000 3677.975 ;
        RECT 0.000 3671.995 3160.600 3673.395 ;
        RECT 0.000 3670.175 3165.000 3671.995 ;
        RECT 0.000 3668.775 3160.600 3670.175 ;
        RECT 0.000 3666.955 3165.000 3668.775 ;
        RECT 0.000 3665.555 3160.600 3666.955 ;
        RECT 0.000 3660.975 3165.000 3665.555 ;
        RECT 0.000 3659.575 3160.600 3660.975 ;
        RECT 0.000 3643.280 3165.000 3659.575 ;
        RECT 0.000 3640.080 9.480 3643.280 ;
        RECT 120.840 3640.080 3042.640 3643.280 ;
        RECT 3155.320 3640.080 3165.000 3643.280 ;
        RECT 0.000 3638.880 3165.000 3640.080 ;
        RECT 0.000 3635.680 9.480 3638.880 ;
        RECT 120.840 3635.680 3042.640 3638.880 ;
        RECT 3155.320 3635.680 3165.000 3638.880 ;
        RECT 0.000 3634.480 3165.000 3635.680 ;
        RECT 0.000 3631.280 9.480 3634.480 ;
        RECT 120.840 3631.280 3042.640 3634.480 ;
        RECT 3155.320 3631.280 3165.000 3634.480 ;
        RECT 0.000 3630.080 3165.000 3631.280 ;
        RECT 0.000 3626.880 9.480 3630.080 ;
        RECT 120.840 3626.880 3047.740 3630.080 ;
        RECT 3155.320 3626.880 3165.000 3630.080 ;
        RECT 0.000 3625.680 3165.000 3626.880 ;
        RECT 0.000 3622.480 9.480 3625.680 ;
        RECT 120.840 3622.480 3042.640 3625.680 ;
        RECT 3155.320 3622.480 3165.000 3625.680 ;
        RECT 0.000 3621.280 3165.000 3622.480 ;
        RECT 0.000 3618.080 9.480 3621.280 ;
        RECT 120.840 3618.080 3042.640 3621.280 ;
        RECT 3155.320 3618.080 3165.000 3621.280 ;
        RECT 0.000 3616.880 3165.000 3618.080 ;
        RECT 0.000 3613.680 9.480 3616.880 ;
        RECT 120.840 3613.680 3042.640 3616.880 ;
        RECT 3155.320 3613.680 3165.000 3616.880 ;
        RECT 0.000 3612.480 3165.000 3613.680 ;
        RECT 0.000 3609.280 9.480 3612.480 ;
        RECT 120.840 3609.280 3042.640 3612.480 ;
        RECT 3155.320 3609.280 3165.000 3612.480 ;
        RECT 0.000 3571.425 3165.000 3609.280 ;
        RECT 4.400 3570.025 3165.000 3571.425 ;
        RECT 0.000 3565.445 3165.000 3570.025 ;
        RECT 4.400 3564.045 3165.000 3565.445 ;
        RECT 0.000 3562.225 3165.000 3564.045 ;
        RECT 4.400 3560.825 3165.000 3562.225 ;
        RECT 0.000 3559.005 3165.000 3560.825 ;
        RECT 4.400 3557.605 3165.000 3559.005 ;
        RECT 0.000 3553.025 3165.000 3557.605 ;
        RECT 4.400 3551.625 3165.000 3553.025 ;
        RECT 0.000 3547.045 3165.000 3551.625 ;
        RECT 4.400 3545.645 3165.000 3547.045 ;
        RECT 0.000 3543.825 3165.000 3545.645 ;
        RECT 4.400 3543.280 3165.000 3543.825 ;
        RECT 4.400 3542.425 9.480 3543.280 ;
        RECT 0.000 3540.605 9.480 3542.425 ;
        RECT 4.400 3540.080 9.480 3540.605 ;
        RECT 120.840 3540.080 3042.640 3543.280 ;
        RECT 3155.320 3540.080 3165.000 3543.280 ;
        RECT 4.400 3539.205 3165.000 3540.080 ;
        RECT 0.000 3538.880 3165.000 3539.205 ;
        RECT 0.000 3537.845 9.480 3538.880 ;
        RECT 4.400 3536.445 9.480 3537.845 ;
        RECT 0.000 3535.680 9.480 3536.445 ;
        RECT 120.840 3535.680 3042.640 3538.880 ;
        RECT 3155.320 3535.680 3165.000 3538.880 ;
        RECT 0.000 3534.480 3165.000 3535.680 ;
        RECT 0.000 3531.280 9.480 3534.480 ;
        RECT 120.840 3531.280 3042.640 3534.480 ;
        RECT 3155.320 3531.280 3165.000 3534.480 ;
        RECT 0.000 3530.080 3165.000 3531.280 ;
        RECT 0.000 3526.880 9.480 3530.080 ;
        RECT 120.840 3526.880 3042.640 3530.080 ;
        RECT 3155.320 3526.880 3165.000 3530.080 ;
        RECT 0.000 3525.680 3165.000 3526.880 ;
        RECT 0.000 3525.425 9.480 3525.680 ;
        RECT 4.400 3524.025 9.480 3525.425 ;
        RECT 0.000 3522.480 9.480 3524.025 ;
        RECT 120.840 3522.480 3042.640 3525.680 ;
        RECT 3155.320 3522.480 3165.000 3525.680 ;
        RECT 0.000 3522.205 3165.000 3522.480 ;
        RECT 4.400 3521.280 3165.000 3522.205 ;
        RECT 4.400 3520.805 9.480 3521.280 ;
        RECT 0.000 3518.985 9.480 3520.805 ;
        RECT 4.400 3518.080 9.480 3518.985 ;
        RECT 120.840 3518.080 3042.640 3521.280 ;
        RECT 3155.320 3518.080 3165.000 3521.280 ;
        RECT 4.400 3517.585 3165.000 3518.080 ;
        RECT 0.000 3516.880 3165.000 3517.585 ;
        RECT 0.000 3516.225 9.480 3516.880 ;
        RECT 4.400 3514.825 9.480 3516.225 ;
        RECT 0.000 3513.680 9.480 3514.825 ;
        RECT 115.740 3513.680 3042.640 3516.880 ;
        RECT 3155.320 3513.680 3165.000 3516.880 ;
        RECT 0.000 3512.480 3165.000 3513.680 ;
        RECT 0.000 3509.280 9.480 3512.480 ;
        RECT 120.840 3509.280 3042.640 3512.480 ;
        RECT 3155.320 3509.280 3165.000 3512.480 ;
        RECT 0.000 3507.025 3165.000 3509.280 ;
        RECT 4.400 3506.815 3165.000 3507.025 ;
        RECT 4.400 3505.625 3160.600 3506.815 ;
        RECT 0.000 3505.415 3160.600 3505.625 ;
        RECT 0.000 3503.805 3165.000 3505.415 ;
        RECT 4.400 3503.595 3165.000 3503.805 ;
        RECT 4.400 3502.405 3160.600 3503.595 ;
        RECT 0.000 3502.195 3160.600 3502.405 ;
        RECT 0.000 3500.585 3165.000 3502.195 ;
        RECT 4.400 3500.375 3165.000 3500.585 ;
        RECT 4.400 3499.185 3160.600 3500.375 ;
        RECT 0.000 3498.975 3160.600 3499.185 ;
        RECT 0.000 3491.175 3165.000 3498.975 ;
        RECT 0.000 3489.775 3160.600 3491.175 ;
        RECT 0.000 3488.415 3165.000 3489.775 ;
        RECT 0.000 3487.015 3160.600 3488.415 ;
        RECT 0.000 3485.195 3165.000 3487.015 ;
        RECT 0.000 3483.795 3160.600 3485.195 ;
        RECT 0.000 3481.975 3165.000 3483.795 ;
        RECT 0.000 3480.575 3160.600 3481.975 ;
        RECT 0.000 3469.555 3165.000 3480.575 ;
        RECT 0.000 3468.155 3160.600 3469.555 ;
        RECT 0.000 3466.795 3165.000 3468.155 ;
        RECT 0.000 3465.395 3160.600 3466.795 ;
        RECT 0.000 3463.575 3165.000 3465.395 ;
        RECT 0.000 3462.175 3160.600 3463.575 ;
        RECT 0.000 3460.355 3165.000 3462.175 ;
        RECT 0.000 3458.955 3160.600 3460.355 ;
        RECT 0.000 3454.375 3165.000 3458.955 ;
        RECT 0.000 3452.975 3160.600 3454.375 ;
        RECT 0.000 3448.395 3165.000 3452.975 ;
        RECT 0.000 3446.995 3160.600 3448.395 ;
        RECT 0.000 3445.175 3165.000 3446.995 ;
        RECT 0.000 3443.775 3160.600 3445.175 ;
        RECT 0.000 3443.280 3165.000 3443.775 ;
        RECT 0.000 3440.080 9.480 3443.280 ;
        RECT 120.840 3440.080 3042.640 3443.280 ;
        RECT 3155.320 3441.955 3165.000 3443.280 ;
        RECT 3155.320 3440.555 3160.600 3441.955 ;
        RECT 3155.320 3440.080 3165.000 3440.555 ;
        RECT 0.000 3438.880 3165.000 3440.080 ;
        RECT 0.000 3435.680 9.480 3438.880 ;
        RECT 120.840 3435.680 3042.640 3438.880 ;
        RECT 3155.320 3435.975 3165.000 3438.880 ;
        RECT 3155.320 3435.680 3160.600 3435.975 ;
        RECT 0.000 3434.575 3160.600 3435.680 ;
        RECT 0.000 3434.480 3165.000 3434.575 ;
        RECT 0.000 3431.280 9.480 3434.480 ;
        RECT 120.840 3431.280 3042.640 3434.480 ;
        RECT 3155.320 3431.280 3165.000 3434.480 ;
        RECT 0.000 3430.080 3165.000 3431.280 ;
        RECT 0.000 3426.880 9.480 3430.080 ;
        RECT 120.840 3426.880 3047.740 3430.080 ;
        RECT 3155.320 3426.880 3165.000 3430.080 ;
        RECT 0.000 3425.680 3165.000 3426.880 ;
        RECT 0.000 3422.480 9.480 3425.680 ;
        RECT 120.840 3422.480 3042.640 3425.680 ;
        RECT 3155.320 3422.480 3165.000 3425.680 ;
        RECT 0.000 3421.280 3165.000 3422.480 ;
        RECT 0.000 3418.080 9.480 3421.280 ;
        RECT 120.840 3418.080 3042.640 3421.280 ;
        RECT 3155.320 3418.080 3165.000 3421.280 ;
        RECT 0.000 3416.880 3165.000 3418.080 ;
        RECT 0.000 3413.680 9.480 3416.880 ;
        RECT 120.840 3413.680 3042.640 3416.880 ;
        RECT 3155.320 3413.680 3165.000 3416.880 ;
        RECT 0.000 3412.480 3165.000 3413.680 ;
        RECT 0.000 3409.280 9.480 3412.480 ;
        RECT 120.840 3409.280 3042.640 3412.480 ;
        RECT 3155.320 3409.280 3165.000 3412.480 ;
        RECT 0.000 3355.425 3165.000 3409.280 ;
        RECT 4.400 3354.025 3165.000 3355.425 ;
        RECT 0.000 3349.445 3165.000 3354.025 ;
        RECT 4.400 3348.045 3165.000 3349.445 ;
        RECT 0.000 3346.225 3165.000 3348.045 ;
        RECT 4.400 3344.825 3165.000 3346.225 ;
        RECT 0.000 3343.280 3165.000 3344.825 ;
        RECT 0.000 3343.005 9.480 3343.280 ;
        RECT 4.400 3341.605 9.480 3343.005 ;
        RECT 0.000 3340.080 9.480 3341.605 ;
        RECT 120.840 3340.080 3042.640 3343.280 ;
        RECT 3155.320 3340.080 3165.000 3343.280 ;
        RECT 0.000 3338.880 3165.000 3340.080 ;
        RECT 0.000 3337.025 9.480 3338.880 ;
        RECT 4.400 3335.680 9.480 3337.025 ;
        RECT 120.840 3335.680 3042.640 3338.880 ;
        RECT 3155.320 3335.680 3165.000 3338.880 ;
        RECT 4.400 3335.625 3165.000 3335.680 ;
        RECT 0.000 3334.480 3165.000 3335.625 ;
        RECT 0.000 3331.280 9.480 3334.480 ;
        RECT 120.840 3331.280 3042.640 3334.480 ;
        RECT 3155.320 3331.280 3165.000 3334.480 ;
        RECT 0.000 3331.045 3165.000 3331.280 ;
        RECT 4.400 3330.080 3165.000 3331.045 ;
        RECT 4.400 3329.645 9.480 3330.080 ;
        RECT 0.000 3327.825 9.480 3329.645 ;
        RECT 4.400 3326.880 9.480 3327.825 ;
        RECT 120.840 3326.880 3042.640 3330.080 ;
        RECT 3155.320 3326.880 3165.000 3330.080 ;
        RECT 4.400 3326.425 3165.000 3326.880 ;
        RECT 0.000 3325.680 3165.000 3326.425 ;
        RECT 0.000 3324.605 9.480 3325.680 ;
        RECT 4.690 3323.205 9.480 3324.605 ;
        RECT 0.000 3322.480 9.480 3323.205 ;
        RECT 120.840 3322.480 3042.640 3325.680 ;
        RECT 3155.320 3322.480 3165.000 3325.680 ;
        RECT 0.000 3321.845 3165.000 3322.480 ;
        RECT 4.400 3321.280 3165.000 3321.845 ;
        RECT 4.400 3320.445 9.480 3321.280 ;
        RECT 0.000 3318.080 9.480 3320.445 ;
        RECT 115.740 3318.080 3042.640 3321.280 ;
        RECT 3155.320 3318.080 3165.000 3321.280 ;
        RECT 0.000 3316.880 3165.000 3318.080 ;
        RECT 0.000 3313.680 9.480 3316.880 ;
        RECT 120.840 3313.680 3042.640 3316.880 ;
        RECT 3155.320 3313.680 3165.000 3316.880 ;
        RECT 0.000 3312.480 3165.000 3313.680 ;
        RECT 0.000 3309.425 9.480 3312.480 ;
        RECT 4.400 3309.280 9.480 3309.425 ;
        RECT 120.840 3309.280 3042.640 3312.480 ;
        RECT 3155.320 3309.280 3165.000 3312.480 ;
        RECT 4.400 3308.025 3165.000 3309.280 ;
        RECT 0.000 3306.205 3165.000 3308.025 ;
        RECT 4.400 3304.805 3165.000 3306.205 ;
        RECT 0.000 3302.985 3165.000 3304.805 ;
        RECT 4.400 3301.585 3165.000 3302.985 ;
        RECT 0.000 3300.225 3165.000 3301.585 ;
        RECT 4.400 3298.825 3165.000 3300.225 ;
        RECT 0.000 3291.025 3165.000 3298.825 ;
        RECT 4.400 3289.625 3165.000 3291.025 ;
        RECT 0.000 3287.805 3165.000 3289.625 ;
        RECT 4.400 3286.405 3165.000 3287.805 ;
        RECT 0.000 3284.585 3165.000 3286.405 ;
        RECT 4.400 3283.185 3165.000 3284.585 ;
        RECT 0.000 3281.815 3165.000 3283.185 ;
        RECT 0.000 3280.415 3160.600 3281.815 ;
        RECT 0.000 3278.595 3165.000 3280.415 ;
        RECT 0.000 3277.195 3160.600 3278.595 ;
        RECT 0.000 3275.375 3165.000 3277.195 ;
        RECT 0.000 3273.975 3160.600 3275.375 ;
        RECT 0.000 3266.175 3165.000 3273.975 ;
        RECT 0.000 3264.775 3160.600 3266.175 ;
        RECT 0.000 3263.415 3165.000 3264.775 ;
        RECT 0.000 3262.015 3160.600 3263.415 ;
        RECT 0.000 3260.195 3165.000 3262.015 ;
        RECT 0.000 3258.795 3160.600 3260.195 ;
        RECT 0.000 3256.975 3165.000 3258.795 ;
        RECT 0.000 3255.575 3160.600 3256.975 ;
        RECT 0.000 3244.555 3165.000 3255.575 ;
        RECT 0.000 3243.280 3160.600 3244.555 ;
        RECT 0.000 3240.080 9.480 3243.280 ;
        RECT 120.840 3240.080 3042.640 3243.280 ;
        RECT 3155.320 3243.155 3160.600 3243.280 ;
        RECT 3155.320 3241.795 3165.000 3243.155 ;
        RECT 3155.320 3240.395 3160.600 3241.795 ;
        RECT 3155.320 3240.080 3165.000 3240.395 ;
        RECT 0.000 3238.880 3165.000 3240.080 ;
        RECT 0.000 3235.680 9.480 3238.880 ;
        RECT 120.840 3235.680 3042.640 3238.880 ;
        RECT 3155.320 3238.575 3165.000 3238.880 ;
        RECT 3155.320 3237.175 3160.600 3238.575 ;
        RECT 3155.320 3235.680 3165.000 3237.175 ;
        RECT 0.000 3235.355 3165.000 3235.680 ;
        RECT 0.000 3234.480 3160.600 3235.355 ;
        RECT 0.000 3231.280 9.480 3234.480 ;
        RECT 120.840 3231.280 3042.640 3234.480 ;
        RECT 3155.320 3233.955 3160.600 3234.480 ;
        RECT 3155.320 3231.280 3165.000 3233.955 ;
        RECT 0.000 3230.080 3165.000 3231.280 ;
        RECT 0.000 3226.880 9.480 3230.080 ;
        RECT 120.840 3226.880 3047.740 3230.080 ;
        RECT 3155.320 3229.375 3165.000 3230.080 ;
        RECT 3155.320 3227.975 3160.600 3229.375 ;
        RECT 3155.320 3226.880 3165.000 3227.975 ;
        RECT 0.000 3225.680 3165.000 3226.880 ;
        RECT 0.000 3222.480 9.480 3225.680 ;
        RECT 120.840 3222.480 3042.640 3225.680 ;
        RECT 3155.320 3223.395 3165.000 3225.680 ;
        RECT 3155.320 3222.480 3160.600 3223.395 ;
        RECT 0.000 3221.995 3160.600 3222.480 ;
        RECT 0.000 3221.280 3165.000 3221.995 ;
        RECT 0.000 3218.080 9.480 3221.280 ;
        RECT 120.840 3218.080 3042.640 3221.280 ;
        RECT 3155.320 3220.175 3165.000 3221.280 ;
        RECT 3155.320 3218.775 3160.600 3220.175 ;
        RECT 3155.320 3218.080 3165.000 3218.775 ;
        RECT 0.000 3216.955 3165.000 3218.080 ;
        RECT 0.000 3216.880 3160.600 3216.955 ;
        RECT 0.000 3213.680 9.480 3216.880 ;
        RECT 120.840 3213.680 3042.640 3216.880 ;
        RECT 3155.320 3215.555 3160.600 3216.880 ;
        RECT 3155.320 3213.680 3165.000 3215.555 ;
        RECT 0.000 3212.480 3165.000 3213.680 ;
        RECT 0.000 3209.280 9.480 3212.480 ;
        RECT 120.840 3209.280 3042.640 3212.480 ;
        RECT 3155.320 3210.975 3165.000 3212.480 ;
        RECT 3155.320 3209.575 3160.600 3210.975 ;
        RECT 3155.320 3209.280 3165.000 3209.575 ;
        RECT 0.000 3143.280 3165.000 3209.280 ;
        RECT 0.000 3140.080 9.480 3143.280 ;
        RECT 120.840 3140.080 3042.640 3143.280 ;
        RECT 3155.320 3140.080 3165.000 3143.280 ;
        RECT 0.000 3139.425 3165.000 3140.080 ;
        RECT 4.400 3138.880 3165.000 3139.425 ;
        RECT 4.400 3138.025 9.480 3138.880 ;
        RECT 0.000 3135.680 9.480 3138.025 ;
        RECT 120.840 3135.680 3042.640 3138.880 ;
        RECT 3155.320 3135.680 3165.000 3138.880 ;
        RECT 0.000 3134.480 3165.000 3135.680 ;
        RECT 0.000 3133.445 9.480 3134.480 ;
        RECT 4.400 3132.045 9.480 3133.445 ;
        RECT 0.000 3131.280 9.480 3132.045 ;
        RECT 120.840 3131.280 3042.640 3134.480 ;
        RECT 3155.320 3131.280 3165.000 3134.480 ;
        RECT 0.000 3130.225 3165.000 3131.280 ;
        RECT 4.400 3130.080 3165.000 3130.225 ;
        RECT 4.400 3128.825 9.480 3130.080 ;
        RECT 0.000 3127.005 9.480 3128.825 ;
        RECT 4.400 3126.880 9.480 3127.005 ;
        RECT 120.840 3126.880 3042.640 3130.080 ;
        RECT 3155.320 3126.880 3165.000 3130.080 ;
        RECT 4.400 3125.680 3165.000 3126.880 ;
        RECT 4.400 3125.605 9.480 3125.680 ;
        RECT 0.000 3122.480 9.480 3125.605 ;
        RECT 115.740 3122.480 3042.640 3125.680 ;
        RECT 3155.320 3122.480 3165.000 3125.680 ;
        RECT 0.000 3121.280 3165.000 3122.480 ;
        RECT 0.000 3121.025 9.480 3121.280 ;
        RECT 4.400 3119.625 9.480 3121.025 ;
        RECT 0.000 3118.080 9.480 3119.625 ;
        RECT 120.840 3118.080 3042.640 3121.280 ;
        RECT 3155.320 3118.080 3165.000 3121.280 ;
        RECT 0.000 3116.880 3165.000 3118.080 ;
        RECT 0.000 3115.045 9.480 3116.880 ;
        RECT 4.400 3113.680 9.480 3115.045 ;
        RECT 120.840 3113.680 3042.640 3116.880 ;
        RECT 3155.320 3113.680 3165.000 3116.880 ;
        RECT 4.400 3113.645 3165.000 3113.680 ;
        RECT 0.000 3112.480 3165.000 3113.645 ;
        RECT 0.000 3111.825 9.480 3112.480 ;
        RECT 4.400 3110.425 9.480 3111.825 ;
        RECT 0.000 3109.280 9.480 3110.425 ;
        RECT 120.840 3109.280 3042.640 3112.480 ;
        RECT 3155.320 3109.280 3165.000 3112.480 ;
        RECT 0.000 3108.605 3165.000 3109.280 ;
        RECT 4.400 3107.205 3165.000 3108.605 ;
        RECT 0.000 3105.845 3165.000 3107.205 ;
        RECT 4.400 3104.445 3165.000 3105.845 ;
        RECT 0.000 3093.425 3165.000 3104.445 ;
        RECT 4.400 3092.025 3165.000 3093.425 ;
        RECT 0.000 3090.205 3165.000 3092.025 ;
        RECT 4.400 3088.805 3165.000 3090.205 ;
        RECT 0.000 3086.985 3165.000 3088.805 ;
        RECT 4.400 3085.585 3165.000 3086.985 ;
        RECT 0.000 3084.225 3165.000 3085.585 ;
        RECT 4.400 3082.825 3165.000 3084.225 ;
        RECT 0.000 3075.025 3165.000 3082.825 ;
        RECT 4.400 3073.625 3165.000 3075.025 ;
        RECT 0.000 3071.805 3165.000 3073.625 ;
        RECT 4.400 3070.405 3165.000 3071.805 ;
        RECT 0.000 3068.585 3165.000 3070.405 ;
        RECT 4.400 3067.185 3165.000 3068.585 ;
        RECT 0.000 3055.815 3165.000 3067.185 ;
        RECT 0.000 3054.415 3160.600 3055.815 ;
        RECT 0.000 3052.595 3165.000 3054.415 ;
        RECT 0.000 3051.195 3160.600 3052.595 ;
        RECT 0.000 3049.375 3165.000 3051.195 ;
        RECT 0.000 3047.975 3160.600 3049.375 ;
        RECT 0.000 3043.280 3165.000 3047.975 ;
        RECT 0.000 3040.080 9.480 3043.280 ;
        RECT 120.840 3040.080 3042.640 3043.280 ;
        RECT 3155.320 3040.175 3165.000 3043.280 ;
        RECT 3155.320 3040.080 3160.600 3040.175 ;
        RECT 0.000 3038.880 3160.600 3040.080 ;
        RECT 0.000 3035.680 9.480 3038.880 ;
        RECT 120.840 3035.680 3042.640 3038.880 ;
        RECT 3155.320 3038.775 3160.600 3038.880 ;
        RECT 3155.320 3037.415 3165.000 3038.775 ;
        RECT 3155.320 3036.015 3160.600 3037.415 ;
        RECT 3155.320 3035.680 3165.000 3036.015 ;
        RECT 0.000 3034.480 3165.000 3035.680 ;
        RECT 0.000 3031.280 9.480 3034.480 ;
        RECT 120.840 3031.280 3047.740 3034.480 ;
        RECT 3155.320 3034.195 3165.000 3034.480 ;
        RECT 3155.320 3032.795 3160.600 3034.195 ;
        RECT 3155.320 3031.280 3165.000 3032.795 ;
        RECT 0.000 3030.975 3165.000 3031.280 ;
        RECT 0.000 3030.080 3160.600 3030.975 ;
        RECT 0.000 3026.880 9.480 3030.080 ;
        RECT 120.840 3026.880 3047.740 3030.080 ;
        RECT 3155.320 3029.575 3160.600 3030.080 ;
        RECT 3155.320 3026.880 3165.000 3029.575 ;
        RECT 0.000 3025.680 3165.000 3026.880 ;
        RECT 0.000 3022.480 9.480 3025.680 ;
        RECT 120.840 3022.480 3042.640 3025.680 ;
        RECT 3155.320 3022.480 3165.000 3025.680 ;
        RECT 0.000 3021.280 3165.000 3022.480 ;
        RECT 0.000 3018.080 9.480 3021.280 ;
        RECT 120.840 3018.080 3042.640 3021.280 ;
        RECT 3155.320 3018.555 3165.000 3021.280 ;
        RECT 3155.320 3018.080 3160.600 3018.555 ;
        RECT 0.000 3017.155 3160.600 3018.080 ;
        RECT 0.000 3016.880 3165.000 3017.155 ;
        RECT 0.000 3013.680 9.480 3016.880 ;
        RECT 120.840 3013.680 3042.640 3016.880 ;
        RECT 3155.320 3015.795 3165.000 3016.880 ;
        RECT 3155.320 3014.395 3160.600 3015.795 ;
        RECT 3155.320 3013.680 3165.000 3014.395 ;
        RECT 0.000 3012.575 3165.000 3013.680 ;
        RECT 0.000 3012.480 3160.600 3012.575 ;
        RECT 0.000 3009.280 9.480 3012.480 ;
        RECT 120.840 3009.280 3042.640 3012.480 ;
        RECT 3155.320 3011.175 3160.600 3012.480 ;
        RECT 3155.320 3009.355 3165.000 3011.175 ;
        RECT 3155.320 3009.280 3160.600 3009.355 ;
        RECT 0.000 3007.955 3160.600 3009.280 ;
        RECT 0.000 3003.375 3165.000 3007.955 ;
        RECT 0.000 3001.975 3160.600 3003.375 ;
        RECT 0.000 2997.395 3165.000 3001.975 ;
        RECT 0.000 2995.995 3160.600 2997.395 ;
        RECT 0.000 2994.175 3165.000 2995.995 ;
        RECT 0.000 2992.775 3160.600 2994.175 ;
        RECT 0.000 2990.955 3165.000 2992.775 ;
        RECT 0.000 2989.555 3160.600 2990.955 ;
        RECT 0.000 2984.975 3165.000 2989.555 ;
        RECT 0.000 2983.575 3160.600 2984.975 ;
        RECT 0.000 2943.280 3165.000 2983.575 ;
        RECT 0.000 2940.080 9.480 2943.280 ;
        RECT 120.840 2940.080 3042.640 2943.280 ;
        RECT 3155.320 2940.080 3165.000 2943.280 ;
        RECT 0.000 2938.880 3165.000 2940.080 ;
        RECT 0.000 2935.680 9.480 2938.880 ;
        RECT 120.840 2935.680 3042.640 2938.880 ;
        RECT 3155.320 2935.680 3165.000 2938.880 ;
        RECT 0.000 2934.480 3165.000 2935.680 ;
        RECT 0.000 2931.280 9.480 2934.480 ;
        RECT 120.840 2931.280 3042.640 2934.480 ;
        RECT 3155.320 2931.280 3165.000 2934.480 ;
        RECT 0.000 2930.080 3165.000 2931.280 ;
        RECT 0.000 2926.880 9.480 2930.080 ;
        RECT 115.740 2926.880 3042.640 2930.080 ;
        RECT 3155.320 2926.880 3165.000 2930.080 ;
        RECT 0.000 2925.680 3165.000 2926.880 ;
        RECT 0.000 2923.425 9.480 2925.680 ;
        RECT 4.400 2922.480 9.480 2923.425 ;
        RECT 120.840 2922.480 3042.640 2925.680 ;
        RECT 3155.320 2922.480 3165.000 2925.680 ;
        RECT 4.400 2922.025 3165.000 2922.480 ;
        RECT 0.000 2921.280 3165.000 2922.025 ;
        RECT 0.000 2918.080 9.480 2921.280 ;
        RECT 120.840 2918.080 3042.640 2921.280 ;
        RECT 3155.320 2918.080 3165.000 2921.280 ;
        RECT 0.000 2917.445 3165.000 2918.080 ;
        RECT 4.400 2916.880 3165.000 2917.445 ;
        RECT 4.400 2916.045 9.480 2916.880 ;
        RECT 0.000 2914.225 9.480 2916.045 ;
        RECT 4.400 2913.680 9.480 2914.225 ;
        RECT 120.840 2913.680 3042.640 2916.880 ;
        RECT 3155.320 2913.680 3165.000 2916.880 ;
        RECT 4.400 2912.825 3165.000 2913.680 ;
        RECT 0.000 2912.480 3165.000 2912.825 ;
        RECT 0.000 2911.005 9.480 2912.480 ;
        RECT 4.400 2909.605 9.480 2911.005 ;
        RECT 0.000 2909.280 9.480 2909.605 ;
        RECT 120.840 2909.280 3042.640 2912.480 ;
        RECT 3155.320 2909.280 3165.000 2912.480 ;
        RECT 0.000 2905.025 3165.000 2909.280 ;
        RECT 4.400 2903.625 3165.000 2905.025 ;
        RECT 0.000 2899.045 3165.000 2903.625 ;
        RECT 4.400 2897.645 3165.000 2899.045 ;
        RECT 0.000 2895.825 3165.000 2897.645 ;
        RECT 4.400 2894.425 3165.000 2895.825 ;
        RECT 0.000 2892.605 3165.000 2894.425 ;
        RECT 4.400 2891.205 3165.000 2892.605 ;
        RECT 0.000 2889.845 3165.000 2891.205 ;
        RECT 4.400 2888.445 3165.000 2889.845 ;
        RECT 0.000 2877.425 3165.000 2888.445 ;
        RECT 4.400 2876.025 3165.000 2877.425 ;
        RECT 0.000 2874.205 3165.000 2876.025 ;
        RECT 4.400 2872.805 3165.000 2874.205 ;
        RECT 0.000 2870.985 3165.000 2872.805 ;
        RECT 4.400 2869.585 3165.000 2870.985 ;
        RECT 0.000 2868.225 3165.000 2869.585 ;
        RECT 4.400 2866.825 3165.000 2868.225 ;
        RECT 0.000 2859.025 3165.000 2866.825 ;
        RECT 4.400 2857.625 3165.000 2859.025 ;
        RECT 0.000 2855.805 3165.000 2857.625 ;
        RECT 4.400 2854.405 3165.000 2855.805 ;
        RECT 0.000 2852.585 3165.000 2854.405 ;
        RECT 4.400 2851.185 3165.000 2852.585 ;
        RECT 0.000 2843.280 3165.000 2851.185 ;
        RECT 0.000 2840.080 9.480 2843.280 ;
        RECT 120.840 2840.080 3042.640 2843.280 ;
        RECT 3155.320 2840.080 3165.000 2843.280 ;
        RECT 0.000 2838.880 3165.000 2840.080 ;
        RECT 0.000 2835.680 9.480 2838.880 ;
        RECT 120.840 2835.680 3042.640 2838.880 ;
        RECT 3155.320 2835.680 3165.000 2838.880 ;
        RECT 0.000 2834.480 3165.000 2835.680 ;
        RECT 0.000 2831.280 9.480 2834.480 ;
        RECT 120.840 2831.280 3047.740 2834.480 ;
        RECT 3155.320 2831.280 3165.000 2834.480 ;
        RECT 0.000 2830.815 3165.000 2831.280 ;
        RECT 0.000 2830.080 3160.600 2830.815 ;
        RECT 0.000 2826.880 9.480 2830.080 ;
        RECT 120.840 2826.880 3042.640 2830.080 ;
        RECT 3155.320 2829.415 3160.600 2830.080 ;
        RECT 3155.320 2827.595 3165.000 2829.415 ;
        RECT 3155.320 2826.880 3160.600 2827.595 ;
        RECT 0.000 2826.195 3160.600 2826.880 ;
        RECT 0.000 2825.680 3165.000 2826.195 ;
        RECT 0.000 2822.480 9.480 2825.680 ;
        RECT 120.840 2822.480 3042.640 2825.680 ;
        RECT 3155.320 2824.375 3165.000 2825.680 ;
        RECT 3155.320 2822.975 3160.600 2824.375 ;
        RECT 3155.320 2822.480 3165.000 2822.975 ;
        RECT 0.000 2821.280 3165.000 2822.480 ;
        RECT 0.000 2818.080 9.480 2821.280 ;
        RECT 120.840 2818.080 3042.640 2821.280 ;
        RECT 3155.320 2818.080 3165.000 2821.280 ;
        RECT 0.000 2816.880 3165.000 2818.080 ;
        RECT 0.000 2813.680 9.480 2816.880 ;
        RECT 120.840 2813.680 3042.640 2816.880 ;
        RECT 3155.320 2815.175 3165.000 2816.880 ;
        RECT 3155.320 2813.775 3160.600 2815.175 ;
        RECT 3155.320 2813.680 3165.000 2813.775 ;
        RECT 0.000 2812.480 3165.000 2813.680 ;
        RECT 0.000 2809.280 9.480 2812.480 ;
        RECT 120.840 2809.280 3042.640 2812.480 ;
        RECT 3155.320 2812.415 3165.000 2812.480 ;
        RECT 3155.320 2811.015 3160.600 2812.415 ;
        RECT 3155.320 2809.280 3165.000 2811.015 ;
        RECT 0.000 2809.195 3165.000 2809.280 ;
        RECT 0.000 2807.795 3160.600 2809.195 ;
        RECT 0.000 2805.975 3165.000 2807.795 ;
        RECT 0.000 2804.575 3160.600 2805.975 ;
        RECT 0.000 2793.555 3165.000 2804.575 ;
        RECT 0.000 2792.155 3160.600 2793.555 ;
        RECT 0.000 2790.795 3165.000 2792.155 ;
        RECT 0.000 2789.395 3160.600 2790.795 ;
        RECT 0.000 2787.575 3165.000 2789.395 ;
        RECT 0.000 2786.175 3160.600 2787.575 ;
        RECT 0.000 2784.355 3165.000 2786.175 ;
        RECT 0.000 2782.955 3160.600 2784.355 ;
        RECT 0.000 2778.375 3165.000 2782.955 ;
        RECT 0.000 2776.975 3160.600 2778.375 ;
        RECT 0.000 2772.395 3165.000 2776.975 ;
        RECT 0.000 2770.995 3160.600 2772.395 ;
        RECT 0.000 2769.175 3165.000 2770.995 ;
        RECT 0.000 2767.775 3160.600 2769.175 ;
        RECT 0.000 2765.955 3165.000 2767.775 ;
        RECT 0.000 2764.555 3160.600 2765.955 ;
        RECT 0.000 2759.975 3165.000 2764.555 ;
        RECT 0.000 2758.575 3160.600 2759.975 ;
        RECT 0.000 2743.280 3165.000 2758.575 ;
        RECT 0.000 2740.080 9.480 2743.280 ;
        RECT 120.840 2740.080 3042.640 2743.280 ;
        RECT 3155.320 2740.080 3165.000 2743.280 ;
        RECT 0.000 2738.880 3165.000 2740.080 ;
        RECT 0.000 2735.680 9.480 2738.880 ;
        RECT 120.840 2735.680 3042.640 2738.880 ;
        RECT 3155.320 2735.680 3165.000 2738.880 ;
        RECT 0.000 2734.480 3165.000 2735.680 ;
        RECT 0.000 2731.280 9.480 2734.480 ;
        RECT 115.740 2731.280 3042.640 2734.480 ;
        RECT 3155.320 2731.280 3165.000 2734.480 ;
        RECT 0.000 2730.080 3165.000 2731.280 ;
        RECT 0.000 2726.880 9.480 2730.080 ;
        RECT 120.840 2726.880 3042.640 2730.080 ;
        RECT 3155.320 2726.880 3165.000 2730.080 ;
        RECT 0.000 2725.680 3165.000 2726.880 ;
        RECT 0.000 2722.480 9.480 2725.680 ;
        RECT 120.840 2722.480 3042.640 2725.680 ;
        RECT 3155.320 2722.480 3165.000 2725.680 ;
        RECT 0.000 2721.280 3165.000 2722.480 ;
        RECT 0.000 2718.080 9.480 2721.280 ;
        RECT 120.840 2718.080 3042.640 2721.280 ;
        RECT 3155.320 2718.080 3165.000 2721.280 ;
        RECT 0.000 2716.880 3165.000 2718.080 ;
        RECT 0.000 2713.680 9.480 2716.880 ;
        RECT 120.840 2713.680 3042.640 2716.880 ;
        RECT 3155.320 2713.680 3165.000 2716.880 ;
        RECT 0.000 2712.480 3165.000 2713.680 ;
        RECT 0.000 2709.280 9.480 2712.480 ;
        RECT 120.840 2709.280 3042.640 2712.480 ;
        RECT 3155.320 2709.280 3165.000 2712.480 ;
        RECT 0.000 2707.425 3165.000 2709.280 ;
        RECT 4.400 2706.025 3165.000 2707.425 ;
        RECT 0.000 2701.445 3165.000 2706.025 ;
        RECT 4.400 2700.045 3165.000 2701.445 ;
        RECT 0.000 2698.225 3165.000 2700.045 ;
        RECT 4.400 2696.825 3165.000 2698.225 ;
        RECT 0.000 2695.005 3165.000 2696.825 ;
        RECT 4.400 2693.605 3165.000 2695.005 ;
        RECT 0.000 2689.025 3165.000 2693.605 ;
        RECT 4.400 2687.625 3165.000 2689.025 ;
        RECT 0.000 2683.045 3165.000 2687.625 ;
        RECT 4.400 2681.645 3165.000 2683.045 ;
        RECT 0.000 2679.825 3165.000 2681.645 ;
        RECT 4.400 2678.425 3165.000 2679.825 ;
        RECT 0.000 2676.605 3165.000 2678.425 ;
        RECT 4.400 2675.205 3165.000 2676.605 ;
        RECT 0.000 2673.845 3165.000 2675.205 ;
        RECT 4.400 2672.445 3165.000 2673.845 ;
        RECT 0.000 2661.425 3165.000 2672.445 ;
        RECT 4.400 2660.025 3165.000 2661.425 ;
        RECT 0.000 2658.205 3165.000 2660.025 ;
        RECT 4.400 2656.805 3165.000 2658.205 ;
        RECT 0.000 2654.985 3165.000 2656.805 ;
        RECT 4.400 2653.585 3165.000 2654.985 ;
        RECT 0.000 2652.225 3165.000 2653.585 ;
        RECT 4.400 2650.825 3165.000 2652.225 ;
        RECT 0.000 2643.280 3165.000 2650.825 ;
        RECT 0.000 2643.025 9.480 2643.280 ;
        RECT 4.400 2641.625 9.480 2643.025 ;
        RECT 0.000 2640.080 9.480 2641.625 ;
        RECT 120.840 2640.080 3042.640 2643.280 ;
        RECT 3155.320 2640.080 3165.000 2643.280 ;
        RECT 0.000 2639.805 3165.000 2640.080 ;
        RECT 4.400 2638.880 3165.000 2639.805 ;
        RECT 4.400 2638.405 9.480 2638.880 ;
        RECT 0.000 2636.585 9.480 2638.405 ;
        RECT 4.400 2635.680 9.480 2636.585 ;
        RECT 120.840 2635.680 3042.640 2638.880 ;
        RECT 3155.320 2635.680 3165.000 2638.880 ;
        RECT 4.400 2635.185 3165.000 2635.680 ;
        RECT 0.000 2634.480 3165.000 2635.185 ;
        RECT 0.000 2631.280 9.480 2634.480 ;
        RECT 120.840 2631.280 3047.740 2634.480 ;
        RECT 3155.320 2631.280 3165.000 2634.480 ;
        RECT 0.000 2630.080 3165.000 2631.280 ;
        RECT 0.000 2626.880 9.480 2630.080 ;
        RECT 120.840 2626.880 3042.640 2630.080 ;
        RECT 3155.320 2626.880 3165.000 2630.080 ;
        RECT 0.000 2625.680 3165.000 2626.880 ;
        RECT 0.000 2622.480 9.480 2625.680 ;
        RECT 120.840 2622.480 3042.640 2625.680 ;
        RECT 3155.320 2622.480 3165.000 2625.680 ;
        RECT 0.000 2621.280 3165.000 2622.480 ;
        RECT 0.000 2618.080 9.480 2621.280 ;
        RECT 120.840 2618.080 3042.640 2621.280 ;
        RECT 3155.320 2618.080 3165.000 2621.280 ;
        RECT 0.000 2616.880 3165.000 2618.080 ;
        RECT 0.000 2613.680 9.480 2616.880 ;
        RECT 120.840 2613.680 3042.640 2616.880 ;
        RECT 3155.320 2613.680 3165.000 2616.880 ;
        RECT 0.000 2612.480 3165.000 2613.680 ;
        RECT 0.000 2609.280 9.480 2612.480 ;
        RECT 120.840 2609.280 3042.640 2612.480 ;
        RECT 3155.320 2609.280 3165.000 2612.480 ;
        RECT 0.000 2604.815 3165.000 2609.280 ;
        RECT 0.000 2603.415 3160.600 2604.815 ;
        RECT 0.000 2601.595 3165.000 2603.415 ;
        RECT 0.000 2600.195 3160.600 2601.595 ;
        RECT 0.000 2598.375 3165.000 2600.195 ;
        RECT 0.000 2596.975 3160.600 2598.375 ;
        RECT 0.000 2589.175 3165.000 2596.975 ;
        RECT 0.000 2587.775 3160.600 2589.175 ;
        RECT 0.000 2586.415 3165.000 2587.775 ;
        RECT 0.000 2585.015 3160.600 2586.415 ;
        RECT 0.000 2583.195 3165.000 2585.015 ;
        RECT 0.000 2581.795 3160.600 2583.195 ;
        RECT 0.000 2579.975 3165.000 2581.795 ;
        RECT 0.000 2578.575 3160.600 2579.975 ;
        RECT 0.000 2567.555 3165.000 2578.575 ;
        RECT 0.000 2566.155 3160.600 2567.555 ;
        RECT 0.000 2564.795 3165.000 2566.155 ;
        RECT 0.000 2563.395 3160.600 2564.795 ;
        RECT 0.000 2561.575 3165.000 2563.395 ;
        RECT 0.000 2560.175 3160.600 2561.575 ;
        RECT 0.000 2558.355 3165.000 2560.175 ;
        RECT 0.000 2556.955 3160.600 2558.355 ;
        RECT 0.000 2552.375 3165.000 2556.955 ;
        RECT 0.000 2550.975 3160.600 2552.375 ;
        RECT 0.000 2546.395 3165.000 2550.975 ;
        RECT 0.000 2544.995 3160.600 2546.395 ;
        RECT 0.000 2543.280 3165.000 2544.995 ;
        RECT 0.000 2540.080 9.480 2543.280 ;
        RECT 120.840 2540.080 3042.640 2543.280 ;
        RECT 3155.320 2543.175 3165.000 2543.280 ;
        RECT 3155.320 2541.775 3160.600 2543.175 ;
        RECT 3155.320 2540.080 3165.000 2541.775 ;
        RECT 0.000 2539.955 3165.000 2540.080 ;
        RECT 0.000 2538.880 3160.600 2539.955 ;
        RECT 0.000 2535.680 9.480 2538.880 ;
        RECT 115.740 2535.680 3042.640 2538.880 ;
        RECT 3155.320 2538.555 3160.600 2538.880 ;
        RECT 3155.320 2535.680 3165.000 2538.555 ;
        RECT 0.000 2534.480 3165.000 2535.680 ;
        RECT 0.000 2531.280 9.480 2534.480 ;
        RECT 120.840 2531.280 3042.640 2534.480 ;
        RECT 3155.320 2533.975 3165.000 2534.480 ;
        RECT 3155.320 2532.575 3160.600 2533.975 ;
        RECT 3155.320 2531.280 3165.000 2532.575 ;
        RECT 0.000 2530.080 3165.000 2531.280 ;
        RECT 0.000 2526.880 9.480 2530.080 ;
        RECT 120.840 2526.880 3042.640 2530.080 ;
        RECT 3155.320 2526.880 3165.000 2530.080 ;
        RECT 0.000 2525.680 3165.000 2526.880 ;
        RECT 0.000 2522.480 9.480 2525.680 ;
        RECT 120.840 2522.480 3042.640 2525.680 ;
        RECT 3155.320 2522.480 3165.000 2525.680 ;
        RECT 0.000 2521.280 3165.000 2522.480 ;
        RECT 0.000 2518.080 9.480 2521.280 ;
        RECT 120.840 2518.080 3042.640 2521.280 ;
        RECT 3155.320 2518.080 3165.000 2521.280 ;
        RECT 0.000 2516.880 3165.000 2518.080 ;
        RECT 0.000 2513.680 9.480 2516.880 ;
        RECT 120.840 2513.680 3042.640 2516.880 ;
        RECT 3155.320 2513.680 3165.000 2516.880 ;
        RECT 0.000 2512.480 3165.000 2513.680 ;
        RECT 0.000 2509.280 9.480 2512.480 ;
        RECT 120.840 2509.280 3042.640 2512.480 ;
        RECT 3155.320 2509.280 3165.000 2512.480 ;
        RECT 0.000 2491.425 3165.000 2509.280 ;
        RECT 4.400 2490.025 3165.000 2491.425 ;
        RECT 0.000 2485.445 3165.000 2490.025 ;
        RECT 4.400 2484.045 3165.000 2485.445 ;
        RECT 0.000 2482.225 3165.000 2484.045 ;
        RECT 4.400 2480.825 3165.000 2482.225 ;
        RECT 0.000 2479.005 3165.000 2480.825 ;
        RECT 4.400 2477.605 3165.000 2479.005 ;
        RECT 0.000 2473.025 3165.000 2477.605 ;
        RECT 4.400 2471.625 3165.000 2473.025 ;
        RECT 0.000 2467.045 3165.000 2471.625 ;
        RECT 4.400 2465.645 3165.000 2467.045 ;
        RECT 0.000 2463.825 3165.000 2465.645 ;
        RECT 4.400 2462.425 3165.000 2463.825 ;
        RECT 0.000 2460.605 3165.000 2462.425 ;
        RECT 4.400 2459.205 3165.000 2460.605 ;
        RECT 0.000 2457.845 3165.000 2459.205 ;
        RECT 4.400 2456.445 3165.000 2457.845 ;
        RECT 0.000 2445.425 3165.000 2456.445 ;
        RECT 4.400 2444.025 3165.000 2445.425 ;
        RECT 0.000 2443.280 3165.000 2444.025 ;
        RECT 0.000 2442.205 9.480 2443.280 ;
        RECT 4.400 2440.805 9.480 2442.205 ;
        RECT 0.000 2440.080 9.480 2440.805 ;
        RECT 120.840 2440.080 3042.640 2443.280 ;
        RECT 3155.320 2440.080 3165.000 2443.280 ;
        RECT 0.000 2438.985 3165.000 2440.080 ;
        RECT 4.400 2438.880 3165.000 2438.985 ;
        RECT 4.400 2437.585 9.480 2438.880 ;
        RECT 0.000 2436.225 9.480 2437.585 ;
        RECT 4.400 2435.680 9.480 2436.225 ;
        RECT 120.840 2435.680 3042.640 2438.880 ;
        RECT 3155.320 2435.680 3165.000 2438.880 ;
        RECT 4.400 2434.825 3165.000 2435.680 ;
        RECT 0.000 2434.480 3165.000 2434.825 ;
        RECT 0.000 2431.280 9.480 2434.480 ;
        RECT 120.840 2431.280 3047.740 2434.480 ;
        RECT 3155.320 2431.280 3165.000 2434.480 ;
        RECT 0.000 2430.080 3165.000 2431.280 ;
        RECT 0.000 2427.025 9.480 2430.080 ;
        RECT 4.400 2426.880 9.480 2427.025 ;
        RECT 120.840 2426.880 3042.640 2430.080 ;
        RECT 3155.320 2426.880 3165.000 2430.080 ;
        RECT 4.400 2425.680 3165.000 2426.880 ;
        RECT 4.400 2425.625 9.480 2425.680 ;
        RECT 0.000 2423.805 9.480 2425.625 ;
        RECT 4.400 2422.480 9.480 2423.805 ;
        RECT 120.840 2422.480 3042.640 2425.680 ;
        RECT 3155.320 2422.480 3165.000 2425.680 ;
        RECT 4.400 2422.405 3165.000 2422.480 ;
        RECT 0.000 2421.280 3165.000 2422.405 ;
        RECT 0.000 2420.585 9.480 2421.280 ;
        RECT 4.400 2419.185 9.480 2420.585 ;
        RECT 0.000 2418.080 9.480 2419.185 ;
        RECT 120.840 2418.080 3042.640 2421.280 ;
        RECT 3155.320 2418.080 3165.000 2421.280 ;
        RECT 0.000 2416.880 3165.000 2418.080 ;
        RECT 0.000 2413.680 9.480 2416.880 ;
        RECT 120.840 2413.680 3042.640 2416.880 ;
        RECT 3155.320 2413.680 3165.000 2416.880 ;
        RECT 0.000 2412.480 3165.000 2413.680 ;
        RECT 0.000 2409.280 9.480 2412.480 ;
        RECT 120.840 2409.280 3042.640 2412.480 ;
        RECT 3155.320 2409.280 3165.000 2412.480 ;
        RECT 0.000 2383.005 3165.000 2409.280 ;
        RECT 0.000 2359.060 3178.020 2383.005 ;
        RECT 0.000 2343.280 3165.000 2359.060 ;
        RECT 0.000 2340.080 9.480 2343.280 ;
        RECT 115.740 2340.080 3042.640 2343.280 ;
        RECT 3155.320 2340.080 3165.000 2343.280 ;
        RECT 0.000 2338.880 3165.000 2340.080 ;
        RECT 0.000 2335.680 9.480 2338.880 ;
        RECT 120.840 2335.680 3042.640 2338.880 ;
        RECT 3155.320 2335.680 3165.000 2338.880 ;
        RECT 0.000 2334.480 3165.000 2335.680 ;
        RECT 0.000 2331.280 9.480 2334.480 ;
        RECT 120.840 2331.280 3042.640 2334.480 ;
        RECT 3155.320 2333.090 3165.000 2334.480 ;
        RECT 3155.320 2331.280 3178.020 2333.090 ;
        RECT 0.000 2330.080 3178.020 2331.280 ;
        RECT 0.000 2326.880 9.480 2330.080 ;
        RECT 120.840 2326.880 3042.640 2330.080 ;
        RECT 3155.320 2326.880 3178.020 2330.080 ;
        RECT 0.000 2325.680 3178.020 2326.880 ;
        RECT 0.000 2322.480 9.480 2325.680 ;
        RECT 120.840 2322.480 3042.640 2325.680 ;
        RECT 3155.320 2322.480 3178.020 2325.680 ;
        RECT 0.000 2321.280 3178.020 2322.480 ;
        RECT 0.000 2318.080 9.480 2321.280 ;
        RECT 120.840 2318.080 3042.640 2321.280 ;
        RECT 3155.320 2318.080 3178.020 2321.280 ;
        RECT 0.000 2316.880 3178.020 2318.080 ;
        RECT 0.000 2313.680 9.480 2316.880 ;
        RECT 120.840 2313.680 3042.640 2316.880 ;
        RECT 3155.320 2313.680 3178.020 2316.880 ;
        RECT 0.000 2312.480 3178.020 2313.680 ;
        RECT 0.000 2309.280 9.480 2312.480 ;
        RECT 120.840 2309.280 3042.640 2312.480 ;
        RECT 3155.320 2309.280 3178.020 2312.480 ;
        RECT 0.000 2309.145 3178.020 2309.280 ;
        RECT 0.000 2278.790 3165.000 2309.145 ;
        RECT -16.080 2254.845 3165.000 2278.790 ;
        RECT 0.000 2243.280 3165.000 2254.845 ;
        RECT 0.000 2240.080 9.480 2243.280 ;
        RECT 120.840 2240.080 3042.640 2243.280 ;
        RECT 3155.320 2240.080 3165.000 2243.280 ;
        RECT 0.000 2238.880 3165.000 2240.080 ;
        RECT 0.000 2235.680 9.480 2238.880 ;
        RECT 120.840 2235.680 3042.640 2238.880 ;
        RECT 3155.320 2235.680 3165.000 2238.880 ;
        RECT 0.000 2234.480 3165.000 2235.680 ;
        RECT 0.000 2231.280 9.480 2234.480 ;
        RECT 120.840 2231.280 3047.740 2234.480 ;
        RECT 3155.320 2231.280 3165.000 2234.480 ;
        RECT 0.000 2230.080 3165.000 2231.280 ;
        RECT 0.000 2228.895 9.480 2230.080 ;
        RECT -16.080 2226.880 9.480 2228.895 ;
        RECT 120.840 2226.880 3042.640 2230.080 ;
        RECT 3155.320 2226.880 3165.000 2230.080 ;
        RECT -16.080 2225.680 3165.000 2226.880 ;
        RECT -16.080 2222.480 9.480 2225.680 ;
        RECT 120.840 2222.480 3042.640 2225.680 ;
        RECT 3155.320 2222.480 3165.000 2225.680 ;
        RECT -16.080 2221.280 3165.000 2222.480 ;
        RECT -16.080 2218.080 9.480 2221.280 ;
        RECT 120.840 2218.080 3042.640 2221.280 ;
        RECT 3155.320 2218.080 3165.000 2221.280 ;
        RECT -16.080 2216.880 3165.000 2218.080 ;
        RECT -16.080 2213.680 9.480 2216.880 ;
        RECT 120.840 2213.680 3042.640 2216.880 ;
        RECT 3155.320 2213.680 3165.000 2216.880 ;
        RECT -16.080 2212.480 3165.000 2213.680 ;
        RECT -16.080 2209.280 9.480 2212.480 ;
        RECT 115.740 2209.280 3042.640 2212.480 ;
        RECT 3155.320 2209.280 3165.000 2212.480 ;
        RECT -16.080 2204.950 3165.000 2209.280 ;
        RECT 0.000 2163.000 3165.000 2204.950 ;
        RECT 0.000 2143.280 3178.020 2163.000 ;
        RECT 0.000 2140.080 9.480 2143.280 ;
        RECT 120.840 2140.080 3042.640 2143.280 ;
        RECT 3155.320 2140.080 3178.020 2143.280 ;
        RECT 0.000 2139.055 3178.020 2140.080 ;
        RECT 0.000 2138.880 3165.000 2139.055 ;
        RECT 0.000 2135.680 9.480 2138.880 ;
        RECT 120.840 2135.680 3042.640 2138.880 ;
        RECT 3155.320 2137.450 3165.000 2138.880 ;
        RECT 3155.320 2135.680 3176.020 2137.450 ;
        RECT 0.000 2134.480 3176.020 2135.680 ;
        RECT 0.000 2131.280 9.480 2134.480 ;
        RECT 120.840 2131.280 3042.640 2134.480 ;
        RECT 3155.320 2131.280 3176.020 2134.480 ;
        RECT 0.000 2130.080 3176.020 2131.280 ;
        RECT 0.000 2126.880 9.480 2130.080 ;
        RECT 120.840 2126.880 3042.640 2130.080 ;
        RECT 3155.320 2126.880 3176.020 2130.080 ;
        RECT 0.000 2125.680 3176.020 2126.880 ;
        RECT 0.000 2122.480 9.480 2125.680 ;
        RECT 120.840 2122.480 3042.640 2125.680 ;
        RECT 3155.320 2122.480 3176.020 2125.680 ;
        RECT 0.000 2121.280 3176.020 2122.480 ;
        RECT 0.000 2118.080 9.480 2121.280 ;
        RECT 120.840 2118.080 3042.640 2121.280 ;
        RECT 3155.320 2118.080 3176.020 2121.280 ;
        RECT 0.000 2116.880 3176.020 2118.080 ;
        RECT 0.000 2113.680 9.480 2116.880 ;
        RECT 120.840 2113.680 3042.640 2116.880 ;
        RECT 3155.320 2114.345 3176.020 2116.880 ;
        RECT 3155.320 2113.680 3165.000 2114.345 ;
        RECT 0.000 2112.745 3165.000 2113.680 ;
        RECT 0.000 2112.480 3178.020 2112.745 ;
        RECT 0.000 2109.280 9.480 2112.480 ;
        RECT 120.840 2109.280 3042.640 2112.480 ;
        RECT 3155.320 2109.280 3178.020 2112.480 ;
        RECT 0.000 2088.800 3178.020 2109.280 ;
        RECT 0.000 2068.200 3165.000 2088.800 ;
        RECT -16.080 2044.255 3165.000 2068.200 ;
        RECT 0.000 2043.280 3165.000 2044.255 ;
        RECT 0.000 2042.650 9.480 2043.280 ;
        RECT -11.080 2040.080 9.480 2042.650 ;
        RECT 120.840 2040.080 3042.640 2043.280 ;
        RECT 3155.320 2040.080 3165.000 2043.280 ;
        RECT -11.080 2038.880 3165.000 2040.080 ;
        RECT -11.080 2035.680 9.480 2038.880 ;
        RECT 120.840 2035.680 3042.640 2038.880 ;
        RECT 3155.320 2035.680 3165.000 2038.880 ;
        RECT -11.080 2034.480 3165.000 2035.680 ;
        RECT -11.080 2031.280 9.480 2034.480 ;
        RECT 120.840 2031.280 3047.740 2034.480 ;
        RECT 3155.320 2031.280 3165.000 2034.480 ;
        RECT -11.080 2030.080 3165.000 2031.280 ;
        RECT -11.080 2026.880 9.480 2030.080 ;
        RECT 120.840 2026.880 3042.640 2030.080 ;
        RECT 3155.320 2026.880 3165.000 2030.080 ;
        RECT -11.080 2025.680 3165.000 2026.880 ;
        RECT -11.080 2022.480 9.480 2025.680 ;
        RECT 120.840 2022.480 3042.640 2025.680 ;
        RECT 3155.320 2022.480 3165.000 2025.680 ;
        RECT -11.080 2021.280 3165.000 2022.480 ;
        RECT -11.080 2019.600 9.480 2021.280 ;
        RECT 0.000 2018.080 9.480 2019.600 ;
        RECT 120.840 2018.080 3042.640 2021.280 ;
        RECT 3155.320 2018.080 3165.000 2021.280 ;
        RECT 0.000 2018.000 3165.000 2018.080 ;
        RECT -16.080 2016.880 3165.000 2018.000 ;
        RECT -16.080 2013.680 9.480 2016.880 ;
        RECT 115.740 2013.680 3042.640 2016.880 ;
        RECT 3155.320 2013.680 3165.000 2016.880 ;
        RECT -16.080 2012.480 3165.000 2013.680 ;
        RECT -16.080 2009.280 9.480 2012.480 ;
        RECT 120.840 2009.280 3042.640 2012.480 ;
        RECT 3155.320 2009.280 3165.000 2012.480 ;
        RECT -16.080 1994.055 3165.000 2009.280 ;
        RECT 0.000 1943.280 3165.000 1994.055 ;
        RECT 0.000 1940.080 9.480 1943.280 ;
        RECT 120.840 1940.080 3042.640 1943.280 ;
        RECT 3155.320 1942.045 3165.000 1943.280 ;
        RECT 3155.320 1940.080 3178.020 1942.045 ;
        RECT 0.000 1938.880 3178.020 1940.080 ;
        RECT 0.000 1935.680 9.480 1938.880 ;
        RECT 120.840 1935.680 3042.640 1938.880 ;
        RECT 3155.320 1935.680 3178.020 1938.880 ;
        RECT 0.000 1934.480 3178.020 1935.680 ;
        RECT 0.000 1931.280 9.480 1934.480 ;
        RECT 120.840 1931.280 3042.640 1934.480 ;
        RECT 3155.320 1931.280 3178.020 1934.480 ;
        RECT 0.000 1930.080 3178.020 1931.280 ;
        RECT 0.000 1926.880 9.480 1930.080 ;
        RECT 120.840 1926.880 3042.640 1930.080 ;
        RECT 3155.320 1926.880 3178.020 1930.080 ;
        RECT 0.000 1925.680 3178.020 1926.880 ;
        RECT 0.000 1922.480 9.480 1925.680 ;
        RECT 120.840 1922.480 3042.640 1925.680 ;
        RECT 3155.320 1922.480 3178.020 1925.680 ;
        RECT 0.000 1921.280 3178.020 1922.480 ;
        RECT 0.000 1918.080 9.480 1921.280 ;
        RECT 120.840 1918.080 3042.640 1921.280 ;
        RECT 3155.320 1918.100 3178.020 1921.280 ;
        RECT 3155.320 1918.080 3165.000 1918.100 ;
        RECT 0.000 1916.880 3165.000 1918.080 ;
        RECT 0.000 1913.680 9.480 1916.880 ;
        RECT 120.840 1913.680 3042.640 1916.880 ;
        RECT 3155.320 1913.680 3165.000 1916.880 ;
        RECT 0.000 1912.480 3165.000 1913.680 ;
        RECT 0.000 1909.280 9.480 1912.480 ;
        RECT 120.840 1909.280 3042.640 1912.480 ;
        RECT 3155.320 1909.280 3165.000 1912.480 ;
        RECT 0.000 1892.130 3165.000 1909.280 ;
        RECT 0.000 1868.185 3178.020 1892.130 ;
        RECT 0.000 1853.425 3165.000 1868.185 ;
        RECT 4.400 1852.025 3165.000 1853.425 ;
        RECT 0.000 1847.445 3165.000 1852.025 ;
        RECT 4.400 1846.045 3165.000 1847.445 ;
        RECT 0.000 1844.225 3165.000 1846.045 ;
        RECT 4.400 1843.280 3165.000 1844.225 ;
        RECT 4.400 1842.825 9.480 1843.280 ;
        RECT 0.000 1841.005 9.480 1842.825 ;
        RECT 4.400 1840.080 9.480 1841.005 ;
        RECT 120.840 1840.080 3042.640 1843.280 ;
        RECT 3155.320 1840.080 3165.000 1843.280 ;
        RECT 4.400 1839.605 3165.000 1840.080 ;
        RECT 0.000 1838.880 3165.000 1839.605 ;
        RECT 0.000 1835.680 9.480 1838.880 ;
        RECT 120.840 1835.680 3047.740 1838.880 ;
        RECT 3155.320 1835.680 3165.000 1838.880 ;
        RECT 0.000 1835.025 3165.000 1835.680 ;
        RECT 4.400 1834.480 3165.000 1835.025 ;
        RECT 4.400 1833.625 9.480 1834.480 ;
        RECT 0.000 1831.280 9.480 1833.625 ;
        RECT 120.840 1831.280 3042.640 1834.480 ;
        RECT 3155.320 1831.280 3165.000 1834.480 ;
        RECT 0.000 1830.080 3165.000 1831.280 ;
        RECT 0.000 1829.045 9.480 1830.080 ;
        RECT 4.400 1827.645 9.480 1829.045 ;
        RECT 0.000 1826.880 9.480 1827.645 ;
        RECT 120.840 1826.880 3042.640 1830.080 ;
        RECT 3155.320 1826.880 3165.000 1830.080 ;
        RECT 0.000 1825.825 3165.000 1826.880 ;
        RECT 4.400 1825.680 3165.000 1825.825 ;
        RECT 4.400 1824.425 9.480 1825.680 ;
        RECT 0.000 1822.605 9.480 1824.425 ;
        RECT 4.400 1822.480 9.480 1822.605 ;
        RECT 120.840 1822.480 3042.640 1825.680 ;
        RECT 3155.320 1822.480 3165.000 1825.680 ;
        RECT 4.400 1821.280 3165.000 1822.480 ;
        RECT 4.400 1821.205 9.480 1821.280 ;
        RECT 0.000 1819.845 9.480 1821.205 ;
        RECT 4.400 1818.445 9.480 1819.845 ;
        RECT 0.000 1818.080 9.480 1818.445 ;
        RECT 115.740 1818.080 3042.640 1821.280 ;
        RECT 3155.320 1818.080 3165.000 1821.280 ;
        RECT 0.000 1816.880 3165.000 1818.080 ;
        RECT 0.000 1813.680 9.480 1816.880 ;
        RECT 120.840 1813.680 3042.640 1816.880 ;
        RECT 3155.320 1813.680 3165.000 1816.880 ;
        RECT 0.000 1812.480 3165.000 1813.680 ;
        RECT 0.000 1809.280 9.480 1812.480 ;
        RECT 120.840 1809.280 3042.640 1812.480 ;
        RECT 3155.320 1809.280 3165.000 1812.480 ;
        RECT 0.000 1807.425 3165.000 1809.280 ;
        RECT 4.400 1806.025 3165.000 1807.425 ;
        RECT 0.000 1804.205 3165.000 1806.025 ;
        RECT 4.400 1802.805 3165.000 1804.205 ;
        RECT 0.000 1800.985 3165.000 1802.805 ;
        RECT 4.400 1799.585 3165.000 1800.985 ;
        RECT 0.000 1798.225 3165.000 1799.585 ;
        RECT 4.400 1796.825 3165.000 1798.225 ;
        RECT 0.000 1789.025 3165.000 1796.825 ;
        RECT 4.400 1787.625 3165.000 1789.025 ;
        RECT 0.000 1785.805 3165.000 1787.625 ;
        RECT 4.400 1784.405 3165.000 1785.805 ;
        RECT 0.000 1782.585 3165.000 1784.405 ;
        RECT 4.400 1781.185 3165.000 1782.585 ;
        RECT 0.000 1743.280 3165.000 1781.185 ;
        RECT 0.000 1740.080 9.480 1743.280 ;
        RECT 120.840 1740.080 3042.640 1743.280 ;
        RECT 3155.320 1740.080 3165.000 1743.280 ;
        RECT 0.000 1738.880 3165.000 1740.080 ;
        RECT 0.000 1735.680 9.480 1738.880 ;
        RECT 120.840 1735.680 3042.640 1738.880 ;
        RECT 3155.320 1735.680 3165.000 1738.880 ;
        RECT 0.000 1734.480 3165.000 1735.680 ;
        RECT 0.000 1731.280 9.480 1734.480 ;
        RECT 120.840 1731.280 3042.640 1734.480 ;
        RECT 3155.320 1731.280 3165.000 1734.480 ;
        RECT 0.000 1730.080 3165.000 1731.280 ;
        RECT 0.000 1726.880 9.480 1730.080 ;
        RECT 120.840 1726.880 3042.640 1730.080 ;
        RECT 3155.320 1726.880 3165.000 1730.080 ;
        RECT 0.000 1725.680 3165.000 1726.880 ;
        RECT 0.000 1722.480 9.480 1725.680 ;
        RECT 120.840 1722.480 3042.640 1725.680 ;
        RECT 3155.320 1722.480 3165.000 1725.680 ;
        RECT 0.000 1721.280 3165.000 1722.480 ;
        RECT 0.000 1718.080 9.480 1721.280 ;
        RECT 120.840 1718.080 3042.640 1721.280 ;
        RECT 3155.320 1718.815 3165.000 1721.280 ;
        RECT 3155.320 1718.080 3160.600 1718.815 ;
        RECT 0.000 1717.415 3160.600 1718.080 ;
        RECT 0.000 1716.880 3165.000 1717.415 ;
        RECT 0.000 1713.680 9.480 1716.880 ;
        RECT 120.840 1713.680 3042.640 1716.880 ;
        RECT 3155.320 1715.595 3165.000 1716.880 ;
        RECT 3155.320 1714.195 3160.600 1715.595 ;
        RECT 3155.320 1713.680 3165.000 1714.195 ;
        RECT 0.000 1712.480 3165.000 1713.680 ;
        RECT 0.000 1709.280 9.480 1712.480 ;
        RECT 120.840 1709.280 3042.640 1712.480 ;
        RECT 3155.320 1712.375 3165.000 1712.480 ;
        RECT 3155.320 1710.975 3160.600 1712.375 ;
        RECT 3155.320 1709.280 3165.000 1710.975 ;
        RECT 0.000 1703.175 3165.000 1709.280 ;
        RECT 0.000 1701.775 3160.600 1703.175 ;
        RECT 0.000 1700.415 3165.000 1701.775 ;
        RECT 0.000 1699.015 3160.600 1700.415 ;
        RECT 0.000 1697.195 3165.000 1699.015 ;
        RECT 0.000 1695.795 3160.600 1697.195 ;
        RECT 0.000 1693.975 3165.000 1695.795 ;
        RECT 0.000 1692.575 3160.600 1693.975 ;
        RECT 0.000 1681.555 3165.000 1692.575 ;
        RECT 0.000 1680.155 3160.600 1681.555 ;
        RECT 0.000 1678.795 3165.000 1680.155 ;
        RECT 0.000 1677.395 3160.600 1678.795 ;
        RECT 0.000 1675.575 3165.000 1677.395 ;
        RECT 0.000 1674.175 3160.600 1675.575 ;
        RECT 0.000 1672.355 3165.000 1674.175 ;
        RECT 0.000 1670.955 3160.600 1672.355 ;
        RECT 0.000 1666.375 3165.000 1670.955 ;
        RECT 0.000 1664.975 3160.600 1666.375 ;
        RECT 0.000 1657.175 3165.000 1664.975 ;
        RECT 0.000 1655.775 3160.600 1657.175 ;
        RECT 0.000 1653.955 3165.000 1655.775 ;
        RECT 0.000 1652.555 3160.600 1653.955 ;
        RECT 0.000 1647.975 3165.000 1652.555 ;
        RECT 0.000 1646.575 3160.600 1647.975 ;
        RECT 0.000 1643.280 3165.000 1646.575 ;
        RECT 0.000 1640.080 9.480 1643.280 ;
        RECT 120.840 1640.080 3042.640 1643.280 ;
        RECT 3155.320 1640.080 3165.000 1643.280 ;
        RECT 0.000 1638.880 3165.000 1640.080 ;
        RECT 0.000 1637.425 9.480 1638.880 ;
        RECT 4.400 1636.025 9.480 1637.425 ;
        RECT 0.000 1635.680 9.480 1636.025 ;
        RECT 120.840 1635.680 3047.740 1638.880 ;
        RECT 3155.320 1635.680 3165.000 1638.880 ;
        RECT 0.000 1634.480 3165.000 1635.680 ;
        RECT 0.000 1631.445 9.480 1634.480 ;
        RECT 4.400 1631.280 9.480 1631.445 ;
        RECT 120.840 1631.280 3042.640 1634.480 ;
        RECT 3155.320 1631.280 3165.000 1634.480 ;
        RECT 4.400 1630.080 3165.000 1631.280 ;
        RECT 4.400 1630.045 9.480 1630.080 ;
        RECT 0.000 1628.225 9.480 1630.045 ;
        RECT 4.400 1626.880 9.480 1628.225 ;
        RECT 120.840 1626.880 3042.640 1630.080 ;
        RECT 3155.320 1626.880 3165.000 1630.080 ;
        RECT 4.400 1626.825 3165.000 1626.880 ;
        RECT 0.000 1625.680 3165.000 1626.825 ;
        RECT 0.000 1625.005 9.480 1625.680 ;
        RECT 4.400 1623.605 9.480 1625.005 ;
        RECT 0.000 1622.480 9.480 1623.605 ;
        RECT 115.740 1622.480 3042.640 1625.680 ;
        RECT 3155.320 1622.480 3165.000 1625.680 ;
        RECT 0.000 1621.280 3165.000 1622.480 ;
        RECT 0.000 1619.025 9.480 1621.280 ;
        RECT 4.400 1618.080 9.480 1619.025 ;
        RECT 120.840 1618.080 3042.640 1621.280 ;
        RECT 3155.320 1618.080 3165.000 1621.280 ;
        RECT 4.400 1617.625 3165.000 1618.080 ;
        RECT 0.000 1616.880 3165.000 1617.625 ;
        RECT 0.000 1613.680 9.480 1616.880 ;
        RECT 120.840 1613.680 3042.640 1616.880 ;
        RECT 3155.320 1613.680 3165.000 1616.880 ;
        RECT 0.000 1613.045 3165.000 1613.680 ;
        RECT 4.400 1612.480 3165.000 1613.045 ;
        RECT 4.400 1611.645 9.480 1612.480 ;
        RECT 0.000 1609.825 9.480 1611.645 ;
        RECT 4.400 1609.280 9.480 1609.825 ;
        RECT 120.840 1609.280 3042.640 1612.480 ;
        RECT 3155.320 1609.280 3165.000 1612.480 ;
        RECT 4.400 1608.425 3165.000 1609.280 ;
        RECT 0.000 1606.605 3165.000 1608.425 ;
        RECT 4.400 1605.205 3165.000 1606.605 ;
        RECT 0.000 1603.845 3165.000 1605.205 ;
        RECT 4.400 1602.445 3165.000 1603.845 ;
        RECT 0.000 1591.425 3165.000 1602.445 ;
        RECT 4.400 1590.025 3165.000 1591.425 ;
        RECT 0.000 1588.205 3165.000 1590.025 ;
        RECT 4.400 1586.805 3165.000 1588.205 ;
        RECT 0.000 1584.985 3165.000 1586.805 ;
        RECT 4.400 1583.585 3165.000 1584.985 ;
        RECT 0.000 1582.225 3165.000 1583.585 ;
        RECT 4.400 1580.825 3165.000 1582.225 ;
        RECT 0.000 1573.025 3165.000 1580.825 ;
        RECT 4.400 1571.625 3165.000 1573.025 ;
        RECT 0.000 1569.805 3165.000 1571.625 ;
        RECT 4.400 1568.405 3165.000 1569.805 ;
        RECT 0.000 1566.585 3165.000 1568.405 ;
        RECT 4.400 1565.185 3165.000 1566.585 ;
        RECT 0.000 1543.280 3165.000 1565.185 ;
        RECT 0.000 1540.080 9.480 1543.280 ;
        RECT 120.840 1540.080 3042.640 1543.280 ;
        RECT 3155.320 1540.080 3165.000 1543.280 ;
        RECT 0.000 1538.880 3165.000 1540.080 ;
        RECT 0.000 1535.680 9.480 1538.880 ;
        RECT 120.840 1535.680 3042.640 1538.880 ;
        RECT 3155.320 1535.680 3165.000 1538.880 ;
        RECT 0.000 1534.480 3165.000 1535.680 ;
        RECT 0.000 1531.280 9.480 1534.480 ;
        RECT 120.840 1531.280 3042.640 1534.480 ;
        RECT 3155.320 1531.280 3165.000 1534.480 ;
        RECT 0.000 1530.080 3165.000 1531.280 ;
        RECT 0.000 1526.880 9.480 1530.080 ;
        RECT 120.840 1526.880 3042.640 1530.080 ;
        RECT 3155.320 1526.880 3165.000 1530.080 ;
        RECT 0.000 1525.680 3165.000 1526.880 ;
        RECT 0.000 1522.480 9.480 1525.680 ;
        RECT 120.840 1522.480 3042.640 1525.680 ;
        RECT 3155.320 1522.480 3165.000 1525.680 ;
        RECT 0.000 1521.280 3165.000 1522.480 ;
        RECT 0.000 1518.080 9.480 1521.280 ;
        RECT 120.840 1518.080 3042.640 1521.280 ;
        RECT 3155.320 1518.080 3165.000 1521.280 ;
        RECT 0.000 1516.880 3165.000 1518.080 ;
        RECT 0.000 1513.680 9.480 1516.880 ;
        RECT 120.840 1513.680 3042.640 1516.880 ;
        RECT 3155.320 1513.680 3165.000 1516.880 ;
        RECT 0.000 1512.480 3165.000 1513.680 ;
        RECT 0.000 1509.280 9.480 1512.480 ;
        RECT 120.840 1509.280 3042.640 1512.480 ;
        RECT 3155.320 1509.280 3165.000 1512.480 ;
        RECT 0.000 1492.815 3165.000 1509.280 ;
        RECT 0.000 1491.415 3160.600 1492.815 ;
        RECT 0.000 1489.595 3165.000 1491.415 ;
        RECT 0.000 1488.195 3160.600 1489.595 ;
        RECT 0.000 1486.375 3165.000 1488.195 ;
        RECT 0.000 1484.975 3160.600 1486.375 ;
        RECT 0.000 1477.175 3165.000 1484.975 ;
        RECT 0.000 1475.775 3160.600 1477.175 ;
        RECT 0.000 1474.415 3165.000 1475.775 ;
        RECT 0.000 1473.015 3160.600 1474.415 ;
        RECT 0.000 1471.195 3165.000 1473.015 ;
        RECT 0.000 1469.795 3160.600 1471.195 ;
        RECT 0.000 1467.975 3165.000 1469.795 ;
        RECT 0.000 1466.575 3160.600 1467.975 ;
        RECT 0.000 1455.555 3165.000 1466.575 ;
        RECT 0.000 1454.155 3160.600 1455.555 ;
        RECT 0.000 1452.795 3165.000 1454.155 ;
        RECT 0.000 1451.395 3160.600 1452.795 ;
        RECT 0.000 1449.575 3165.000 1451.395 ;
        RECT 0.000 1448.175 3160.600 1449.575 ;
        RECT 0.000 1446.355 3165.000 1448.175 ;
        RECT 0.000 1444.955 3160.600 1446.355 ;
        RECT 0.000 1443.280 3165.000 1444.955 ;
        RECT 0.000 1440.080 9.480 1443.280 ;
        RECT 120.840 1440.080 3042.640 1443.280 ;
        RECT 3155.320 1440.375 3165.000 1443.280 ;
        RECT 3155.320 1440.080 3160.600 1440.375 ;
        RECT 0.000 1438.975 3160.600 1440.080 ;
        RECT 0.000 1438.880 3165.000 1438.975 ;
        RECT 0.000 1435.680 9.480 1438.880 ;
        RECT 120.840 1435.680 3047.740 1438.880 ;
        RECT 3155.320 1435.680 3165.000 1438.880 ;
        RECT 0.000 1434.480 3165.000 1435.680 ;
        RECT 0.000 1431.280 9.480 1434.480 ;
        RECT 120.840 1431.280 3042.640 1434.480 ;
        RECT 3155.320 1431.280 3165.000 1434.480 ;
        RECT 0.000 1431.175 3165.000 1431.280 ;
        RECT 0.000 1430.080 3160.600 1431.175 ;
        RECT 0.000 1426.880 9.480 1430.080 ;
        RECT 115.740 1426.880 3042.640 1430.080 ;
        RECT 3155.320 1429.775 3160.600 1430.080 ;
        RECT 3155.320 1427.955 3165.000 1429.775 ;
        RECT 3155.320 1426.880 3160.600 1427.955 ;
        RECT 0.000 1426.555 3160.600 1426.880 ;
        RECT 0.000 1425.680 3165.000 1426.555 ;
        RECT 0.000 1422.480 9.480 1425.680 ;
        RECT 120.840 1422.480 3042.640 1425.680 ;
        RECT 3155.320 1422.480 3165.000 1425.680 ;
        RECT 0.000 1421.975 3165.000 1422.480 ;
        RECT 0.000 1421.425 3160.600 1421.975 ;
        RECT 4.400 1421.280 3160.600 1421.425 ;
        RECT 4.400 1420.025 9.480 1421.280 ;
        RECT 0.000 1418.080 9.480 1420.025 ;
        RECT 120.840 1418.080 3042.640 1421.280 ;
        RECT 3155.320 1420.575 3160.600 1421.280 ;
        RECT 3155.320 1418.080 3165.000 1420.575 ;
        RECT 0.000 1416.880 3165.000 1418.080 ;
        RECT 0.000 1415.445 9.480 1416.880 ;
        RECT 4.400 1414.045 9.480 1415.445 ;
        RECT 0.000 1413.680 9.480 1414.045 ;
        RECT 120.840 1413.680 3042.640 1416.880 ;
        RECT 3155.320 1413.680 3165.000 1416.880 ;
        RECT 0.000 1412.480 3165.000 1413.680 ;
        RECT 0.000 1412.225 9.480 1412.480 ;
        RECT 4.400 1410.825 9.480 1412.225 ;
        RECT 0.000 1409.280 9.480 1410.825 ;
        RECT 120.840 1409.280 3042.640 1412.480 ;
        RECT 3155.320 1409.280 3165.000 1412.480 ;
        RECT 0.000 1409.005 3165.000 1409.280 ;
        RECT 4.400 1407.605 3165.000 1409.005 ;
        RECT 0.000 1403.025 3165.000 1407.605 ;
        RECT 4.400 1401.625 3165.000 1403.025 ;
        RECT 0.000 1397.045 3165.000 1401.625 ;
        RECT 4.400 1395.645 3165.000 1397.045 ;
        RECT 0.000 1393.825 3165.000 1395.645 ;
        RECT 4.400 1392.425 3165.000 1393.825 ;
        RECT 0.000 1390.605 3165.000 1392.425 ;
        RECT 4.400 1389.205 3165.000 1390.605 ;
        RECT 0.000 1387.845 3165.000 1389.205 ;
        RECT 4.400 1386.445 3165.000 1387.845 ;
        RECT 0.000 1375.425 3165.000 1386.445 ;
        RECT 4.400 1374.025 3165.000 1375.425 ;
        RECT 0.000 1372.205 3165.000 1374.025 ;
        RECT 4.400 1370.805 3165.000 1372.205 ;
        RECT 0.000 1368.985 3165.000 1370.805 ;
        RECT 4.400 1367.585 3165.000 1368.985 ;
        RECT 0.000 1366.225 3165.000 1367.585 ;
        RECT 4.400 1364.825 3165.000 1366.225 ;
        RECT 0.000 1357.025 3165.000 1364.825 ;
        RECT 4.400 1355.625 3165.000 1357.025 ;
        RECT 0.000 1353.805 3165.000 1355.625 ;
        RECT 4.400 1352.405 3165.000 1353.805 ;
        RECT 0.000 1350.585 3165.000 1352.405 ;
        RECT 4.400 1349.185 3165.000 1350.585 ;
        RECT 0.000 1343.280 3165.000 1349.185 ;
        RECT 0.000 1340.080 9.480 1343.280 ;
        RECT 120.840 1340.080 3042.640 1343.280 ;
        RECT 3155.320 1340.080 3165.000 1343.280 ;
        RECT 0.000 1338.880 3165.000 1340.080 ;
        RECT 0.000 1335.680 9.480 1338.880 ;
        RECT 120.840 1335.680 3042.640 1338.880 ;
        RECT 3155.320 1335.680 3165.000 1338.880 ;
        RECT 0.000 1334.480 3165.000 1335.680 ;
        RECT 0.000 1331.280 9.480 1334.480 ;
        RECT 120.840 1331.280 3042.640 1334.480 ;
        RECT 3155.320 1331.280 3165.000 1334.480 ;
        RECT 0.000 1330.080 3165.000 1331.280 ;
        RECT 0.000 1326.880 9.480 1330.080 ;
        RECT 120.840 1326.880 3042.640 1330.080 ;
        RECT 3155.320 1326.880 3165.000 1330.080 ;
        RECT 0.000 1325.680 3165.000 1326.880 ;
        RECT 0.000 1322.480 9.480 1325.680 ;
        RECT 120.840 1322.480 3042.640 1325.680 ;
        RECT 3155.320 1322.480 3165.000 1325.680 ;
        RECT 0.000 1321.280 3165.000 1322.480 ;
        RECT 0.000 1318.080 9.480 1321.280 ;
        RECT 120.840 1318.080 3042.640 1321.280 ;
        RECT 3155.320 1318.080 3165.000 1321.280 ;
        RECT 0.000 1316.880 3165.000 1318.080 ;
        RECT 0.000 1313.680 9.480 1316.880 ;
        RECT 120.840 1313.680 3042.640 1316.880 ;
        RECT 3155.320 1313.680 3165.000 1316.880 ;
        RECT 0.000 1312.480 3165.000 1313.680 ;
        RECT 0.000 1309.280 9.480 1312.480 ;
        RECT 120.840 1309.280 3042.640 1312.480 ;
        RECT 3155.320 1309.280 3165.000 1312.480 ;
        RECT 0.000 1267.815 3165.000 1309.280 ;
        RECT 0.000 1266.415 3160.600 1267.815 ;
        RECT 0.000 1264.595 3165.000 1266.415 ;
        RECT 0.000 1263.195 3160.600 1264.595 ;
        RECT 0.000 1261.375 3165.000 1263.195 ;
        RECT 0.000 1259.975 3160.600 1261.375 ;
        RECT 0.000 1252.175 3165.000 1259.975 ;
        RECT 0.000 1250.775 3160.600 1252.175 ;
        RECT 0.000 1249.415 3165.000 1250.775 ;
        RECT 0.000 1248.015 3160.600 1249.415 ;
        RECT 0.000 1246.195 3165.000 1248.015 ;
        RECT 0.000 1244.795 3160.600 1246.195 ;
        RECT 0.000 1243.280 3165.000 1244.795 ;
        RECT 0.000 1240.080 9.480 1243.280 ;
        RECT 120.840 1240.080 3042.640 1243.280 ;
        RECT 3155.320 1242.975 3165.000 1243.280 ;
        RECT 3155.320 1241.575 3160.600 1242.975 ;
        RECT 3155.320 1240.080 3165.000 1241.575 ;
        RECT 0.000 1238.880 3165.000 1240.080 ;
        RECT 0.000 1235.680 9.480 1238.880 ;
        RECT 120.840 1235.680 3047.740 1238.880 ;
        RECT 3155.320 1235.680 3165.000 1238.880 ;
        RECT 0.000 1234.480 3165.000 1235.680 ;
        RECT 0.000 1231.280 9.480 1234.480 ;
        RECT 115.740 1231.280 3042.640 1234.480 ;
        RECT 3155.320 1231.280 3165.000 1234.480 ;
        RECT 0.000 1230.555 3165.000 1231.280 ;
        RECT 0.000 1230.080 3160.600 1230.555 ;
        RECT 0.000 1226.880 9.480 1230.080 ;
        RECT 120.840 1226.880 3042.640 1230.080 ;
        RECT 3155.320 1229.155 3160.600 1230.080 ;
        RECT 3155.320 1227.795 3165.000 1229.155 ;
        RECT 3155.320 1226.880 3160.600 1227.795 ;
        RECT 0.000 1226.395 3160.600 1226.880 ;
        RECT 0.000 1225.680 3165.000 1226.395 ;
        RECT 0.000 1222.480 9.480 1225.680 ;
        RECT 120.840 1222.480 3042.640 1225.680 ;
        RECT 3155.320 1224.575 3165.000 1225.680 ;
        RECT 3155.320 1223.175 3160.600 1224.575 ;
        RECT 3155.320 1222.480 3165.000 1223.175 ;
        RECT 0.000 1221.355 3165.000 1222.480 ;
        RECT 0.000 1221.280 3160.600 1221.355 ;
        RECT 0.000 1218.080 9.480 1221.280 ;
        RECT 120.840 1218.080 3042.640 1221.280 ;
        RECT 3155.320 1219.955 3160.600 1221.280 ;
        RECT 3155.320 1218.080 3165.000 1219.955 ;
        RECT 0.000 1216.880 3165.000 1218.080 ;
        RECT 0.000 1213.680 9.480 1216.880 ;
        RECT 120.840 1213.680 3042.640 1216.880 ;
        RECT 3155.320 1215.375 3165.000 1216.880 ;
        RECT 3155.320 1213.975 3160.600 1215.375 ;
        RECT 3155.320 1213.680 3165.000 1213.975 ;
        RECT 0.000 1212.480 3165.000 1213.680 ;
        RECT 0.000 1209.280 9.480 1212.480 ;
        RECT 120.840 1209.280 3042.640 1212.480 ;
        RECT 3155.320 1209.280 3165.000 1212.480 ;
        RECT 0.000 1206.175 3165.000 1209.280 ;
        RECT 0.000 1205.425 3160.600 1206.175 ;
        RECT 4.400 1204.775 3160.600 1205.425 ;
        RECT 4.400 1204.025 3165.000 1204.775 ;
        RECT 0.000 1202.955 3165.000 1204.025 ;
        RECT 0.000 1201.555 3160.600 1202.955 ;
        RECT 0.000 1199.445 3165.000 1201.555 ;
        RECT 4.400 1198.045 3165.000 1199.445 ;
        RECT 0.000 1196.975 3165.000 1198.045 ;
        RECT 0.000 1196.225 3160.600 1196.975 ;
        RECT 4.400 1195.575 3160.600 1196.225 ;
        RECT 4.400 1194.825 3165.000 1195.575 ;
        RECT 0.000 1193.005 3165.000 1194.825 ;
        RECT 4.400 1191.605 3165.000 1193.005 ;
        RECT 0.000 1187.025 3165.000 1191.605 ;
        RECT 4.400 1185.625 3165.000 1187.025 ;
        RECT 0.000 1181.045 3165.000 1185.625 ;
        RECT 4.400 1179.645 3165.000 1181.045 ;
        RECT 0.000 1177.825 3165.000 1179.645 ;
        RECT 4.400 1176.425 3165.000 1177.825 ;
        RECT 0.000 1174.605 3165.000 1176.425 ;
        RECT 4.400 1173.205 3165.000 1174.605 ;
        RECT 0.000 1171.845 3165.000 1173.205 ;
        RECT 4.400 1170.445 3165.000 1171.845 ;
        RECT 0.000 1159.425 3165.000 1170.445 ;
        RECT 4.400 1158.025 3165.000 1159.425 ;
        RECT 0.000 1156.205 3165.000 1158.025 ;
        RECT 4.400 1154.805 3165.000 1156.205 ;
        RECT 0.000 1152.985 3165.000 1154.805 ;
        RECT 4.400 1151.585 3165.000 1152.985 ;
        RECT 0.000 1150.225 3165.000 1151.585 ;
        RECT 4.400 1148.825 3165.000 1150.225 ;
        RECT 0.000 1141.025 3165.000 1148.825 ;
        RECT 4.400 1139.625 3165.000 1141.025 ;
        RECT 0.000 1137.805 3165.000 1139.625 ;
        RECT 4.400 1136.405 3165.000 1137.805 ;
        RECT 0.000 1134.585 3165.000 1136.405 ;
        RECT 4.400 1133.185 3165.000 1134.585 ;
        RECT 0.000 1042.815 3165.000 1133.185 ;
        RECT 0.000 1041.415 3160.600 1042.815 ;
        RECT 0.000 1039.595 3165.000 1041.415 ;
        RECT 0.000 1038.195 3160.600 1039.595 ;
        RECT 0.000 1036.375 3165.000 1038.195 ;
        RECT 0.000 1034.975 3160.600 1036.375 ;
        RECT 0.000 1027.175 3165.000 1034.975 ;
        RECT 0.000 1025.775 3160.600 1027.175 ;
        RECT 0.000 1024.415 3165.000 1025.775 ;
        RECT 0.000 1023.015 3160.600 1024.415 ;
        RECT 0.000 1021.195 3165.000 1023.015 ;
        RECT 0.000 1019.795 3160.600 1021.195 ;
        RECT 0.000 1017.975 3165.000 1019.795 ;
        RECT 0.000 1016.575 3160.600 1017.975 ;
        RECT 0.000 1005.555 3165.000 1016.575 ;
        RECT 0.000 1004.155 3160.600 1005.555 ;
        RECT 0.000 1002.795 3165.000 1004.155 ;
        RECT 0.000 1001.395 3160.600 1002.795 ;
        RECT 0.000 999.575 3165.000 1001.395 ;
        RECT 0.000 998.175 3160.600 999.575 ;
        RECT 0.000 996.355 3165.000 998.175 ;
        RECT 0.000 994.955 3160.600 996.355 ;
        RECT 0.000 990.375 3165.000 994.955 ;
        RECT 0.000 989.425 3160.600 990.375 ;
        RECT 4.400 988.975 3160.600 989.425 ;
        RECT 4.400 988.025 3165.000 988.975 ;
        RECT 0.000 983.445 3165.000 988.025 ;
        RECT 4.400 982.045 3165.000 983.445 ;
        RECT 0.000 981.175 3165.000 982.045 ;
        RECT 0.000 980.225 3160.600 981.175 ;
        RECT 4.400 979.775 3160.600 980.225 ;
        RECT 4.400 978.825 3165.000 979.775 ;
        RECT 0.000 977.955 3165.000 978.825 ;
        RECT 0.000 976.555 3160.600 977.955 ;
        RECT 0.000 971.975 3165.000 976.555 ;
        RECT 0.000 971.025 3160.600 971.975 ;
        RECT 4.400 970.575 3160.600 971.025 ;
        RECT 4.400 969.625 3165.000 970.575 ;
        RECT 0.000 965.045 3165.000 969.625 ;
        RECT 4.400 963.645 3165.000 965.045 ;
        RECT 0.000 961.825 3165.000 963.645 ;
        RECT 4.400 960.425 3165.000 961.825 ;
        RECT 0.000 958.605 3165.000 960.425 ;
        RECT 4.400 957.205 3165.000 958.605 ;
        RECT 0.000 955.845 3165.000 957.205 ;
        RECT 4.400 954.445 3165.000 955.845 ;
        RECT 0.000 943.425 3165.000 954.445 ;
        RECT 4.400 942.025 3165.000 943.425 ;
        RECT 0.000 940.205 3165.000 942.025 ;
        RECT 4.400 938.805 3165.000 940.205 ;
        RECT 0.000 936.985 3165.000 938.805 ;
        RECT 4.400 935.585 3165.000 936.985 ;
        RECT 0.000 934.225 3165.000 935.585 ;
        RECT 4.400 932.825 3165.000 934.225 ;
        RECT 0.000 925.025 3165.000 932.825 ;
        RECT 4.400 923.625 3165.000 925.025 ;
        RECT 0.000 921.805 3165.000 923.625 ;
        RECT 4.400 920.405 3165.000 921.805 ;
        RECT 0.000 918.585 3165.000 920.405 ;
        RECT 4.400 917.185 3165.000 918.585 ;
        RECT 0.000 816.815 3165.000 917.185 ;
        RECT 0.000 815.415 3160.600 816.815 ;
        RECT 0.000 813.595 3165.000 815.415 ;
        RECT 0.000 812.195 3160.600 813.595 ;
        RECT 0.000 810.375 3165.000 812.195 ;
        RECT 0.000 808.975 3160.600 810.375 ;
        RECT 0.000 801.175 3165.000 808.975 ;
        RECT 0.000 799.775 3160.600 801.175 ;
        RECT 0.000 798.415 3165.000 799.775 ;
        RECT 0.000 797.015 3160.600 798.415 ;
        RECT 0.000 795.195 3165.000 797.015 ;
        RECT 0.000 793.795 3160.600 795.195 ;
        RECT 0.000 791.975 3165.000 793.795 ;
        RECT 0.000 790.575 3160.600 791.975 ;
        RECT 0.000 779.555 3165.000 790.575 ;
        RECT 0.000 778.155 3160.600 779.555 ;
        RECT 0.000 776.795 3165.000 778.155 ;
        RECT 0.000 775.395 3160.600 776.795 ;
        RECT 0.000 773.575 3165.000 775.395 ;
        RECT 0.000 773.425 3160.600 773.575 ;
        RECT 4.400 772.175 3160.600 773.425 ;
        RECT 4.400 772.025 3165.000 772.175 ;
        RECT 0.000 770.355 3165.000 772.025 ;
        RECT 0.000 768.955 3160.600 770.355 ;
        RECT 0.000 767.445 3165.000 768.955 ;
        RECT 4.400 766.045 3165.000 767.445 ;
        RECT 0.000 764.375 3165.000 766.045 ;
        RECT 0.000 764.225 3160.600 764.375 ;
        RECT 4.400 762.975 3160.600 764.225 ;
        RECT 4.400 762.825 3165.000 762.975 ;
        RECT 0.000 755.175 3165.000 762.825 ;
        RECT 0.000 755.025 3160.600 755.175 ;
        RECT 4.400 753.775 3160.600 755.025 ;
        RECT 4.400 753.625 3165.000 753.775 ;
        RECT 0.000 751.955 3165.000 753.625 ;
        RECT 0.000 750.555 3160.600 751.955 ;
        RECT 0.000 749.045 3165.000 750.555 ;
        RECT 4.400 747.645 3165.000 749.045 ;
        RECT 0.000 745.975 3165.000 747.645 ;
        RECT 0.000 745.825 3160.600 745.975 ;
        RECT 4.400 744.575 3160.600 745.825 ;
        RECT 4.400 744.425 3165.000 744.575 ;
        RECT 0.000 742.605 3165.000 744.425 ;
        RECT 4.400 741.205 3165.000 742.605 ;
        RECT 0.000 739.845 3165.000 741.205 ;
        RECT 4.400 738.445 3165.000 739.845 ;
        RECT 0.000 727.425 3165.000 738.445 ;
        RECT 4.400 726.025 3165.000 727.425 ;
        RECT 0.000 724.205 3165.000 726.025 ;
        RECT 4.400 722.805 3165.000 724.205 ;
        RECT 0.000 720.985 3165.000 722.805 ;
        RECT 4.400 719.585 3165.000 720.985 ;
        RECT 0.000 718.225 3165.000 719.585 ;
        RECT 4.400 716.825 3165.000 718.225 ;
        RECT 0.000 709.025 3165.000 716.825 ;
        RECT 4.400 707.625 3165.000 709.025 ;
        RECT 0.000 705.805 3165.000 707.625 ;
        RECT 4.690 704.405 3165.000 705.805 ;
        RECT 0.000 702.585 3165.000 704.405 ;
        RECT 4.400 701.185 3165.000 702.585 ;
        RECT 0.000 591.815 3165.000 701.185 ;
        RECT 0.000 590.415 3160.600 591.815 ;
        RECT 0.000 588.595 3165.000 590.415 ;
        RECT 0.000 587.195 3160.600 588.595 ;
        RECT 0.000 585.375 3165.000 587.195 ;
        RECT 0.000 583.975 3160.600 585.375 ;
        RECT 0.000 576.175 3165.000 583.975 ;
        RECT 0.000 574.775 3160.600 576.175 ;
        RECT 0.000 573.415 3165.000 574.775 ;
        RECT 0.000 572.015 3160.600 573.415 ;
        RECT 0.000 570.195 3165.000 572.015 ;
        RECT 0.000 568.795 3160.600 570.195 ;
        RECT 0.000 566.975 3165.000 568.795 ;
        RECT 0.000 565.575 3160.600 566.975 ;
        RECT 0.000 554.555 3165.000 565.575 ;
        RECT 0.000 553.155 3160.600 554.555 ;
        RECT 0.000 551.795 3165.000 553.155 ;
        RECT 0.000 550.395 3160.600 551.795 ;
        RECT 0.000 548.575 3165.000 550.395 ;
        RECT 0.000 547.175 3160.600 548.575 ;
        RECT 0.000 545.355 3165.000 547.175 ;
        RECT 0.000 543.955 3160.600 545.355 ;
        RECT 0.000 539.375 3165.000 543.955 ;
        RECT 0.000 537.975 3160.600 539.375 ;
        RECT 0.000 530.175 3165.000 537.975 ;
        RECT 0.000 528.775 3160.600 530.175 ;
        RECT 0.000 526.955 3165.000 528.775 ;
        RECT 0.000 525.555 3160.600 526.955 ;
        RECT 0.000 520.975 3165.000 525.555 ;
        RECT 0.000 519.575 3160.600 520.975 ;
        RECT 0.000 365.815 3165.000 519.575 ;
        RECT 0.000 364.415 3160.600 365.815 ;
        RECT 0.000 362.595 3165.000 364.415 ;
        RECT 0.000 361.195 3160.600 362.595 ;
        RECT 0.000 359.375 3165.000 361.195 ;
        RECT 0.000 357.975 3160.600 359.375 ;
        RECT 0.000 350.175 3165.000 357.975 ;
        RECT 0.000 348.775 3160.600 350.175 ;
        RECT 0.000 347.415 3165.000 348.775 ;
        RECT 0.000 346.015 3160.600 347.415 ;
        RECT 0.000 344.195 3165.000 346.015 ;
        RECT 0.000 342.795 3160.600 344.195 ;
        RECT 0.000 340.975 3165.000 342.795 ;
        RECT 0.000 339.575 3160.600 340.975 ;
        RECT 0.000 328.555 3165.000 339.575 ;
        RECT 0.000 327.155 3160.600 328.555 ;
        RECT 0.000 325.795 3165.000 327.155 ;
        RECT 0.000 324.395 3160.600 325.795 ;
        RECT 0.000 322.575 3165.000 324.395 ;
        RECT 0.000 321.175 3160.600 322.575 ;
        RECT 0.000 319.355 3165.000 321.175 ;
        RECT 0.000 317.955 3160.600 319.355 ;
        RECT 0.000 313.375 3165.000 317.955 ;
        RECT 0.000 311.975 3160.600 313.375 ;
        RECT 0.000 304.175 3165.000 311.975 ;
        RECT 0.000 302.775 3160.600 304.175 ;
        RECT 0.000 300.955 3165.000 302.775 ;
        RECT 0.000 299.555 3160.600 300.955 ;
        RECT 0.000 294.975 3165.000 299.555 ;
        RECT 0.000 293.575 3160.600 294.975 ;
        RECT 0.000 204.200 3165.000 293.575 ;
        RECT -16.080 180.255 3165.000 204.200 ;
        RECT 0.000 154.000 3165.000 180.255 ;
        RECT -16.080 130.055 3165.000 154.000 ;
        RECT 0.000 0.000 3165.000 130.055 ;
        RECT 878.500 -31.255 896.510 -0.675 ;
        RECT 994.715 -14.690 1018.745 -0.110 ;
        RECT 1044.970 -14.690 1069.000 -0.110 ;
        RECT 1075.025 -40.985 1088.745 -0.675 ;
      LAYER met4 ;
        RECT 2666.935 4767.000 2690.965 4772.410 ;
        RECT 2716.840 4767.000 2740.870 4772.410 ;
        RECT 0.000 4755.200 3165.000 4767.000 ;
        RECT 0.000 4424.200 10.520 4755.200 ;
        RECT -9.290 4400.255 10.520 4424.200 ;
        RECT 0.000 4398.650 10.520 4400.255 ;
        RECT -9.290 4375.600 10.520 4398.650 ;
        RECT 0.000 4374.000 10.520 4375.600 ;
        RECT -9.290 4350.055 10.520 4374.000 ;
        RECT 0.000 4001.790 10.520 4350.055 ;
        RECT -9.290 3977.845 10.520 4001.790 ;
        RECT 0.000 3951.590 10.520 3977.845 ;
        RECT -9.290 3927.945 10.520 3951.590 ;
        RECT 0.000 2278.790 10.520 3927.945 ;
        RECT -9.290 2254.845 10.520 2278.790 ;
        RECT 0.000 2228.590 10.520 2254.845 ;
        RECT -9.290 2204.945 10.520 2228.590 ;
        RECT 0.000 2068.200 10.520 2204.945 ;
        RECT -9.290 2044.255 10.520 2068.200 ;
        RECT 0.000 2042.650 10.520 2044.255 ;
        RECT -9.290 2019.600 10.520 2042.650 ;
        RECT 0.000 2018.000 10.520 2019.600 ;
        RECT -9.290 1994.055 10.520 2018.000 ;
        RECT 0.000 204.200 10.520 1994.055 ;
        RECT -9.290 180.255 10.520 204.200 ;
        RECT 0.000 154.000 10.520 180.255 ;
        RECT -9.290 130.055 10.520 154.000 ;
        RECT 0.000 10.240 10.520 130.055 ;
        RECT 16.320 10.240 16.520 4755.200 ;
        RECT 22.320 10.240 22.520 4755.200 ;
        RECT 28.320 10.240 28.520 4755.200 ;
        RECT 34.320 10.240 34.520 4755.200 ;
        RECT 40.320 10.240 40.520 4755.200 ;
        RECT 46.320 10.240 46.520 4755.200 ;
        RECT 52.320 10.240 52.520 4755.200 ;
        RECT 58.320 10.240 58.520 4755.200 ;
        RECT 64.320 10.240 64.520 4755.200 ;
        RECT 70.320 10.240 70.520 4755.200 ;
        RECT 73.320 10.240 73.520 4755.200 ;
        RECT 76.320 4630.950 123.520 4755.200 ;
        RECT 130.720 4630.950 131.120 4755.200 ;
        RECT 138.320 4630.950 223.520 4755.200 ;
        RECT 230.720 4630.950 231.120 4755.200 ;
        RECT 238.320 4630.950 255.640 4755.200 ;
        RECT 262.840 4630.950 263.240 4755.200 ;
        RECT 270.440 4630.950 323.520 4755.200 ;
        RECT 330.720 4630.950 331.120 4755.200 ;
        RECT 338.320 4630.950 423.520 4755.200 ;
        RECT 430.720 4630.950 431.120 4755.200 ;
        RECT 438.320 4630.950 523.520 4755.200 ;
        RECT 530.720 4630.950 531.120 4755.200 ;
        RECT 538.320 4630.950 555.640 4755.200 ;
        RECT 562.840 4630.950 563.240 4755.200 ;
        RECT 570.440 4630.950 623.520 4755.200 ;
        RECT 630.720 4630.950 631.120 4755.200 ;
        RECT 638.320 4630.950 723.520 4755.200 ;
        RECT 730.720 4630.950 731.120 4755.200 ;
        RECT 738.320 4630.950 823.520 4755.200 ;
        RECT 830.720 4630.950 831.120 4755.200 ;
        RECT 838.320 4630.950 850.320 4755.200 ;
        RECT 855.920 4630.950 858.320 4755.200 ;
        RECT 863.920 4630.950 900.320 4755.200 ;
        RECT 905.920 4630.950 908.320 4755.200 ;
        RECT 913.920 4630.950 923.520 4755.200 ;
        RECT 930.720 4630.950 931.120 4755.200 ;
        RECT 938.320 4630.950 955.640 4755.200 ;
        RECT 962.840 4630.950 963.240 4755.200 ;
        RECT 970.440 4630.950 1023.520 4755.200 ;
        RECT 1030.720 4630.950 1031.120 4755.200 ;
        RECT 1038.320 4630.950 1123.520 4755.200 ;
        RECT 1130.720 4630.950 1131.120 4755.200 ;
        RECT 1138.320 4630.950 1155.640 4755.200 ;
        RECT 1162.840 4630.950 1163.240 4755.200 ;
        RECT 1170.440 4630.950 1223.520 4755.200 ;
        RECT 1230.720 4630.950 1231.120 4755.200 ;
        RECT 1238.320 4630.950 1275.320 4755.200 ;
        RECT 1280.920 4630.950 1283.320 4755.200 ;
        RECT 1288.920 4630.950 1323.520 4755.200 ;
        RECT 1330.720 4630.950 1331.120 4755.200 ;
        RECT 1338.320 4630.950 1375.320 4755.200 ;
        RECT 1380.920 4630.950 1383.320 4755.200 ;
        RECT 1388.920 4630.950 1423.520 4755.200 ;
        RECT 1430.720 4630.950 1431.120 4755.200 ;
        RECT 1438.320 4630.950 1455.640 4755.200 ;
        RECT 1462.840 4630.950 1463.240 4755.200 ;
        RECT 1470.440 4630.950 1475.320 4755.200 ;
        RECT 1480.920 4630.950 1483.320 4755.200 ;
        RECT 1488.920 4630.950 1523.520 4755.200 ;
        RECT 1530.720 4630.950 1531.120 4755.200 ;
        RECT 1538.320 4630.950 1623.520 4755.200 ;
        RECT 1630.720 4630.950 1631.120 4755.200 ;
        RECT 1638.320 4630.950 1723.520 4755.200 ;
        RECT 1730.720 4630.950 1731.120 4755.200 ;
        RECT 1738.320 4630.950 1755.640 4755.200 ;
        RECT 1762.840 4630.950 1763.240 4755.200 ;
        RECT 1770.440 4630.950 1823.520 4755.200 ;
        RECT 1830.720 4630.950 1831.120 4755.200 ;
        RECT 1838.320 4630.950 1843.320 4755.200 ;
        RECT 1848.920 4630.950 1851.320 4755.200 ;
        RECT 1856.920 4630.950 1859.320 4755.200 ;
        RECT 1864.920 4630.950 1867.320 4755.200 ;
        RECT 1872.920 4630.950 1883.320 4755.200 ;
        RECT 1888.920 4630.950 1891.320 4755.200 ;
        RECT 1896.920 4630.950 1899.320 4755.200 ;
        RECT 1904.920 4630.950 1907.320 4755.200 ;
        RECT 1912.920 4630.950 1923.520 4755.200 ;
        RECT 1930.720 4630.950 1931.120 4755.200 ;
        RECT 1938.320 4630.950 2023.520 4755.200 ;
        RECT 2030.720 4630.950 2031.120 4755.200 ;
        RECT 2038.320 4630.950 2055.640 4755.200 ;
        RECT 2062.840 4630.950 2063.240 4755.200 ;
        RECT 2070.440 4630.950 2123.520 4755.200 ;
        RECT 2130.720 4630.950 2131.120 4755.200 ;
        RECT 2138.320 4630.950 2223.520 4755.200 ;
        RECT 2230.720 4630.950 2231.120 4755.200 ;
        RECT 2238.320 4630.950 2323.520 4755.200 ;
        RECT 2330.720 4630.950 2331.120 4755.200 ;
        RECT 2338.320 4630.950 2355.640 4755.200 ;
        RECT 2362.840 4630.950 2363.240 4755.200 ;
        RECT 2370.440 4630.950 2423.520 4755.200 ;
        RECT 2430.720 4630.950 2431.120 4755.200 ;
        RECT 2438.320 4630.950 2523.520 4755.200 ;
        RECT 2530.720 4630.950 2531.120 4755.200 ;
        RECT 2538.320 4630.950 2623.520 4755.200 ;
        RECT 2630.720 4630.950 2631.120 4755.200 ;
        RECT 2638.320 4630.950 2755.640 4755.200 ;
        RECT 2762.840 4630.950 2763.240 4755.200 ;
        RECT 2770.440 4630.950 2823.520 4755.200 ;
        RECT 2830.720 4630.950 2831.120 4755.200 ;
        RECT 2838.320 4630.950 2923.520 4755.200 ;
        RECT 2930.720 4630.950 2931.120 4755.200 ;
        RECT 2938.320 4630.950 2967.975 4755.200 ;
        RECT 76.320 4630.850 2967.975 4630.950 ;
        RECT 2970.375 4630.850 2990.355 4755.200 ;
        RECT 2992.755 4630.950 3023.520 4755.200 ;
        RECT 3030.720 4630.950 3031.120 4755.200 ;
        RECT 3038.320 4630.950 3086.780 4755.200 ;
        RECT 2992.755 4630.850 3086.780 4630.950 ;
        RECT 76.320 1032.830 3086.780 4630.850 ;
        RECT 76.320 1032.730 2967.975 1032.830 ;
        RECT 76.320 835.105 123.520 1032.730 ;
        RECT 130.720 835.105 131.120 1032.730 ;
        RECT 138.320 835.105 223.520 1032.730 ;
        RECT 230.720 835.105 231.120 1032.730 ;
        RECT 238.320 850.560 255.640 1032.730 ;
        RECT 262.840 850.560 263.240 1032.730 ;
        RECT 270.440 850.560 323.520 1032.730 ;
        RECT 238.320 835.105 323.520 850.560 ;
        RECT 330.720 835.105 331.120 1032.730 ;
        RECT 338.320 835.105 423.520 1032.730 ;
        RECT 430.720 835.105 431.120 1032.730 ;
        RECT 438.320 835.105 523.520 1032.730 ;
        RECT 530.720 835.105 531.120 1032.730 ;
        RECT 538.320 850.560 555.640 1032.730 ;
        RECT 562.840 850.560 563.240 1032.730 ;
        RECT 570.440 850.560 623.520 1032.730 ;
        RECT 538.320 835.105 623.520 850.560 ;
        RECT 630.720 835.105 631.120 1032.730 ;
        RECT 638.320 835.105 723.520 1032.730 ;
        RECT 730.720 835.105 731.120 1032.730 ;
        RECT 738.320 835.105 823.520 1032.730 ;
        RECT 830.720 835.105 831.120 1032.730 ;
        RECT 838.320 850.560 850.320 1032.730 ;
        RECT 855.920 850.560 858.320 1032.730 ;
        RECT 838.320 835.105 858.320 850.560 ;
        RECT 863.920 850.560 900.320 1032.730 ;
        RECT 905.920 850.560 908.320 1032.730 ;
        RECT 863.920 835.105 908.320 850.560 ;
        RECT 913.920 835.105 923.520 1032.730 ;
        RECT 930.720 835.105 931.120 1032.730 ;
        RECT 938.320 850.560 955.640 1032.730 ;
        RECT 962.840 850.560 963.240 1032.730 ;
        RECT 970.440 850.560 1023.520 1032.730 ;
        RECT 938.320 835.105 1023.520 850.560 ;
        RECT 1030.720 835.105 1031.120 1032.730 ;
        RECT 1038.320 835.105 1123.520 1032.730 ;
        RECT 1130.720 835.105 1131.120 1032.730 ;
        RECT 1138.320 850.560 1155.640 1032.730 ;
        RECT 1162.840 850.560 1163.240 1032.730 ;
        RECT 1170.440 850.560 1223.520 1032.730 ;
        RECT 1138.320 835.105 1223.520 850.560 ;
        RECT 1230.720 835.105 1231.120 1032.730 ;
        RECT 1238.320 835.105 1275.320 1032.730 ;
        RECT 1280.920 835.105 1283.320 1032.730 ;
        RECT 1288.920 835.105 1323.520 1032.730 ;
        RECT 1330.720 835.105 1331.120 1032.730 ;
        RECT 1338.320 835.105 1375.320 1032.730 ;
        RECT 1380.920 835.105 1383.320 1032.730 ;
        RECT 1388.920 835.105 1423.520 1032.730 ;
        RECT 1430.720 835.105 1431.120 1032.730 ;
        RECT 1438.320 850.560 1455.640 1032.730 ;
        RECT 1462.840 850.560 1463.240 1032.730 ;
        RECT 1470.440 850.560 1475.320 1032.730 ;
        RECT 1438.320 835.105 1475.320 850.560 ;
        RECT 1480.920 835.105 1483.320 1032.730 ;
        RECT 1488.920 835.105 1523.520 1032.730 ;
        RECT 1530.720 835.105 1531.120 1032.730 ;
        RECT 1538.320 835.105 1623.520 1032.730 ;
        RECT 1630.720 835.105 1631.120 1032.730 ;
        RECT 1638.320 835.105 1723.520 1032.730 ;
        RECT 1730.720 835.105 1731.120 1032.730 ;
        RECT 1738.320 850.560 1755.640 1032.730 ;
        RECT 1762.840 850.560 1763.240 1032.730 ;
        RECT 1770.440 850.560 1823.520 1032.730 ;
        RECT 1738.320 835.105 1823.520 850.560 ;
        RECT 1830.720 835.105 1831.120 1032.730 ;
        RECT 1838.320 835.105 1843.320 1032.730 ;
        RECT 1848.920 850.560 1851.320 1032.730 ;
        RECT 1856.920 850.560 1859.320 1032.730 ;
        RECT 1848.920 835.105 1859.320 850.560 ;
        RECT 1864.920 850.560 1867.320 1032.730 ;
        RECT 1872.920 850.560 1883.320 1032.730 ;
        RECT 1864.920 835.105 1883.320 850.560 ;
        RECT 1888.920 835.105 1891.320 1032.730 ;
        RECT 1896.920 835.105 1899.320 1032.730 ;
        RECT 1904.920 850.560 1907.320 1032.730 ;
        RECT 1912.920 850.560 1923.520 1032.730 ;
        RECT 1904.920 835.105 1923.520 850.560 ;
        RECT 1930.720 835.105 1931.120 1032.730 ;
        RECT 1938.320 835.105 2023.520 1032.730 ;
        RECT 2030.720 835.105 2031.120 1032.730 ;
        RECT 2038.320 850.560 2055.640 1032.730 ;
        RECT 2062.840 850.560 2063.240 1032.730 ;
        RECT 2070.440 850.560 2123.520 1032.730 ;
        RECT 2038.320 835.105 2123.520 850.560 ;
        RECT 2130.720 835.105 2131.120 1032.730 ;
        RECT 2138.320 835.105 2223.520 1032.730 ;
        RECT 2230.720 835.105 2231.120 1032.730 ;
        RECT 2238.320 835.105 2323.520 1032.730 ;
        RECT 2330.720 835.105 2331.120 1032.730 ;
        RECT 2338.320 850.560 2355.640 1032.730 ;
        RECT 2362.840 850.560 2363.240 1032.730 ;
        RECT 2370.440 850.560 2423.520 1032.730 ;
        RECT 2338.320 835.105 2423.520 850.560 ;
        RECT 2430.720 835.105 2431.120 1032.730 ;
        RECT 2438.320 835.105 2523.520 1032.730 ;
        RECT 2530.720 835.105 2531.120 1032.730 ;
        RECT 2538.320 835.105 2623.520 1032.730 ;
        RECT 76.320 114.415 2623.520 835.105 ;
        RECT 76.320 10.240 123.520 114.415 ;
        RECT 130.720 10.240 131.120 114.415 ;
        RECT 138.320 10.240 223.520 114.415 ;
        RECT 230.720 10.240 231.120 114.415 ;
        RECT 238.320 108.480 323.520 114.415 ;
        RECT 238.320 10.240 255.640 108.480 ;
        RECT 262.840 10.240 263.240 108.480 ;
        RECT 270.440 10.240 323.520 108.480 ;
        RECT 330.720 10.240 331.120 114.415 ;
        RECT 338.320 10.240 423.520 114.415 ;
        RECT 430.720 10.240 431.120 114.415 ;
        RECT 438.320 10.240 523.520 114.415 ;
        RECT 530.720 10.240 531.120 114.415 ;
        RECT 538.320 108.480 623.520 114.415 ;
        RECT 538.320 10.240 555.640 108.480 ;
        RECT 562.840 10.240 563.240 108.480 ;
        RECT 570.440 10.240 623.520 108.480 ;
        RECT 630.720 10.240 631.120 114.415 ;
        RECT 638.320 10.240 723.520 114.415 ;
        RECT 730.720 10.240 731.120 114.415 ;
        RECT 738.320 10.240 823.520 114.415 ;
        RECT 830.720 10.240 831.120 114.415 ;
        RECT 838.320 108.480 858.320 114.415 ;
        RECT 838.320 10.240 850.320 108.480 ;
        RECT 855.920 10.240 858.320 108.480 ;
        RECT 863.920 108.480 908.320 114.415 ;
        RECT 863.920 10.240 900.320 108.480 ;
        RECT 905.920 10.240 908.320 108.480 ;
        RECT 913.920 10.240 923.520 114.415 ;
        RECT 930.720 10.240 931.120 114.415 ;
        RECT 938.320 108.480 1123.520 114.415 ;
        RECT 938.320 10.240 955.640 108.480 ;
        RECT 962.840 10.240 963.240 108.480 ;
        RECT 970.440 10.240 1123.520 108.480 ;
        RECT 1130.720 10.240 1131.120 114.415 ;
        RECT 1138.320 108.480 1223.520 114.415 ;
        RECT 1138.320 10.240 1155.640 108.480 ;
        RECT 1162.840 10.240 1163.240 108.480 ;
        RECT 1170.440 10.240 1223.520 108.480 ;
        RECT 1230.720 10.240 1231.120 114.415 ;
        RECT 1238.320 10.240 1275.320 114.415 ;
        RECT 1280.920 10.240 1283.320 114.415 ;
        RECT 1288.920 10.240 1323.520 114.415 ;
        RECT 1330.720 10.240 1331.120 114.415 ;
        RECT 1338.320 10.240 1375.320 114.415 ;
        RECT 1380.920 10.240 1383.320 114.415 ;
        RECT 1388.920 10.240 1423.520 114.415 ;
        RECT 1430.720 10.240 1431.120 114.415 ;
        RECT 1438.320 108.480 1475.320 114.415 ;
        RECT 1438.320 10.240 1455.640 108.480 ;
        RECT 1462.840 10.240 1463.240 108.480 ;
        RECT 1470.440 10.240 1475.320 108.480 ;
        RECT 1480.920 10.240 1483.320 114.415 ;
        RECT 1488.920 10.240 1523.520 114.415 ;
        RECT 1530.720 10.240 1531.120 114.415 ;
        RECT 1538.320 10.240 1623.520 114.415 ;
        RECT 1630.720 10.240 1631.120 114.415 ;
        RECT 1638.320 10.240 1723.520 114.415 ;
        RECT 1730.720 10.240 1731.120 114.415 ;
        RECT 1738.320 108.480 1823.520 114.415 ;
        RECT 1738.320 10.240 1755.640 108.480 ;
        RECT 1762.840 10.240 1763.240 108.480 ;
        RECT 1770.440 10.240 1823.520 108.480 ;
        RECT 1830.720 10.240 1831.120 114.415 ;
        RECT 1838.320 10.240 1843.320 114.415 ;
        RECT 1848.920 108.480 1859.320 114.415 ;
        RECT 1848.920 10.240 1851.320 108.480 ;
        RECT 1856.920 10.240 1859.320 108.480 ;
        RECT 1864.920 108.480 1883.320 114.415 ;
        RECT 1864.920 10.240 1867.320 108.480 ;
        RECT 1872.920 10.240 1883.320 108.480 ;
        RECT 1888.920 10.240 1891.320 114.415 ;
        RECT 1896.920 10.240 1899.320 114.415 ;
        RECT 1904.920 108.480 1923.520 114.415 ;
        RECT 1904.920 10.240 1907.320 108.480 ;
        RECT 1912.920 10.240 1923.520 108.480 ;
        RECT 1930.720 10.240 1931.120 114.415 ;
        RECT 1938.320 10.240 2023.520 114.415 ;
        RECT 2030.720 10.240 2031.120 114.415 ;
        RECT 2038.320 108.480 2123.520 114.415 ;
        RECT 2038.320 10.240 2055.640 108.480 ;
        RECT 2062.840 10.240 2063.240 108.480 ;
        RECT 2070.440 10.240 2123.520 108.480 ;
        RECT 2130.720 10.240 2131.120 114.415 ;
        RECT 2138.320 10.240 2223.520 114.415 ;
        RECT 2230.720 10.240 2231.120 114.415 ;
        RECT 2238.320 10.240 2323.520 114.415 ;
        RECT 2330.720 10.240 2331.120 114.415 ;
        RECT 2338.320 108.480 2423.520 114.415 ;
        RECT 2338.320 10.240 2355.640 108.480 ;
        RECT 2362.840 10.240 2363.240 108.480 ;
        RECT 2370.440 10.240 2423.520 108.480 ;
        RECT 2430.720 10.240 2431.120 114.415 ;
        RECT 2438.320 10.240 2523.520 114.415 ;
        RECT 2530.720 10.240 2531.120 114.415 ;
        RECT 2538.320 10.240 2623.520 114.415 ;
        RECT 2630.720 10.240 2631.120 1032.730 ;
        RECT 2638.320 10.240 2648.320 1032.730 ;
        RECT 2653.920 10.240 2655.120 1032.730 ;
        RECT 2660.720 939.420 2723.520 1032.730 ;
        RECT 2730.720 939.420 2731.120 1032.730 ;
        RECT 2738.320 939.420 2755.640 1032.730 ;
        RECT 2762.840 939.420 2763.240 1032.730 ;
        RECT 2660.720 904.100 2763.240 939.420 ;
        RECT 2660.720 797.420 2723.520 904.100 ;
        RECT 2730.720 797.420 2731.120 904.100 ;
        RECT 2660.720 793.305 2731.120 797.420 ;
        RECT 2738.320 797.420 2755.640 904.100 ;
        RECT 2762.840 797.420 2763.240 904.100 ;
        RECT 2770.440 960.800 2823.520 1032.730 ;
        RECT 2770.440 886.080 2776.880 960.800 ;
        RECT 2782.680 886.080 2783.320 960.800 ;
        RECT 2789.120 939.420 2823.520 960.800 ;
        RECT 2830.720 939.420 2831.120 1032.730 ;
        RECT 2838.320 939.420 2923.520 1032.730 ;
        RECT 2789.120 904.100 2923.520 939.420 ;
        RECT 2789.120 886.080 2823.520 904.100 ;
        RECT 2770.440 797.420 2823.520 886.080 ;
        RECT 2738.320 793.305 2823.520 797.420 ;
        RECT 2830.720 793.305 2831.120 904.100 ;
        RECT 2838.320 793.305 2923.520 904.100 ;
        RECT 2930.720 793.305 2931.120 1032.730 ;
        RECT 2938.320 793.305 2967.975 1032.730 ;
        RECT 2660.720 793.205 2967.975 793.305 ;
        RECT 2970.375 793.205 2990.355 1032.830 ;
        RECT 2992.755 1032.730 3086.780 1032.830 ;
        RECT 2992.755 793.305 3023.520 1032.730 ;
        RECT 3030.720 797.420 3031.120 1032.730 ;
        RECT 3038.320 797.420 3086.780 1032.730 ;
        RECT 3030.720 793.305 3086.780 797.420 ;
        RECT 2992.755 793.205 3086.780 793.305 ;
        RECT 2660.720 269.915 3086.780 793.205 ;
        RECT 2660.720 269.815 2967.975 269.915 ;
        RECT 2660.720 267.060 2731.120 269.815 ;
        RECT 2660.720 10.240 2723.520 267.060 ;
        RECT 2730.720 10.240 2731.120 267.060 ;
        RECT 2738.320 267.060 2823.520 269.815 ;
        RECT 2738.320 10.240 2755.640 267.060 ;
        RECT 2762.840 10.240 2763.240 267.060 ;
        RECT 2770.440 103.220 2823.520 267.060 ;
        RECT 2830.720 103.220 2831.120 269.815 ;
        RECT 2838.320 103.220 2923.520 269.815 ;
        RECT 2770.440 10.240 2923.520 103.220 ;
        RECT 2930.720 10.240 2931.120 269.815 ;
        RECT 2938.320 10.240 2967.975 269.815 ;
        RECT 2970.375 10.240 2990.355 269.915 ;
        RECT 2992.755 269.815 3086.780 269.915 ;
        RECT 2992.755 10.240 3023.520 269.815 ;
        RECT 3030.720 267.060 3086.780 269.815 ;
        RECT 3030.720 10.240 3031.120 267.060 ;
        RECT 3038.320 10.240 3086.780 267.060 ;
        RECT 3089.580 10.240 3089.780 4755.200 ;
        RECT 3092.580 10.240 3092.780 4755.200 ;
        RECT 3098.580 10.240 3098.780 4755.200 ;
        RECT 3104.580 10.240 3104.780 4755.200 ;
        RECT 3110.580 10.240 3110.780 4755.200 ;
        RECT 3116.580 10.240 3116.780 4755.200 ;
        RECT 3122.580 10.240 3122.780 4755.200 ;
        RECT 3128.580 10.240 3128.780 4755.200 ;
        RECT 3134.580 10.240 3134.780 4755.200 ;
        RECT 3140.580 10.240 3140.780 4755.200 ;
        RECT 3146.580 10.240 3146.780 4755.200 ;
        RECT 3152.580 4402.000 3165.000 4755.200 ;
        RECT 3152.580 4378.055 3171.230 4402.000 ;
        RECT 3152.580 4376.450 3165.000 4378.055 ;
        RECT 3152.580 4353.345 3171.230 4376.450 ;
        RECT 3152.580 4351.745 3165.000 4353.345 ;
        RECT 3152.580 4327.800 3171.230 4351.745 ;
        RECT 3152.580 3956.005 3165.000 4327.800 ;
        RECT 3152.580 3932.060 3171.230 3956.005 ;
        RECT 3152.580 3906.090 3165.000 3932.060 ;
        RECT 3152.580 3882.145 3171.230 3906.090 ;
        RECT 3152.580 2383.005 3165.000 3882.145 ;
        RECT 3152.580 2359.060 3171.230 2383.005 ;
        RECT 3152.580 2333.090 3165.000 2359.060 ;
        RECT 3152.580 2309.145 3171.230 2333.090 ;
        RECT 3152.580 2163.000 3165.000 2309.145 ;
        RECT 3152.580 2139.055 3171.230 2163.000 ;
        RECT 3152.580 2137.450 3165.000 2139.055 ;
        RECT 3152.580 2114.345 3171.230 2137.450 ;
        RECT 3152.580 2112.745 3165.000 2114.345 ;
        RECT 3152.580 2088.800 3171.230 2112.745 ;
        RECT 3152.580 1942.045 3165.000 2088.800 ;
        RECT 3152.580 1918.100 3171.230 1942.045 ;
        RECT 3152.580 1892.130 3165.000 1918.100 ;
        RECT 3152.580 1868.185 3171.230 1892.130 ;
        RECT 3152.580 10.240 3165.000 1868.185 ;
        RECT 0.000 0.000 3165.000 10.240 ;
        RECT 878.500 -9.685 896.510 0.000 ;
        RECT 994.715 -9.120 1018.745 0.000 ;
        RECT 1044.970 -9.120 1069.000 0.000 ;
        RECT 1075.025 -9.685 1088.745 0.000 ;
        RECT 1075.025 -40.985 1088.745 -36.425 ;
      LAYER met5 ;
        RECT 0.000 4629.480 3165.000 4629.950 ;
        RECT 0.000 4611.080 8.280 4629.480 ;
        RECT 75.510 4620.680 3087.590 4629.480 ;
        RECT 77.520 4611.080 3085.580 4620.680 ;
        RECT 3156.520 4611.080 3165.000 4629.480 ;
        RECT 0.000 4529.480 3165.000 4611.080 ;
        RECT 0.000 4511.080 8.280 4529.480 ;
        RECT 77.520 4520.680 3086.580 4529.480 ;
        RECT 77.520 4511.080 3085.580 4520.680 ;
        RECT 3156.520 4511.080 3165.000 4529.480 ;
        RECT 0.000 4429.480 3165.000 4511.080 ;
        RECT 0.000 4424.200 3086.580 4429.480 ;
        RECT -9.290 4420.680 3086.580 4424.200 ;
        RECT -9.290 4411.080 3085.580 4420.680 ;
        RECT 3156.520 4411.080 3165.000 4429.480 ;
        RECT -9.290 4402.000 3165.000 4411.080 ;
        RECT -9.290 4400.250 3171.230 4402.000 ;
        RECT 0.000 4398.650 3171.230 4400.250 ;
        RECT -9.290 4378.050 3171.230 4398.650 ;
        RECT -9.290 4376.450 3165.000 4378.050 ;
        RECT -9.290 4375.600 3171.230 4376.450 ;
        RECT 0.000 4374.000 3171.230 4375.600 ;
        RECT -9.290 4353.345 3171.230 4374.000 ;
        RECT -9.290 4351.745 3165.000 4353.345 ;
        RECT -9.290 4350.050 3171.230 4351.745 ;
        RECT 0.000 4329.480 3171.230 4350.050 ;
        RECT 0.000 4311.080 8.280 4329.480 ;
        RECT 77.520 4327.795 3171.230 4329.480 ;
        RECT 77.520 4320.680 3165.000 4327.795 ;
        RECT 77.520 4311.080 3085.580 4320.680 ;
        RECT 3156.520 4311.080 3165.000 4320.680 ;
        RECT 0.000 4229.480 3165.000 4311.080 ;
        RECT 0.000 4211.080 8.280 4229.480 ;
        RECT 77.520 4220.680 3086.580 4229.480 ;
        RECT 77.520 4211.080 3085.580 4220.680 ;
        RECT 3156.520 4211.080 3165.000 4229.480 ;
        RECT 0.000 4129.480 3165.000 4211.080 ;
        RECT 0.000 4111.080 8.280 4129.480 ;
        RECT 77.520 4120.680 3086.580 4129.480 ;
        RECT 77.520 4111.080 3085.580 4120.680 ;
        RECT 3156.520 4111.080 3165.000 4129.480 ;
        RECT 0.000 4029.480 3165.000 4111.080 ;
        RECT 0.000 4011.080 8.280 4029.480 ;
        RECT 77.520 4020.680 3086.580 4029.480 ;
        RECT 77.520 4011.080 3085.580 4020.680 ;
        RECT 3156.520 4011.080 3165.000 4029.480 ;
        RECT 0.000 4001.790 3165.000 4011.080 ;
        RECT -9.290 3977.840 3165.000 4001.790 ;
        RECT 0.000 3956.005 3165.000 3977.840 ;
        RECT 0.000 3951.895 3171.230 3956.005 ;
        RECT -9.290 3932.055 3171.230 3951.895 ;
        RECT -9.290 3927.945 3165.000 3932.055 ;
        RECT 0.000 3906.090 3165.000 3927.945 ;
        RECT 0.000 3882.140 3171.230 3906.090 ;
        RECT 0.000 3829.480 3165.000 3882.140 ;
        RECT 0.000 3811.080 8.280 3829.480 ;
        RECT 77.520 3820.680 3086.580 3829.480 ;
        RECT 77.520 3811.080 3085.580 3820.680 ;
        RECT 3156.520 3811.080 3165.000 3829.480 ;
        RECT 0.000 3729.480 3165.000 3811.080 ;
        RECT 0.000 3711.080 8.280 3729.480 ;
        RECT 77.520 3720.680 3086.580 3729.480 ;
        RECT 77.520 3711.080 3085.580 3720.680 ;
        RECT 3156.520 3711.080 3165.000 3729.480 ;
        RECT 0.000 3629.480 3165.000 3711.080 ;
        RECT 0.000 3611.080 8.280 3629.480 ;
        RECT 77.520 3620.680 3086.580 3629.480 ;
        RECT 77.520 3611.080 3085.580 3620.680 ;
        RECT 3156.520 3611.080 3165.000 3629.480 ;
        RECT 0.000 3529.480 3165.000 3611.080 ;
        RECT 0.000 3511.080 8.280 3529.480 ;
        RECT 77.520 3520.680 3086.580 3529.480 ;
        RECT 77.520 3511.080 3085.580 3520.680 ;
        RECT 3156.520 3511.080 3165.000 3529.480 ;
        RECT 0.000 3429.480 3165.000 3511.080 ;
        RECT 0.000 3411.080 8.280 3429.480 ;
        RECT 77.520 3420.680 3086.580 3429.480 ;
        RECT 77.520 3411.080 3085.580 3420.680 ;
        RECT 3156.520 3411.080 3165.000 3429.480 ;
        RECT 0.000 3329.480 3165.000 3411.080 ;
        RECT 0.000 3311.080 8.280 3329.480 ;
        RECT 77.520 3320.680 3086.580 3329.480 ;
        RECT 77.520 3311.080 3085.580 3320.680 ;
        RECT 3156.520 3311.080 3165.000 3329.480 ;
        RECT 0.000 3229.480 3165.000 3311.080 ;
        RECT 0.000 3211.080 8.280 3229.480 ;
        RECT 77.520 3220.680 3086.580 3229.480 ;
        RECT 77.520 3211.080 3085.580 3220.680 ;
        RECT 3156.520 3211.080 3165.000 3229.480 ;
        RECT 0.000 3129.480 3165.000 3211.080 ;
        RECT 0.000 3111.080 8.280 3129.480 ;
        RECT 77.520 3120.680 3086.580 3129.480 ;
        RECT 77.520 3111.080 3085.580 3120.680 ;
        RECT 3156.520 3111.080 3165.000 3129.480 ;
        RECT 0.000 3029.480 3165.000 3111.080 ;
        RECT 0.000 3011.080 8.280 3029.480 ;
        RECT 77.520 3020.680 3086.580 3029.480 ;
        RECT 77.520 3011.080 3085.580 3020.680 ;
        RECT 3156.520 3011.080 3165.000 3029.480 ;
        RECT 0.000 2929.480 3165.000 3011.080 ;
        RECT 0.000 2911.080 8.280 2929.480 ;
        RECT 77.520 2920.680 3086.580 2929.480 ;
        RECT 77.520 2911.080 3085.580 2920.680 ;
        RECT 3156.520 2911.080 3165.000 2929.480 ;
        RECT 0.000 2829.480 3165.000 2911.080 ;
        RECT 0.000 2811.080 8.280 2829.480 ;
        RECT 77.520 2820.680 3086.580 2829.480 ;
        RECT 77.520 2811.080 3085.580 2820.680 ;
        RECT 3156.520 2811.080 3165.000 2829.480 ;
        RECT 0.000 2729.480 3165.000 2811.080 ;
        RECT 0.000 2711.080 8.280 2729.480 ;
        RECT 77.520 2720.680 3086.580 2729.480 ;
        RECT 77.520 2711.080 3085.580 2720.680 ;
        RECT 3156.520 2711.080 3165.000 2729.480 ;
        RECT 0.000 2629.480 3165.000 2711.080 ;
        RECT 0.000 2611.080 8.280 2629.480 ;
        RECT 77.520 2620.680 3086.580 2629.480 ;
        RECT 77.520 2611.080 3085.580 2620.680 ;
        RECT 3156.520 2611.080 3165.000 2629.480 ;
        RECT 0.000 2529.480 3165.000 2611.080 ;
        RECT 0.000 2511.080 8.280 2529.480 ;
        RECT 77.520 2520.680 3086.580 2529.480 ;
        RECT 77.520 2511.080 3085.580 2520.680 ;
        RECT 3156.520 2511.080 3165.000 2529.480 ;
        RECT 0.000 2429.480 3165.000 2511.080 ;
        RECT 0.000 2411.080 8.280 2429.480 ;
        RECT 77.520 2420.680 3086.580 2429.480 ;
        RECT 77.520 2411.080 3085.580 2420.680 ;
        RECT 3156.520 2411.080 3165.000 2429.480 ;
        RECT 0.000 2383.005 3165.000 2411.080 ;
        RECT 0.000 2359.055 3171.230 2383.005 ;
        RECT 0.000 2333.090 3165.000 2359.055 ;
        RECT 0.000 2329.480 3171.230 2333.090 ;
        RECT 0.000 2311.080 8.280 2329.480 ;
        RECT 77.520 2311.080 3171.230 2329.480 ;
        RECT 0.000 2309.140 3171.230 2311.080 ;
        RECT 0.000 2278.790 3165.000 2309.140 ;
        RECT -9.290 2254.840 3165.000 2278.790 ;
        RECT 0.000 2229.480 3165.000 2254.840 ;
        RECT 0.000 2228.895 3086.580 2229.480 ;
        RECT -9.290 2220.680 3086.580 2228.895 ;
        RECT -9.290 2211.080 3085.580 2220.680 ;
        RECT 3156.520 2211.080 3165.000 2229.480 ;
        RECT -9.290 2204.945 3165.000 2211.080 ;
        RECT 0.000 2163.000 3165.000 2204.945 ;
        RECT 0.000 2139.050 3171.230 2163.000 ;
        RECT 0.000 2137.450 3165.000 2139.050 ;
        RECT 0.000 2129.480 3171.230 2137.450 ;
        RECT 0.000 2111.080 8.280 2129.480 ;
        RECT 77.520 2114.345 3171.230 2129.480 ;
        RECT 77.520 2112.745 3165.000 2114.345 ;
        RECT 77.520 2111.080 3171.230 2112.745 ;
        RECT 0.000 2088.795 3171.230 2111.080 ;
        RECT 0.000 2068.200 3165.000 2088.795 ;
        RECT -9.290 2044.250 3165.000 2068.200 ;
        RECT 0.000 2042.650 3165.000 2044.250 ;
        RECT -9.290 2029.480 3165.000 2042.650 ;
        RECT -9.290 2020.680 3086.580 2029.480 ;
        RECT -9.290 2019.600 3085.580 2020.680 ;
        RECT 0.000 2018.000 3085.580 2019.600 ;
        RECT -9.290 2011.080 3085.580 2018.000 ;
        RECT 3156.520 2011.080 3165.000 2029.480 ;
        RECT -9.290 1994.050 3165.000 2011.080 ;
        RECT 0.000 1942.045 3165.000 1994.050 ;
        RECT 0.000 1929.480 3171.230 1942.045 ;
        RECT 0.000 1911.080 8.280 1929.480 ;
        RECT 77.520 1918.095 3171.230 1929.480 ;
        RECT 77.520 1911.080 3165.000 1918.095 ;
        RECT 0.000 1892.130 3165.000 1911.080 ;
        RECT 0.000 1868.180 3171.230 1892.130 ;
        RECT 0.000 1829.480 3165.000 1868.180 ;
        RECT 0.000 1811.080 8.280 1829.480 ;
        RECT 77.520 1820.680 3086.580 1829.480 ;
        RECT 77.520 1811.080 3085.580 1820.680 ;
        RECT 3156.520 1811.080 3165.000 1829.480 ;
        RECT 0.000 1729.480 3165.000 1811.080 ;
        RECT 0.000 1711.080 8.280 1729.480 ;
        RECT 77.520 1720.680 3086.580 1729.480 ;
        RECT 77.520 1711.080 3085.580 1720.680 ;
        RECT 3156.520 1711.080 3165.000 1729.480 ;
        RECT 0.000 1629.480 3165.000 1711.080 ;
        RECT 0.000 1611.080 8.280 1629.480 ;
        RECT 77.520 1620.680 3086.580 1629.480 ;
        RECT 77.520 1611.080 3085.580 1620.680 ;
        RECT 3156.520 1611.080 3165.000 1629.480 ;
        RECT 0.000 1529.480 3165.000 1611.080 ;
        RECT 0.000 1511.080 8.280 1529.480 ;
        RECT 77.520 1520.680 3086.580 1529.480 ;
        RECT 77.520 1511.080 3085.580 1520.680 ;
        RECT 3156.520 1511.080 3165.000 1529.480 ;
        RECT 0.000 1429.480 3165.000 1511.080 ;
        RECT 0.000 1411.080 8.280 1429.480 ;
        RECT 77.520 1420.680 3086.580 1429.480 ;
        RECT 77.520 1411.080 3085.580 1420.680 ;
        RECT 3156.520 1411.080 3165.000 1429.480 ;
        RECT 0.000 1329.480 3165.000 1411.080 ;
        RECT 0.000 1311.080 8.280 1329.480 ;
        RECT 77.520 1320.680 3086.580 1329.480 ;
        RECT 77.520 1311.080 3085.580 1320.680 ;
        RECT 3156.520 1311.080 3165.000 1329.480 ;
        RECT 0.000 1229.480 3165.000 1311.080 ;
        RECT 0.000 1211.080 8.280 1229.480 ;
        RECT 77.520 1220.680 3086.580 1229.480 ;
        RECT 77.520 1211.080 3085.580 1220.680 ;
        RECT 3156.520 1211.080 3165.000 1229.480 ;
        RECT 0.000 1129.480 3165.000 1211.080 ;
        RECT 0.000 1111.080 8.280 1129.480 ;
        RECT 77.520 1120.680 3086.580 1129.480 ;
        RECT 77.520 1111.080 3085.580 1120.680 ;
        RECT 3156.520 1111.080 3165.000 1129.480 ;
        RECT 0.000 1029.480 3165.000 1111.080 ;
        RECT 0.000 1011.080 8.280 1029.480 ;
        RECT 3156.520 1011.080 3165.000 1029.480 ;
        RECT 0.000 985.800 3165.000 1011.080 ;
        RECT 0.000 951.400 8.280 985.800 ;
        RECT 3156.520 951.400 3165.000 985.800 ;
        RECT 0.000 929.480 3165.000 951.400 ;
        RECT 0.000 911.080 8.280 929.480 ;
        RECT 3156.520 911.080 3165.000 929.480 ;
        RECT 0.000 906.780 3165.000 911.080 ;
        RECT 0.000 851.180 8.280 906.780 ;
        RECT 3156.520 851.180 3165.000 906.780 ;
        RECT 0.000 829.480 3165.000 851.180 ;
        RECT 0.000 811.080 8.280 829.480 ;
        RECT 556.860 811.080 2601.300 819.880 ;
        RECT 3156.520 811.080 3165.000 829.480 ;
        RECT 0.000 729.480 3165.000 811.080 ;
        RECT 0.000 711.080 8.280 729.480 ;
        RECT 556.860 711.080 2601.300 729.480 ;
        RECT 3156.520 711.080 3165.000 729.480 ;
        RECT 0.000 629.480 3165.000 711.080 ;
        RECT 0.000 611.080 8.280 629.480 ;
        RECT 556.860 611.080 2601.300 629.480 ;
        RECT 3156.520 611.080 3165.000 629.480 ;
        RECT 0.000 529.480 3165.000 611.080 ;
        RECT 0.000 511.080 8.280 529.480 ;
        RECT 556.860 511.080 2601.300 529.480 ;
        RECT 3156.520 511.080 3165.000 529.480 ;
        RECT 0.000 429.480 3165.000 511.080 ;
        RECT 0.000 411.080 8.280 429.480 ;
        RECT 556.860 411.080 2601.300 429.480 ;
        RECT 3156.520 411.080 3165.000 429.480 ;
        RECT 0.000 329.480 3165.000 411.080 ;
        RECT 0.000 311.080 8.280 329.480 ;
        RECT 556.860 311.080 2601.300 329.480 ;
        RECT 3156.520 311.080 3165.000 329.480 ;
        RECT 0.000 229.480 3165.000 311.080 ;
        RECT 0.000 211.080 8.280 229.480 ;
        RECT 556.860 211.080 2601.300 229.480 ;
        RECT 3156.520 211.080 3165.000 229.480 ;
        RECT 0.000 204.200 3165.000 211.080 ;
        RECT -9.290 180.250 3165.000 204.200 ;
        RECT 0.000 167.980 3165.000 180.250 ;
        RECT 0.000 158.780 2601.300 167.980 ;
        RECT 2722.055 158.780 3165.000 167.980 ;
        RECT 0.000 154.000 2612.860 158.780 ;
        RECT -9.290 150.780 2612.860 154.000 ;
        RECT 2682.965 150.780 3165.000 158.780 ;
        RECT -9.290 133.980 3165.000 150.780 ;
        RECT -9.290 130.050 120.000 133.980 ;
        RECT 0.000 116.780 120.000 130.050 ;
        RECT 2682.965 116.780 3165.000 133.980 ;
        RECT 0.000 109.580 3165.000 116.780 ;
  END
END caravel_core
END LIBRARY

