* NGSPICE file created from gpio_control_block.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VPWR X VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VPWR X VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VPWR X VNB VPB
X0 a_244_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X1 VPWR a_244_47# a_355_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X2 X a_355_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_244_47# a_355_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X6 X a_355_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_244_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VPWR X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_791_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR RESET_B a_941_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1415_315# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_791_47# a_941_21# a_647_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VGND a_1415_315# a_1363_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1340_413# a_27_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_473_413# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_1555_47# a_941_21# a_1415_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VPWR a_1415_315# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1256_413# a_193_47# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_581_47# a_27_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_647_21# a_473_413# a_791_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_647_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_941_21# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 a_557_413# a_193_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_473_413# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_891_329# a_473_413# a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q_N a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND RESET_B a_941_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_647_21# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1112_329# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 VGND a_647_21# a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_1415_315# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VPWR a_941_21# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VPWR a_1415_315# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1363_47# a_193_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1159_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1672_329# a_1256_413# a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1256_413# a_27_47# a_1159_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 a_1415_315# a_1256_413# a_1555_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VPWR Z VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X21 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X26 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X32 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VPWR X VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_logic1 gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_4_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VPWR X VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VPWR Z VNB VPB
X0 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_116_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X14 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_301_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_301_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_116_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X31 VGND A a_116_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X33 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X36 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
X_200_ _200_/A vssd vccd _201_/A vssd vccd sky130_fd_sc_hd__buf_1
X_131_ _131_/A vssd vccd _131_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_114_ _114_/A vssd vccd _114_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 user_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput31 _205_/X vssd vccd pad_gpio_outenb vssd vccd sky130_fd_sc_hd__buf_2
X_130_ _136_/A _132_/B vssd vccd _131_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_113_ _187_/A _113_/B vssd vccd _114_/A vssd vccd sky130_fd_sc_hd__or2_1
XFILLER_0_58 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput32 _212_/Q vssd vccd pad_gpio_slow_sel vssd vccd sky130_fd_sc_hd__buf_2
Xoutput21 _220_/Q vssd vccd pad_gpio_ana_en vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_6 user_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_189_ _189_/A _189_/B vssd vccd _190_/A vssd vccd sky130_fd_sc_hd__or2_1
Xhold10 _226_/D vssd vccd _211_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_112_ _202_/A vssd vccd _187_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_7 serial_data_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput33 _213_/Q vssd vccd pad_gpio_vtrip_sel vssd vccd sky130_fd_sc_hd__buf_2
Xoutput22 _222_/Q vssd vccd pad_gpio_ana_pol vssd vccd sky130_fd_sc_hd__buf_2
X_188_ _188_/A vssd vccd _188_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_111_ _111_/A vssd vccd _111_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold11 _224_/D vssd vccd _210_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput34 _202_/X vssd vccd resetn_out vssd vccd sky130_fd_sc_hd__buf_2
Xoutput23 _221_/Q vssd vccd pad_gpio_ana_sel vssd vccd sky130_fd_sc_hd__buf_2
X_187_ _187_/A _189_/A vssd vccd _188_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_110_ _136_/A _113_/B vssd vccd _111_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold12 _230_/D vssd vccd _221_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput24 _217_/Q vssd vccd pad_gpio_dm[0] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput35 _203_/X vssd vccd serial_clock_out vssd vccd sky130_fd_sc_hd__clkbuf_1
X_186_ _186_/A vssd vccd _186_/X vssd vccd sky130_fd_sc_hd__buf_1
X_169_ _169_/A _171_/B vssd vccd _170_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold13 _233_/D vssd vccd hold1/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput36 _199_/X vssd vccd serial_data_out vssd vccd sky130_fd_sc_hd__buf_2
Xoutput25 _218_/Q vssd vccd pad_gpio_dm[1] vssd vccd sky130_fd_sc_hd__buf_2
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_185_ _185_/A vssd vccd _186_/A vssd vccd sky130_fd_sc_hd__buf_1
X_168_ _168_/A vssd vccd _168_/X vssd vccd sky130_fd_sc_hd__buf_1
Xhold14 _231_/D vssd vccd _222_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput37 _204_/X vssd vccd serial_load_out vssd vccd sky130_fd_sc_hd__clkbuf_1
Xoutput26 _219_/Q vssd vccd pad_gpio_dm[2] vssd vccd sky130_fd_sc_hd__buf_2
X_184_ _184_/A vssd vccd _184_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_167_ _173_/A vssd vccd _168_/A vssd vccd sky130_fd_sc_hd__buf_1
Xhold15 _232_/D vssd vccd hold4/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_219_ _129_/X hold8/X _133_/X _131_/X vssd vccd _219_/Q _219_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
Xoutput27 _211_/Q vssd vccd pad_gpio_holdover vssd vccd sky130_fd_sc_hd__buf_2
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_183_ _183_/A _183_/B vssd vccd _184_/A vssd vccd sky130_fd_sc_hd__or2_1
X_166_ _166_/A vssd vccd _166_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_235_ _203_/A _235_/D _202_/A vssd vccd hold8/A vssd vccd sky130_fd_sc_hd__dfrtp_1
Xoutput28 _215_/Q vssd vccd pad_gpio_ib_mode_sel vssd vccd sky130_fd_sc_hd__buf_2
Xhold16 _228_/D vssd vccd hold2/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_149_ _149_/A vssd vccd _149_/X vssd vccd sky130_fd_sc_hd__buf_1
X_218_ _135_/X hold5/X _139_/X _137_/X vssd vccd _218_/Q _218_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_182_ _182_/A vssd vccd _182_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_148_ _173_/A vssd vccd _149_/A vssd vccd sky130_fd_sc_hd__buf_1
X_165_ _183_/A _165_/B vssd vccd _166_/A vssd vccd sky130_fd_sc_hd__or2_1
X_217_ _141_/X hold6/X _146_/X _144_/X vssd vccd _217_/Q _206_/A0 vssd vccd sky130_fd_sc_hd__dfbbn_1
X_234_ _203_/A _234_/D _202_/A vssd vccd _235_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xhold17 _234_/D vssd vccd hold6/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput29 _214_/Q vssd vccd pad_gpio_inenb vssd vccd sky130_fd_sc_hd__buf_2
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_181_ _187_/A _183_/B vssd vccd _182_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_164_ _164_/A vssd vccd _164_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_233_ _203_/A _233_/D _202_/A vssd vccd _234_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xhold18 _225_/D vssd vccd hold3/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_216_ _149_/X hold3/X _153_/X _151_/X vssd vccd _216_/Q _216_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_147_ _147_/A vssd vccd _173_/A vssd vccd sky130_fd_sc_hd__buf_1
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_180_ _180_/A vssd vccd _180_/X vssd vccd sky130_fd_sc_hd__buf_1
X_232_ _203_/A _232_/D _202_/A vssd vccd _233_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_163_ _169_/A _165_/B vssd vccd _164_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold19 _235_/D vssd vccd hold5/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_146_ _146_/A vssd vccd _146_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_215_ _155_/X hold2/X _160_/X _157_/X vssd vccd _215_/Q _215_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_129_ _129_/A vssd vccd _129_/X vssd vccd sky130_fd_sc_hd__buf_1
X_231_ _231_/CLK _231_/D _202_/A vssd vccd _232_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_162_ _162_/A vssd vccd _162_/X vssd vccd sky130_fd_sc_hd__buf_1
X_145_ _152_/A _145_/B vssd vccd _146_/A vssd vccd sky130_fd_sc_hd__or2_1
X_214_ _162_/X hold7/X _166_/X _164_/X vssd vccd _214_/Q _214_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
Xinput1 gpio_defaults[0] vssd vccd _189_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_128_ _140_/A vssd vccd _129_/A vssd vccd sky130_fd_sc_hd__buf_1
X_161_ _173_/A vssd vccd _162_/A vssd vccd sky130_fd_sc_hd__buf_1
X_230_ _231_/CLK _230_/D _202_/A vssd vccd _231_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xinput2 gpio_defaults[10] vssd vccd _145_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xgpio_in_buf _197_/Y gpio_in_buf/TE vssd vccd user_gpio_in vssd vccd sky130_fd_sc_hd__einvp_8
X_144_ _144_/A vssd vccd _144_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_213_ _168_/X hold1/X _172_/X _170_/X vssd vccd _213_/Q _213_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_127_ _127_/A vssd vccd _127_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_212_ _174_/X hold4/X _178_/X _176_/X vssd vccd _212_/Q _212_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_143_ _169_/A _145_/B vssd vccd _144_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_160_ _160_/A vssd vccd _160_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput3 gpio_defaults[11] vssd vccd _138_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_126_ _152_/A _126_/B vssd vccd _127_/A vssd vccd sky130_fd_sc_hd__or2_1
X_109_ _189_/B vssd vccd _136_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput4 gpio_defaults[12] vssd vccd _132_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_211_ _180_/X _211_/D _184_/X _182_/X vssd vccd _211_/Q _211_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_125_ _189_/B vssd vccd _152_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_142_ _189_/B vssd vccd _169_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_108_ _202_/A vssd vccd _189_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_210_ _186_/X _210_/D _190_/X _188_/X vssd vccd _210_/Q _210_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_141_ _141_/A vssd vccd _141_/X vssd vccd sky130_fd_sc_hd__buf_1
Xinput5 gpio_defaults[1] vssd vccd _152_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vccd _203_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
X_124_ _124_/A vssd vccd _124_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_115__1 serial_load vssd vccd _200_/A vssd vccd sky130_fd_sc_hd__inv_2
X_140_ _140_/A vssd vccd _141_/A vssd vccd sky130_fd_sc_hd__buf_1
Xinput6 gpio_defaults[2] vssd vccd _183_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput20 user_gpio_out vssd vccd _208_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
X_123_ _136_/A _126_/B vssd vccd _124_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_115__2 serial_load vssd vccd _185_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput7 gpio_defaults[3] vssd vccd _165_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_199_ _199_/A vssd vccd _199_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput10 gpio_defaults[6] vssd vccd _119_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_122_ _122_/A vssd vccd _122_/X vssd vccd sky130_fd_sc_hd__buf_1
X_115__3 serial_load vssd vccd _179_/A vssd vccd sky130_fd_sc_hd__inv_2
X_198_ one hold8/A vssd vccd _199_/A vssd vccd sky130_fd_sc_hd__and2_1
Xinput8 gpio_defaults[4] vssd vccd _159_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput11 gpio_defaults[7] vssd vccd _113_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_121_ _140_/A vssd vccd _122_/A vssd vccd sky130_fd_sc_hd__buf_1
X_115__4 serial_load vssd vccd _147_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput9 gpio_defaults[5] vssd vccd _126_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput12 gpio_defaults[8] vssd vccd _177_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_120_ _120_/A vssd vccd _120_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_197_ _209_/A vssd vccd _197_/Y vssd vccd sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd vccd hold1/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_115__5 serial_load vssd vccd _116_/A vssd vccd sky130_fd_sc_hd__inv_2
X_196_ _196_/A vssd vccd _206_/S vssd vccd sky130_fd_sc_hd__clkbuf_1
X_179_ _179_/A vssd vccd _180_/A vssd vccd sky130_fd_sc_hd__buf_1
Xinput13 gpio_defaults[9] vssd vccd _171_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold2 hold2/A vssd vccd hold2/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
X_195_ _219_/Q _218_/Q vssd vccd _196_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xinput14 mgmt_gpio_oeb vssd vccd _207_/S vssd vccd sky130_fd_sc_hd__clkbuf_1
X_178_ _178_/A vssd vccd _178_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold3 hold3/A vssd vccd hold3/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_30 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_194_ _194_/A vssd vccd _194_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_177_ _183_/A _177_/B vssd vccd _178_/A vssd vccd sky130_fd_sc_hd__or2_1
Xinput15 mgmt_gpio_out vssd vccd _207_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold4 hold4/A vssd vccd hold4/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_229_ _231_/CLK hold9/A _202_/A vssd vccd _230_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
XPHY_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_193_ _216_/Q _207_/S vssd vccd _194_/A vssd vccd sky130_fd_sc_hd__and2_1
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_176_ _176_/A vssd vccd _176_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_159_ _183_/A _159_/B vssd vccd _160_/A vssd vccd sky130_fd_sc_hd__or2_1
X_228_ _231_/CLK _228_/D _202_/A vssd vccd hold9/A vssd vccd sky130_fd_sc_hd__dfrtp_1
Xinput16 pad_gpio_in vssd vccd _209_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold5 hold5/A vssd vccd hold5/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_32 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_192_ _192_/A vssd vccd _192_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput17 resetn vssd vccd _202_/A vssd vccd sky130_fd_sc_hd__buf_6
X_175_ _187_/A _177_/B vssd vccd _176_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_158_ _189_/B vssd vccd _183_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold6 hold6/A vssd vccd hold6/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_227_ _231_/CLK hold7/A _202_/A vssd vccd _228_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vccd _231_/CLK vssd vccd sky130_fd_sc_hd__clkbuf_2
XPHY_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vccd clkbuf_0_serial_clock/X vssd vccd sky130_fd_sc_hd__clkbuf_16
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_191_ _214_/Q _216_/Q vssd vccd _192_/A vssd vccd sky130_fd_sc_hd__or2b_1
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_174_ _174_/A vssd vccd _174_/X vssd vccd sky130_fd_sc_hd__buf_1
X_226_ _231_/CLK _226_/D _202_/A vssd vccd hold7/A vssd vccd sky130_fd_sc_hd__dfrtp_1
X_157_ _157_/A vssd vccd _157_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput18 serial_data_in vssd vccd _223_/D vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold7 hold7/A vssd vccd hold7/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_209_ _209_/A _192_/X vssd vccd mgmt_gpio_in vssd vccd sky130_fd_sc_hd__ebufn_8
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_173_ _173_/A vssd vccd _174_/A vssd vccd sky130_fd_sc_hd__buf_1
XPHY_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_190_ _190_/A vssd vccd _190_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput19 user_gpio_oeb vssd vccd _205_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
X_225_ _231_/CLK _225_/D _202_/A vssd vccd _226_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_156_ _169_/A _159_/B vssd vccd _157_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold8 hold8/A vssd vccd hold8/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_208_ _208_/A0 _207_/X _210_/Q vssd vccd _208_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_139_ _139_/A vssd vccd _139_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_172_ _172_/A vssd vccd _172_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_224_ _231_/CLK _224_/D _202_/A vssd vccd _225_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_155_ _155_/A vssd vccd _155_/X vssd vccd sky130_fd_sc_hd__buf_1
X_207_ _207_/A0 _206_/X _207_/S vssd vccd _207_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_138_ _152_/A _138_/B vssd vccd _139_/A vssd vccd sky130_fd_sc_hd__or2_1
Xhold9 hold9/A vssd vccd hold9/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_171_ _183_/A _171_/B vssd vccd _172_/A vssd vccd sky130_fd_sc_hd__or2_1
XPHY_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_223_ _203_/A _223_/D _202_/A vssd vccd _224_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_154_ _173_/A vssd vccd _155_/A vssd vccd sky130_fd_sc_hd__buf_1
X_206_ _206_/A0 _207_/A0 _206_/S vssd vccd _206_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_137_ _137_/A vssd vccd _137_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_170_ _170_/A vssd vccd _170_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_153_ _153_/A vssd vccd _153_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_205_ _205_/A0 _194_/X _210_/Q vssd vccd _205_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_222_ _201_/X _222_/D _114_/X _111_/X vssd vccd _222_/Q _222_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_136_ _136_/A _138_/B vssd vccd _137_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_119_ _187_/A _119_/B vssd vccd _120_/A vssd vccd sky130_fd_sc_hd__or2_1
XPHY_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_0 mgmt_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_152_ _152_/A _152_/B vssd vccd _153_/A vssd vccd sky130_fd_sc_hd__or2_1
X_221_ _140_/A _221_/D _120_/X _118_/X vssd vccd _221_/Q _221_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_204_ serial_load vssd vccd _204_/X vssd vccd sky130_fd_sc_hd__buf_2
X_118_ _118_/A vssd vccd _118_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_135_ _135_/A vssd vccd _135_/X vssd vccd sky130_fd_sc_hd__buf_1
XPHY_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1 mgmt_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_203_ _203_/A vssd vccd _203_/X vssd vccd sky130_fd_sc_hd__buf_2
X_151_ _151_/A vssd vccd _151_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_134_ _140_/A vssd vccd _135_/A vssd vccd sky130_fd_sc_hd__buf_1
X_220_ _122_/X hold9/X _127_/X _124_/X vssd vccd _220_/Q _220_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_117_ _136_/A _119_/B vssd vccd _118_/A vssd vccd sky130_fd_sc_hd__or2b_1
XPHY_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2 one vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_150_ _169_/A _152_/B vssd vccd _151_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_133_ _133_/A vssd vccd _133_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_202_ _202_/A vssd vccd _202_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_116_ _116_/A vssd vccd _140_/A vssd vccd sky130_fd_sc_hd__buf_1
XANTENNA_3 one vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_132_ _152_/A _132_/B vssd vccd _133_/A vssd vccd sky130_fd_sc_hd__or2_1
X_201_ _201_/A vssd vccd _201_/X vssd vccd sky130_fd_sc_hd__buf_1
Xoutput30 _208_/X vssd vccd pad_gpio_out vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_4 pad_gpio_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
.ends

