magic
tech sky130A
magscale 1 2
timestamp 1636033645
<< viali >>
rect 1041 1853 1075 1887
<< metal1 >>
rect 0 2746 1380 2768
rect 0 2694 78 2746
rect 130 2694 142 2746
rect 194 2694 206 2746
rect 258 2694 270 2746
rect 322 2694 1380 2746
rect 0 2672 1380 2694
rect 0 2202 1380 2224
rect 0 2150 818 2202
rect 870 2150 882 2202
rect 934 2150 946 2202
rect 998 2150 1010 2202
rect 1062 2150 1380 2202
rect 0 2128 1380 2150
rect 474 1844 480 1896
rect 532 1884 538 1896
rect 1029 1887 1087 1893
rect 1029 1884 1041 1887
rect 532 1856 1041 1884
rect 532 1844 538 1856
rect 1029 1853 1041 1856
rect 1075 1853 1087 1887
rect 1029 1847 1087 1853
rect 0 1658 1380 1680
rect 0 1606 78 1658
rect 130 1606 142 1658
rect 194 1606 206 1658
rect 258 1606 270 1658
rect 322 1606 1380 1658
rect 0 1584 1380 1606
rect 0 1114 1380 1136
rect 0 1062 818 1114
rect 870 1062 882 1114
rect 934 1062 946 1114
rect 998 1062 1010 1114
rect 1062 1062 1380 1114
rect 0 1040 1380 1062
rect 0 570 1380 592
rect 0 518 78 570
rect 130 518 142 570
rect 194 518 206 570
rect 258 518 270 570
rect 322 518 1380 570
rect 0 496 1380 518
rect 0 26 1380 48
rect 0 -26 818 26
rect 870 -26 882 26
rect 934 -26 946 26
rect 998 -26 1010 26
rect 1062 -26 1380 26
rect 0 -48 1380 -26
<< via1 >>
rect 78 2694 130 2746
rect 142 2694 194 2746
rect 206 2694 258 2746
rect 270 2694 322 2746
rect 818 2150 870 2202
rect 882 2150 934 2202
rect 946 2150 998 2202
rect 1010 2150 1062 2202
rect 480 1844 532 1896
rect 78 1606 130 1658
rect 142 1606 194 1658
rect 206 1606 258 1658
rect 270 1606 322 1658
rect 818 1062 870 1114
rect 882 1062 934 1114
rect 946 1062 998 1114
rect 1010 1062 1062 1114
rect 78 518 130 570
rect 142 518 194 570
rect 206 518 258 570
rect 270 518 322 570
rect 818 -26 870 26
rect 882 -26 934 26
rect 946 -26 998 26
rect 1010 -26 1062 26
<< metal2 >>
rect 78 2748 322 2768
rect 78 2746 92 2748
rect 148 2746 172 2748
rect 228 2746 252 2748
rect 308 2746 322 2748
rect 78 2692 92 2694
rect 148 2692 172 2694
rect 228 2692 252 2694
rect 308 2692 322 2694
rect 78 2672 322 2692
rect 818 2204 1062 2224
rect 818 2202 832 2204
rect 888 2202 912 2204
rect 968 2202 992 2204
rect 1048 2202 1062 2204
rect 818 2148 832 2150
rect 888 2148 912 2150
rect 968 2148 992 2150
rect 1048 2148 1062 2150
rect 818 2128 1062 2148
rect 480 1896 532 1902
rect 480 1838 532 1844
rect 492 1737 520 1838
rect 478 1728 534 1737
rect 78 1660 322 1680
rect 478 1663 534 1672
rect 78 1658 92 1660
rect 148 1658 172 1660
rect 228 1658 252 1660
rect 308 1658 322 1660
rect 78 1604 92 1606
rect 148 1604 172 1606
rect 228 1604 252 1606
rect 308 1604 322 1606
rect 78 1584 322 1604
rect 818 1116 1062 1136
rect 818 1114 832 1116
rect 888 1114 912 1116
rect 968 1114 992 1116
rect 1048 1114 1062 1116
rect 818 1060 832 1062
rect 888 1060 912 1062
rect 968 1060 992 1062
rect 1048 1060 1062 1062
rect 818 1040 1062 1060
rect 78 572 322 592
rect 78 570 92 572
rect 148 570 172 572
rect 228 570 252 572
rect 308 570 322 572
rect 78 516 92 518
rect 148 516 172 518
rect 228 516 252 518
rect 308 516 322 518
rect 78 496 322 516
rect 818 28 1062 48
rect 818 26 832 28
rect 888 26 912 28
rect 968 26 992 28
rect 1048 26 1062 28
rect 818 -28 832 -26
rect 888 -28 912 -26
rect 968 -28 992 -26
rect 1048 -28 1062 -26
rect 818 -48 1062 -28
<< via2 >>
rect 92 2746 148 2748
rect 172 2746 228 2748
rect 252 2746 308 2748
rect 92 2694 130 2746
rect 130 2694 142 2746
rect 142 2694 148 2746
rect 172 2694 194 2746
rect 194 2694 206 2746
rect 206 2694 228 2746
rect 252 2694 258 2746
rect 258 2694 270 2746
rect 270 2694 308 2746
rect 92 2692 148 2694
rect 172 2692 228 2694
rect 252 2692 308 2694
rect 832 2202 888 2204
rect 912 2202 968 2204
rect 992 2202 1048 2204
rect 832 2150 870 2202
rect 870 2150 882 2202
rect 882 2150 888 2202
rect 912 2150 934 2202
rect 934 2150 946 2202
rect 946 2150 968 2202
rect 992 2150 998 2202
rect 998 2150 1010 2202
rect 1010 2150 1048 2202
rect 832 2148 888 2150
rect 912 2148 968 2150
rect 992 2148 1048 2150
rect 478 1672 534 1728
rect 92 1658 148 1660
rect 172 1658 228 1660
rect 252 1658 308 1660
rect 92 1606 130 1658
rect 130 1606 142 1658
rect 142 1606 148 1658
rect 172 1606 194 1658
rect 194 1606 206 1658
rect 206 1606 228 1658
rect 252 1606 258 1658
rect 258 1606 270 1658
rect 270 1606 308 1658
rect 92 1604 148 1606
rect 172 1604 228 1606
rect 252 1604 308 1606
rect 832 1114 888 1116
rect 912 1114 968 1116
rect 992 1114 1048 1116
rect 832 1062 870 1114
rect 870 1062 882 1114
rect 882 1062 888 1114
rect 912 1062 934 1114
rect 934 1062 946 1114
rect 946 1062 968 1114
rect 992 1062 998 1114
rect 998 1062 1010 1114
rect 1010 1062 1048 1114
rect 832 1060 888 1062
rect 912 1060 968 1062
rect 992 1060 1048 1062
rect 92 570 148 572
rect 172 570 228 572
rect 252 570 308 572
rect 92 518 130 570
rect 130 518 142 570
rect 142 518 148 570
rect 172 518 194 570
rect 194 518 206 570
rect 206 518 228 570
rect 252 518 258 570
rect 258 518 270 570
rect 270 518 308 570
rect 92 516 148 518
rect 172 516 228 518
rect 252 516 308 518
rect 832 26 888 28
rect 912 26 968 28
rect 992 26 1048 28
rect 832 -26 870 26
rect 870 -26 882 26
rect 882 -26 888 26
rect 912 -26 934 26
rect 934 -26 946 26
rect 946 -26 968 26
rect 992 -26 998 26
rect 998 -26 1010 26
rect 1010 -26 1048 26
rect 832 -28 888 -26
rect 912 -28 968 -26
rect 992 -28 1048 -26
<< metal3 >>
rect 60 2752 340 2753
rect 60 2688 88 2752
rect 152 2688 168 2752
rect 232 2688 248 2752
rect 312 2688 340 2752
rect 60 2687 340 2688
rect 800 2208 1080 2209
rect 800 2144 828 2208
rect 892 2144 908 2208
rect 972 2144 988 2208
rect 1052 2144 1080 2208
rect 800 2143 1080 2144
rect 473 1730 539 1733
rect 600 1730 1400 1760
rect 473 1728 1400 1730
rect 473 1672 478 1728
rect 534 1672 1400 1728
rect 473 1670 1400 1672
rect 473 1667 539 1670
rect 60 1664 340 1665
rect 60 1600 88 1664
rect 152 1600 168 1664
rect 232 1600 248 1664
rect 312 1600 340 1664
rect 600 1640 1400 1670
rect 60 1599 340 1600
rect 800 1120 1080 1121
rect 800 1056 828 1120
rect 892 1056 908 1120
rect 972 1056 988 1120
rect 1052 1056 1080 1120
rect 800 1055 1080 1056
rect 60 576 340 577
rect 60 512 88 576
rect 152 512 168 576
rect 232 512 248 576
rect 312 512 340 576
rect 60 511 340 512
rect 800 32 1080 33
rect 800 -32 828 32
rect 892 -32 908 32
rect 972 -32 988 32
rect 1052 -32 1080 32
rect 800 -33 1080 -32
<< via3 >>
rect 88 2748 152 2752
rect 88 2692 92 2748
rect 92 2692 148 2748
rect 148 2692 152 2748
rect 88 2688 152 2692
rect 168 2748 232 2752
rect 168 2692 172 2748
rect 172 2692 228 2748
rect 228 2692 232 2748
rect 168 2688 232 2692
rect 248 2748 312 2752
rect 248 2692 252 2748
rect 252 2692 308 2748
rect 308 2692 312 2748
rect 248 2688 312 2692
rect 828 2204 892 2208
rect 828 2148 832 2204
rect 832 2148 888 2204
rect 888 2148 892 2204
rect 828 2144 892 2148
rect 908 2204 972 2208
rect 908 2148 912 2204
rect 912 2148 968 2204
rect 968 2148 972 2204
rect 908 2144 972 2148
rect 988 2204 1052 2208
rect 988 2148 992 2204
rect 992 2148 1048 2204
rect 1048 2148 1052 2204
rect 988 2144 1052 2148
rect 88 1660 152 1664
rect 88 1604 92 1660
rect 92 1604 148 1660
rect 148 1604 152 1660
rect 88 1600 152 1604
rect 168 1660 232 1664
rect 168 1604 172 1660
rect 172 1604 228 1660
rect 228 1604 232 1660
rect 168 1600 232 1604
rect 248 1660 312 1664
rect 248 1604 252 1660
rect 252 1604 308 1660
rect 308 1604 312 1660
rect 248 1600 312 1604
rect 828 1116 892 1120
rect 828 1060 832 1116
rect 832 1060 888 1116
rect 888 1060 892 1116
rect 828 1056 892 1060
rect 908 1116 972 1120
rect 908 1060 912 1116
rect 912 1060 968 1116
rect 968 1060 972 1116
rect 908 1056 972 1060
rect 988 1116 1052 1120
rect 988 1060 992 1116
rect 992 1060 1048 1116
rect 1048 1060 1052 1116
rect 988 1056 1052 1060
rect 88 572 152 576
rect 88 516 92 572
rect 92 516 148 572
rect 148 516 152 572
rect 88 512 152 516
rect 168 572 232 576
rect 168 516 172 572
rect 172 516 228 572
rect 228 516 232 572
rect 168 512 232 516
rect 248 572 312 576
rect 248 516 252 572
rect 252 516 308 572
rect 308 516 312 572
rect 248 512 312 516
rect 828 28 892 32
rect 828 -28 832 28
rect 832 -28 888 28
rect 888 -28 892 28
rect 828 -32 892 -28
rect 908 28 972 32
rect 908 -28 912 28
rect 912 -28 968 28
rect 968 -28 972 28
rect 908 -32 972 -28
rect 988 28 1052 32
rect 988 -28 992 28
rect 992 -28 1048 28
rect 1048 -28 1052 28
rect 988 -32 1052 -28
<< metal4 >>
rect 60 2752 340 2768
rect 60 2688 88 2752
rect 152 2688 168 2752
rect 232 2688 248 2752
rect 312 2688 340 2752
rect 60 1664 340 2688
rect 60 1600 88 1664
rect 152 1600 168 1664
rect 232 1600 248 1664
rect 312 1600 340 1664
rect 60 576 340 1600
rect 60 512 88 576
rect 152 512 168 576
rect 232 512 248 576
rect 312 512 340 576
rect 60 -48 340 512
rect 800 2208 1080 2768
rect 800 2144 828 2208
rect 892 2144 908 2208
rect 972 2144 988 2208
rect 1052 2144 1080 2208
rect 800 1120 1080 2144
rect 800 1056 828 1120
rect 892 1056 908 1120
rect 972 1056 988 1120
rect 1052 1056 1080 1120
rect 800 32 1080 1056
rect 800 -32 828 32
rect 892 -32 908 32
rect 972 -32 988 32
rect 1052 -32 1080 32
rect 800 -48 1080 -32
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635271187
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 644 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 276 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 736 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 1380 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 1380 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1635271187
transform 1 0 1012 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp 1635271187
transform 1 0 828 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 276 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1635271187
transform 1 0 276 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1635271187
transform 1 0 644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp 1635271187
transform 1 0 828 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635271187
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_11
timestamp 1635271187
transform 1 0 736 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 276 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1635271187
transform 1 0 276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1635271187
transform 1 0 644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp 1635271187
transform 1 0 828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1635271187
transform 1 0 736 0 1 2176
box -38 -48 130 592
<< labels >>
rlabel metal3 s 600 1640 1400 1760 6 gpio_logic1
port 0 nsew signal tristate
rlabel metal4 s 60 -48 340 2768 6 vccd1
port 1 nsew power input
rlabel metal4 s 800 -48 1080 2768 6 vssd1
port 2 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 1400 3200
<< end >>
