* NGSPICE file created from gpio_defaults_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

.subckt gpio_defaults_block VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
Xgpio_default_value\[8\] VGND VGND VPWR VPWR gpio_default_value\[8\]/HI gpio_defaults[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgpio_default_value\[6\] VGND VGND VPWR VPWR gpio_default_value\[6\]/HI gpio_defaults[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[4\] VGND VGND VPWR VPWR gpio_default_value\[4\]/HI gpio_defaults[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[2\] VGND VGND VPWR VPWR gpio_default_value\[2\]/HI gpio_defaults[2]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[12\] VGND VGND VPWR VPWR gpio_default_value\[12\]/HI gpio_defaults[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgpio_default_value\[0\] VGND VGND VPWR VPWR gpio_default_value\[0\]/HI gpio_defaults[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[10\] VGND VGND VPWR VPWR gpio_defaults[10] gpio_default_value\[10\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[9\] VGND VGND VPWR VPWR gpio_default_value\[9\]/HI gpio_defaults[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgpio_default_value\[7\] VGND VGND VPWR VPWR gpio_default_value\[7\]/HI gpio_defaults[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_default_value\[5\] VGND VGND VPWR VPWR gpio_default_value\[5\]/HI gpio_defaults[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgpio_default_value\[3\] VGND VGND VPWR VPWR gpio_default_value\[3\]/HI gpio_defaults[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[1\] VGND VGND VPWR VPWR gpio_defaults[1] gpio_default_value\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[11\] VGND VGND VPWR VPWR gpio_default_value\[11\]/HI gpio_defaults[11]
+ sky130_fd_sc_hd__conb_1
.ends

