magic
tech sky130A
magscale 1 2
timestamp 1637412622
<< obsli1 >>
rect 1104 2159 58880 107729
<< obsm1 >>
rect 14 2128 60044 107976
<< metal2 >>
rect 202 109390 258 110190
rect 662 109390 718 110190
rect 1122 109390 1178 110190
rect 1582 109390 1638 110190
rect 2042 109390 2098 110190
rect 2502 109390 2558 110190
rect 2962 109390 3018 110190
rect 3422 109390 3478 110190
rect 3882 109390 3938 110190
rect 4342 109390 4398 110190
rect 4802 109390 4858 110190
rect 5262 109390 5318 110190
rect 5722 109390 5778 110190
rect 6182 109390 6238 110190
rect 6642 109390 6698 110190
rect 7102 109390 7158 110190
rect 7562 109390 7618 110190
rect 8114 109390 8170 110190
rect 8574 109390 8630 110190
rect 9034 109390 9090 110190
rect 9494 109390 9550 110190
rect 9954 109390 10010 110190
rect 10414 109390 10470 110190
rect 10874 109390 10930 110190
rect 11334 109390 11390 110190
rect 11794 109390 11850 110190
rect 12254 109390 12310 110190
rect 12714 109390 12770 110190
rect 13174 109390 13230 110190
rect 13634 109390 13690 110190
rect 14094 109390 14150 110190
rect 14554 109390 14610 110190
rect 15014 109390 15070 110190
rect 15566 109390 15622 110190
rect 16026 109390 16082 110190
rect 16486 109390 16542 110190
rect 16946 109390 17002 110190
rect 17406 109390 17462 110190
rect 17866 109390 17922 110190
rect 18326 109390 18382 110190
rect 18786 109390 18842 110190
rect 19246 109390 19302 110190
rect 19706 109390 19762 110190
rect 20166 109390 20222 110190
rect 20626 109390 20682 110190
rect 21086 109390 21142 110190
rect 21546 109390 21602 110190
rect 22006 109390 22062 110190
rect 22466 109390 22522 110190
rect 23018 109390 23074 110190
rect 23478 109390 23534 110190
rect 23938 109390 23994 110190
rect 24398 109390 24454 110190
rect 24858 109390 24914 110190
rect 25318 109390 25374 110190
rect 25778 109390 25834 110190
rect 26238 109390 26294 110190
rect 26698 109390 26754 110190
rect 27158 109390 27214 110190
rect 27618 109390 27674 110190
rect 28078 109390 28134 110190
rect 28538 109390 28594 110190
rect 28998 109390 29054 110190
rect 29458 109390 29514 110190
rect 29918 109390 29974 110190
rect 30470 109390 30526 110190
rect 30930 109390 30986 110190
rect 31390 109390 31446 110190
rect 31850 109390 31906 110190
rect 32310 109390 32366 110190
rect 32770 109390 32826 110190
rect 33230 109390 33286 110190
rect 33690 109390 33746 110190
rect 34150 109390 34206 110190
rect 34610 109390 34666 110190
rect 35070 109390 35126 110190
rect 35530 109390 35586 110190
rect 35990 109390 36046 110190
rect 36450 109390 36506 110190
rect 36910 109390 36966 110190
rect 37370 109390 37426 110190
rect 37922 109390 37978 110190
rect 38382 109390 38438 110190
rect 38842 109390 38898 110190
rect 39302 109390 39358 110190
rect 39762 109390 39818 110190
rect 40222 109390 40278 110190
rect 40682 109390 40738 110190
rect 41142 109390 41198 110190
rect 41602 109390 41658 110190
rect 42062 109390 42118 110190
rect 42522 109390 42578 110190
rect 42982 109390 43038 110190
rect 43442 109390 43498 110190
rect 43902 109390 43958 110190
rect 44362 109390 44418 110190
rect 44822 109390 44878 110190
rect 45374 109390 45430 110190
rect 45834 109390 45890 110190
rect 46294 109390 46350 110190
rect 46754 109390 46810 110190
rect 47214 109390 47270 110190
rect 47674 109390 47730 110190
rect 48134 109390 48190 110190
rect 48594 109390 48650 110190
rect 49054 109390 49110 110190
rect 49514 109390 49570 110190
rect 49974 109390 50030 110190
rect 50434 109390 50490 110190
rect 50894 109390 50950 110190
rect 51354 109390 51410 110190
rect 51814 109390 51870 110190
rect 52274 109390 52330 110190
rect 52826 109390 52882 110190
rect 53286 109390 53342 110190
rect 53746 109390 53802 110190
rect 54206 109390 54262 110190
rect 54666 109390 54722 110190
rect 55126 109390 55182 110190
rect 55586 109390 55642 110190
rect 56046 109390 56102 110190
rect 56506 109390 56562 110190
rect 56966 109390 57022 110190
rect 57426 109390 57482 110190
rect 57886 109390 57942 110190
rect 58346 109390 58402 110190
rect 58806 109390 58862 110190
rect 59266 109390 59322 110190
rect 59726 109390 59782 110190
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2226 0 2282 800
rect 2870 0 2926 800
rect 3514 0 3570 800
rect 4158 0 4214 800
rect 4802 0 4858 800
rect 5446 0 5502 800
rect 6090 0 6146 800
rect 6734 0 6790 800
rect 7470 0 7526 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9402 0 9458 800
rect 10046 0 10102 800
rect 10690 0 10746 800
rect 11334 0 11390 800
rect 11978 0 12034 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14646 0 14702 800
rect 15290 0 15346 800
rect 15934 0 15990 800
rect 16578 0 16634 800
rect 17222 0 17278 800
rect 17866 0 17922 800
rect 18510 0 18566 800
rect 19154 0 19210 800
rect 19798 0 19854 800
rect 20534 0 20590 800
rect 21178 0 21234 800
rect 21822 0 21878 800
rect 22466 0 22522 800
rect 23110 0 23166 800
rect 23754 0 23810 800
rect 24398 0 24454 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34242 0 34298 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36174 0 36230 800
rect 36818 0 36874 800
rect 37462 0 37518 800
rect 38106 0 38162 800
rect 38750 0 38806 800
rect 39394 0 39450 800
rect 40038 0 40094 800
rect 40774 0 40830 800
rect 41418 0 41474 800
rect 42062 0 42118 800
rect 42706 0 42762 800
rect 43350 0 43406 800
rect 43994 0 44050 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46570 0 46626 800
rect 47306 0 47362 800
rect 47950 0 48006 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53838 0 53894 800
rect 54482 0 54538 800
rect 55126 0 55182 800
rect 55770 0 55826 800
rect 56414 0 56470 800
rect 57058 0 57114 800
rect 57702 0 57758 800
rect 58346 0 58402 800
rect 58990 0 59046 800
rect 59634 0 59690 800
<< obsm2 >>
rect 20 109334 146 109426
rect 314 109334 606 109426
rect 774 109334 1066 109426
rect 1234 109334 1526 109426
rect 1694 109334 1986 109426
rect 2154 109334 2446 109426
rect 2614 109334 2906 109426
rect 3074 109334 3366 109426
rect 3534 109334 3826 109426
rect 3994 109334 4286 109426
rect 4454 109334 4746 109426
rect 4914 109334 5206 109426
rect 5374 109334 5666 109426
rect 5834 109334 6126 109426
rect 6294 109334 6586 109426
rect 6754 109334 7046 109426
rect 7214 109334 7506 109426
rect 7674 109334 8058 109426
rect 8226 109334 8518 109426
rect 8686 109334 8978 109426
rect 9146 109334 9438 109426
rect 9606 109334 9898 109426
rect 10066 109334 10358 109426
rect 10526 109334 10818 109426
rect 10986 109334 11278 109426
rect 11446 109334 11738 109426
rect 11906 109334 12198 109426
rect 12366 109334 12658 109426
rect 12826 109334 13118 109426
rect 13286 109334 13578 109426
rect 13746 109334 14038 109426
rect 14206 109334 14498 109426
rect 14666 109334 14958 109426
rect 15126 109334 15510 109426
rect 15678 109334 15970 109426
rect 16138 109334 16430 109426
rect 16598 109334 16890 109426
rect 17058 109334 17350 109426
rect 17518 109334 17810 109426
rect 17978 109334 18270 109426
rect 18438 109334 18730 109426
rect 18898 109334 19190 109426
rect 19358 109334 19650 109426
rect 19818 109334 20110 109426
rect 20278 109334 20570 109426
rect 20738 109334 21030 109426
rect 21198 109334 21490 109426
rect 21658 109334 21950 109426
rect 22118 109334 22410 109426
rect 22578 109334 22962 109426
rect 23130 109334 23422 109426
rect 23590 109334 23882 109426
rect 24050 109334 24342 109426
rect 24510 109334 24802 109426
rect 24970 109334 25262 109426
rect 25430 109334 25722 109426
rect 25890 109334 26182 109426
rect 26350 109334 26642 109426
rect 26810 109334 27102 109426
rect 27270 109334 27562 109426
rect 27730 109334 28022 109426
rect 28190 109334 28482 109426
rect 28650 109334 28942 109426
rect 29110 109334 29402 109426
rect 29570 109334 29862 109426
rect 30030 109334 30414 109426
rect 30582 109334 30874 109426
rect 31042 109334 31334 109426
rect 31502 109334 31794 109426
rect 31962 109334 32254 109426
rect 32422 109334 32714 109426
rect 32882 109334 33174 109426
rect 33342 109334 33634 109426
rect 33802 109334 34094 109426
rect 34262 109334 34554 109426
rect 34722 109334 35014 109426
rect 35182 109334 35474 109426
rect 35642 109334 35934 109426
rect 36102 109334 36394 109426
rect 36562 109334 36854 109426
rect 37022 109334 37314 109426
rect 37482 109334 37866 109426
rect 38034 109334 38326 109426
rect 38494 109334 38786 109426
rect 38954 109334 39246 109426
rect 39414 109334 39706 109426
rect 39874 109334 40166 109426
rect 40334 109334 40626 109426
rect 40794 109334 41086 109426
rect 41254 109334 41546 109426
rect 41714 109334 42006 109426
rect 42174 109334 42466 109426
rect 42634 109334 42926 109426
rect 43094 109334 43386 109426
rect 43554 109334 43846 109426
rect 44014 109334 44306 109426
rect 44474 109334 44766 109426
rect 44934 109334 45318 109426
rect 45486 109334 45778 109426
rect 45946 109334 46238 109426
rect 46406 109334 46698 109426
rect 46866 109334 47158 109426
rect 47326 109334 47618 109426
rect 47786 109334 48078 109426
rect 48246 109334 48538 109426
rect 48706 109334 48998 109426
rect 49166 109334 49458 109426
rect 49626 109334 49918 109426
rect 50086 109334 50378 109426
rect 50546 109334 50838 109426
rect 51006 109334 51298 109426
rect 51466 109334 51758 109426
rect 51926 109334 52218 109426
rect 52386 109334 52770 109426
rect 52938 109334 53230 109426
rect 53398 109334 53690 109426
rect 53858 109334 54150 109426
rect 54318 109334 54610 109426
rect 54778 109334 55070 109426
rect 55238 109334 55530 109426
rect 55698 109334 55990 109426
rect 56158 109334 56450 109426
rect 56618 109334 56910 109426
rect 57078 109334 57370 109426
rect 57538 109334 57830 109426
rect 57998 109334 58290 109426
rect 58458 109334 58750 109426
rect 58918 109334 59210 109426
rect 59378 109334 59670 109426
rect 59838 109334 60044 109426
rect 20 856 60044 109334
rect 20 800 238 856
rect 406 800 882 856
rect 1050 800 1526 856
rect 1694 800 2170 856
rect 2338 800 2814 856
rect 2982 800 3458 856
rect 3626 800 4102 856
rect 4270 800 4746 856
rect 4914 800 5390 856
rect 5558 800 6034 856
rect 6202 800 6678 856
rect 6846 800 7414 856
rect 7582 800 8058 856
rect 8226 800 8702 856
rect 8870 800 9346 856
rect 9514 800 9990 856
rect 10158 800 10634 856
rect 10802 800 11278 856
rect 11446 800 11922 856
rect 12090 800 12566 856
rect 12734 800 13210 856
rect 13378 800 13946 856
rect 14114 800 14590 856
rect 14758 800 15234 856
rect 15402 800 15878 856
rect 16046 800 16522 856
rect 16690 800 17166 856
rect 17334 800 17810 856
rect 17978 800 18454 856
rect 18622 800 19098 856
rect 19266 800 19742 856
rect 19910 800 20478 856
rect 20646 800 21122 856
rect 21290 800 21766 856
rect 21934 800 22410 856
rect 22578 800 23054 856
rect 23222 800 23698 856
rect 23866 800 24342 856
rect 24510 800 24986 856
rect 25154 800 25630 856
rect 25798 800 26274 856
rect 26442 800 27010 856
rect 27178 800 27654 856
rect 27822 800 28298 856
rect 28466 800 28942 856
rect 29110 800 29586 856
rect 29754 800 30230 856
rect 30398 800 30874 856
rect 31042 800 31518 856
rect 31686 800 32162 856
rect 32330 800 32806 856
rect 32974 800 33450 856
rect 33618 800 34186 856
rect 34354 800 34830 856
rect 34998 800 35474 856
rect 35642 800 36118 856
rect 36286 800 36762 856
rect 36930 800 37406 856
rect 37574 800 38050 856
rect 38218 800 38694 856
rect 38862 800 39338 856
rect 39506 800 39982 856
rect 40150 800 40718 856
rect 40886 800 41362 856
rect 41530 800 42006 856
rect 42174 800 42650 856
rect 42818 800 43294 856
rect 43462 800 43938 856
rect 44106 800 44582 856
rect 44750 800 45226 856
rect 45394 800 45870 856
rect 46038 800 46514 856
rect 46682 800 47250 856
rect 47418 800 47894 856
rect 48062 800 48538 856
rect 48706 800 49182 856
rect 49350 800 49826 856
rect 49994 800 50470 856
rect 50638 800 51114 856
rect 51282 800 51758 856
rect 51926 800 52402 856
rect 52570 800 53046 856
rect 53214 800 53782 856
rect 53950 800 54426 856
rect 54594 800 55070 856
rect 55238 800 55714 856
rect 55882 800 56358 856
rect 56526 800 57002 856
rect 57170 800 57646 856
rect 57814 800 58290 856
rect 58458 800 58934 856
rect 59102 800 59578 856
rect 59746 800 60044 856
<< metal3 >>
rect 0 109488 800 109608
rect 59246 109216 60046 109336
rect 0 108536 800 108656
rect 0 107448 800 107568
rect 59246 107584 60046 107704
rect 0 106496 800 106616
rect 59246 105816 60046 105936
rect 0 105408 800 105528
rect 0 104456 800 104576
rect 59246 104184 60046 104304
rect 0 103368 800 103488
rect 0 102416 800 102536
rect 59246 102416 60046 102536
rect 0 101328 800 101448
rect 59246 100784 60046 100904
rect 0 100376 800 100496
rect 0 99288 800 99408
rect 59246 99016 60046 99136
rect 0 98336 800 98456
rect 0 97248 800 97368
rect 59246 97384 60046 97504
rect 0 96296 800 96416
rect 59246 95616 60046 95736
rect 0 95208 800 95328
rect 0 94256 800 94376
rect 59246 93984 60046 94104
rect 0 93168 800 93288
rect 0 92216 800 92336
rect 59246 92216 60046 92336
rect 0 91128 800 91248
rect 59246 90584 60046 90704
rect 0 90176 800 90296
rect 0 89088 800 89208
rect 59246 88952 60046 89072
rect 0 88136 800 88256
rect 0 87048 800 87168
rect 59246 87184 60046 87304
rect 0 86096 800 86216
rect 59246 85552 60046 85672
rect 0 85008 800 85128
rect 0 84056 800 84176
rect 59246 83784 60046 83904
rect 0 82968 800 83088
rect 0 82016 800 82136
rect 59246 82152 60046 82272
rect 0 80928 800 81048
rect 59246 80384 60046 80504
rect 0 79976 800 80096
rect 0 78888 800 79008
rect 59246 78752 60046 78872
rect 0 77936 800 78056
rect 0 76848 800 76968
rect 59246 76984 60046 77104
rect 0 75896 800 76016
rect 59246 75352 60046 75472
rect 0 74808 800 74928
rect 0 73856 800 73976
rect 59246 73584 60046 73704
rect 0 72768 800 72888
rect 0 71816 800 71936
rect 59246 71952 60046 72072
rect 0 70728 800 70848
rect 59246 70184 60046 70304
rect 0 69776 800 69896
rect 0 68688 800 68808
rect 59246 68552 60046 68672
rect 0 67736 800 67856
rect 59246 66920 60046 67040
rect 0 66648 800 66768
rect 0 65696 800 65816
rect 59246 65152 60046 65272
rect 0 64608 800 64728
rect 0 63656 800 63776
rect 59246 63520 60046 63640
rect 0 62568 800 62688
rect 0 61616 800 61736
rect 59246 61752 60046 61872
rect 0 60528 800 60648
rect 59246 60120 60046 60240
rect 0 59576 800 59696
rect 0 58488 800 58608
rect 59246 58352 60046 58472
rect 0 57536 800 57656
rect 59246 56720 60046 56840
rect 0 56448 800 56568
rect 0 55496 800 55616
rect 59246 54952 60046 55072
rect 0 54408 800 54528
rect 0 53456 800 53576
rect 59246 53320 60046 53440
rect 0 52368 800 52488
rect 0 51416 800 51536
rect 59246 51552 60046 51672
rect 0 50328 800 50448
rect 59246 49920 60046 50040
rect 0 49376 800 49496
rect 0 48288 800 48408
rect 59246 48152 60046 48272
rect 0 47336 800 47456
rect 59246 46520 60046 46640
rect 0 46248 800 46368
rect 0 45296 800 45416
rect 59246 44888 60046 45008
rect 0 44208 800 44328
rect 0 43256 800 43376
rect 59246 43120 60046 43240
rect 0 42168 800 42288
rect 59246 41488 60046 41608
rect 0 41216 800 41336
rect 0 40128 800 40248
rect 59246 39720 60046 39840
rect 0 39176 800 39296
rect 0 38088 800 38208
rect 59246 38088 60046 38208
rect 0 37136 800 37256
rect 59246 36320 60046 36440
rect 0 36048 800 36168
rect 0 35096 800 35216
rect 59246 34688 60046 34808
rect 0 34008 800 34128
rect 0 33056 800 33176
rect 59246 32920 60046 33040
rect 0 31968 800 32088
rect 59246 31288 60046 31408
rect 0 31016 800 31136
rect 0 29928 800 30048
rect 59246 29520 60046 29640
rect 0 28976 800 29096
rect 0 27888 800 28008
rect 59246 27888 60046 28008
rect 0 26936 800 27056
rect 59246 26120 60046 26240
rect 0 25848 800 25968
rect 0 24896 800 25016
rect 59246 24488 60046 24608
rect 0 23808 800 23928
rect 0 22856 800 22976
rect 59246 22856 60046 22976
rect 0 21768 800 21888
rect 59246 21088 60046 21208
rect 0 20816 800 20936
rect 0 19728 800 19848
rect 59246 19456 60046 19576
rect 0 18776 800 18896
rect 0 17688 800 17808
rect 59246 17688 60046 17808
rect 0 16736 800 16856
rect 59246 16056 60046 16176
rect 0 15648 800 15768
rect 0 14696 800 14816
rect 59246 14288 60046 14408
rect 0 13608 800 13728
rect 0 12656 800 12776
rect 59246 12656 60046 12776
rect 0 11568 800 11688
rect 59246 10888 60046 11008
rect 0 10616 800 10736
rect 0 9528 800 9648
rect 59246 9256 60046 9376
rect 0 8576 800 8696
rect 0 7488 800 7608
rect 59246 7488 60046 7608
rect 0 6536 800 6656
rect 59246 5856 60046 5976
rect 0 5448 800 5568
rect 0 4496 800 4616
rect 59246 4088 60046 4208
rect 0 3408 800 3528
rect 0 2456 800 2576
rect 59246 2456 60046 2576
rect 0 1368 800 1488
rect 59246 824 60046 944
rect 0 416 800 536
<< obsm3 >>
rect 880 109416 60016 109578
rect 880 109408 59166 109416
rect 381 109136 59166 109408
rect 381 108736 60016 109136
rect 880 108456 60016 108736
rect 381 107784 60016 108456
rect 381 107648 59166 107784
rect 880 107504 59166 107648
rect 880 107368 60016 107504
rect 381 106696 60016 107368
rect 880 106416 60016 106696
rect 381 106016 60016 106416
rect 381 105736 59166 106016
rect 381 105608 60016 105736
rect 880 105328 60016 105608
rect 381 104656 60016 105328
rect 880 104384 60016 104656
rect 880 104376 59166 104384
rect 381 104104 59166 104376
rect 381 103568 60016 104104
rect 880 103288 60016 103568
rect 381 102616 60016 103288
rect 880 102336 59166 102616
rect 381 101528 60016 102336
rect 880 101248 60016 101528
rect 381 100984 60016 101248
rect 381 100704 59166 100984
rect 381 100576 60016 100704
rect 880 100296 60016 100576
rect 381 99488 60016 100296
rect 880 99216 60016 99488
rect 880 99208 59166 99216
rect 381 98936 59166 99208
rect 381 98536 60016 98936
rect 880 98256 60016 98536
rect 381 97584 60016 98256
rect 381 97448 59166 97584
rect 880 97304 59166 97448
rect 880 97168 60016 97304
rect 381 96496 60016 97168
rect 880 96216 60016 96496
rect 381 95816 60016 96216
rect 381 95536 59166 95816
rect 381 95408 60016 95536
rect 880 95128 60016 95408
rect 381 94456 60016 95128
rect 880 94184 60016 94456
rect 880 94176 59166 94184
rect 381 93904 59166 94176
rect 381 93368 60016 93904
rect 880 93088 60016 93368
rect 381 92416 60016 93088
rect 880 92136 59166 92416
rect 381 91328 60016 92136
rect 880 91048 60016 91328
rect 381 90784 60016 91048
rect 381 90504 59166 90784
rect 381 90376 60016 90504
rect 880 90096 60016 90376
rect 381 89288 60016 90096
rect 880 89152 60016 89288
rect 880 89008 59166 89152
rect 381 88872 59166 89008
rect 381 88336 60016 88872
rect 880 88056 60016 88336
rect 381 87384 60016 88056
rect 381 87248 59166 87384
rect 880 87104 59166 87248
rect 880 86968 60016 87104
rect 381 86296 60016 86968
rect 880 86016 60016 86296
rect 381 85752 60016 86016
rect 381 85472 59166 85752
rect 381 85208 60016 85472
rect 880 84928 60016 85208
rect 381 84256 60016 84928
rect 880 83984 60016 84256
rect 880 83976 59166 83984
rect 381 83704 59166 83976
rect 381 83168 60016 83704
rect 880 82888 60016 83168
rect 381 82352 60016 82888
rect 381 82216 59166 82352
rect 880 82072 59166 82216
rect 880 81936 60016 82072
rect 381 81128 60016 81936
rect 880 80848 60016 81128
rect 381 80584 60016 80848
rect 381 80304 59166 80584
rect 381 80176 60016 80304
rect 880 79896 60016 80176
rect 381 79088 60016 79896
rect 880 78952 60016 79088
rect 880 78808 59166 78952
rect 381 78672 59166 78808
rect 381 78136 60016 78672
rect 880 77856 60016 78136
rect 381 77184 60016 77856
rect 381 77048 59166 77184
rect 880 76904 59166 77048
rect 880 76768 60016 76904
rect 381 76096 60016 76768
rect 880 75816 60016 76096
rect 381 75552 60016 75816
rect 381 75272 59166 75552
rect 381 75008 60016 75272
rect 880 74728 60016 75008
rect 381 74056 60016 74728
rect 880 73784 60016 74056
rect 880 73776 59166 73784
rect 381 73504 59166 73776
rect 381 72968 60016 73504
rect 880 72688 60016 72968
rect 381 72152 60016 72688
rect 381 72016 59166 72152
rect 880 71872 59166 72016
rect 880 71736 60016 71872
rect 381 70928 60016 71736
rect 880 70648 60016 70928
rect 381 70384 60016 70648
rect 381 70104 59166 70384
rect 381 69976 60016 70104
rect 880 69696 60016 69976
rect 381 68888 60016 69696
rect 880 68752 60016 68888
rect 880 68608 59166 68752
rect 381 68472 59166 68608
rect 381 67936 60016 68472
rect 880 67656 60016 67936
rect 381 67120 60016 67656
rect 381 66848 59166 67120
rect 880 66840 59166 66848
rect 880 66568 60016 66840
rect 381 65896 60016 66568
rect 880 65616 60016 65896
rect 381 65352 60016 65616
rect 381 65072 59166 65352
rect 381 64808 60016 65072
rect 880 64528 60016 64808
rect 381 63856 60016 64528
rect 880 63720 60016 63856
rect 880 63576 59166 63720
rect 381 63440 59166 63576
rect 381 62768 60016 63440
rect 880 62488 60016 62768
rect 381 61952 60016 62488
rect 381 61816 59166 61952
rect 880 61672 59166 61816
rect 880 61536 60016 61672
rect 381 60728 60016 61536
rect 880 60448 60016 60728
rect 381 60320 60016 60448
rect 381 60040 59166 60320
rect 381 59776 60016 60040
rect 880 59496 60016 59776
rect 381 58688 60016 59496
rect 880 58552 60016 58688
rect 880 58408 59166 58552
rect 381 58272 59166 58408
rect 381 57736 60016 58272
rect 880 57456 60016 57736
rect 381 56920 60016 57456
rect 381 56648 59166 56920
rect 880 56640 59166 56648
rect 880 56368 60016 56640
rect 381 55696 60016 56368
rect 880 55416 60016 55696
rect 381 55152 60016 55416
rect 381 54872 59166 55152
rect 381 54608 60016 54872
rect 880 54328 60016 54608
rect 381 53656 60016 54328
rect 880 53520 60016 53656
rect 880 53376 59166 53520
rect 381 53240 59166 53376
rect 381 52568 60016 53240
rect 880 52288 60016 52568
rect 381 51752 60016 52288
rect 381 51616 59166 51752
rect 880 51472 59166 51616
rect 880 51336 60016 51472
rect 381 50528 60016 51336
rect 880 50248 60016 50528
rect 381 50120 60016 50248
rect 381 49840 59166 50120
rect 381 49576 60016 49840
rect 880 49296 60016 49576
rect 381 48488 60016 49296
rect 880 48352 60016 48488
rect 880 48208 59166 48352
rect 381 48072 59166 48208
rect 381 47536 60016 48072
rect 880 47256 60016 47536
rect 381 46720 60016 47256
rect 381 46448 59166 46720
rect 880 46440 59166 46448
rect 880 46168 60016 46440
rect 381 45496 60016 46168
rect 880 45216 60016 45496
rect 381 45088 60016 45216
rect 381 44808 59166 45088
rect 381 44408 60016 44808
rect 880 44128 60016 44408
rect 381 43456 60016 44128
rect 880 43320 60016 43456
rect 880 43176 59166 43320
rect 381 43040 59166 43176
rect 381 42368 60016 43040
rect 880 42088 60016 42368
rect 381 41688 60016 42088
rect 381 41416 59166 41688
rect 880 41408 59166 41416
rect 880 41136 60016 41408
rect 381 40328 60016 41136
rect 880 40048 60016 40328
rect 381 39920 60016 40048
rect 381 39640 59166 39920
rect 381 39376 60016 39640
rect 880 39096 60016 39376
rect 381 38288 60016 39096
rect 880 38008 59166 38288
rect 381 37336 60016 38008
rect 880 37056 60016 37336
rect 381 36520 60016 37056
rect 381 36248 59166 36520
rect 880 36240 59166 36248
rect 880 35968 60016 36240
rect 381 35296 60016 35968
rect 880 35016 60016 35296
rect 381 34888 60016 35016
rect 381 34608 59166 34888
rect 381 34208 60016 34608
rect 880 33928 60016 34208
rect 381 33256 60016 33928
rect 880 33120 60016 33256
rect 880 32976 59166 33120
rect 381 32840 59166 32976
rect 381 32168 60016 32840
rect 880 31888 60016 32168
rect 381 31488 60016 31888
rect 381 31216 59166 31488
rect 880 31208 59166 31216
rect 880 30936 60016 31208
rect 381 30128 60016 30936
rect 880 29848 60016 30128
rect 381 29720 60016 29848
rect 381 29440 59166 29720
rect 381 29176 60016 29440
rect 880 28896 60016 29176
rect 381 28088 60016 28896
rect 880 27808 59166 28088
rect 381 27136 60016 27808
rect 880 26856 60016 27136
rect 381 26320 60016 26856
rect 381 26048 59166 26320
rect 880 26040 59166 26048
rect 880 25768 60016 26040
rect 381 25096 60016 25768
rect 880 24816 60016 25096
rect 381 24688 60016 24816
rect 381 24408 59166 24688
rect 381 24008 60016 24408
rect 880 23728 60016 24008
rect 381 23056 60016 23728
rect 880 22776 59166 23056
rect 381 21968 60016 22776
rect 880 21688 60016 21968
rect 381 21288 60016 21688
rect 381 21016 59166 21288
rect 880 21008 59166 21016
rect 880 20736 60016 21008
rect 381 19928 60016 20736
rect 880 19656 60016 19928
rect 880 19648 59166 19656
rect 381 19376 59166 19648
rect 381 18976 60016 19376
rect 880 18696 60016 18976
rect 381 17888 60016 18696
rect 880 17608 59166 17888
rect 381 16936 60016 17608
rect 880 16656 60016 16936
rect 381 16256 60016 16656
rect 381 15976 59166 16256
rect 381 15848 60016 15976
rect 880 15568 60016 15848
rect 381 14896 60016 15568
rect 880 14616 60016 14896
rect 381 14488 60016 14616
rect 381 14208 59166 14488
rect 381 13808 60016 14208
rect 880 13528 60016 13808
rect 381 12856 60016 13528
rect 880 12576 59166 12856
rect 381 11768 60016 12576
rect 880 11488 60016 11768
rect 381 11088 60016 11488
rect 381 10816 59166 11088
rect 880 10808 59166 10816
rect 880 10536 60016 10808
rect 381 9728 60016 10536
rect 880 9456 60016 9728
rect 880 9448 59166 9456
rect 381 9176 59166 9448
rect 381 8776 60016 9176
rect 880 8496 60016 8776
rect 381 7688 60016 8496
rect 880 7408 59166 7688
rect 381 6736 60016 7408
rect 880 6456 60016 6736
rect 381 6056 60016 6456
rect 381 5776 59166 6056
rect 381 5648 60016 5776
rect 880 5368 60016 5648
rect 381 4696 60016 5368
rect 880 4416 60016 4696
rect 381 4288 60016 4416
rect 381 4008 59166 4288
rect 381 3608 60016 4008
rect 880 3328 60016 3608
rect 381 2656 60016 3328
rect 880 2376 59166 2656
rect 381 1568 60016 2376
rect 880 1288 60016 1568
rect 381 1024 60016 1288
rect 381 744 59166 1024
rect 381 616 60016 744
rect 880 446 60016 616
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
<< obsm4 >>
rect 1163 3299 4128 106589
rect 4608 3299 19488 106589
rect 19968 3299 34848 106589
rect 35328 3299 50208 106589
rect 50688 3299 59925 106589
<< metal5 >>
rect 1104 97206 58880 97526
rect 1104 81888 58880 82208
rect 1104 66570 58880 66890
rect 1104 51252 58880 51572
rect 1104 35934 58880 36254
rect 1104 20616 58880 20936
rect 1104 5298 58880 5618
<< obsm5 >>
rect 3244 38940 28036 39260
<< labels >>
rlabel metal5 s 1104 20616 58880 20936 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 51252 58880 51572 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 81888 58880 82208 6 VGND
port 1 nsew ground input
rlabel metal4 s 19568 2128 19888 107760 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 107760 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 5298 58880 5618 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 35934 58880 36254 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 66570 58880 66890 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 97206 58880 97526 6 VPWR
port 2 nsew power input
rlabel metal4 s 4208 2128 4528 107760 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 107760 6 VPWR
port 2 nsew power input
rlabel metal3 s 0 43256 800 43376 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 59246 9256 60046 9376 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 59246 60120 60046 60240 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 59246 65152 60046 65272 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 59246 70184 60046 70304 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 59246 75352 60046 75472 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 59246 80384 60046 80504 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 59246 85552 60046 85672 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 59246 90584 60046 90704 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 59246 95616 60046 95736 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 59246 100784 60046 100904 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 59246 105816 60046 105936 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 59246 14288 60046 14408 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal2 s 35070 109390 35126 110190 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal2 s 36450 109390 36506 110190 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal2 s 37922 109390 37978 110190 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal2 s 39302 109390 39358 110190 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal2 s 40682 109390 40738 110190 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal2 s 42062 109390 42118 110190 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal2 s 43442 109390 43498 110190 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal2 s 44822 109390 44878 110190 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal2 s 46294 109390 46350 110190 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal2 s 47674 109390 47730 110190 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 59246 19456 60046 19576 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal2 s 49054 109390 49110 110190 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal2 s 50434 109390 50490 110190 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal2 s 51814 109390 51870 110190 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal2 s 53286 109390 53342 110190 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal2 s 54666 109390 54722 110190 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal2 s 56046 109390 56102 110190 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal2 s 57426 109390 57482 110190 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal2 s 58806 109390 58862 110190 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 59246 24488 60046 24608 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 59246 29520 60046 29640 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 59246 34688 60046 34808 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 59246 39720 60046 39840 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 59246 44888 60046 45008 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 59246 49920 60046 50040 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 59246 54952 60046 55072 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 59246 10888 60046 11008 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 59246 61752 60046 61872 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 59246 66920 60046 67040 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 59246 71952 60046 72072 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 59246 76984 60046 77104 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 59246 82152 60046 82272 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 59246 87184 60046 87304 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 59246 92216 60046 92336 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 59246 97384 60046 97504 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 59246 102416 60046 102536 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 59246 107584 60046 107704 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 59246 16056 60046 16176 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal2 s 35530 109390 35586 110190 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal2 s 36910 109390 36966 110190 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal2 s 38382 109390 38438 110190 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal2 s 39762 109390 39818 110190 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal2 s 41142 109390 41198 110190 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal2 s 42522 109390 42578 110190 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal2 s 43902 109390 43958 110190 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal2 s 45374 109390 45430 110190 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal2 s 46754 109390 46810 110190 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal2 s 48134 109390 48190 110190 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 59246 21088 60046 21208 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal2 s 49514 109390 49570 110190 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal2 s 50894 109390 50950 110190 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal2 s 52274 109390 52330 110190 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal2 s 53746 109390 53802 110190 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal2 s 55126 109390 55182 110190 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal2 s 56506 109390 56562 110190 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal2 s 57886 109390 57942 110190 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal2 s 59266 109390 59322 110190 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 59246 26120 60046 26240 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 59246 31288 60046 31408 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 59246 36320 60046 36440 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 59246 41488 60046 41608 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 59246 46520 60046 46640 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 59246 51552 60046 51672 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 59246 56720 60046 56840 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 59246 12656 60046 12776 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 59246 63520 60046 63640 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 59246 68552 60046 68672 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 59246 73584 60046 73704 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 59246 78752 60046 78872 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 59246 83784 60046 83904 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 59246 88952 60046 89072 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 59246 93984 60046 94104 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 59246 99016 60046 99136 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 59246 104184 60046 104304 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 59246 109216 60046 109336 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 59246 17688 60046 17808 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal2 s 35990 109390 36046 110190 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal2 s 37370 109390 37426 110190 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal2 s 38842 109390 38898 110190 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal2 s 40222 109390 40278 110190 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal2 s 41602 109390 41658 110190 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal2 s 42982 109390 43038 110190 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal2 s 44362 109390 44418 110190 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal2 s 45834 109390 45890 110190 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal2 s 47214 109390 47270 110190 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal2 s 48594 109390 48650 110190 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 59246 22856 60046 22976 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal2 s 49974 109390 50030 110190 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal2 s 51354 109390 51410 110190 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal2 s 52826 109390 52882 110190 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal2 s 54206 109390 54262 110190 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal2 s 55586 109390 55642 110190 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal2 s 56966 109390 57022 110190 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal2 s 58346 109390 58402 110190 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal2 s 59726 109390 59782 110190 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 59246 27888 60046 28008 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 59246 32920 60046 33040 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 59246 38088 60046 38208 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 59246 43120 60046 43240 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 59246 48152 60046 48272 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 59246 53320 60046 53440 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 59246 58352 60046 58472 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 294 0 350 800 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 938 0 994 800 6 pad_flash_clk_oeb
port 157 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 pad_flash_csb_oeb
port 159 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 pad_flash_io0_ieb
port 162 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 pad_flash_io0_oeb
port 163 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 pad_flash_io1_ieb
port 166 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 pad_flash_io1_oeb
port 167 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 porb
port 208 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 pwr_ctrl_out[0]
port 209 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 pwr_ctrl_out[1]
port 210 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 pwr_ctrl_out[2]
port 211 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 pwr_ctrl_out[3]
port 212 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 qspi_enabled
port 213 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 reset
port 214 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 ser_rx
port 215 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 ser_tx
port 216 nsew signal input
rlabel metal3 s 59246 824 60046 944 6 serial_clock
port 217 nsew signal output
rlabel metal3 s 59246 5856 60046 5976 6 serial_data_1
port 218 nsew signal output
rlabel metal3 s 59246 7488 60046 7608 6 serial_data_2
port 219 nsew signal output
rlabel metal3 s 59246 4088 60046 4208 6 serial_load
port 220 nsew signal output
rlabel metal3 s 59246 2456 60046 2576 6 serial_resetn
port 221 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 spi_csb
port 222 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 spi_enabled
port 223 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 spi_sck
port 224 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 spi_sdi
port 225 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 spi_sdo
port 226 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 spi_sdoenb
port 227 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 spimemio_flash_clk
port 228 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 spimemio_flash_csb
port 229 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 spimemio_flash_io0_di
port 230 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 spimemio_flash_io0_do
port 231 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 spimemio_flash_io0_oeb
port 232 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 spimemio_flash_io1_di
port 233 nsew signal output
rlabel metal3 s 0 102416 800 102536 6 spimemio_flash_io1_do
port 234 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 spimemio_flash_io1_oeb
port 235 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 spimemio_flash_io2_di
port 236 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 spimemio_flash_io2_do
port 237 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 spimemio_flash_io2_oeb
port 238 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 spimemio_flash_io3_di
port 239 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 spimemio_flash_io3_do
port 240 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 spimemio_flash_io3_oeb
port 241 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 sram_ro_addr[0]
port 242 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 sram_ro_addr[1]
port 243 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 sram_ro_addr[2]
port 244 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 sram_ro_addr[3]
port 245 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 sram_ro_addr[4]
port 246 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 sram_ro_addr[5]
port 247 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 sram_ro_addr[6]
port 248 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 sram_ro_addr[7]
port 249 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 sram_ro_clk
port 250 nsew signal output
rlabel metal3 s 0 416 800 536 6 sram_ro_csb
port 251 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 sram_ro_data[0]
port 252 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 sram_ro_data[10]
port 253 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 sram_ro_data[11]
port 254 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 sram_ro_data[12]
port 255 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 sram_ro_data[13]
port 256 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 sram_ro_data[14]
port 257 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 sram_ro_data[15]
port 258 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 sram_ro_data[16]
port 259 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 sram_ro_data[17]
port 260 nsew signal input
rlabel metal3 s 0 28976 800 29096 6 sram_ro_data[18]
port 261 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 sram_ro_data[19]
port 262 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 sram_ro_data[1]
port 263 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 sram_ro_data[20]
port 264 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 sram_ro_data[21]
port 265 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 sram_ro_data[22]
port 266 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 sram_ro_data[23]
port 267 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 sram_ro_data[24]
port 268 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 sram_ro_data[25]
port 269 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 sram_ro_data[26]
port 270 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 sram_ro_data[27]
port 271 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 sram_ro_data[28]
port 272 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 sram_ro_data[29]
port 273 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 sram_ro_data[2]
port 274 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 sram_ro_data[30]
port 275 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 sram_ro_data[31]
port 276 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 sram_ro_data[3]
port 277 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 sram_ro_data[4]
port 278 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 sram_ro_data[5]
port 279 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 sram_ro_data[6]
port 280 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 sram_ro_data[7]
port 281 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 sram_ro_data[8]
port 282 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 sram_ro_data[9]
port 283 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 trap
port 284 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 uart_enabled
port 285 nsew signal input
rlabel metal2 s 32770 109390 32826 110190 6 user_clock
port 286 nsew signal input
rlabel metal2 s 33230 109390 33286 110190 6 usr1_vcc_pwrgood
port 287 nsew signal input
rlabel metal2 s 34150 109390 34206 110190 6 usr1_vdd_pwrgood
port 288 nsew signal input
rlabel metal2 s 33690 109390 33746 110190 6 usr2_vcc_pwrgood
port 289 nsew signal input
rlabel metal2 s 34610 109390 34666 110190 6 usr2_vdd_pwrgood
port 290 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 wb_ack_o
port 291 nsew signal output
rlabel metal2 s 202 109390 258 110190 6 wb_adr_i[0]
port 292 nsew signal input
rlabel metal2 s 4802 109390 4858 110190 6 wb_adr_i[10]
port 293 nsew signal input
rlabel metal2 s 5262 109390 5318 110190 6 wb_adr_i[11]
port 294 nsew signal input
rlabel metal2 s 5722 109390 5778 110190 6 wb_adr_i[12]
port 295 nsew signal input
rlabel metal2 s 6182 109390 6238 110190 6 wb_adr_i[13]
port 296 nsew signal input
rlabel metal2 s 6642 109390 6698 110190 6 wb_adr_i[14]
port 297 nsew signal input
rlabel metal2 s 7102 109390 7158 110190 6 wb_adr_i[15]
port 298 nsew signal input
rlabel metal2 s 7562 109390 7618 110190 6 wb_adr_i[16]
port 299 nsew signal input
rlabel metal2 s 8114 109390 8170 110190 6 wb_adr_i[17]
port 300 nsew signal input
rlabel metal2 s 8574 109390 8630 110190 6 wb_adr_i[18]
port 301 nsew signal input
rlabel metal2 s 9034 109390 9090 110190 6 wb_adr_i[19]
port 302 nsew signal input
rlabel metal2 s 662 109390 718 110190 6 wb_adr_i[1]
port 303 nsew signal input
rlabel metal2 s 9494 109390 9550 110190 6 wb_adr_i[20]
port 304 nsew signal input
rlabel metal2 s 9954 109390 10010 110190 6 wb_adr_i[21]
port 305 nsew signal input
rlabel metal2 s 10414 109390 10470 110190 6 wb_adr_i[22]
port 306 nsew signal input
rlabel metal2 s 10874 109390 10930 110190 6 wb_adr_i[23]
port 307 nsew signal input
rlabel metal2 s 11334 109390 11390 110190 6 wb_adr_i[24]
port 308 nsew signal input
rlabel metal2 s 11794 109390 11850 110190 6 wb_adr_i[25]
port 309 nsew signal input
rlabel metal2 s 12254 109390 12310 110190 6 wb_adr_i[26]
port 310 nsew signal input
rlabel metal2 s 12714 109390 12770 110190 6 wb_adr_i[27]
port 311 nsew signal input
rlabel metal2 s 13174 109390 13230 110190 6 wb_adr_i[28]
port 312 nsew signal input
rlabel metal2 s 13634 109390 13690 110190 6 wb_adr_i[29]
port 313 nsew signal input
rlabel metal2 s 1122 109390 1178 110190 6 wb_adr_i[2]
port 314 nsew signal input
rlabel metal2 s 14094 109390 14150 110190 6 wb_adr_i[30]
port 315 nsew signal input
rlabel metal2 s 14554 109390 14610 110190 6 wb_adr_i[31]
port 316 nsew signal input
rlabel metal2 s 1582 109390 1638 110190 6 wb_adr_i[3]
port 317 nsew signal input
rlabel metal2 s 2042 109390 2098 110190 6 wb_adr_i[4]
port 318 nsew signal input
rlabel metal2 s 2502 109390 2558 110190 6 wb_adr_i[5]
port 319 nsew signal input
rlabel metal2 s 2962 109390 3018 110190 6 wb_adr_i[6]
port 320 nsew signal input
rlabel metal2 s 3422 109390 3478 110190 6 wb_adr_i[7]
port 321 nsew signal input
rlabel metal2 s 3882 109390 3938 110190 6 wb_adr_i[8]
port 322 nsew signal input
rlabel metal2 s 4342 109390 4398 110190 6 wb_adr_i[9]
port 323 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wb_clk_i
port 324 nsew signal input
rlabel metal2 s 32310 109390 32366 110190 6 wb_cyc_i
port 325 nsew signal input
rlabel metal2 s 15014 109390 15070 110190 6 wb_dat_i[0]
port 326 nsew signal input
rlabel metal2 s 19706 109390 19762 110190 6 wb_dat_i[10]
port 327 nsew signal input
rlabel metal2 s 20166 109390 20222 110190 6 wb_dat_i[11]
port 328 nsew signal input
rlabel metal2 s 20626 109390 20682 110190 6 wb_dat_i[12]
port 329 nsew signal input
rlabel metal2 s 21086 109390 21142 110190 6 wb_dat_i[13]
port 330 nsew signal input
rlabel metal2 s 21546 109390 21602 110190 6 wb_dat_i[14]
port 331 nsew signal input
rlabel metal2 s 22006 109390 22062 110190 6 wb_dat_i[15]
port 332 nsew signal input
rlabel metal2 s 22466 109390 22522 110190 6 wb_dat_i[16]
port 333 nsew signal input
rlabel metal2 s 23018 109390 23074 110190 6 wb_dat_i[17]
port 334 nsew signal input
rlabel metal2 s 23478 109390 23534 110190 6 wb_dat_i[18]
port 335 nsew signal input
rlabel metal2 s 23938 109390 23994 110190 6 wb_dat_i[19]
port 336 nsew signal input
rlabel metal2 s 15566 109390 15622 110190 6 wb_dat_i[1]
port 337 nsew signal input
rlabel metal2 s 24398 109390 24454 110190 6 wb_dat_i[20]
port 338 nsew signal input
rlabel metal2 s 24858 109390 24914 110190 6 wb_dat_i[21]
port 339 nsew signal input
rlabel metal2 s 25318 109390 25374 110190 6 wb_dat_i[22]
port 340 nsew signal input
rlabel metal2 s 25778 109390 25834 110190 6 wb_dat_i[23]
port 341 nsew signal input
rlabel metal2 s 26238 109390 26294 110190 6 wb_dat_i[24]
port 342 nsew signal input
rlabel metal2 s 26698 109390 26754 110190 6 wb_dat_i[25]
port 343 nsew signal input
rlabel metal2 s 27158 109390 27214 110190 6 wb_dat_i[26]
port 344 nsew signal input
rlabel metal2 s 27618 109390 27674 110190 6 wb_dat_i[27]
port 345 nsew signal input
rlabel metal2 s 28078 109390 28134 110190 6 wb_dat_i[28]
port 346 nsew signal input
rlabel metal2 s 28538 109390 28594 110190 6 wb_dat_i[29]
port 347 nsew signal input
rlabel metal2 s 16026 109390 16082 110190 6 wb_dat_i[2]
port 348 nsew signal input
rlabel metal2 s 28998 109390 29054 110190 6 wb_dat_i[30]
port 349 nsew signal input
rlabel metal2 s 29458 109390 29514 110190 6 wb_dat_i[31]
port 350 nsew signal input
rlabel metal2 s 16486 109390 16542 110190 6 wb_dat_i[3]
port 351 nsew signal input
rlabel metal2 s 16946 109390 17002 110190 6 wb_dat_i[4]
port 352 nsew signal input
rlabel metal2 s 17406 109390 17462 110190 6 wb_dat_i[5]
port 353 nsew signal input
rlabel metal2 s 17866 109390 17922 110190 6 wb_dat_i[6]
port 354 nsew signal input
rlabel metal2 s 18326 109390 18382 110190 6 wb_dat_i[7]
port 355 nsew signal input
rlabel metal2 s 18786 109390 18842 110190 6 wb_dat_i[8]
port 356 nsew signal input
rlabel metal2 s 19246 109390 19302 110190 6 wb_dat_i[9]
port 357 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wb_dat_o[0]
port 358 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 wb_dat_o[10]
port 359 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_dat_o[11]
port 360 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 wb_dat_o[12]
port 361 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 wb_dat_o[13]
port 362 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 wb_dat_o[14]
port 363 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 wb_dat_o[15]
port 364 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 wb_dat_o[16]
port 365 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 wb_dat_o[17]
port 366 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 wb_dat_o[18]
port 367 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 wb_dat_o[19]
port 368 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 wb_dat_o[1]
port 369 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 wb_dat_o[20]
port 370 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 wb_dat_o[21]
port 371 nsew signal output
rlabel metal3 s 0 86096 800 86216 6 wb_dat_o[22]
port 372 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 wb_dat_o[23]
port 373 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 wb_dat_o[24]
port 374 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 wb_dat_o[25]
port 375 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 wb_dat_o[26]
port 376 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 wb_dat_o[27]
port 377 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 wb_dat_o[28]
port 378 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 wb_dat_o[29]
port 379 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 wb_dat_o[2]
port 380 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 wb_dat_o[30]
port 381 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 wb_dat_o[31]
port 382 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 wb_dat_o[3]
port 383 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 wb_dat_o[4]
port 384 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 wb_dat_o[5]
port 385 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 wb_dat_o[6]
port 386 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 wb_dat_o[7]
port 387 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 wb_dat_o[8]
port 388 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 wb_dat_o[9]
port 389 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wb_rstn_i
port 390 nsew signal input
rlabel metal2 s 29918 109390 29974 110190 6 wb_sel_i[0]
port 391 nsew signal input
rlabel metal2 s 30470 109390 30526 110190 6 wb_sel_i[1]
port 392 nsew signal input
rlabel metal2 s 30930 109390 30986 110190 6 wb_sel_i[2]
port 393 nsew signal input
rlabel metal2 s 31390 109390 31446 110190 6 wb_sel_i[3]
port 394 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 wb_stb_i
port 395 nsew signal input
rlabel metal2 s 31850 109390 31906 110190 6 wb_we_i
port 396 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60046 110190
string LEFview TRUE
string GDS_FILE /home/ma/ef/caravel_openframe/openlane/housekeeping/runs/housekeeping/results/magic/housekeeping.gds
string GDS_END 22580570
string GDS_START 1111786
<< end >>

