* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s15_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XANTENNA__6209__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5530__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3691__A2 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2978_A _7073_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6914_ _6994_/CLK _6914_/D fanout462/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3443__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6845_ _7017_/CLK _6845_/D fanout461/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6776_ _3958_/A1 _6776_/D _6428_/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtn_1
X_3988_ _3988_/A _5220_/C VGND VGND VPWR VPWR _3999_/S sky130_fd_sc_hd__and2_4
XFILLER_167_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5727_ _5727_/A _5727_/B _5727_/C _5727_/D VGND VGND VPWR VPWR _5727_/Y sky130_fd_sc_hd__nor4_1
XFILLER_163_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5658_ _5689_/A _5686_/B _5689_/C VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__and3b_4
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4609_ _5100_/C _4609_/B _4609_/C _4609_/D VGND VGND VPWR VPWR _4614_/B sky130_fd_sc_hd__and4_1
XFILLER_117_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _6490_/Q _6492_/Q VGND VGND VPWR VPWR _5589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold340 hold340/A VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold351 hold351/A VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold373 hold373/A VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold384 hold384/A VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5006__A _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5120__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 hold32/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 hold69/X VGND VGND VPWR VPWR _3998_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5440__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3682__A2 _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1062 _3249_/X VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input127_A wb_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1073 _3269_/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1084 hold66/X VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _6754_/Q VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1980_A _6585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6081__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3434__A2 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input92_A spimemio_flash_io3_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5895__B1 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3370__A1 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7201__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5350__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4960_ _4552_/B _5033_/B _4782_/X VGND VGND VPWR VPWR _4961_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3911_ _5643_/A _3911_/B VGND VGND VPWR VPWR _3912_/B sky130_fd_sc_hd__and2b_1
X_4891_ _5114_/A _5102_/A _5130_/A _5103_/A VGND VGND VPWR VPWR _4892_/D sky130_fd_sc_hd__and4_1
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6630_ _6794_/CLK _6630_/D fanout434/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_4
X_3842_ _3182_/Y _3846_/S _3840_/B _3842_/C1 VGND VGND VPWR VPWR _3842_/X sky130_fd_sc_hd__o211a_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6561_ _7184_/CLK _6561_/D VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfxtp_1
X_3773_ input93/X _5226_/A _5207_/A _5254_/A _6845_/Q VGND VGND VPWR VPWR _3773_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2461_A _6569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5512_ _5512_/A0 _5575_/A1 _5514_/S VGND VGND VPWR VPWR _5512_/X sky130_fd_sc_hd__mux2_1
X_6492_ _7179_/CLK _6492_/D fanout446/X VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5443_ _5443_/A _5533_/B VGND VGND VPWR VPWR _5451_/S sky130_fd_sc_hd__and2_4
XFILLER_161_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5525__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5886__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5374_ _5374_/A0 _5563_/A1 _5379_/S VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7113_ _7137_/CLK _7113_/D fanout466/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3361__A1 _6852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4325_ hold168/X _5527_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7044_ _7139_/CLK hold72/X fanout471/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_4
X_4256_ _4256_/A _5533_/B VGND VGND VPWR VPWR _4261_/S sky130_fd_sc_hd__and2_4
XFILLER_68_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3207_ _7096_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4187_ _4187_/A0 _5277_/A1 _4187_/S VGND VGND VPWR VPWR _4187_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout377_A hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4861__B2 _4714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6924__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3416__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5810__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6091__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1394_A _6807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6828_ _6828_/CLK hold49/X _6411_/A VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6759_ _6761_/CLK _6759_/D _6416_/A VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6118__B2 _6985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5435__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3744__A _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5877__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 hold170/A VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold192 _4059_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6266__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4852__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3407__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4907__A2 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6109__A1 _7088_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6109__B2 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5345__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4110_ _3675_/Y hold998/A _4115_/S VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__mux2_1
X_5090_ _4950_/X _4769_/Y _5090_/C _5090_/D VGND VGND VPWR VPWR _5137_/B sky130_fd_sc_hd__and4bb_1
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1809 hold252/X VGND VGND VPWR VPWR _5495_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6293__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4041_ hold602/X _5584_/A1 _4056_/C VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3646__A2 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6045__B1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5992_ _6014_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _5992_/X sky130_fd_sc_hd__and3_4
XFILLER_52_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4943_ _4462_/Y _4938_/X _4791_/C VGND VGND VPWR VPWR _5151_/C sky130_fd_sc_hd__o21a_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ _4500_/Y _4652_/Y _4873_/Y VGND VGND VPWR VPWR _4875_/D sky130_fd_sc_hd__o21a_1
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ _6746_/CLK _6613_/D _6416_/A VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_2
X_3825_ _3253_/A _3824_/X _3835_/S VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6544_ _7191_/CLK _6544_/D VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3756_ _6973_/Q _5398_/A _5434_/A _7005_/Q _3755_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5763__B _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6475_ _6733_/CLK _6475_/D fanout433/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3687_ _7134_/Q _3295_/Y _5175_/A _6783_/Q _3685_/X VGND VGND VPWR VPWR _3694_/A
+ sky130_fd_sc_hd__a221o_1
X_5426_ _5426_/A0 _5561_/A1 _5433_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
Xoutput220 _7216_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7226_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
XFILLER_133_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput242 _7208_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput253 _3961_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
XFILLER_114_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5357_ _5357_/A0 _5537_/A1 _5361_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
Xoutput264 _6786_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput275 _6476_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput286 _6802_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput297 _6804_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
X_4308_ _4308_/A0 _5195_/A1 _4309_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5288_ _5288_/A0 _5567_/A1 _5289_/S VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5087__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6284__B1 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7027_ _7082_/CLK _7027_/D fanout464/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_4
X_4239_ _5244_/A0 _5577_/A1 _5236_/C VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3637__A2 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6036__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7126__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3573__B2 _6710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input55_A mgmt_gpio_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6894__SET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6275__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3628__A2 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6027__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output309_A _3965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3800__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3610_ _7024_/Q _5452_/A _5398_/A _6976_/Q _3609_/X VGND VGND VPWR VPWR _3614_/C
+ sky130_fd_sc_hd__a221o_1
X_4590_ _4638_/A _4590_/B VGND VGND VPWR VPWR _4590_/Y sky130_fd_sc_hd__nand2_8
XFILLER_190_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3564__A1 _7088_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3541_ _6799_/Q _3319_/Y _4140_/A _6593_/Q VGND VGND VPWR VPWR _3541_/X sky130_fd_sc_hd__a22o_4
XANTENNA__3564__B2 _6617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold906 hold906/A VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold917 hold917/A VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold928 hold928/A VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold939 hold939/A VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6260_ _6723_/Q _5978_/X _5995_/X _6600_/Q _6259_/X VGND VGND VPWR VPWR _6263_/C
+ sky130_fd_sc_hd__a221o_1
X_3472_ _6985_/Q _5407_/A _4292_/A _6726_/Q _3471_/X VGND VGND VPWR VPWR _3481_/B
+ sky130_fd_sc_hd__a221o_1
X_5211_ hold24/X _5569_/B VGND VGND VPWR VPWR _5217_/S sky130_fd_sc_hd__and2_4
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6191_ _6490_/Q _6191_/A2 _5649_/Y VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2307 _6857_/Q VGND VGND VPWR VPWR hold744/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5142_ _4688_/A _4995_/B _5023_/C _5141_/X _4815_/X VGND VGND VPWR VPWR _5143_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold2318 _5427_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2329 hold600/X VGND VGND VPWR VPWR _5584_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1606 _5348_/X VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1617 _7092_/Q VGND VGND VPWR VPWR hold389/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1628 _5280_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5073_ _4776_/A _5073_/B _5073_/C _5100_/B VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__and4b_1
XFILLER_38_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1639 hold294/X VGND VGND VPWR VPWR _4293_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3619__A2 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4816__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4816__B2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4024_ _6514_/Q hold39/X _4047_/C VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ _6017_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _5976_/B sky130_fd_sc_hd__and3_4
XANTENNA__5241__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _4633_/B _4698_/Y _4702_/Y _4616_/B _4616_/A VGND VGND VPWR VPWR _4931_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4857_ _4917_/D _4857_/B _4857_/C VGND VGND VPWR VPWR _4857_/Y sky130_fd_sc_hd__nand3_1
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ _3814_/B _6468_/Q _6469_/Q VGND VGND VPWR VPWR _3811_/B sky130_fd_sc_hd__and3b_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4788_ _4947_/A _4698_/Y _4531_/B VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6527_ _6803_/CLK _6527_/D fanout442/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3555__B2 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3739_ _3738_/X _3739_/A1 _3739_/S VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6458_ _3958_/A1 _6458_/D _6408_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5409_ _5409_/A0 _5562_/A1 _5415_/S VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6389_ _4222_/B _3189_/Y _4220_/B _6388_/X _6387_/X VGND VGND VPWR VPWR _7204_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6257__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2830 hold935/X VGND VGND VPWR VPWR _4228_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2841 _7058_/Q VGND VGND VPWR VPWR hold957/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2852 _3424_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2863 _6679_/Q VGND VGND VPWR VPWR _3918_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2874 _6242_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2885 _7161_/Q VGND VGND VPWR VPWR _5750_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2896 _7202_/Q VGND VGND VPWR VPWR _6384_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6009__B1 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5480__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5232__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4064__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5783__A2 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3546__B2 _7009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7145__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output259_A _6794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6248__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4239__S _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5471__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2005_A _6740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5578__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5223__A1 _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _5760_/A _5760_/B _5760_/C VGND VGND VPWR VPWR _5760_/Y sky130_fd_sc_hd__nor3_4
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5774__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4711_ _4826_/A _4730_/B VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__nand2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5691_ _7077_/Q _5689_/X _5690_/X _5683_/X VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4642_ _4640_/Y _4857_/B VGND VGND VPWR VPWR _4642_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4573_ _4811_/B _4607_/B VGND VGND VPWR VPWR _4757_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold703 hold703/A VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap422 _4677_/A VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__clkbuf_2
Xhold714 hold714/A VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6312_ _6587_/Q _5989_/X _6309_/X _6311_/X VGND VGND VPWR VPWR _6313_/C sky130_fd_sc_hd__a211oi_1
X_3524_ _7089_/Q _5524_/A _4262_/A _6701_/Q VGND VGND VPWR VPWR _3524_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold736 hold736/A VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold747 hold747/A VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6768__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold758 hold758/A VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6243_ _6595_/Q _5991_/X _6018_/X _6718_/Q VGND VGND VPWR VPWR _6243_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _7074_/Q _5506_/A _5434_/A _7010_/Q VGND VGND VPWR VPWR _3455_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6174_ _7059_/Q _5990_/X _5998_/X _6891_/Q _6173_/X VGND VGND VPWR VPWR _6179_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2104 hold804/X VGND VGND VPWR VPWR _4338_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2115 _6716_/Q VGND VGND VPWR VPWR hold837/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3386_ _6448_/Q _6656_/Q VGND VGND VPWR VPWR _3739_/S sky130_fd_sc_hd__nand2_8
Xhold2126 _7086_/Q VGND VGND VPWR VPWR hold551/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5125_ _5139_/B _5125_/B _5125_/C VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__and3_1
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2137 _5313_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1403 _7139_/Q VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2148 _6479_/Q VGND VGND VPWR VPWR hold731/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1414 _7049_/Q VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2159 _4279_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1425 _3978_/X VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1436 hold254/X VGND VGND VPWR VPWR _5463_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1447 _6959_/Q VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5056_ _4610_/A _4693_/B _4508_/B VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__o21ai_1
Xhold1458 _5327_/X VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1469 _5432_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5462__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4007_ hold233/X wire371/X _4008_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout457_A _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5488__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5214__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5958_ _6756_/Q _5681_/X _5956_/X _5957_/X VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5765__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__B2 _6782_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4909_ _4633_/B _4688_/A _4872_/A _4889_/B VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__o211a_1
X_5889_ _6693_/Q _5658_/X _5664_/X _6758_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3528__B2 _6889_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6190__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7168__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1641_A _6631_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input157_A wb_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4567__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4059__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__buf_12
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2660 hold664/X VGND VGND VPWR VPWR _4175_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2671 _6745_/Q VGND VGND VPWR VPWR hold797/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__buf_2
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2682 _6727_/Q VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2693 _6577_/Q VGND VGND VPWR VPWR hold788/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5453__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1970 _6523_/Q VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1981 hold528/X VGND VGND VPWR VPWR _4136_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input18_A mask_rev_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1992 _6501_/Q VGND VGND VPWR VPWR hold887/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _3950_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5398__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5205__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5756__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3767__A1 _6803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3767__B2 _7021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6181__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4192__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _3543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5141__B1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6685__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5444__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _6936_/CLK _6930_/D fanout463/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3455__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6861_ _7101_/CLK _6861_/D fanout450/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_6_csclk _6549_/CLK VGND VGND VPWR VPWR _6756_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5812_ _6914_/Q _5670_/X _5685_/X _7074_/Q VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__a22o_1
X_6792_ _6793_/CLK _6792_/D fanout434/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5747__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5743_ _6855_/Q _5651_/X _5653_/X _6847_/Q VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5528__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5674_ _5689_/A _5679_/B _5688_/C VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__and3b_4
XFILLER_136_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4625_ _4625_/A _4625_/B VGND VGND VPWR VPWR _4625_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6172__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold500 hold500/A VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4183__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4556_ _4921_/A _4554_/X _4556_/C _5136_/A VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__and4bb_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold522 _4058_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold533 hold533/A VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold544 _4238_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3507_ _3535_/A _3523_/B VGND VGND VPWR VPWR _4182_/A sky130_fd_sc_hd__nor2_8
XFILLER_116_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold555 hold555/A VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold566 hold566/A VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4487_ _4595_/B _4488_/B VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__and2_4
Xhold577 _4046_/X VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold588 hold588/A VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6226_ _6535_/Q _5983_/X _6005_/X _6692_/Q VGND VGND VPWR VPWR _6226_/X sky130_fd_sc_hd__a22o_1
X_3438_ input49/X _4047_/C _5560_/A _7122_/Q VGND VGND VPWR VPWR _3438_/X sky130_fd_sc_hd__a22o_1
Xhold599 hold599/A VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5683__B2 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6157_ _7122_/Q _5978_/X _5995_/X _6922_/Q _6156_/X VGND VGND VPWR VPWR _6163_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1200 hold242/X VGND VGND VPWR VPWR _5437_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _7004_/Q _5425_/A _3310_/Y input19/X _3358_/X VGND VGND VPWR VPWR _3369_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1211 hold1211/A VGND VGND VPWR VPWR _5235_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1222_A _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1222 _7044_/Q VGND VGND VPWR VPWR _5478_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5125_/B sky130_fd_sc_hd__and3_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1233 _6968_/Q VGND VGND VPWR VPWR hold383/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6088_ _6088_/A _6088_/B _6088_/C _6088_/D VGND VGND VPWR VPWR _6089_/D sky130_fd_sc_hd__nor4_1
Xhold1244 _6848_/Q VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1255 _7038_/Q VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5435__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1266 hold124/X VGND VGND VPWR VPWR _5320_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _5285_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5039_ _5026_/B _4719_/B _4771_/X VGND VGND VPWR VPWR _5039_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3446__B1 _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1288 hold126/X VGND VGND VPWR VPWR _5419_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1299 _5267_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3997__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1591_A _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5738__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3749__B2 input98/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5438__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4174__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5910__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _3893_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6371_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6377_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_4
XFILLER_64_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5426__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2490 hold971/X VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3437__B1 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5202__A _5202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5348__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6154__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4410_ _4719_/A _4590_/B VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__and2_4
XANTENNA__4165__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5390_ _5390_/A0 _5534_/A1 _5397_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5901__A2 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4341_ _3890_/Y _4340_/Y _4395_/A VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__o21a_2
XFILLER_172_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7060_ _7130_/CLK _7060_/D fanout462/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4272_ hold67/X hold43/X _4273_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6011_ _6002_/X _6011_/B VGND VGND VPWR VPWR _6313_/D sky130_fd_sc_hd__nand2b_4
X_3223_ _6968_/Q VGND VGND VPWR VPWR _5763_/A sky130_fd_sc_hd__inv_2
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4000__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5417__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7148__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6090__A1 _6839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3979__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6913_ _6967_/CLK _6913_/D fanout465/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6844_ _7084_/CLK _6844_/D fanout447/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3987_ _3987_/A0 _5189_/A1 _3987_/S VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6775_ _3958_/A1 _6775_/D _6427_/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5726_ _6990_/Q _5929_/B _5688_/X _6886_/Q _5725_/X VGND VGND VPWR VPWR _5727_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3600__B1 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5657_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5689_/C sky130_fd_sc_hd__and2_4
XANTENNA__6145__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4156__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4608_ _4570_/A _4564_/Y _4574_/A _4495_/B VGND VGND VPWR VPWR _4609_/D sky130_fd_sc_hd__a211o_1
X_5588_ _6816_/Q _6489_/Q _3197_/Y _5588_/B1 _5587_/X VGND VGND VPWR VPWR _5588_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_190_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold341 hold341/A VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4539_ _4621_/A _4972_/A VGND VGND VPWR VPWR _4539_/Y sky130_fd_sc_hd__nand2_2
Xhold352 _4061_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold363 hold363/A VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 hold396/A VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ _6956_/Q _5997_/X _6012_/X _7004_/Q VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__a22o_1
X_7189_ _7194_/CLK _7189_/D VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5120__A3 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1030 hold3/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _6441_/Q VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5408__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _3998_/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _3648_/B VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3419__B1 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1074 _3272_/Y VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5959__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1085 _6768_/Q VGND VGND VPWR VPWR _5167_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1096 hold180/X VGND VGND VPWR VPWR _4331_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1973_A _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input85_A spimemio_flash_io0_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6136__A2 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4147__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7013__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3370__A2 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output241_A _3931_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6733_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3910_ _7142_/Q _7143_/Q _7144_/Q _7145_/Q VGND VGND VPWR VPWR _3911_/B sky130_fd_sc_hd__and4bb_1
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _4464_/Y _4601_/A _4601_/B _4581_/X VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__a211o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3841_ _3841_/A _3841_/B VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__xnor2_1
XFILLER_158_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3772_ _6579_/Q _4128_/A _4212_/A _6649_/Q _3771_/X VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a221o_1
X_6560_ _7191_/CLK _6560_/D VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ hold99/X hold95/X _5514_/S VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6491_ _7180_/CLK _6491_/D fanout446/X VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6127__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4138__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5442_ _5442_/A0 _5577_/A1 _5442_/S VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5886__B2 _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5373_ hold596/X _5562_/A1 _5379_/S VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2621_A _6796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7072_/CLK sky130_fd_sc_hd__clkbuf_16
X_7112_ _7112_/CLK _7112_/D fanout473/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_4
X_4324_ _4324_/A0 _5238_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3361__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7043_ _7136_/CLK _7043_/D fanout471/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4255_ _4255_/A0 _5189_/A1 _4255_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5541__S _5541_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3206_ _7104_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4186_ _4186_/A0 _5233_/A1 _4187_/S VGND VGND VPWR VPWR _4186_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6992_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4861__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _6549_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_55_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3996__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4613__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6827_ _6828_/CLK _6827_/D _6411_/A VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6758_ _6830_/CLK _6758_/D _6407_/A VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5709_ _5729_/A0 _5649_/Y _5707_/Y _5708_/X VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__a22o_1
XANTENNA__6118__A2 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6689_ _6701_/CLK _6689_/D fanout436/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_hold1554_A _6452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3888__B1 _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold171 hold171/A VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5451__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7232__A _7232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4301__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4852__A2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6634__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6109__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output289_A _6481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3591__A2 _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4540__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5361__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6293__A1 _6617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4040_ _4040_/A0 _4039_/X _4046_/S VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6293__B2 _6582_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6045__A1 _7054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6045__B2 _6950_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5991_ _6017_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__and3_4
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _5026_/B _5033_/A VGND VGND VPWR VPWR _5032_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4873_ _4988_/A _4607_/B _4526_/X VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2571_A _6804_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6612_ _6756_/CLK _6612_/D fanout441/X VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_4
X_3824_ _3254_/X _3253_/Y _3827_/B VGND VGND VPWR VPWR _3824_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3755_ _6861_/Q _5272_/A _3521_/Y _6535_/Q VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__a22o_1
X_6543_ _7194_/CLK _6543_/D VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5536__S _5541_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3582__A2 _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6474_ _6733_/CLK _6474_/D fanout433/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfstp_4
X_3686_ _3686_/A _3686_/B VGND VGND VPWR VPWR _5175_/A sky130_fd_sc_hd__nor2_4
XFILLER_173_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5425_ _5425_/A _5578_/B VGND VGND VPWR VPWR _5433_/S sky130_fd_sc_hd__and2_4
Xoutput210 _3233_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput221 _7217_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_160_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 _7227_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7209_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
XFILLER_133_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput254 _7231_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ _5356_/A0 _5527_/A1 _5361_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6787_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput276 _6477_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_160_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput287 _6487_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
X_4307_ _4307_/A0 _5194_/A1 _4309_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _6805_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XANTENNA__4676__A _4751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5287_ _5287_/A0 _5575_/A1 _5289_/S VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5271__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6284__A1 _6689_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4238_ _4238_/A0 _4237_/X _4240_/S VGND VGND VPWR VPWR _4238_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6284__B2 _6739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7026_ _7072_/CLK _7026_/D fanout464/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _4169_/A0 _5448_/A1 _4169_/S VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold1302_A _6713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6036__A1 _7133_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3270__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5446__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3573__A2 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input48_A mgmt_gpio_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3730__C1 _3729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout470 input75/X VGND VGND VPWR VPWR fanout470/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_5__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6027__A1 _6901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6027__B2 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5786__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5210__A _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5356__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3564__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3540_ _3544_/A _3550_/B VGND VGND VPWR VPWR _4140_/A sky130_fd_sc_hd__nor2_8
Xhold907 hold907/A VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold918 hold918/A VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3471_ _6841_/Q _5245_/A _5178_/A _6788_/Q VGND VGND VPWR VPWR _3471_/X sky130_fd_sc_hd__a22o_4
Xhold929 hold929/A VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5210_ _5220_/C _5210_/B VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__and2_1
X_6190_ _6843_/Q _6339_/B _6189_/Y _6166_/S VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5710__B1 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5141_ _5011_/A _4590_/Y _4676_/Y VGND VGND VPWR VPWR _5141_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2308 hold744/X VGND VGND VPWR VPWR _5268_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2319 _7101_/Q VGND VGND VPWR VPWR hold832/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1607 _6980_/Q VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5072_ _5135_/A _5102_/C _5072_/C _5135_/C VGND VGND VPWR VPWR _5074_/C sky130_fd_sc_hd__and4_1
Xhold1618 hold389/X VGND VGND VPWR VPWR _5532_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1629 _6819_/Q VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4816__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4023_ _4023_/A0 _4022_/X _4029_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3965__A_N _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5777__B1 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5974_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6019_/C sky130_fd_sc_hd__nor2_8
XFILLER_80_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3252__A1 _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4925_ _4925_/A _5052_/B _4925_/C VGND VGND VPWR VPWR _4925_/X sky130_fd_sc_hd__and3_1
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4638_/Y _4662_/Y _5073_/B VGND VGND VPWR VPWR _4856_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3807_ _3903_/A _3807_/B VGND VGND VPWR VPWR _3814_/B sky130_fd_sc_hd__and2_2
X_4787_ _4411_/Y _4683_/A _4664_/Y _4509_/Y VGND VGND VPWR VPWR _5034_/B sky130_fd_sc_hd__o31a_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5266__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout402_A hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6526_ _6803_/CLK _6526_/D fanout442/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3555__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3738_ _6774_/Q _3737_/Y _3738_/S VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6457_ _3958_/A1 _6457_/D _6407_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3669_ _7111_/Q _5551_/A hold57/A _6571_/Q VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1252_A _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5408_ _5408_/A0 _5561_/A1 _5415_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5701__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6388_ _6682_/Q hold7/A _6355_/Y VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__o21ba_1
XFILLER_88_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5339_ _5339_/A0 _5537_/A1 _5343_/S VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6257__A1 _6708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2820 hold945/X VGND VGND VPWR VPWR _5269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1517_A _6851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2831 _6660_/Q VGND VGND VPWR VPWR hold967/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2842 hold957/X VGND VGND VPWR VPWR _5494_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2853 _6777_/Q VGND VGND VPWR VPWR _3618_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2864 _6683_/Q VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4807__A2 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2875 hold26/A VGND VGND VPWR VPWR _3829_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7009_ _7137_/CLK _7009_/D fanout466/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2886 _7173_/Q VGND VGND VPWR VPWR _6066_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2897 _7169_/Q VGND VGND VPWR VPWR _5925_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5768__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input102_A wb_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3794__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6193__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3546__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4710_ _4710_/A _5150_/C VGND VGND VPWR VPWR _4832_/C sky130_fd_sc_hd__nand2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A2 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6910__SET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5690_ _6989_/Q _5929_/B _5670_/X _6909_/Q VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6973__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4641_ _4498_/X _4499_/Y _4500_/Y _4501_/X VGND VGND VPWR VPWR _4857_/B sky130_fd_sc_hd__o211a_1
XANTENNA__6184__B1 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4734__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4572_ _4637_/B _4823_/A VGND VGND VPWR VPWR _4572_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5931__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold704 hold704/A VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6311_ _6652_/Q _5996_/X _6012_/X _6750_/Q _6310_/X VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap423 _4677_/A VGND VGND VPWR VPWR _4751_/C sky130_fd_sc_hd__clkbuf_2
Xhold715 hold715/A VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3523_ _3550_/A _3523_/B VGND VGND VPWR VPWR _4262_/A sky130_fd_sc_hd__nor2_8
Xhold726 hold726/A VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold737 hold737/A VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold748 hold748/A VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6242_ _6266_/A0 _6241_/X _6342_/S VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3454_ _7050_/Q hold16/A _5245_/A _6842_/Q _3436_/X VGND VGND VPWR VPWR _3460_/A
+ sky130_fd_sc_hd__a221o_1
Xhold759 hold759/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6173_ _6907_/Q _5985_/X _6018_/X _6971_/Q VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__a22o_1
X_3385_ _3385_/A _3385_/B VGND VGND VPWR VPWR _3385_/Y sky130_fd_sc_hd__nand2_8
Xhold2105 _4338_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2116 hold837/X VGND VGND VPWR VPWR _4285_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2127 hold551/X VGND VGND VPWR VPWR _5526_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2138 _7014_/Q VGND VGND VPWR VPWR hold545/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5124_ _4636_/X _5124_/B _5124_/C _5136_/A VGND VGND VPWR VPWR _5125_/C sky130_fd_sc_hd__and4b_1
Xhold1404 hold215/X VGND VGND VPWR VPWR _5585_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2149 hold731/X VGND VGND VPWR VPWR _4001_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1415 hold339/X VGND VGND VPWR VPWR _5484_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1426 hold274/X VGND VGND VPWR VPWR hold1426/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1437 _5463_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5055_ _4570_/D _4523_/Y _4931_/B _5054_/X VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__o211a_2
Xhold1448 hold224/X VGND VGND VPWR VPWR _5383_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1459 _6583_/Q VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4006_ hold226/X wire375/X _4008_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5957_ _6613_/Q _5660_/X _5669_/X _6653_/Q VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4908_ _4636_/X _5127_/B _5127_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__and3b_1
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3776__A2 _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ _6595_/Q _5670_/X _5685_/X _6770_/Q VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4839_ _4917_/A _4643_/C _4504_/X VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6175__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1467_A _7003_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _6512_/CLK _6509_/D fanout473/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3700__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2650 _6772_/Q VGND VGND VPWR VPWR hold703/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2661 _4175_/X VGND VGND VPWR VPWR hold665/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2672 hold797/X VGND VGND VPWR VPWR _4320_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__clkbuf_4
Xhold2683 hold697/X VGND VGND VPWR VPWR _4299_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2694 hold788/X VGND VGND VPWR VPWR _4126_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1960 _5519_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1971 hold292/X VGND VGND VPWR VPWR _4063_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4583__B _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1982 _4136_/X VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1993 hold887/X VGND VGND VPWR VPWR _4032_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3767__A2 _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5913__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 _3697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5141__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5692__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2115_A _6716_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6860_ _7091_/CLK _6860_/D fanout452/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5811_ _6954_/Q _5672_/X _5679_/X _6906_/Q _5810_/X VGND VGND VPWR VPWR _5811_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6791_ _6793_/CLK _6791_/D fanout434/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3758__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5742_ _6879_/Q _5667_/X _5682_/X _7039_/Q VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6157__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5673_ _5685_/A _5684_/B _5676_/B VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4624_ _4569_/C _4655_/A _4901_/B _4622_/X _5098_/A VGND VGND VPWR VPWR _4624_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_191_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold501 hold501/A VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4555_ _5026_/B _4948_/A _4392_/X VGND VGND VPWR VPWR _4556_/C sky130_fd_sc_hd__a21oi_1
XFILLER_144_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5544__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold523 hold523/A VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold545 hold545/A VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3506_ _6598_/Q _4146_/A _4122_/A _6578_/Q VGND VGND VPWR VPWR _3506_/X sky130_fd_sc_hd__a22o_1
Xhold556 hold556/A VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4486_ _4486_/A _4486_/B VGND VGND VPWR VPWR _4569_/C sky130_fd_sc_hd__nand2_4
Xhold567 hold567/A VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold578 hold578/A VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6225_ _6742_/Q _6014_/X _6219_/X _6224_/X VGND VGND VPWR VPWR _6230_/A sky130_fd_sc_hd__a211o_1
XFILLER_104_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold589 hold589/A VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3437_ input31/X _3307_/Y _3988_/A _6476_/Q VGND VGND VPWR VPWR _3437_/X sky130_fd_sc_hd__a22o_4
XANTENNA__5683__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3368_/A _3368_/B _3368_/C _3368_/D VGND VGND VPWR VPWR _3385_/A sky130_fd_sc_hd__nor4_4
X_6156_ _7106_/Q _6008_/X _6016_/X _7042_/Q VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__a22o_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1201 _5437_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1212 _5235_/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1223 _5478_/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5107_ _5107_/A _5107_/B _5107_/C VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__and3_1
Xhold1234 hold383/X VGND VGND VPWR VPWR _5393_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6087_ _7135_/Q _5977_/X _5984_/X _7095_/Q _6086_/X VGND VGND VPWR VPWR _6088_/D
+ sky130_fd_sc_hd__a221o_1
X_3299_ _3346_/A _3726_/A VGND VGND VPWR VPWR _5254_/A sky130_fd_sc_hd__nor2_8
Xhold1245 hold384/X VGND VGND VPWR VPWR _5258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1256 _6992_/Q VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1267 _5320_/X VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5038_ _4769_/Y _5038_/B _5038_/C VGND VGND VPWR VPWR _5043_/A sky130_fd_sc_hd__and3b_1
XFILLER_26_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1278 _6888_/Q VGND VGND VPWR VPWR hold369/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3446__A1 _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1289 _5419_/X VGND VGND VPWR VPWR hold127/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3446__B2 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5199__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6989_ _7094_/CLK _6989_/D fanout450/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6148__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6778__CLK_N _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5454__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3382__B1 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4578__B _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6320__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__buf_8
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4637_/D sky130_fd_sc_hd__buf_12
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6362_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input30_A mask_rev_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6364_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6368_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6355_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold2480 hold868/X VGND VGND VPWR VPWR _3987_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2491 _6623_/Q VGND VGND VPWR VPWR hold674/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5202__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1790 _7192_/Q VGND VGND VPWR VPWR hold992/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4937__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5872__B _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5364__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2065_A _6846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__B1 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4340_ _4649_/C _4649_/D VGND VGND VPWR VPWR _4340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4271_ _4271_/A0 _5581_/A1 _4273_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6311__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6010_ _6010_/A _6010_/B _6010_/C VGND VGND VPWR VPWR _6011_/B sky130_fd_sc_hd__nor3_2
X_3222_ _6976_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__3676__A1 _3675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6090__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7158__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6912_ _6994_/CLK _6912_/D fanout462/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4009__A _4009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _7084_/CLK _6843_/D fanout447/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5539__S _5541_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ _3958_/A1 _6774_/D _6426_/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtn_1
X_3986_ _3986_/A0 _7199_/Q _3998_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5050__B1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5725_ _6854_/Q _5651_/X _5684_/X _6926_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5656_ _5689_/A _5676_/B _5689_/B VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__and3_4
XFILLER_136_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ _4988_/A _4607_/B VGND VGND VPWR VPWR _4754_/D sky130_fd_sc_hd__nand2_1
XFILLER_191_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5587_ _5610_/A _3915_/Y _6492_/Q VGND VGND VPWR VPWR _5587_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5274__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold320 hold320/A VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3364__B1 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold331 hold331/A VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4538_ _4724_/C _4621_/A VGND VGND VPWR VPWR _4894_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold353 hold353/A VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold364 hold364/A VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold375 _5550_/X VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6302__B1 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4469_ _4917_/A _4469_/B VGND VGND VPWR VPWR _4568_/A sky130_fd_sc_hd__nor2_4
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold397 hold397/A VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6208_ _7092_/Q _5638_/X _5992_/X _6964_/Q _6207_/X VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a221o_1
X_7188_ _7194_/CLK _7188_/D VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6120_/X _6139_/B _6139_/C VGND VGND VPWR VPWR _6139_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1020 _5223_/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1031 _7047_/Q VGND VGND VPWR VPWR _5482_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 hold93/X VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 hold70/X VGND VGND VPWR VPWR hold1053/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3419__A1 _7003_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1064 hold23/X VGND VGND VPWR VPWR _3726_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1075 _3294_/Y VGND VGND VPWR VPWR _3686_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1086 _3257_/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _4331_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6081__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5449__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5592__A1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input78_A spi_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5895__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6493__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_csclk _6549_/CLK VGND VGND VPWR VPWR _6760_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3658__A1 _6596_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4855__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6072__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5359__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3840_ _3840_/A _3840_/B VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5583__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3771_ _6644_/Q _4206_/A _4328_/A _6752_/Q VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3594__B1 _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5510_ _5510_/A0 _5537_/A1 _5514_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6490_ _7179_/CLK _6490_/D fanout447/X VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5441_ _5441_/A0 _5567_/A1 _5442_/S VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5886__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5372_ hold771/X _5561_/A1 _5379_/S VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__mux2_1
X_7111_ _7133_/CLK _7111_/D fanout469/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_4
X_4323_ _4323_/A0 _5543_/A1 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7042_ _7139_/CLK _7042_/D fanout471/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ _4254_/A0 _5195_/A1 _4255_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3649__A1 _6734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3649__B2 _6818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4846__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _7112_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4185_ _4185_/A0 _5581_/A1 _4187_/S VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4074__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5810__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5269__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6826_ _6826_/CLK _6826_/D _6407_/A VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5574__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6757_ _6760_/CLK _6757_/D _6407_/A VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_4
X_3969_ _3969_/A _3969_/B VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_77_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3585__B1 _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5708_ _5692_/X _5697_/X _5706_/X _5647_/Y VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__o31a_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6688_ _6701_/CLK _6688_/D fanout436/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5639_ _5639_/A _5639_/B VGND VGND VPWR VPWR _5639_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6401__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5877__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold150 hold150/A VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold161 hold161/A VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold172 hold172/A VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold194 hold194/A VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A wb_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5801__A2 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5565__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3576__B1 _5202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6674__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5868__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6293__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6045__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5990_ _6014_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__and3_4
XFILLER_18_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4941_ _4729_/A _4691_/Y _4935_/X _4477_/Y _4534_/Y VGND VGND VPWR VPWR _4963_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4872_ _4872_/A _5046_/A _4872_/C _4872_/D VGND VGND VPWR VPWR _4875_/C sky130_fd_sc_hd__and4_1
X_6611_ _6746_/CLK _6611_/D _6416_/A VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5556__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3823_ hold26/A _3826_/B VGND VGND VPWR VPWR _3827_/B sky130_fd_sc_hd__and2_1
XFILLER_20_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7155__SET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__B1 _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6542_ _7194_/CLK _6542_/D VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfxtp_1
X_3754_ _6989_/Q _5416_/A hold16/A _7045_/Q _3753_/X VGND VGND VPWR VPWR _3759_/B
+ sky130_fd_sc_hd__a221o_1
X_6473_ _6486_/CLK _6473_/D fanout433/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfstp_4
X_3685_ _6758_/Q _4334_/A _4176_/A _6620_/Q VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2731_A _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5424_ _5424_/A0 _5568_/A1 _5424_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
Xoutput200 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
XFILLER_173_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput211 _3232_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _3945_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7207_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
Xoutput244 _7210_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
XFILLER_161_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5355_ _5355_/A0 _5571_/A1 _5361_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
Xoutput255 _3963_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5552__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput266 _6788_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _6478_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
X_4306_ _4306_/A0 _5193_/A1 _4309_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
Xoutput288 _6488_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput299 _6806_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
X_5286_ _5286_/A0 _5448_/A1 _5289_/S VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7025_ _7135_/CLK _7025_/D fanout466/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6284__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4237_ _5243_/A0 wire371/X _4237_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout382_A _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4295__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A0 _5233_/A1 _4169_/S VGND VGND VPWR VPWR _4168_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7194_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6036__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7132__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4099_ _3803_/Y hold970/A _4106_/S VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5547__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6809_ _6809_/CLK _6809_/D fanout433/X VGND VGND VPWR VPWR _7206_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6809_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5462__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3730__B1 _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6275__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout460 fanout461/X VGND VGND VPWR VPWR fanout460/X sky130_fd_sc_hd__buf_12
Xfanout471 fanout472/X VGND VGND VPWR VPWR fanout471/X sky130_fd_sc_hd__buf_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6027__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3797__B1 _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6855__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5538__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4210__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold908 hold908/A VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold919 hold919/A VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3470_ hold15/X hold23/X VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__nor2_8
XFILLER_155_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5710__A1 _6998_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5372__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5140_ _5140_/A _5140_/B _5140_/C VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__and3_1
XANTENNA__3721__B1 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2309 _5268_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5071_ _5135_/C VGND VGND VPWR VPWR _5071_/Y sky130_fd_sc_hd__inv_2
Xhold1608 hold367/X VGND VGND VPWR VPWR _5406_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1619 _5532_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4277__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4022_ hold883/X _5583_/A1 _4047_/C VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5973_ _6015_/B _6008_/A _6018_/B VGND VGND VPWR VPWR _5973_/X sky130_fd_sc_hd__and3_4
XANTENNA__5777__B2 _6865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4924_ _4924_/A _4924_/B _4924_/C _5046_/B VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__and4_1
XFILLER_178_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5529__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4855_ _4570_/D _4655_/A _4590_/Y _4674_/Y VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__o22a_1
XANTENNA__5547__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3806_ _6657_/Q _6656_/Q VGND VGND VPWR VPWR _3807_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4201__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4786_ _4729_/A _4698_/Y _5095_/A VGND VGND VPWR VPWR _4786_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _6735_/CLK _6525_/D fanout442/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_4
X_3737_ _3737_/A _3737_/B VGND VGND VPWR VPWR _3737_/Y sky130_fd_sc_hd__nand2_8
XFILLER_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6456_ _3958_/A1 _6456_/D _6406_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_4
X_3668_ _6473_/Q _3988_/A _4262_/A _6699_/Q _3667_/X VGND VGND VPWR VPWR _3673_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5407_ _5407_/A _5578_/B VGND VGND VPWR VPWR _5415_/S sky130_fd_sc_hd__and2_4
XANTENNA__5701__A1 _6981_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6387_ _6686_/Q _6357_/A _6358_/A _6386_/Y VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5701__B2 _7021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5282__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3599_ _7072_/Q _5506_/A _4065_/A _6528_/Q _3598_/X VGND VGND VPWR VPWR _3604_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3712__B1 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A0 _5572_/A1 _5343_/S VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__mux2_1
Xhold2810 hold715/X VGND VGND VPWR VPWR _5522_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6257__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2821 _5269_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2832 hold967/X VGND VGND VPWR VPWR _4226_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_125_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2843 _5494_/X VGND VGND VPWR VPWR hold958/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5269_ _5269_/A0 _5575_/A1 _5271_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2854 _3618_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_7008_ _7133_/CLK _7008_/D fanout468/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2865 _6677_/Q VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2876 _7197_/Q VGND VGND VPWR VPWR _6369_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2887 _6656_/Q VGND VGND VPWR VPWR _3928_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2898 _6449_/Q VGND VGND VPWR VPWR _3858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5768__A1 _6944_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1879_A _7056_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3779__B1 _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4440__A1 _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4991__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5457__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6193__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6193__B2 _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input60_A mgmt_gpio_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5192__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6248__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4259__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5759__A1 _6888_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5367__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4640_ _4341_/X _4640_/B VGND VGND VPWR VPWR _4640_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4571_ _4988_/A _4808_/B VGND VGND VPWR VPWR _4823_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5931__A1 _6533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5931__B2 _6587_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6310_ _6637_/Q _5994_/X _6018_/X _6720_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
X_3522_ _6945_/Q _5362_/A _3521_/Y _6539_/Q _3520_/X VGND VGND VPWR VPWR _3529_/B
+ sky130_fd_sc_hd__a221o_1
Xhold705 hold705/A VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap424 _4726_/B VGND VGND VPWR VPWR _4732_/B sky130_fd_sc_hd__clkbuf_2
Xhold716 hold716/A VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold727 hold727/A VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold738 hold738/A VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6241_ _7180_/Q _6240_/X _6341_/S VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3453_ _6930_/Q _5344_/A _5515_/A _7082_/Q _3452_/X VGND VGND VPWR VPWR _3461_/B
+ sky130_fd_sc_hd__a221oi_1
XFILLER_115_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5695__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2527_A _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6172_ _6915_/Q _5991_/X _5996_/X _7051_/Q _6171_/X VGND VGND VPWR VPWR _6179_/A
+ sky130_fd_sc_hd__a221o_1
X_3384_ _3384_/A _3384_/B _3383_/Y VGND VGND VPWR VPWR _3385_/B sky130_fd_sc_hd__nor3b_4
Xhold2106 _6482_/Q VGND VGND VPWR VPWR hold723/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2117 _4285_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5123_ _5123_/A _5123_/B _5123_/C _5123_/D VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__and4_1
Xhold2128 _5526_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2139 hold545/X VGND VGND VPWR VPWR _5445_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1405 _7078_/Q VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1416 _5484_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1427 hold1427/A VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1438 _6838_/Q VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5054_ _4638_/Y _4698_/Y _4689_/Y _5063_/B VGND VGND VPWR VPWR _5054_/X sky130_fd_sc_hd__o211a_1
XFILLER_38_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1449 _5383_/X VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4005_ hold857/X _5189_/A1 _4008_/S VGND VGND VPWR VPWR _4005_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5956_ _6573_/Q _5674_/X _5680_/X _6711_/Q VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ _4907_/A1 _5139_/A _4906_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__5785__B _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5887_ _6635_/Q _5671_/X _5886_/X VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3630__C1 _3389_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5277__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4838_ _4917_/C _4838_/B VGND VGND VPWR VPWR _4857_/C sky130_fd_sc_hd__nor2_1
XANTENNA__6175__B2 _6875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5922__A1 _6586_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4769_ _5011_/A _4729_/A _4514_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__a21oi_1
X_6508_ _7106_/CLK _6508_/D fanout472/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6439_ net399_2/A _6439_/D _6394_/X VGND VGND VPWR VPWR _6439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__buf_2
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2640 _5503_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2651 hold703/X VGND VGND VPWR VPWR _5173_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2662 _6960_/Q VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__buf_8
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2673 _4320_/X VGND VGND VPWR VPWR hold798/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__buf_2
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4110__A0 _3675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2684 _4299_/X VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1950 _5366_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2695 _4126_/X VGND VGND VPWR VPWR hold789/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1961 _6964_/Q VGND VGND VPWR VPWR hold344/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1996_A _7118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1972 _6877_/Q VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1983 _7016_/Q VGND VGND VPWR VPWR hold813/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1994 _4032_/X VGND VGND VPWR VPWR hold888/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3240__1 net399_2/A VGND VGND VPWR VPWR _6436_/CLK sky130_fd_sc_hd__inv_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3767__A3 hold47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4091__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 _3748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output264_A _6786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5141__A2 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4101__A0 _3675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3455__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5810_ _6938_/Q _5659_/X _5687_/X _6922_/Q VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _6793_/CLK _6790_/D fanout434/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5741_ _6911_/Q _5670_/X _5685_/X _7071_/Q VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _5685_/A _5689_/B _5689_/C VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__and3b_4
X_4623_ _4625_/A _4971_/A VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ _4637_/B _4590_/B _5033_/A _4959_/A _4553_/Y VGND VGND VPWR VPWR _4554_/X
+ sky130_fd_sc_hd__a311o_1
Xhold502 hold502/A VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold513 hold513/A VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold524 hold524/A VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3505_ _3544_/A _3553_/B VGND VGND VPWR VPWR _4122_/A sky130_fd_sc_hd__nor2_4
Xhold535 hold535/A VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold546 hold546/A VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4485_ _4486_/A _4485_/B _4568_/A VGND VGND VPWR VPWR _4621_/A sky130_fd_sc_hd__and3_2
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold568 hold568/A VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold579 hold579/A VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6224_ _6589_/Q _5985_/X _5994_/X _6634_/Q _6218_/X VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a221o_1
X_3436_ _6850_/Q _5254_/A _3431_/Y _7233_/A VGND VGND VPWR VPWR _3436_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5236__A_N _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6155_ _7130_/Q _5973_/X _5988_/X _6874_/Q _6154_/X VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _6972_/Q _5389_/A _5308_/A _6900_/Q _3366_/X VGND VGND VPWR VPWR _3368_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1202 _7229_/A VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5106_ _4569_/A _4523_/Y _4583_/B _4688_/C _4871_/A VGND VGND VPWR VPWR _5107_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _6935_/Q VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _6806_/Q VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6086_ _6927_/Q _5982_/X _5987_/X _7111_/Q VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__a22o_1
Xhold1235 _5393_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3298_ hold79/X hold14/X VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__nand2_8
Xhold1246 _7110_/Q VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6093__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1257 hold395/X VGND VGND VPWR VPWR _5420_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5037_ _5117_/C _5151_/B _5037_/C VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__and3_1
XFILLER_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout462_A fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1268 _6879_/Q VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1279 hold369/X VGND VGND VPWR VPWR _5303_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3446__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5840__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6988_ _7082_/CLK _6988_/D fanout464/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3603__C1 _3602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5939_ _6551_/Q _5673_/X _5937_/X _5938_/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6404__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input162_A wb_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4345_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4649_/B sky130_fd_sc_hd__buf_12
XFILLER_163_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6367_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6373_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6380_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6356_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2470 _7132_/Q VGND VGND VPWR VPWR hold419/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2481 _3987_/X VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input23_A mask_rev_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6084__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4086__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2492 hold674/X VGND VGND VPWR VPWR _4181_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3437__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5831__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1780 hold434/X VGND VGND VPWR VPWR hold1780/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1791 hold992/X VGND VGND VPWR VPWR hold480/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4937__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3954__A _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5898__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3373__B2 _3973_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A0 _5580_/A1 _4273_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3221_ _6984_/Q VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6075__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5822__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6911_ _6967_/CLK _6911_/D fanout465/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4009__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6842_ _7084_/CLK _6842_/D fanout447/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6773_ _6809_/CLK _6773_/D fanout433/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfrtp_4
X_3985_ _3985_/A0 _5195_/A1 _3987_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _7046_/Q _5669_/X _5680_/X _6958_/Q _5723_/X VGND VGND VPWR VPWR _5727_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3600__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5655_ _5689_/A _5679_/B _5687_/C VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__and3_4
XANTENNA__5555__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5889__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4606_ _4625_/A _4611_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nand2_2
X_5586_ hold92/X hold71/X _5586_/S VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3364__A1 _6996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold321 hold321/A VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4537_ _4601_/A _4570_/C _4535_/X _4536_/Y VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3364__B2 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold332 hold332/A VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold365 hold365/A VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6302__A1 _6607_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4468_ _4638_/B _4488_/B VGND VGND VPWR VPWR _4601_/A sky130_fd_sc_hd__nand2_8
XANTENNA__6302__B2 _6710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold387 hold387/A VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold398 hold398/A VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6207_ _7100_/Q _5984_/X _6015_/X _7020_/Q VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__a22o_1
X_3419_ _7003_/Q _5425_/A _5506_/A _7075_/Q VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7187_ _7194_/CLK _7187_/D VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfxtp_1
X_4399_ _4637_/D _4574_/A VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__and2b_4
XANTENNA__3667__A2 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6131_/X _6133_/X _6138_/C _6339_/B VGND VGND VPWR VPWR _6139_/C sky130_fd_sc_hd__and4bb_2
Xhold1010 hold41/X VGND VGND VPWR VPWR _3984_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1021 hold11/X VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _5482_/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _3986_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 hold1054/A VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6069_ _6911_/Q _5991_/X _6018_/X _6967_/Q VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _5212_/X VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3419__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 _3295_/Y VGND VGND VPWR VPWR _5578_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5813__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 hold54/X VGND VGND VPWR VPWR _3259_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 _6646_/Q VGND VGND VPWR VPWR hold188/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5465__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3658__A2 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6057__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5804__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5280__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _3770_/A _3770_/B _3770_/C VGND VGND VPWR VPWR _3803_/A sky130_fd_sc_hd__and3_2
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3594__A1 _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5375__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5440_ _5440_/A0 _5575_/A1 _5442_/S VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5371_/A _5578_/B VGND VGND VPWR VPWR _5379_/S sky130_fd_sc_hd__and2_4
X_7110_ _7124_/CLK _7110_/D fanout467/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfstp_2
X_4322_ _4322_/A _5533_/B VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__and2_4
XFILLER_113_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6296__B1 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold31_A hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7041_ _7137_/CLK _7041_/D fanout466/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
X_4253_ _4253_/A0 _5194_/A1 _4255_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3649__A2 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3204_ _7120_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__4846__B2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4184_ _4184_/A0 _5238_/A1 _4187_/S VGND VGND VPWR VPWR _4184_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6048__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5271__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6825_ _7125_/CLK _6825_/D fanout468/X VGND VGND VPWR VPWR _7230_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_51_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6220__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3968_ _3968_/A _3975_/B VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__and2_1
X_6756_ _6756_/CLK _6756_/D fanout454/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3585__A1 _6572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5707_ _6837_/Q _5707_/B VGND VGND VPWR VPWR _5707_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__3585__B2 _6607_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6687_ _6701_/CLK _6687_/D fanout436/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_4
X_3899_ _4345_/A _4345_/B _3899_/C _3899_/D VGND VGND VPWR VPWR _3900_/D sky130_fd_sc_hd__and4bb_2
XANTENNA__5285__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1275_A _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5638_ _6014_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__and3_4
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5569_ _5569_/A _5569_/B VGND VGND VPWR VPWR _5577_/S sky130_fd_sc_hd__and2_4
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3888__A2 _6434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold140 _5311_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold173 hold173/A VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold195 hold195/A VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1707_A _6901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A wb_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6211__B1 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input90_A spimemio_flash_io2_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3576__A1 _6944_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3576__B2 _6807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5195__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7148__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6643__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6278__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5253__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4940_ _4462_/Y _4935_/X _4796_/A VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__o21a_1
XFILLER_33_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4871_ _4871_/A _4871_/B _4871_/C _4871_/D VGND VGND VPWR VPWR _4872_/D sky130_fd_sc_hd__and4_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6202__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _6745_/CLK _6610_/D fanout441/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
X_3822_ hold52/A hold19/A _3834_/S VGND VGND VPWR VPWR _3826_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_21_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3567__A1 _6888_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6541_ _7194_/CLK _6541_/D VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6821_/Q _5226_/A _5226_/B _3315_/Y input34/X VGND VGND VPWR VPWR _3753_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3567__B2 _6582_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2557_A _7021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6472_ _6486_/CLK _6472_/D fanout433/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_173_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ _3684_/A _3684_/B _3684_/C VGND VGND VPWR VPWR _3704_/A sky130_fd_sc_hd__nor3_1
XFILLER_146_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ _5423_/A0 _5549_/A1 _5424_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
Xoutput201 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput223 _7218_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
XFILLER_161_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput234 _7228_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ _5354_/A0 _5534_/A1 _5361_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput245 _3942_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_99_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput256 _3963_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _6782_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
XANTENNA__6269__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4305_ _4305_/A0 _5237_/A1 _4309_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput278 _6795_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
X_5285_ _5285_/A0 _5537_/A1 _5289_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
Xoutput289 _6481_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_87_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7024_ _7133_/CLK _7024_/D fanout468/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4236_ _4236_/A0 _4235_/X _4240_/S VGND VGND VPWR VPWR _4236_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5492__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4167_ _4167_/A0 _5581_/A1 _4169_/S VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4098_ _6678_/Q _6346_/B VGND VGND VPWR VPWR _4106_/S sky130_fd_sc_hd__nand2_8
XANTENNA__5244__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk _6549_/CLK VGND VGND VPWR VPWR _6830_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6808_ _6826_/CLK _6808_/D _6407_/A VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_1
X_6739_ _6803_/CLK _6739_/D fanout449/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6412__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3730__B2 _6785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3263__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout450 fanout454/X VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__buf_12
XFILLER_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout461 fanout465/X VGND VGND VPWR VPWR fanout461/X sky130_fd_sc_hd__buf_12
XANTENNA__5483__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout472 fanout473/X VGND VGND VPWR VPWR fanout472/X sky130_fd_sc_hd__buf_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3494__B1 _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5786__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3797__A1 _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output294_A _6486_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5219__A _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _5237_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3962__A _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5710__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3721__B2 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2138_A _7014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5070_ _4476_/X _4568_/Y _4920_/B _4972_/Y VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__o211a_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 _5406_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5474__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4021_ _4021_/A0 _4020_/X _4029_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5972_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6018_/B sky130_fd_sc_hd__nor2_4
XFILLER_53_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5777__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3202__A _7136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3788__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3788__B2 _6525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4923_ _4633_/B _4691_/Y _4846_/X _4894_/B VGND VGND VPWR VPWR _5052_/B sky130_fd_sc_hd__o211a_1
XFILLER_33_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4569_/A _4655_/A _4590_/Y _4688_/C VGND VGND VPWR VPWR _4871_/B sky130_fd_sc_hd__o22a_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3805_ _3805_/A1 _3739_/S _3803_/Y _3804_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__a22o_1
X_4785_ _4718_/A _4463_/B _4570_/D _4691_/Y _4947_/A VGND VGND VPWR VPWR _4785_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6524_ _7106_/CLK hold83/X fanout472/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
X_3736_ _3707_/X _3736_/B _3736_/C _3736_/D VGND VGND VPWR VPWR _3737_/B sky130_fd_sc_hd__and4b_4
XFILLER_174_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3667_ _6855_/Q _5263_/A _4334_/A _6759_/Q VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__a22o_1
X_6455_ _3940_/A1 _6455_/D _6405_/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5563__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5406_ _5406_/A0 _5577_/A1 _5406_/S VGND VGND VPWR VPWR _5406_/X sky130_fd_sc_hd__mux2_1
X_6386_ _3969_/A _6356_/Y _6358_/Y _3967_/A VGND VGND VPWR VPWR _6386_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__5701__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3598_ _7048_/Q hold16/A _5169_/A _6772_/Q VGND VGND VPWR VPWR _3598_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6651__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ _5337_/A0 _5580_/A1 _5343_/S VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2800 _5314_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2811 _5522_/X VGND VGND VPWR VPWR hold716/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2822 _7010_/Q VGND VGND VPWR VPWR hold956/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5268_ _5268_/A0 _5448_/A1 _5271_/S VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__mux2_1
Xhold2833 _6994_/Q VGND VGND VPWR VPWR hold951/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5465__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2844 _7090_/Q VGND VGND VPWR VPWR hold959/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2855 _6775_/Q VGND VGND VPWR VPWR _3739_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4219_ _6682_/Q _4220_/B VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__and2b_4
X_7007_ _7135_/CLK _7007_/D fanout466/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2866 _7175_/Q VGND VGND VPWR VPWR _6116_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2877 _7166_/Q VGND VGND VPWR VPWR _5859_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5199_ _5199_/A0 _5577_/A1 _5199_/S VGND VGND VPWR VPWR _5199_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3476__B1 _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2888 _6655_/Q VGND VGND VPWR VPWR _3920_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2899 _7200_/Q VGND VGND VPWR VPWR _6378_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5217__A1 _5228_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5768__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6193__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3400__B1 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5940__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3951__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5473__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4597__B _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A mgmt_gpio_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4089__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5456__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5208__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5759__A2 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3957__A _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6184__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4195__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ _4570_/A _4570_/B _4570_/C _4570_/D VGND VGND VPWR VPWR _4570_/X sky130_fd_sc_hd__and4_1
XANTENNA__5931__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3521_ hold56/X _3533_/B VGND VGND VPWR VPWR _3521_/Y sky130_fd_sc_hd__nor2_8
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap425 _4808_/A VGND VGND VPWR VPWR _4726_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5383__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold717 hold717/A VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold728 hold728/A VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6240_ _6525_/Q _6339_/B _6239_/X VGND VGND VPWR VPWR _6240_/X sky130_fd_sc_hd__o21ba_1
XFILLER_170_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3452_ _6866_/Q _5272_/A _5389_/A _6970_/Q _3451_/X VGND VGND VPWR VPWR _3452_/X
+ sky130_fd_sc_hd__a221o_1
Xhold739 hold739/A VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5695__A1 _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7027_/Q _5971_/X _6014_/X _6995_/Q VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__a22o_1
X_3383_ _3383_/A _3383_/B _3383_/C _3383_/D VGND VGND VPWR VPWR _3383_/Y sky130_fd_sc_hd__nor4_1
XANTENNA_hold2422_A _6643_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2107 hold723/X VGND VGND VPWR VPWR _4004_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5122_ _4491_/Y _4523_/Y _4583_/B _4676_/Y _4872_/C VGND VGND VPWR VPWR _5123_/D
+ sky130_fd_sc_hd__o221a_1
Xhold2118 _7121_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2129 _7005_/Q VGND VGND VPWR VPWR hold750/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5447__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1406 hold263/X VGND VGND VPWR VPWR _5517_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1417 _6805_/Q VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5053_ _5112_/B _5121_/C _5112_/C _5107_/B VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__and4_1
Xhold1428 _5399_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1439 hold265/X VGND VGND VPWR VPWR _5247_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3458__B1 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4004_ _4004_/A0 _5195_/A1 _4008_/S VGND VGND VPWR VPWR _4004_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5955_ _6696_/Q _5658_/X _5664_/X _6761_/Q VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5558__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _4906_/A _4906_/B _4906_/C _4906_/D VGND VGND VPWR VPWR _4906_/X sky130_fd_sc_hd__and4_1
XANTENNA__3630__B1 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5886_ _6748_/Q _5666_/X _5689_/X _6625_/Q VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6746__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4837_ _5114_/A _4837_/B VGND VGND VPWR VPWR _5044_/B sky130_fd_sc_hd__and2_1
XANTENNA__6175__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4186__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4768_ _5033_/A _4955_/D VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5922__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3933__A1 input92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6507_ _7106_/CLK _6507_/D fanout472/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_1
X_3719_ _6902_/Q _5317_/A _5281_/A _6870_/Q VGND VGND VPWR VPWR _3719_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5293__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4699_ _4710_/A _4702_/B VGND VGND VPWR VPWR _4699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ net399_2/A _6438_/D _6393_/X VGND VGND VPWR VPWR _6438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6369_ _6368_/X _6369_/A1 _6384_/S VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3697__B1 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1522_A _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6977_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5438__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2630 hold737/X VGND VGND VPWR VPWR _5468_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__buf_4
Xhold2641 _7225_/A VGND VGND VPWR VPWR hold822/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2652 _5173_/X VGND VGND VPWR VPWR hold704/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2663 hold833/X VGND VGND VPWR VPWR _5384_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2674 _6873_/Q VGND VGND VPWR VPWR hold689/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2685 _6866_/Q VGND VGND VPWR VPWR hold946/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1940 hold289/X VGND VGND VPWR VPWR _5378_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1951 _6515_/Q VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2696 _6769_/Q VGND VGND VPWR VPWR hold672/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__buf_6
Xhold1962 hold344/X VGND VGND VPWR VPWR _5388_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7099_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1973 _6878_/Q VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1984 hold813/X VGND VGND VPWR VPWR _5447_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1995 hold888/X VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5976__B _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5468__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__B1 _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4716__A3 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5913__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 _3769_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output257_A _6792_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7204__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5378__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5740_ _7063_/Q _5671_/X _5733_/X _5735_/X _5739_/X VGND VGND VPWR VPWR _5740_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_188_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3612__B1 _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5671_ _5689_/A _5679_/B _5689_/C VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__and3_4
XANTENNA__6157__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6213__D _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4622_ _4894_/B _4622_/B _4622_/C _5052_/A VGND VGND VPWR VPWR _4622_/X sky130_fd_sc_hd__and4_1
XFILLER_129_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ _4514_/Y _4526_/X _4553_/C _5090_/C VGND VGND VPWR VPWR _4553_/Y sky130_fd_sc_hd__nand4bb_1
XFILLER_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold503 hold503/A VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5407__A _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold525 hold525/A VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3504_ hold56/X _3549_/B VGND VGND VPWR VPWR _4146_/A sky130_fd_sc_hd__nor2_4
Xhold536 hold536/A VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4484_ _4607_/B _4611_/A VGND VGND VPWR VPWR _4531_/B sky130_fd_sc_hd__nand2_2
Xhold547 hold547/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold558 hold558/A VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3435_ input17/X _3310_/Y _4000_/A _6484_/Q VGND VGND VPWR VPWR _3435_/X sky130_fd_sc_hd__a22o_4
X_6223_ _6702_/Q _5977_/X _5984_/X _6614_/Q _6222_/X VGND VGND VPWR VPWR _6238_/B
+ sky130_fd_sc_hd__a221o_4
Xhold569 hold569/A VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6962_/Q _5992_/X _6012_/X _7002_/Q _6153_/X VGND VGND VPWR VPWR _6154_/X
+ sky130_fd_sc_hd__a221o_1
X_3366_ _7140_/Q _3295_/Y _5335_/A _6924_/Q VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__a22o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1203 hold73/X VGND VGND VPWR VPWR _4249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5105_ _5101_/X _5135_/D _5062_/A _5071_/Y VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__a211o_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 hold235/X VGND VGND VPWR VPWR _5356_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6085_ _6863_/Q _5999_/X _6019_/X _6983_/Q _6084_/X VGND VGND VPWR VPWR _6088_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1225 hold243/X VGND VGND VPWR VPWR _5205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3297_ hold13/X hold46/A VGND VGND VPWR VPWR _3297_/Y sky130_fd_sc_hd__nor2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 _7076_/Q VGND VGND VPWR VPWR _5514_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5036_ _4812_/A _4724_/C _5033_/A VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__o21ai_1
Xhold1247 hold138/X VGND VGND VPWR VPWR _5553_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6093__B2 _7080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1258 _5420_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1269 hold132/X VGND VGND VPWR VPWR _5293_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5840__B2 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout455_A _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5796__B _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6987_ _7082_/CLK _6987_/D fanout464/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5288__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3603__B1 _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5938_ _6612_/Q _5660_/X _5669_/X _6652_/Q VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5869_ _5869_/A _5869_/B _5869_/C VGND VGND VPWR VPWR _5869_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__6148__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4159__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5317__A _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3382__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4221__A _6678_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7181__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6320__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4331__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input155_A wb_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4345_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6370_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6376_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3271__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2460 _5225_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6382_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6358_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2471 hold419/X VGND VGND VPWR VPWR _5577_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6084__B2 _7015_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2482 _7133_/Q VGND VGND VPWR VPWR hold854/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2493 _4181_/X VGND VGND VPWR VPWR hold675/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1770 hold978/X VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5831__A1 _6851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input16_A mask_rev_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1781 _6568_/Q VGND VGND VPWR VPWR hold983/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1792 hold480/X VGND VGND VPWR VPWR hold1792/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5198__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3373__A2 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6311__A2 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3970__A _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3220_ _6992_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_141_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4873__A2 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7185_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6075__A1 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6075__B2 _6887_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2218_A _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4086__A0 _3675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5822__A1 _6963_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6910_ _7126_/CLK _6910_/D fanout453/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6841_ _7073_/CLK _6841_/D fanout444/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6772_ _6803_/CLK _6772_/D fanout442/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_4
X_3984_ _3984_/A0 _7198_/Q _3998_/S VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3210__A _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5050__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5723_ _7014_/Q _5664_/X _5668_/X _7054_/Q VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2754_A _6795_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5654_ _7148_/Q _7149_/Q VGND VGND VPWR VPWR _5687_/C sky130_fd_sc_hd__and2b_4
XFILLER_190_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4605_ _4580_/Y _4969_/B _4584_/Y _4604_/X VGND VGND VPWR VPWR _4609_/C sky130_fd_sc_hd__a31o_1
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5585_ _5585_/A0 wire371/X _5586_/S VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 hold300/A VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold311 hold311/A VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3364__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4536_ _4607_/B _4562_/A VGND VGND VPWR VPWR _4536_/Y sky130_fd_sc_hd__nand2_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7197__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold333 hold333/A VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold344 hold344/A VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold355 hold355/A VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4467_ _4638_/B _4488_/B VGND VGND VPWR VPWR _4934_/B sky130_fd_sc_hd__and2_4
XANTENNA__5571__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6302__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold377 hold377/A VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold388 hold388/A VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4313__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6206_ _7052_/Q _5996_/X _6005_/X _6948_/Q _6205_/X VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a221o_1
X_3418_ _6923_/Q _5335_/A _5353_/A _6939_/Q _3417_/X VGND VGND VPWR VPWR _3421_/C
+ sky130_fd_sc_hd__a221o_1
X_4398_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4495_/B sky130_fd_sc_hd__nand2_8
X_7186_ _7203_/CLK _7186_/D _4107_/B VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input8_A mask_rev_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 _4109_/A1 VGND VGND VPWR VPWR hold1877/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6137_ _7041_/Q _6016_/X _6134_/X _6136_/X VGND VGND VPWR VPWR _6138_/C sky130_fd_sc_hd__a211oi_1
X_3349_ _3349_/A hold15/X VGND VGND VPWR VPWR _5407_/A sky130_fd_sc_hd__nor2_8
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1011 _3984_/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1022 _6462_/Q VGND VGND VPWR VPWR _3840_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1033 hold18/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_133_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 hold94/X VGND VGND VPWR VPWR hold1044/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6068_ _6855_/Q _5983_/X _6005_/X _6943_/Q VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__a22o_1
Xhold1055 _5559_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1066 _6617_/Q VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _5578_/X VGND VGND VPWR VPWR _5586_/S sky130_fd_sc_hd__clkdlybuf4s50_2
X_5019_ _4826_/B _4990_/Y _5018_/X _4683_/A VGND VGND VPWR VPWR _5022_/C sky130_fd_sc_hd__o2bb2a_1
Xhold1088 _3259_/X VGND VGND VPWR VPWR _3284_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 hold188/X VGND VGND VPWR VPWR _4209_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6415__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3266__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5481__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4855__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2290 _5448_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5804__B2 _7018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3594__A2 _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5370_ _5370_/A0 _5568_/A1 _5370_/S VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4321_ _4321_/A0 _5448_/A1 _4321_/S VGND VGND VPWR VPWR _4321_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5391__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6296__A1 _6715_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7040_ _7136_/CLK _7040_/D fanout467/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_4
X_4252_ _4252_/A0 _5193_/A1 _4255_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6296__B2 _6642_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3203_ _7128_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4846__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold24_A hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4183_ _4183_/A0 _5543_/A1 _4187_/S VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3205__A _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6048__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6048__B2 _6942_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6824_ _6826_/CLK _6824_/D _6407_/A VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _6756_/CLK _6755_/D fanout441/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_4
X_3967_ _3967_/A _3969_/B VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5566__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5706_ _6973_/Q _5660_/X _5699_/X _5701_/X _5705_/X VGND VGND VPWR VPWR _5706_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3585__A2 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6686_ _3950_/A1 _6686_/D _4107_/B VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3898_ _3898_/A _3898_/B _3898_/C VGND VGND VPWR VPWR _3899_/D sky130_fd_sc_hd__and3_1
XFILLER_12_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5637_ _5637_/A _7156_/Q VGND VGND VPWR VPWR _6019_/B sky130_fd_sc_hd__nor2_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5731__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5568_ _5568_/A0 _5568_/A1 _5568_/S VGND VGND VPWR VPWR _5568_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold141 hold141/A VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4519_ _4637_/D _4522_/B VGND VGND VPWR VPWR _4917_/D sky130_fd_sc_hd__nor2_8
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold152 hold152/A VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5499_ _5499_/A0 _5571_/A1 _5505_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold163 hold163/A VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold174 _7197_/Q VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__A1 _6452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold185 _4050_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold196 hold196/A VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7169_ _7184_/CLK _7169_/D fanout443/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5798__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A wb_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6211__A1 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5476__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3576__A2 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4773__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input83_A spimemio_flash_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5722__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6278__B2 _6532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5789__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _4870_/A _4870_/B _4870_/C _4870_/D VGND VGND VPWR VPWR _4871_/D sky130_fd_sc_hd__and4_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6202__B2 _6852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3821_ hold60/A _6462_/Q _6461_/Q _6460_/Q VGND VGND VPWR VPWR _3834_/S sky130_fd_sc_hd__and4_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5386__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3567__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6540_ _7194_/CLK _6540_/D VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5961__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3752_ _6909_/Q _5326_/A _4316_/A _6742_/Q _3751_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6471_ _6486_/CLK _6471_/D fanout433/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfstp_2
X_3683_ input12/X _3310_/Y _5169_/A _6770_/Q _3682_/X VGND VGND VPWR VPWR _3684_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2452_A _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5422_ _5422_/A0 _5575_/A1 _5424_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5713__B1 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _3205_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
XFILLER_145_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput213 _3946_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput224 _7219_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
XFILLER_99_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput235 _7229_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
X_5353_ _5353_/A _5533_/B VGND VGND VPWR VPWR _5361_/S sky130_fd_sc_hd__and2_4
Xoutput246 _7211_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
Xoutput257 _6792_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A _5220_/C VGND VGND VPWR VPWR _4309_/S sky130_fd_sc_hd__and2_2
Xoutput268 _6789_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
XANTENNA__6269__B2 _6719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput279 _6796_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_99_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5284_ _5284_/A0 _5572_/A1 _5289_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4819__A2 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7023_ _7125_/CLK _7023_/D fanout468/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4235_ _5242_/A0 wire375/X _5236_/C VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4166_ _4166_/A0 _5238_/A1 _4169_/S VGND VGND VPWR VPWR _4166_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4097_ _4097_/A0 _5277_/A1 _4097_/S VGND VGND VPWR VPWR _4097_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout368_A wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6611__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6807_ _6815_/CLK _6807_/D fanout443/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _5010_/B _4999_/B _5139_/B _4999_/D VGND VGND VPWR VPWR _5000_/B sky130_fd_sc_hd__and4_1
XANTENNA__5296__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6738_ _6803_/CLK _6738_/D fanout449/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5952__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6669_ _7125_/CLK _6669_/D fanout468/X VGND VGND VPWR VPWR _7223_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5704__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5180__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3730__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout440 fanout454/X VGND VGND VPWR VPWR fanout440/X sky130_fd_sc_hd__buf_12
Xfanout451 fanout453/X VGND VGND VPWR VPWR fanout451/X sky130_fd_sc_hd__buf_12
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout462 fanout465/X VGND VGND VPWR VPWR fanout462/X sky130_fd_sc_hd__buf_12
Xfanout473 input75/X VGND VGND VPWR VPWR fanout473/X sky130_fd_sc_hd__buf_12
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3494__A1 input30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3494__B2 _6643_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4994__A1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3797__A2 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6196__B1 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5943__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3962__B _3962_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5171__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3721__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6120__B1 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4020_ _6512_/Q _5537_/A1 _4047_/C VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2033_A _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3485__B2 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5971_ _6015_/B _6014_/A _6019_/B VGND VGND VPWR VPWR _5971_/X sky130_fd_sc_hd__and3_4
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3788__A2 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4922_ _4922_/A _4922_/B _4922_/C VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__and3_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4510_/A _4655_/A _4590_/Y _4995_/A VGND VGND VPWR VPWR _4924_/C sky130_fd_sc_hd__o22a_1
XFILLER_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3804_ _6448_/Q _6656_/Q _3857_/B VGND VGND VPWR VPWR _3804_/X sky130_fd_sc_hd__and3_1
XANTENNA__5934__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4784_ _4466_/A _4477_/Y _4510_/B _4736_/Y _4407_/Y VGND VGND VPWR VPWR _4784_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_165_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6523_ _7106_/CLK _6523_/D fanout472/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3735_ _3735_/A _3735_/B _3735_/C _3735_/D VGND VGND VPWR VPWR _3736_/D sky130_fd_sc_hd__nor4_1
XFILLER_118_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6454_ _6733_/CLK _6454_/D fanout433/X VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_4
X_3666_ _7127_/Q _5569_/A _5344_/A _6927_/Q _3665_/X VGND VGND VPWR VPWR _3673_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5698__C1 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5405_ _5405_/A0 _5549_/A1 _5406_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6385_ _3184_/Y _3189_/Y _6385_/A3 _4836_/A _4222_/Y VGND VGND VPWR VPWR _7203_/D
+ sky130_fd_sc_hd__a41o_2
X_3597_ _6474_/Q _3988_/A _4322_/A _6750_/Q _3596_/X VGND VGND VPWR VPWR _3604_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5336_ hold786/X _5561_/A1 _5343_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2801 _6821_/Q VGND VGND VPWR VPWR hold913/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2812 _6867_/Q VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6111__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5267_ _5267_/A0 _5303_/A1 _5271_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
Xhold2823 hold956/X VGND VGND VPWR VPWR _5440_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2834 hold951/X VGND VGND VPWR VPWR _5422_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7006_ _7078_/CLK _7006_/D fanout445/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfstp_1
Xhold2845 hold959/X VGND VGND VPWR VPWR _5530_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4218_ _6684_/Q _6685_/Q _6686_/Q VGND VGND VPWR VPWR _4218_/Y sky130_fd_sc_hd__nor3_4
Xhold2856 _3739_/X VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2867 _6092_/X VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2878 _5838_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5198_ _5198_/A0 _5549_/A1 _5199_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2889 _3920_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4195__S _4199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4149_ _4149_/A0 _5527_/A1 _4151_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3779__A2 hold64/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6178__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6423__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3400__A1 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3400__B2 _6843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4878__B _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6350__A0 _3616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input46_A mgmt_gpio_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_64_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3957__B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4134__A _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5916__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5392__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6655__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3520_ _7137_/Q _3295_/Y _5290_/A _6881_/Q VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap415 _4700_/B VGND VGND VPWR VPWR _4698_/C sky130_fd_sc_hd__clkbuf_2
Xhold707 hold707/A VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap426 _4580_/A VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__clkbuf_2
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold729 hold729/A VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3451_ _6978_/Q _5398_/A _5524_/A _7090_/Q _3450_/X VGND VGND VPWR VPWR _3451_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5695__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3382_ _6932_/Q _5344_/A _5263_/A _6860_/Q _3381_/X VGND VGND VPWR VPWR _3383_/D
+ sky130_fd_sc_hd__a221o_1
X_6170_ _7099_/Q _5984_/X _5997_/X _6955_/Q _6169_/X VGND VGND VPWR VPWR _6170_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk _6549_/CLK VGND VGND VPWR VPWR _6826_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5121_/A _5121_/B _5121_/C _5121_/D VGND VGND VPWR VPWR _5121_/X sky130_fd_sc_hd__and4_2
Xhold2108 _4004_/X VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2119 hold783/X VGND VGND VPWR VPWR _5565_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1407 _5517_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1418 hold255/X VGND VGND VPWR VPWR _5204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5052_ _5052_/A _5052_/B _5052_/C VGND VGND VPWR VPWR _5107_/B sky130_fd_sc_hd__and3_1
Xhold1429 _7224_/A VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4003_ hold513/X _5194_/A1 _4008_/S VGND VGND VPWR VPWR _4003_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3213__A _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5954_ _6583_/Q _5688_/X _5952_/X _5953_/X VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__a211o_1
XFILLER_179_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4905_ _4601_/A _4523_/Y _4491_/Y VGND VGND VPWR VPWR _4905_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5885_ _3200_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5885_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3630__A1 _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3630__B2 _6791_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4836_ _4836_/A _4836_/B VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5907__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5383__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4767_ _4767_/A _4880_/B VGND VGND VPWR VPWR _4933_/C sky130_fd_sc_hd__and2_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5574__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6506_ _7086_/CLK _6506_/D fanout467/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3394__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_A hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3718_ _6815_/Q hold24/A _3431_/Y input62/X _3717_/X VGND VGND VPWR VPWR _3725_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4698_ _4712_/A _4712_/B _4698_/C VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nand3_4
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6437_ _3958_/A1 _6437_/D _6392_/X VGND VGND VPWR VPWR _6437_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6332__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3649_ _6734_/Q _4304_/A _3648_/Y _6818_/Q VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6368_ _6684_/Q _6368_/A2 _6368_/B1 _4218_/Y _6367_/X VGND VGND VPWR VPWR _6368_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3697__A1 _7086_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3697__B2 _7038_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5319_ hold589/X _5562_/A1 _5325_/S VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__mux2_1
X_6299_ _6538_/Q _5983_/X _5993_/X _6622_/Q _6298_/X VGND VGND VPWR VPWR _6304_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2620 _4198_/X VGND VGND VPWR VPWR hold779/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1515_A _6852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2631 _5468_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__buf_12
Xhold2642 hold822/X VGND VGND VPWR VPWR _4245_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2653 _6610_/Q VGND VGND VPWR VPWR hold535/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2664 _5384_/X VGND VGND VPWR VPWR hold834/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__buf_12
Xhold1930 _5342_/X VGND VGND VPWR VPWR hold284/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2675 hold689/X VGND VGND VPWR VPWR _5286_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2686 hold946/X VGND VGND VPWR VPWR _5278_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1941 _5378_/X VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1952 hold280/X VGND VGND VPWR VPWR _4054_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2697 hold672/X VGND VGND VPWR VPWR _5170_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1963 _5388_/X VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1974 hold507/X VGND VGND VPWR VPWR _5292_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1985 _5447_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1996 _7118_/Q VGND VGND VPWR VPWR hold564/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input100_A wb_adr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3621__A1 _6786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3269__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6678__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5374__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5484__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _3765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6323__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4885__B1 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3860__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3612__A1 _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B2 _6592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5685_/A _5686_/B _5687_/C VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__and3b_4
XFILLER_175_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4621_ _4621_/A _5048_/A VGND VGND VPWR VPWR _5052_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5365__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5394__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3376__B1 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ _5009_/A _4552_/B VGND VGND VPWR VPWR _5090_/C sky130_fd_sc_hd__nand2_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3503_ _6583_/Q _4128_/A _4334_/A _6761_/Q _3502_/X VGND VGND VPWR VPWR _3515_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5407__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4483_ _4486_/A _4483_/B VGND VGND VPWR VPWR _4570_/D sky130_fd_sc_hd__nand2_8
XFILLER_171_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold537 hold537/A VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3208__A _7088_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold548 hold548/A VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold559 hold559/A VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6222_ _6604_/Q _5982_/X _5987_/X _6727_/Q VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3434_ input8/X _3315_/Y _3336_/Y input25/X VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__a22o_4
XANTENNA__3679__A1 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3679__B2 _6713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6954_/Q _5997_/X _6004_/X _6882_/Q VGND VGND VPWR VPWR _6153_/X sky130_fd_sc_hd__a22o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _6980_/Q _5398_/A _3315_/Y input10/X _3362_/X VGND VGND VPWR VPWR _3368_/C
+ sky130_fd_sc_hd__a221o_2
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _4976_/B _4976_/A _5104_/C _5104_/D VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__and4bb_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _4249_/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _7087_/Q _5638_/X _6015_/X _7015_/Q VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__a22o_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _5356_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3296_ _3338_/A _3354_/B VGND VGND VPWR VPWR _5344_/A sky130_fd_sc_hd__nor2_8
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _5205_/X VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1237 _5514_/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6093__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5035_ _4683_/A _5029_/X _4961_/D _4529_/B VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__o211a_1
Xhold1248 _5553_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1259 _6937_/Q VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5840__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6986_ _7112_/CLK _6986_/D fanout473/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout448_A fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5937_ _6572_/Q _5674_/X _5680_/X _6710_/Q VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3603__B2 _6453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6967__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5868_ _6752_/Q _5681_/X _5865_/X _5867_/X VGND VGND VPWR VPWR _5869_/C sky130_fd_sc_hd__a211o_1
XANTENNA__6002__C1 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4819_ _4658_/A _4633_/B _4683_/A _4727_/Y _4818_/X VGND VGND VPWR VPWR _4820_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5356__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5799_ _6850_/Q _5653_/X _5662_/X _6898_/Q _5798_/X VGND VGND VPWR VPWR _5799_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1465_A _6811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3367__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5317__B _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6305__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1632_A _6532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4344_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4649_/D sky130_fd_sc_hd__clkbuf_4
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4637_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input148_A wb_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6374_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6379_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2450 hold835/X VGND VGND VPWR VPWR _5457_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6371_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2461 _6569_/Q VGND VGND VPWR VPWR hold881/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6357_/A sky130_fd_sc_hd__clkbuf_2
Xhold2472 _5577_/X VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6084__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4095__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2483 _6861_/Q VGND VGND VPWR VPWR hold917/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2494 _6747_/Q VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1760 _6555_/Q VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1771 hold426/X VGND VGND VPWR VPWR hold1771/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5831__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1782 hold983/X VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1793 _6578_/Q VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5347__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3358__B1 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5898__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6075__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5822__A2 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6840_ _7084_/CLK _6840_/D fanout447/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5586__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6771_ _6809_/CLK _6771_/D fanout442/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfstp_4
X_3983_ _3983_/A0 _5194_/A1 _3987_/S VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2482_A _7133_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5722_ _6902_/Q _5679_/X _5685_/X _7070_/Q _5721_/X VGND VGND VPWR VPWR _5727_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3597__B1 _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7017_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5338__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5653_ _5685_/A _5676_/B _5686_/B VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__and3b_4
XFILLER_191_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4604_ _4580_/Y _4581_/X _4598_/A VGND VGND VPWR VPWR _4604_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5889__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4322__A _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5584_ _5584_/A0 _5584_/A1 _5586_/S VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4010__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7106_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_191_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ _4463_/B _4570_/D _4533_/X _4534_/Y _4893_/A VGND VGND VPWR VPWR _4535_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold301 hold301/A VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4561__A2 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold312 hold312/A VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold323 hold323/A VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold334 _4060_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold345 hold345/A VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4466_ _4466_/A VGND VGND VPWR VPWR _4765_/B sky130_fd_sc_hd__inv_2
Xhold356 hold356/A VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold367 hold367/A VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold378 hold378/A VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold389 hold389/A VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6205_ _7012_/Q _5993_/X _5994_/X _7068_/Q VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__a22o_1
X_3417_ input41/X _4056_/C _5308_/A _6899_/Q VGND VGND VPWR VPWR _3417_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5510__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7185_ _7185_/CLK _7185_/D fanout443/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_1
X_4397_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4523_/A sky130_fd_sc_hd__and2_4
XANTENNA_fanout398_A hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _7049_/Q _5996_/X _6012_/X _7001_/Q _6135_/X VGND VGND VPWR VPWR _6136_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _6884_/Q _5290_/A _5434_/A _7012_/Q VGND VGND VPWR VPWR _3348_/X sky130_fd_sc_hd__a22o_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1001 _4088_/A1 VGND VGND VPWR VPWR hold1839/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1012 hold42/X VGND VGND VPWR VPWR hold1012/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _3265_/X VGND VGND VPWR VPWR _3266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1034 _7204_/Q VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6067_ _6067_/A1 _6342_/S _6065_/X _6066_/X VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__o22a_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3277_/B hold63/A VGND VGND VPWR VPWR _3279_/Y sky130_fd_sc_hd__nand2b_1
Xhold1045 hold1045/A VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _6572_/Q VGND VGND VPWR VPWR _4120_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1067 hold50/X VGND VGND VPWR VPWR _4174_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5018_ _4664_/Y _5011_/X _4736_/Y VGND VGND VPWR VPWR _5018_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5813__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1078 _5586_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _3295_/A VGND VGND VPWR VPWR _3356_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5577__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6969_ _6969_/CLK hold98/X fanout450/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold1582_A _6739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3588__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5329__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6730__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4001__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3760__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5501__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold890 hold890/A VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6057__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4068__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2280 _6598_/Q VGND VGND VPWR VPWR hold932/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2291 _6589_/Q VGND VGND VPWR VPWR hold752/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5804__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1590 _5375_/X VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5568__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4320_ _4320_/A0 _5233_/A1 _4321_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6296__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4251_ _4251_/A0 _5237_/A1 _4255_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3202_ _7136_/Q VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
X_4182_ _4182_/A hold9/A VGND VGND VPWR VPWR _4187_/S sky130_fd_sc_hd__and2_4
XANTENNA__6048__A2 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold17_A hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4059__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3221__A _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5559__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6823_ _6826_/CLK _6823_/D _6407_/A VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6220__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6754_ _6761_/CLK _6754_/D _6416_/A VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4231__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3966_ _6456_/Q _3966_/B VGND VGND VPWR VPWR _3966_/X sky130_fd_sc_hd__and2b_4
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5705_ _6845_/Q _5653_/X _5702_/X _5704_/X VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__a211o_1
X_6685_ _3950_/A1 _6685_/D _4107_/B VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_4
X_3897_ _4344_/C _4344_/D _4343_/A _4343_/B VGND VGND VPWR VPWR _3898_/C sky130_fd_sc_hd__nor4_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ _5634_/B _5635_/Y _5639_/B VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__a21oi_1
XFILLER_176_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ _5567_/A0 _5567_/A1 _5568_/S VGND VGND VPWR VPWR _5567_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold1163_A _7023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3742__B1 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__clkbuf_2
X_4518_ _4615_/B _4972_/A VGND VGND VPWR VPWR _5063_/A sky130_fd_sc_hd__nand2_1
Xhold131 _5257_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold142 hold142/A VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold153 hold153/A VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5498_ _5498_/A0 _5534_/A1 _5505_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold175 hold175/A VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4198__S _4199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6287__A2 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4449_ _4457_/A _4671_/A VGND VGND VPWR VPWR _4450_/B sky130_fd_sc_hd__nor2_1
Xhold186 hold186/A VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold197 hold197/A VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7168_ _7185_/CLK _7168_/D fanout443/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _7089_/Q _5638_/X _5998_/X _6889_/Q _6118_/X VGND VGND VPWR VPWR _6119_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7099_ _7099_/CLK _7099_/D fanout471/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5798__B2 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6911__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6211__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4773__A2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input76_A qspi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5492__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3733__B1 _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7088__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6278__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4289__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4828__A3 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6202__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3820_ _3846_/S VGND VGND VPWR VPWR _3835_/S sky130_fd_sc_hd__inv_2
XFILLER_32_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4213__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3751_ _6614_/Q _4170_/A _4176_/A _6619_/Q VGND VGND VPWR VPWR _3751_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_59_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _3958_/A1 _6470_/D _6420_/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3682_ _6738_/Q _4310_/A _4274_/A _6708_/Q VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5421_ _5421_/A0 _5529_/A1 _5424_/S VGND VGND VPWR VPWR _5421_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5713__A1 _6894_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput203 _3935_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XANTENNA__3724__B1 _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5352_ _5352_/A0 _5577_/A1 _5352_/S VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput214 _3939_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
Xoutput225 _7220_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput236 _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _3941_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput258 _6793_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
XANTENNA__6269__A2 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4303_ _4303_/A0 _5448_/A1 hold65/X VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
Xoutput269 _6790_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5283_ _5283_/A0 _5562_/A1 _5289_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3216__A _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4819__A3 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7022_ _7124_/CLK _7022_/D fanout467/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfstp_2
X_4234_ _4234_/A0 _4233_/X _4240_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4165_ _4165_/A0 _5561_/A1 _4169_/S VGND VGND VPWR VPWR _4165_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4096_ _4096_/A0 _5233_/A1 _4097_/S VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6561__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5577__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _6815_/CLK _6806_/D fanout443/X VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout430_A _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4204__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4998_ _4658_/A _4633_/B _4683_/A _4727_/Y _4885_/X VGND VGND VPWR VPWR _4999_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ _6508_/Q user_clock _6819_/Q VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__mux2_1
X_6737_ _6809_/CLK _6737_/D fanout442/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6668_ _7125_/CLK _6668_/D fanout468/X VGND VGND VPWR VPWR _7222_/A sky130_fd_sc_hd__dfrtp_1
X_5619_ _5685_/A _5639_/A VGND VGND VPWR VPWR _5619_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5704__A1 _6957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6599_ _7045_/CLK _6599_/D fanout444/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3715__B1 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout430 _6430_/B VGND VGND VPWR VPWR _6433_/B sky130_fd_sc_hd__buf_6
XFILLER_132_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout441 fanout454/X VGND VGND VPWR VPWR fanout441/X sky130_fd_sc_hd__buf_12
Xfanout452 fanout453/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__buf_12
Xfanout463 fanout464/X VGND VGND VPWR VPWR fanout463/X sky130_fd_sc_hd__buf_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout474 _6346_/B VGND VGND VPWR VPWR _4107_/B sky130_fd_sc_hd__buf_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3494__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input130_A wb_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5487__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5943__A1 _6735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5943__B2 _6592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output182_A _5763_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3706__B1 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3485__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5970_ _5970_/A1 _6342_/S _5968_/X _5969_/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__o22a_1
XFILLER_92_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4921_ _4921_/A _4921_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5397__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4852_ _4638_/Y _4688_/C _4625_/Y VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__o21a_1
XFILLER_166_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3803_ _3803_/A _3803_/B VGND VGND VPWR VPWR _3803_/Y sky130_fd_sc_hd__nand2_8
X_4783_ _4384_/A _4658_/A _4417_/B _4986_/C VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__o31a_2
X_6522_ _7086_/CLK _6522_/D fanout467/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3734_ input35/X _3315_/Y _5434_/A _7006_/Q _3733_/X VGND VGND VPWR VPWR _3735_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6453_ _6809_/CLK _6453_/D fanout433/X VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_4
X_3665_ _6895_/Q _5308_/A _4250_/A _6689_/Q VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5698__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5404_ _5404_/A0 _5575_/A1 _5406_/S VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__mux2_1
X_6384_ _6383_/X _6384_/A1 _6384_/S VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3596_ _7032_/Q _5461_/A _4200_/A _6642_/Q VGND VGND VPWR VPWR _3596_/X sky130_fd_sc_hd__a22o_1
X_5335_ _5335_/A _5578_/B VGND VGND VPWR VPWR _5343_/S sky130_fd_sc_hd__and2_4
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2802 hold913/X VGND VGND VPWR VPWR _5227_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5266_ _5266_/A0 _5581_/A1 _5271_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
Xhold2813 hold656/X VGND VGND VPWR VPWR _5279_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6111__B2 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2824 _6970_/Q VGND VGND VPWR VPWR hold950/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7005_ _7045_/CLK _7005_/D fanout444/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfstp_2
Xhold2835 _5422_/X VGND VGND VPWR VPWR hold952/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4217_ _4217_/A0 _5448_/A1 _4217_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
Xhold2846 _6922_/Q VGND VGND VPWR VPWR hold964/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout380_A hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2857 _6774_/Q VGND VGND VPWR VPWR _3805_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5197_ hold210/X wire375/X _5199_/S VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__mux2_1
Xhold2868 _7163_/Q VGND VGND VPWR VPWR _5794_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3476__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2879 _7182_/Q VGND VGND VPWR VPWR _6291_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5870__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4148_ _4148_/A0 _5238_/A1 _4151_/S VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4079_ _4079_/A0 _5238_/A1 _4082_/S VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3779__A3 _5220_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6178__A1 _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6457__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4113__A0 _3462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input39_A mgmt_gpio_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5861__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A1 _6641_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__B2 _6631_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4134__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3973__B _3973_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap416 _4738_/B VGND VGND VPWR VPWR _4700_/B sky130_fd_sc_hd__clkbuf_2
Xhold708 hold708/A VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold719 _4057_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3450_ _7058_/Q _5488_/A hold24/A _3428_/X VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3381_ _6868_/Q _5272_/A _5380_/A _6964_/Q VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2143_A _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5120_ _4402_/Y _4523_/Y _4583_/B _4642_/Y _4839_/X VGND VGND VPWR VPWR _5121_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2109 _6782_/Q VGND VGND VPWR VPWR hold666/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4104__A0 _3462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5051_ _4583_/B _4688_/B _4691_/Y _4638_/Y _4622_/C VGND VGND VPWR VPWR _5052_/C
+ sky130_fd_sc_hd__o221a_1
Xhold1408 _6913_/Q VGND VGND VPWR VPWR hold392/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1419 _5204_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3458__A2 _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4002_ _4002_/A0 _5193_/A1 _4008_/S VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5852__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5953_ _6534_/Q _5653_/X _5662_/X _6588_/Q _5951_/X VGND VGND VPWR VPWR _5953_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4904_ _4879_/X _4892_/X _4903_/X _4561_/X VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__a31o_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5884_ _6605_/Q _5684_/X _5686_/X _6620_/Q VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3630__A2 _5184_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4835_ _5114_/B _4834_/X _4716_/Y VGND VGND VPWR VPWR _4836_/B sky130_fd_sc_hd__a21oi_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4766_ _4735_/Y _4765_/Y _4407_/Y VGND VGND VPWR VPWR _4791_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _7106_/CLK _6505_/D fanout472/X VGND VGND VPWR VPWR _7213_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3394__B2 input27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3717_ _6728_/Q _3509_/Y _4065_/A _6526_/Q VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4712_/A _4712_/B _4698_/C VGND VGND VPWR VPWR _4702_/B sky130_fd_sc_hd__and3_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1076_A _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6332__A1 _6726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3648_ _3648_/A _3648_/B VGND VGND VPWR VPWR _3648_/Y sky130_fd_sc_hd__nor2_2
X_6436_ _6436_/CLK _6436_/D _3882_/X VGND VGND VPWR VPWR _6436_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_134_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6367_ _6686_/Q _6367_/A2 _6367_/B1 _6685_/Q VGND VGND VPWR VPWR _6367_/X sky130_fd_sc_hd__a22o_1
X_3579_ _6864_/Q _5272_/A _4122_/A _6577_/Q _3565_/X VGND VGND VPWR VPWR _3580_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3697__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5318_ hold620/X _5561_/A1 _5325_/S VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__mux2_1
X_6298_ _6572_/Q _5988_/X _6014_/X _6745_/Q VGND VGND VPWR VPWR _6298_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2610 hold927/X VGND VGND VPWR VPWR _4291_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2621 _6796_/Q VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5249_ _5249_/A0 _5303_/A1 _5253_/S VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__mux2_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__clkbuf_2
Xhold2632 _6574_/Q VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2643 _4245_/X VGND VGND VPWR VPWR hold823/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2654 hold535/X VGND VGND VPWR VPWR _4166_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__buf_4
Xhold1920 _4021_/X VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2665 _6803_/Q VGND VGND VPWR VPWR hold741/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5843__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1931 _6835_/Q VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1508_A _6865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2676 _5286_/X VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1942 _6480_/Q VGND VGND VPWR VPWR hold514/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2687 _5278_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__clkbuf_16
Xhold2698 _5170_/X VGND VGND VPWR VPWR hold673/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1953 _6536_/Q VGND VGND VPWR VPWR hold556/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1964 _7191_/Q VGND VGND VPWR VPWR _6351_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1975 _7040_/Q VGND VGND VPWR VPWR hold871/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1986 _6600_/Q VGND VGND VPWR VPWR hold517/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1997 hold564/X VGND VGND VPWR VPWR _5562_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__A2 _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6020__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6323__A1 _6539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3688__A2 _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6496__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6087__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5834__B1 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3612__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4620_ _4625_/A _4621_/A VGND VGND VPWR VPWR _4622_/C sky130_fd_sc_hd__nand2_1
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3376__A1 _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3376__B2 _6478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4551_ _4601_/A _4491_/Y _4548_/X _5138_/A _4550_/Y VGND VGND VPWR VPWR _4553_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3502_ _7001_/Q _5425_/A _5461_/A _7033_/Q VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 hold505/A VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4482_ _4486_/A _4485_/B _4564_/B VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__and3_1
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold527 hold527/A VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold538 hold538/A VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7094__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6221_ _6548_/Q _5999_/X _6019_/X _6732_/Q _6220_/X VGND VGND VPWR VPWR _6238_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3433_ _7042_/Q _3325_/Y hold31/A _7098_/Q VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold47_A hold47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3679__A2 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A _6152_/B _6152_/C VGND VGND VPWR VPWR _6164_/C sky130_fd_sc_hd__nor3_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3364_ _6996_/Q _5416_/A _3325_/Y _7044_/Q _3361_/X VGND VGND VPWR VPWR _3368_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6078__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5103_ _5103_/A _5103_/B _5103_/C VGND VGND VPWR VPWR _5104_/D sky130_fd_sc_hd__and3_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6895_/Q _5989_/X _6013_/X _7079_/Q _6082_/X VGND VGND VPWR VPWR _6088_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1205 _7103_/Q VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3295_/A _3686_/A VGND VGND VPWR VPWR _3295_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__3224__A _6720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1216 _6887_/Q VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1227 _6524_/Q VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5034_ _5034_/A _5034_/B _5034_/C _5034_/D VGND VGND VPWR VPWR _5117_/C sky130_fd_sc_hd__and4_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1238 _6896_/Q VGND VGND VPWR VPWR hold356/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1249 _6976_/Q VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ _7001_/CLK _6985_/D fanout466/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5936_ _6695_/Q _5658_/X _5664_/X _6760_/Q VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ _6697_/Q _5672_/X _5680_/X _6707_/Q _5866_/X VGND VGND VPWR VPWR _5867_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4818_ _4818_/A _4818_/B _5080_/A VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__and3_1
XANTENNA__4013__C1 _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5798_ _6882_/Q _5667_/X _5682_/X _7042_/Q VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4749_ _4804_/A _4686_/X _4748_/X VGND VGND VPWR VPWR _4749_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6419_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
XANTENNA__4867__A1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6429__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6069__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4649_/C sky130_fd_sc_hd__buf_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4701_/A sky130_fd_sc_hd__buf_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6377_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2440 _6593_/Q VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2451 _5457_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6383_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6373_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2462 hold881/X VGND VGND VPWR VPWR _4117_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2473 _7061_/Q VGND VGND VPWR VPWR hold911/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput169 wb_stb_i VGND VGND VPWR VPWR _3893_/D sky130_fd_sc_hd__buf_4
XFILLER_57_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2484 hold917/X VGND VGND VPWR VPWR _5273_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1750 _4289_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2495 hold710/X VGND VGND VPWR VPWR _4323_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5292__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1761 hold977/X VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1772 _6906_/Q VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1783 hold432/X VGND VGND VPWR VPWR hold1783/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1794 hold406/X VGND VGND VPWR VPWR _4127_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6164__B _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_csclk _6549_/CLK VGND VGND VPWR VPWR _6752_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5495__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output262_A _6784_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5524__A _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6339__B _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5283__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5035__A1 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6232__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3982_ _3982_/A0 hold174/X _3998_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
X_6770_ _6809_/CLK _6770_/D fanout433/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3597__A1 _6474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5721_ _6910_/Q _5670_/X _5678_/B _6966_/Q _5707_/B VGND VGND VPWR VPWR _5721_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5652_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5686_/B sky130_fd_sc_hd__and2b_4
XFILLER_176_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _4981_/A _4917_/D VGND VGND VPWR VPWR _4616_/B sky130_fd_sc_hd__nand2_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5583_ _5583_/A0 _5583_/A1 _5586_/S VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4322__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3219__A _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4534_ _4562_/A _4972_/A VGND VGND VPWR VPWR _4534_/Y sky130_fd_sc_hd__nand2_2
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 hold313/A VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6299__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold324 hold324/A VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4465_ _4363_/B _4465_/B VGND VGND VPWR VPWR _4466_/A sky130_fd_sc_hd__nand2b_4
Xhold346 hold346/A VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold357 hold357/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5434__A _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _6204_/A _6204_/B _6204_/C _6204_/D VGND VGND VPWR VPWR _6214_/B sky130_fd_sc_hd__nor4_1
X_3416_ _7027_/Q _5452_/A _5254_/A _6851_/Q _3415_/X VGND VGND VPWR VPWR _3421_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7184_ _7184_/CLK _7184_/D fanout443/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_1
X_4396_ _4513_/A _5009_/A _4580_/A _4652_/A VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__and4_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6135_ _7065_/Q _5994_/X _6018_/X _6969_/Q VGND VGND VPWR VPWR _6135_/X sky130_fd_sc_hd__a22o_1
X_3347_ _3347_/A _3686_/A VGND VGND VPWR VPWR _5434_/A sky130_fd_sc_hd__nor2_8
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _4112_/A1 VGND VGND VPWR VPWR hold1866/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1013 hold1013/A VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6066_ _6490_/Q _6066_/A2 _5649_/Y VGND VGND VPWR VPWR _6066_/X sky130_fd_sc_hd__a21o_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1024 _3266_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1035 hold7/X VGND VGND VPWR VPWR _3976_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3278_ hold62/X hold21/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__nor2_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5274__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1046 _5511_/X VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 _4120_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5017_ _4691_/Y _4995_/B _5016_/X _4818_/B VGND VGND VPWR VPWR _5080_/B sky130_fd_sc_hd__o211a_1
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1068 _4174_/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1079 _6607_/Q VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6968_ _6994_/CLK _6968_/D fanout462/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3588__A1 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3588__B2 input23/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5919_ _6532_/Q _5653_/X _5918_/X VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4785__B1 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6899_ _6996_/CLK _6899_/D fanout463/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5734__C1 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5344__A _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input160_A wb_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold880 hold880/A VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold891 hold891/A VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2270 hold615/X VGND VGND VPWR VPWR _4148_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input21_A mask_rev_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5265__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2281 hold932/X VGND VGND VPWR VPWR _4151_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2292 hold752/X VGND VGND VPWR VPWR _4141_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1580 hold353/X VGND VGND VPWR VPWR _5289_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1591 _6918_/Q VGND VGND VPWR VPWR _5337_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5017__A1 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3579__A1 _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5740__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5254__A _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4250_ _4250_/A _5220_/C VGND VGND VPWR VPWR _4255_/S sky130_fd_sc_hd__and2_2
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3201_ _6719_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4181_ _4181_/A0 _5448_/A1 _4181_/S VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_55_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5256__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5008__A1 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6205__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6822_ _7073_/CLK _6822_/D fanout443/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_1
X_6753_ _6753_/CLK _6753_/D fanout454/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3965_ _6457_/Q _3965_/B VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__and2b_4
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5704_ _6957_/Q _5680_/X _5686_/X _7005_/Q _5703_/X VGND VGND VPWR VPWR _5704_/X
+ sky130_fd_sc_hd__a221o_1
X_3896_ _4343_/C _4343_/D _3896_/C VGND VGND VPWR VPWR _3898_/B sky130_fd_sc_hd__nor3_1
X_6684_ _3950_/A1 _6684_/D _4107_/B VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3990__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A _5639_/A VGND VGND VPWR VPWR _5635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5566_ _5566_/A0 _5584_/A1 _5568_/S VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5731__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold110 hold110/A VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3742__A1 _7053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold121 hold121/A VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4517_ _4812_/A _4948_/A VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__and2_1
XANTENNA__3742__B2 _6569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold132 hold132/A VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5497_ _5497_/A _5533_/B VGND VGND VPWR VPWR _5505_/S sky130_fd_sc_hd__and2_4
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold154 hold154/A VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold165 _4119_/X VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold176 hold176/A VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4448_ _4714_/B VGND VGND VPWR VPWR _4671_/A sky130_fd_sc_hd__inv_2
XANTENNA__7150__SET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold187 hold187/A VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold198 hold198/A VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5495__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4379_ _5001_/A _4717_/A _4717_/B VGND VGND VPWR VPWR _4811_/B sky130_fd_sc_hd__and3_4
X_7167_ _7180_/CLK _7167_/D fanout446/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _6849_/Q _6007_/X _6019_/X _6985_/Q VGND VGND VPWR VPWR _6118_/X sky130_fd_sc_hd__a22o_1
X_7098_ _7139_/CLK _7098_/D fanout471/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5247__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6958_/Q _5992_/X _6019_/X _6982_/Q _6048_/X VGND VGND VPWR VPWR _6054_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5798__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3981__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5722__A2 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3733__B2 _6585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input69_A mgmt_gpio_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5486__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5238__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5789__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5946__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5410__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _3750_/A _3750_/B _3750_/C _3750_/D VGND VGND VPWR VPWR _3770_/A sky130_fd_sc_hd__nor4_1
XFILLER_13_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5961__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3681_ _6926_/Q _5344_/A _5290_/A _6878_/Q _3680_/X VGND VGND VPWR VPWR _3684_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2173_A _6474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5420_ _5420_/A0 _5537_/A1 _5424_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5713__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput204 _3934_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _5351_/A0 _5549_/A1 _5352_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
Xoutput215 _7212_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
Xoutput226 _7221_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput237 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2438_A _6483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput248 _3959_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_5_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4302_ _4302_/A0 hold43/X hold65/X VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _6794_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_5282_ hold679/X _5579_/A1 _5289_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5477__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7021_ _7134_/CLK _7021_/D fanout469/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfstp_4
X_4233_ _4233_/A0 hold95/X _5236_/C VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3931__S _3934_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4164_ _4164_/A hold9/A VGND VGND VPWR VPWR _4169_/S sky130_fd_sc_hd__and2_2
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4095_ _4095_/A0 _5527_/A1 _4097_/S VGND VGND VPWR VPWR _4095_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4328__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3232__A _6904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4047__B _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3660__B1 _5202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _6815_/CLK _6805_/D fanout443/X VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4997_ _4997_/A _5104_/C VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__and2_2
XANTENNA__5401__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ _6736_/CLK _6736_/D fanout436/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3948_ _3239_/Y input2/X input1/X VGND VGND VPWR VPWR _3948_/X sky130_fd_sc_hd__mux2_8
XANTENNA__5952__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6667_ _7091_/CLK _6667_/D fanout452/X VGND VGND VPWR VPWR _7211_/A sky130_fd_sc_hd__dfrtp_1
X_3879_ _3879_/A _3879_/B VGND VGND VPWR VPWR _3879_/X sky130_fd_sc_hd__and2_1
XANTENNA_hold1273_A _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5618_ _5620_/S _5617_/X _5611_/Y VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__o21a_1
XANTENNA__5704__A2 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6598_ _6835_/CLK _6598_/D fanout435/X VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3715__A1 _6950_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3715__B2 _7054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5549_ _5549_/A0 _5549_/A1 _5550_/S VGND VGND VPWR VPWR _5549_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1538_A _7099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7179_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5468__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7219_ _7219_/A VGND VGND VPWR VPWR _7219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout431 _6430_/B VGND VGND VPWR VPWR _6423_/B sky130_fd_sc_hd__buf_8
XFILLER_59_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout442 fanout449/X VGND VGND VPWR VPWR fanout442/X sky130_fd_sc_hd__buf_12
Xfanout453 fanout454/X VGND VGND VPWR VPWR fanout453/X sky130_fd_sc_hd__buf_8
Xfanout464 fanout465/X VGND VGND VPWR VPWR fanout464/X sky130_fd_sc_hd__buf_12
XFILLER_101_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout475 input164/X VGND VGND VPWR VPWR _6346_/B sky130_fd_sc_hd__buf_12
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input123_A wb_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6196__A2 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__B1 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5943__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4701__A _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3706__B2 _6570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output175_A _3948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5459__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7161__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6120__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4131__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4920_ _5114_/A _4920_/B _5114_/B VGND VGND VPWR VPWR _4929_/B sky130_fd_sc_hd__and3_1
XFILLER_80_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4851_ _4917_/D _5048_/B VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__nand2_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6187__A2 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4198__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3802_ _3774_/X _3802_/B _3802_/C _3802_/D VGND VGND VPWR VPWR _3803_/B sky130_fd_sc_hd__and4b_2
X_4782_ _4552_/B _4955_/D _4396_/X VGND VGND VPWR VPWR _4782_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5934__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6521_ _7106_/CLK _6521_/D fanout472/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3945__A1 _3966_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ _6480_/Q _4000_/A _4134_/A _6585_/Q VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__a22o_2
X_6452_ _6809_/CLK _6452_/D fanout433/X VGND VGND VPWR VPWR _6452_/Q sky130_fd_sc_hd__dfstp_4
X_3664_ _3664_/A _3664_/B _3664_/C VGND VGND VPWR VPWR _3674_/C sky130_fd_sc_hd__nor3_1
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5403_ _5403_/A0 _5529_/A1 _5406_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6383_ _6684_/Q _6383_/A2 _6383_/B1 _4218_/Y _6382_/X VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a221o_1
X_3595_ _3595_/A _3595_/B _3595_/C _3595_/D VGND VGND VPWR VPWR _3615_/A sky130_fd_sc_hd__nor4_1
XANTENNA__3227__A _6944_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5334_ _5334_/A0 _5577_/A1 _5334_/S VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2803 _5227_/X VGND VGND VPWR VPWR hold914/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6111__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5265_ _5265_/A0 _5562_/A1 _5271_/S VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2814 _5279_/X VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2825 hold950/X VGND VGND VPWR VPWR _5395_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7004_ _7139_/CLK _7004_/D fanout471/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2836 _6549_/Q VGND VGND VPWR VPWR hold940/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4216_ _4216_/A0 _5233_/A1 _4217_/S VGND VGND VPWR VPWR _4216_/X sky130_fd_sc_hd__mux2_1
X_5196_ _5196_/A0 _5277_/A1 _5199_/S VGND VGND VPWR VPWR _5196_/X sky130_fd_sc_hd__mux2_1
Xhold2847 hold964/X VGND VGND VPWR VPWR _5341_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2858 _6779_/Q VGND VGND VPWR VPWR _3464_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2869 _5773_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4147_ _4147_/A0 _5543_/A1 _4151_/S VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout373_A wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1119_A _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4078_ _4078_/A0 _5543_/A1 _4082_/S VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3633__B1 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6178__A2 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4189__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6719_ _6786_/CLK _6719_/D fanout435/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7184__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5861__B2 _6604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5498__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3624__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output292_A _6484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap417 _4712_/C VGND VGND VPWR VPWR _4738_/B sky130_fd_sc_hd__clkbuf_2
Xhold709 hold709/A VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap428 _4389_/Y VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3380_ _6956_/Q _3291_/Y _4047_/C input51/X _3379_/X VGND VGND VPWR VPWR _3383_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5050_ _4510_/A _4523_/Y _4583_/B _4995_/A _4859_/X VGND VGND VPWR VPWR _5112_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 hold392/X VGND VGND VPWR VPWR _5331_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4001_ _4001_/A0 _5237_/A1 _4008_/S VGND VGND VPWR VPWR _4001_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5952_ _6578_/Q _5667_/X _5682_/X _6454_/Q VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4903_ _5155_/A _4903_/B _4903_/C _4903_/D VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__and4_1
X_5883_ _6688_/Q _5659_/X _5687_/X _6600_/Q VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4834_ _4834_/A _4834_/B _4834_/C VGND VGND VPWR VPWR _4834_/X sky130_fd_sc_hd__and3_1
XFILLER_21_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5907__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4765_ _4955_/C _4765_/B _4972_/A VGND VGND VPWR VPWR _4765_/Y sky130_fd_sc_hd__nand3_2
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ _6936_/CLK _6504_/D fanout463/X VGND VGND VPWR VPWR _7212_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3394__A2 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3716_ _3716_/A _3716_/B _3716_/C _3716_/D VGND VGND VPWR VPWR _3736_/B sky130_fd_sc_hd__nor4_1
X_4696_ _4990_/B _4691_/Y _4692_/X _4694_/Y _4922_/B VGND VGND VPWR VPWR _4703_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _3958_/A1 _6435_/D _6391_/X VGND VGND VPWR VPWR _6435_/Q sky130_fd_sc_hd__dfrtp_4
X_3647_ input5/X _3315_/Y _4310_/A _6739_/Q _3646_/X VGND VGND VPWR VPWR _3655_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6332__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1069_A _6710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6366_ _6365_/X _6366_/A1 _6384_/S VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__mux2_1
X_3578_ _6872_/Q _5281_/A _5389_/A _6968_/Q _3577_/X VGND VGND VPWR VPWR _3580_/C
+ sky130_fd_sc_hd__a221o_2
X_5317_ _5317_/A _5317_/B VGND VGND VPWR VPWR _5325_/S sky130_fd_sc_hd__and2_4
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6297_ _6612_/Q _5976_/B _5995_/X _6602_/Q _6296_/X VGND VGND VPWR VPWR _6304_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2600 _6808_/Q VGND VGND VPWR VPWR hold681/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__A1 _6904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2611 _4291_/X VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B2 _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2622 hold508/X VGND VGND VPWR VPWR _5193_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__buf_8
X_5248_ _5248_/A0 _5527_/A1 _5253_/S VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
Xhold2633 hold713/X VGND VGND VPWR VPWR _4123_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2644 _6798_/Q VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1910 _7012_/Q VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2655 _4166_/X VGND VGND VPWR VPWR hold536/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkbuf_4
Xhold1921 hold585/X VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2666 hold741/X VGND VGND VPWR VPWR _5201_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1932 hold316/X VGND VGND VPWR VPWR _5243_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2677 _6731_/Q VGND VGND VPWR VPWR hold670/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5179_ _5179_/A0 _5237_/A1 _5183_/S VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__mux2_1
Xhold1943 hold514/X VGND VGND VPWR VPWR _4002_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2688 _6649_/Q VGND VGND VPWR VPWR hold695/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1403_A _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1954 hold556/X VGND VGND VPWR VPWR _4079_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2699 _6746_/Q VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1965 hold1965/A VGND VGND VPWR VPWR hold488/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1976 hold871/X VGND VGND VPWR VPWR _5474_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1987 hold517/X VGND VGND VPWR VPWR _4154_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1998 _5562_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3606__B1 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6316__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6020__B2 _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6323__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A mgmt_gpio_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5834__A1 _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output305_A _3392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6063__D _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3376__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4550_ _4972_/A _4628_/A VGND VGND VPWR VPWR _4550_/Y sky130_fd_sc_hd__nand2_2
XFILLER_184_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3501_ _3553_/A _3523_/B VGND VGND VPWR VPWR _4334_/A sky130_fd_sc_hd__nor2_4
XFILLER_171_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold506 hold506/A VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4481_ _4724_/C _4562_/A VGND VGND VPWR VPWR _4893_/A sky130_fd_sc_hd__nand2_1
Xhold517 hold517/A VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold528 hold528/A VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold539 hold539/A VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6220_ _6752_/Q _5638_/X _6015_/X _6757_/Q VGND VGND VPWR VPWR _6220_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4325__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3432_ _7138_/Q _3295_/Y _4241_/A input57/X VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _7034_/Q _5986_/X _5998_/X _6890_/Q _6150_/X VGND VGND VPWR VPWR _6152_/C
+ sky130_fd_sc_hd__a221o_1
X_3363_ _7052_/Q hold16/A _5407_/A _6988_/Q _3359_/X VGND VGND VPWR VPWR _3368_/A
+ sky130_fd_sc_hd__a221o_2
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6078__A1 _6959_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5102_ _5102_/A _5102_/B _5102_/C VGND VGND VPWR VPWR _5103_/C sky130_fd_sc_hd__and3_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4100__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4089__A0 _3462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6935_/Q _5980_/X _6017_/X _7071_/Q VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__a22o_1
X_3294_ hold79/X _3430_/A VGND VGND VPWR VPWR _3294_/Y sky130_fd_sc_hd__nand2_8
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 hold237/X VGND VGND VPWR VPWR _5545_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A1 _6955_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1217 hold249/X VGND VGND VPWR VPWR _5302_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1228 hold82/X VGND VGND VPWR VPWR _4064_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5033_ _5033_/A _5033_/B VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__nand2_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1239 hold356/X VGND VGND VPWR VPWR _5312_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6447__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6984_ _7112_/CLK _6984_/D fanout473/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5935_ _6637_/Q _5671_/X _5931_/X _5933_/X _5934_/X VGND VGND VPWR VPWR _5935_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5866_ _6609_/Q _5660_/X _5669_/X _6649_/Q VGND VGND VPWR VPWR _5866_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4817_ _4917_/A _4672_/Y _4812_/Y _4815_/X _5010_/A VGND VGND VPWR VPWR _4820_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_178_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ _3242_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4071__A _5220_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3367__A2 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4748_ _4637_/C _4719_/A _4686_/X _4747_/Y VGND VGND VPWR VPWR _4748_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5761__B1 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4679_ _5009_/B _4826_/A VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__6305__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6418_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4867__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6349_ _3675_/Y hold994/A _6354_/S VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4344_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3896_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__clkbuf_16
Xhold2430 _6487_/Q VGND VGND VPWR VPWR hold920/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4619__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2441 hold867/X VGND VGND VPWR VPWR _4145_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6361_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2452 _7125_/Q VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6376_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2463 _4117_/X VGND VGND VPWR VPWR hold882/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2474 hold911/X VGND VGND VPWR VPWR _5498_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1740 _6603_/Q VGND VGND VPWR VPWR hold327/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2485 _5273_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2496 _4323_/X VGND VGND VPWR VPWR hold711/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1751 _6540_/Q VGND VGND VPWR VPWR hold975/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1762 hold430/X VGND VGND VPWR VPWR hold1762/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1773 hold633/X VGND VGND VPWR VPWR _5323_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1784 _6624_/Q VGND VGND VPWR VPWR hold702/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1795 _4127_/X VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A wb_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3358__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5752__B1 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4307__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5524__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6232__A1 _6707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3981_ _3981_/A0 _5193_/A1 _3987_/S VGND VGND VPWR VPWR _3981_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5720_ _6974_/Q _5660_/X _5686_/X _7006_/Q _5719_/X VGND VGND VPWR VPWR _5727_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3597__A2 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4794__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5651_ _5685_/A _5676_/B _5689_/B VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__and3b_4
XANTENNA__4603__B _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4602_ _4581_/X _4602_/B VGND VGND VPWR VPWR _4602_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5743__B1 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5582_ _5582_/A0 _5582_/A1 _5586_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4533_ _5034_/A _4533_/B _4533_/C _4533_/D VGND VGND VPWR VPWR _4533_/X sky130_fd_sc_hd__and4_1
XFILLER_117_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3934__S _3934_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold303 hold303/A VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold314 hold314/A VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2635_A _6843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold325 hold325/A VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4464_ _4576_/A _4488_/B VGND VGND VPWR VPWR _4464_/Y sky130_fd_sc_hd__nand2_4
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold347 hold347/A VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold358 hold358/A VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5434__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6203_ _7036_/Q _5986_/X _5988_/X _6876_/Q _6202_/X VGND VGND VPWR VPWR _6204_/D
+ sky130_fd_sc_hd__a221o_1
X_3415_ _7043_/Q _3325_/Y _5407_/A _6987_/Q VGND VGND VPWR VPWR _3415_/X sky130_fd_sc_hd__a22o_1
X_7183_ _7184_/CLK _7183_/D fanout449/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_1
X_4395_ _4395_/A _4650_/B VGND VGND VPWR VPWR _4652_/A sky130_fd_sc_hd__nor2_4
XANTENNA__3235__A _6880_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7097_/Q _5984_/X _6013_/X _7081_/Q VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a22o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3346_ _3346_/A _3686_/A VGND VGND VPWR VPWR _5290_/A sky130_fd_sc_hd__nor2_8
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1003 _6351_/A1 VGND VGND VPWR VPWR hold1965/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _5564_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6838_/Q _6339_/B _6064_/Y _6341_/S VGND VGND VPWR VPWR _6065_/X sky130_fd_sc_hd__o211a_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ hold21/X _3277_/B VGND VGND VPWR VPWR _3290_/B sky130_fd_sc_hd__nor2_2
Xhold1025 _3297_/Y VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1036 _3976_/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 _6889_/Q VGND VGND VPWR VPWR hold100/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5016_ _5011_/A _4590_/Y _4688_/B VGND VGND VPWR VPWR _5016_/X sky130_fd_sc_hd__a21o_1
Xhold1058 _7081_/Q VGND VGND VPWR VPWR hold103/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1069 _6710_/Q VGND VGND VPWR VPWR _4278_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout453_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/CLK _6967_/D fanout465/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5918_ _6576_/Q _5667_/X _5682_/X _6452_/Q VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3588__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4785__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6898_ _6996_/CLK _6898_/D fanout462/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5849_ _7028_/Q _5663_/X _5843_/X _5844_/X _5848_/X VGND VGND VPWR VPWR _5849_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_158_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7104__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4537__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5734__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3760__A2 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5344__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold870 hold870/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold881 hold881/A VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold892 hold892/A VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input153_A wb_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2260 _5186_/X VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2271 _4148_/X VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2282 _4151_/X VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2293 _4141_/X VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6762__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1570 _6947_/Q VGND VGND VPWR VPWR hold315/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input14_A mask_rev_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1581 _5289_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1592 _5337_/X VGND VGND VPWR VPWR hold121/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3579__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4528__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4528__B2 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5725__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3751__A2 _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6827__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_max_cap349_A _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5254__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6150__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ _6718_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3503__A2 _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4180_ _4180_/A0 _5233_/A1 _4181_/S VGND VGND VPWR VPWR _4180_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7157__477 VGND VGND VPWR VPWR _7157_/D _7157__477/LO sky130_fd_sc_hd__conb_1
XFILLER_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6821_ _6821_/CLK _6821_/D fanout449/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ _6752_/CLK _6752_/D fanout440/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5964__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3964_ input85/X _3879_/B _6457_/Q VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__mux2_2
X_5703_ _6861_/Q _5673_/X _5687_/X _6917_/Q VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6683_ _7203_/CLK _6683_/D _4107_/B VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_4
X_3895_ _4345_/C _4345_/D _4344_/A _4344_/B VGND VGND VPWR VPWR _3899_/C sky130_fd_sc_hd__nor4_1
XFILLER_149_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5634_ _5637_/A _5634_/B VGND VGND VPWR VPWR _5639_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5716__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5192__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5565_ _5565_/A0 _5583_/A1 _5568_/S VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 hold100/A VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4516_ _4596_/A _4955_/D VGND VGND VPWR VPWR _4767_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3742__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold111 hold111/A VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold122 hold122/A VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ _5496_/A0 _5568_/A1 _5496_/S VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__mux2_1
Xhold133 _5293_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold144 hold144/A VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 hold155/A VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4447_ _4663_/D _4447_/B VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__and2b_4
Xhold166 hold166/A VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold188 hold188/A VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold199 hold199/A VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7166_ _7180_/CLK _7166_/D fanout446/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4378_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__and2b_4
XFILLER_98_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_csclk _6549_/CLK VGND VGND VPWR VPWR _6753_/CLK sky130_fd_sc_hd__clkbuf_16
X_6117_ _6141_/A1 _6116_/X _6342_/S VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__mux2_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A mask_rev_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3430_/A _3390_/B VGND VGND VPWR VPWR _3648_/A sky130_fd_sc_hd__nand2_8
X_7097_ _7137_/CLK _7097_/D fanout469/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6048_ _6878_/Q _6004_/X _6005_/X _6942_/Q VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5955__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5183__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3733__A2 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6132__B1 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4694__B1 _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2090 _4214_/X VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6199__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6658__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3680_ _6580_/Q _4128_/A _4304_/A _6733_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5174__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3724__A2 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5350_ _5350_/A0 _5575_/A1 _5352_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
Xoutput205 _3933_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6661__RESET_B fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 _7213_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7222_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
Xoutput238 _7230_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
X_4301_ _4301_/A0 _5581_/A1 hold65/X VGND VGND VPWR VPWR _4301_/X sky130_fd_sc_hd__mux2_1
Xoutput249 _3956_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
XFILLER_142_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6123__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5281_ _5281_/A _5578_/B VGND VGND VPWR VPWR _5289_/S sky130_fd_sc_hd__and2_4
XFILLER_141_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2333_A _6720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7020_ _7108_/CLK _7020_/D fanout451/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4232_ _4232_/A0 _4231_/X _4240_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4163_ _4163_/A0 _5448_/A1 _4163_/S VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4094_ _4094_/A0 _5238_/A1 _4097_/S VGND VGND VPWR VPWR _4094_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4328__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4047__C _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3660__B2 _6806_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6804_ _6815_/CLK _6804_/D fanout443/X VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5937__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4996_ _4691_/B _4990_/Y _5081_/B VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__a21oi_1
X_6735_ _6735_/CLK _6735_/D fanout442/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _3238_/Y _6436_/Q _6430_/B VGND VGND VPWR VPWR _3947_/X sky130_fd_sc_hd__mux2_4
XANTENNA__3412__A1 _6963_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6666_ _6835_/CLK _6666_/D _3959_/B VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_4
X_3878_ _3879_/B hold4/A _3878_/S VGND VGND VPWR VPWR _6438_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5617_ _7148_/Q _5613_/B _7149_/Q VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__o21a_1
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6597_ _6752_/CLK _6597_/D fanout440/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3715__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5548_ _5548_/A0 _5584_/A1 _5550_/S VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5479_ hold16/X _5569_/B VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__and2_4
X_7218_ _7218_/A VGND VGND VPWR VPWR _7218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout410 _6166_/S VGND VGND VPWR VPWR _6341_/S sky130_fd_sc_hd__buf_12
XFILLER_120_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout432 _3881_/Y VGND VGND VPWR VPWR _6430_/B sky130_fd_sc_hd__buf_12
Xfanout443 fanout449/X VGND VGND VPWR VPWR fanout443/X sky130_fd_sc_hd__buf_12
X_7149_ _7179_/CLK _7149_/D fanout448/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout454 input75/X VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__buf_12
XFILLER_171_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout465 input75/X VGND VGND VPWR VPWR fanout465/X sky130_fd_sc_hd__buf_12
Xfanout476 _4637_/C VGND VGND VPWR VPWR _4574_/A sky130_fd_sc_hd__buf_12
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A wb_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A1 _6887_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5928__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__B2 _6477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input81_A spi_sdo VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6353__A0 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3706__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6105__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5816__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3642__A1 _6724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3642__B2 _6532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4402_/Y _4570_/C _4638_/Y _4674_/Y VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__o22a_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6041__C1 _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3801_ _3801_/A _3801_/B _3801_/C _3801_/D VGND VGND VPWR VPWR _3802_/D sky130_fd_sc_hd__nor4_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4368_/A _4477_/Y _4729_/A _4550_/Y VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__o31a_1
X_6520_ _6936_/CLK _6520_/D fanout463/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_1
X_3732_ input21/X _3336_/Y _4200_/A _6640_/Q _3731_/X VGND VGND VPWR VPWR _3735_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5707__B _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6451_ _6733_/CLK _6451_/D fanout433/X VGND VGND VPWR VPWR _6451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3663_ _6919_/Q _5335_/A _3660_/X _3662_/X VGND VGND VPWR VPWR _3664_/C sky130_fd_sc_hd__a211o_1
XANTENNA__4611__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5698__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5402_ _5402_/A0 _5537_/A1 _5406_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4103__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6382_ _6686_/Q _6382_/A2 _6382_/B1 _6685_/Q VGND VGND VPWR VPWR _6382_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3594_ _6787_/Q _5178_/A _4182_/A _6627_/Q _3593_/X VGND VGND VPWR VPWR _3595_/D
+ sky130_fd_sc_hd__a221o_1
X_5333_ _5333_/A0 _5549_/A1 _5334_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5264_ _5264_/A0 _5561_/A1 _5271_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
Xhold2804 _6939_/Q VGND VGND VPWR VPWR hold647/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7003_ _7139_/CLK _7003_/D fanout471/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2815 _6978_/Q VGND VGND VPWR VPWR hold953/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2826 _5395_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4215_ hold155/X _5581_/A1 _4217_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
Xhold2837 hold940/X VGND VGND VPWR VPWR _4094_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5195_ _5195_/A0 _5195_/A1 _5199_/S VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__mux2_1
Xhold2848 _5341_/X VGND VGND VPWR VPWR hold965/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2859 _3464_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5870__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4146_ _4146_/A _5533_/B VGND VGND VPWR VPWR _4151_/S sky130_fd_sc_hd__and2_2
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ _4077_/A _5533_/B VGND VGND VPWR VPWR _4082_/S sky130_fd_sc_hd__and2_2
XANTENNA_fanout366_A hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5386__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4979_ _4510_/A _4570_/C _4564_/Y _4968_/Y VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__a31o_1
XFILLER_11_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3397__B1 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6718_ _6786_/CLK _6718_/D fanout435/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6512__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6649_ _6745_/CLK _6649_/D fanout441/X VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__6335__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4521__B _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5310__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5861__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5377__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6326__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output285_A _6801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap418 _4751_/C VGND VGND VPWR VPWR _4712_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_183_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5301__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2031_A _6771_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4000_ _4000_/A _5220_/C VGND VGND VPWR VPWR _4008_/S sky130_fd_sc_hd__and2_4
XANTENNA__5852__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5951_ _6598_/Q _5670_/X _5685_/X _6773_/Q VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _4902_/A _5073_/C _5063_/C _5098_/B VGND VGND VPWR VPWR _4903_/D sky130_fd_sc_hd__and4_1
X_5882_ _5903_/A1 _5881_/X _6342_/S VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _4683_/A _4832_/X _5127_/B _5104_/C _5021_/A VGND VGND VPWR VPWR _4834_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5368__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2665_A _6803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3379__B1 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4764_ _5150_/A _4764_/B VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__nand2_1
X_6503_ _6936_/CLK _6503_/D fanout463/X VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfrtp_1
X_3715_ _6950_/Q _3291_/Y _5488_/A _7054_/Q _3714_/X VGND VGND VPWR VPWR _3716_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4695_ _4826_/A _4719_/B VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__nand2_2
XANTENNA__3238__A _6848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6434_ _3547_/A1 _6434_/D _6390_/X VGND VGND VPWR VPWR _6434_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_134_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3646_ _6983_/Q _5407_/A hold24/A _6812_/Q VGND VGND VPWR VPWR _3646_/X sky130_fd_sc_hd__a22o_1
X_6365_ _6686_/Q _6365_/A2 _6365_/B1 _6685_/Q _6364_/X VGND VGND VPWR VPWR _6365_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5540__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3577_ _7136_/Q _3295_/Y _5542_/A _7104_/Q VGND VGND VPWR VPWR _3577_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3551__B1 _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5316_ _5316_/A0 _5568_/A1 _5316_/S VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6296_ _6715_/Q _5973_/X _5986_/X _6642_/Q VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__a22o_1
Xhold2601 hold681/X VGND VGND VPWR VPWR _5208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2612 _6770_/Q VGND VGND VPWR VPWR hold502/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5247_ _5247_/A0 _5571_/A1 _5253_/S VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2623 _5193_/X VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__buf_12
Xhold2634 _4123_/X VGND VGND VPWR VPWR hold714/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2645 hold699/X VGND VGND VPWR VPWR _5195_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1900 _6620_/Q VGND VGND VPWR VPWR hold529/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1911 hold360/X VGND VGND VPWR VPWR _5442_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2656 _6695_/Q VGND VGND VPWR VPWR hold859/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5843__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__buf_8
Xhold1922 _6453_/Q VGND VGND VPWR VPWR hold669/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2667 _5201_/X VGND VGND VPWR VPWR hold742/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5178_ _5178_/A _5220_/C VGND VGND VPWR VPWR _5183_/S sky130_fd_sc_hd__and2_2
Xhold1933 _6580_/Q VGND VGND VPWR VPWR hold546/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2678 hold670/X VGND VGND VPWR VPWR _4303_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1944 _4002_/X VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2689 hold695/X VGND VGND VPWR VPWR _4213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1955 _6963_/Q VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4129_ _4129_/A0 _5543_/A1 _4133_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__mux2_1
Xhold1966 hold488/X VGND VGND VPWR VPWR hold1966/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1977 _6738_/Q VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1988 _4154_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1999 _7032_/Q VGND VGND VPWR VPWR hold827/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3606__A1 _6840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6764__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7151__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6020__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4031__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6308__B1 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3790__B1 _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5531__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A mgmt_gpio_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6087__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5834__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3845__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5302__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4270__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4022__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3500_ _3544_/A _3523_/B VGND VGND VPWR VPWR _4128_/A sky130_fd_sc_hd__nor2_4
XANTENNA__3781__B1 _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _4486_/A _4491_/B VGND VGND VPWR VPWR _4570_/C sky130_fd_sc_hd__nand2_4
XFILLER_116_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold518 hold518/A VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3431_ _3563_/A _3523_/B VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__nor2_8
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5522__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6150_ _6978_/Q _5976_/B _5993_/X _7010_/Q VGND VGND VPWR VPWR _6150_/X sky130_fd_sc_hd__a22o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _7060_/Q _5488_/A _5497_/A _7068_/Q VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__a22o_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6078__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5101_ _5131_/A _5131_/B _5101_/C VGND VGND VPWR VPWR _5101_/X sky130_fd_sc_hd__and3_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7119_/Q _5978_/X _5995_/X _6919_/Q _6080_/X VGND VGND VPWR VPWR _6088_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3293_ _3343_/A _3563_/A VGND VGND VPWR VPWR _3293_/Y sky130_fd_sc_hd__nor2_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _6841_/Q VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2413_A _6604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5032_ _5032_/A _5032_/B _5032_/C VGND VGND VPWR VPWR _5086_/A sky130_fd_sc_hd__and3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1218 _5302_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1229 _6516_/Q VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6983_ _7086_/CLK _6983_/D fanout467/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6250__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5934_ _6750_/Q _5666_/X _5689_/X _6627_/Q VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4261__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5865_ _6569_/Q _5674_/X _5687_/X _6599_/Q VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4816_ _4729_/A _4688_/B _4688_/C _4583_/B VGND VGND VPWR VPWR _5080_/A sky130_fd_sc_hd__o22a_1
X_5796_ _6994_/Q _5929_/B VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__and2_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ _4415_/B _4714_/Y _4746_/Y VGND VGND VPWR VPWR _4747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4071__B _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5761__A1 _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5761__B2 _6952_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3772__B1 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4678_ _4638_/Y _4674_/Y _4676_/Y _4633_/B _5049_/A VGND VGND VPWR VPWR _4678_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6417_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5513__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3629_ _6601_/Q _4152_/A _4164_/A _6611_/Q _3628_/X VGND VGND VPWR VPWR _3636_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3524__B1 _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6348_ _3737_/Y hold996/A _6354_/S VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6069__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4344_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6279_ _6279_/A _6279_/B _6279_/C _6279_/D VGND VGND VPWR VPWR _6289_/B sky130_fd_sc_hd__nor4_2
XFILLER_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR _3898_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2420 hold905/X VGND VGND VPWR VPWR _4287_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4447_/B sky130_fd_sc_hd__clkbuf_16
Xhold2431 hold920/X VGND VGND VPWR VPWR _4010_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6382_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2442 _4145_/X VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6365_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2453 hold866/X VGND VGND VPWR VPWR _5570_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2464 _6985_/Q VGND VGND VPWR VPWR hold802/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2475 _5498_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1730 hold989/X VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2486 _7001_/Q VGND VGND VPWR VPWR hold803/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1741 hold327/X VGND VGND VPWR VPWR _4157_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1752 hold975/X VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2497 _7129_/Q VGND VGND VPWR VPWR hold838/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1763 _6627_/Q VGND VGND VPWR VPWR hold821/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1774 _5323_/X VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1785 hold702/X VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1796 _6552_/Q VGND VGND VPWR VPWR hold403/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1882_A _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4252__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4262__A _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4004__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5752__A1 _7056_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5752__B2 _7088_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5504__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5807__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7197__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6232__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3980_ _3980_/A0 hold119/X _3998_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_2
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4243__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4794__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5650_ _7146_/Q _7147_/Q VGND VGND VPWR VPWR _5689_/B sky130_fd_sc_hd__and2b_4
XFILLER_31_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4601_ _4601_/A _4601_/B VGND VGND VPWR VPWR _4602_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5581_ _5581_/A0 _5581_/A1 _5586_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4546__A2 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2363_A _7018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3754__B1 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4532_ _4607_/B _4934_/B _4981_/A VGND VGND VPWR VPWR _4533_/D sky130_fd_sc_hd__o21ai_1
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6299__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold315 hold315/A VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4463_ _4718_/A _4463_/B VGND VGND VPWR VPWR _4607_/B sky130_fd_sc_hd__nor2_8
Xhold337 _5244_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2530_A _6528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold348 hold348/A VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6202_ _6860_/Q _5983_/X _6007_/X _6852_/Q VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4111__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3414_ _6875_/Q _5281_/A _5389_/A _6971_/Q _3413_/X VGND VGND VPWR VPWR _3421_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7182_ _7184_/CLK _7182_/D fanout449/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_1
X_4394_ _4394_/A _4650_/B VGND VGND VPWR VPWR _4394_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6133_ _7025_/Q _5971_/X _5990_/X _7057_/Q _6132_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3354_/B hold15/X VGND VGND VPWR VPWR _5335_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3950__S _6818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _4233_/A0 VGND VGND VPWR VPWR hold1143/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6064_ _6045_/X _6064_/B _6064_/C VGND VGND VPWR VPWR _6064_/Y sky130_fd_sc_hd__nand3b_2
Xhold1015 _6439_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3276_ _3276_/A hold55/X VGND VGND VPWR VPWR _3277_/B sky130_fd_sc_hd__nand2_1
Xhold1026 _3298_/Y VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__buf_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _4702_/B _4990_/Y _5014_/X _4822_/Y VGND VGND VPWR VPWR _5015_/X sky130_fd_sc_hd__a211o_1
Xhold1037 hold8/X VGND VGND VPWR VPWR _5317_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1048 hold100/X VGND VGND VPWR VPWR _5304_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1059 hold103/X VGND VGND VPWR VPWR _5520_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout446_A fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6966_ _7061_/CLK _6966_/D fanout450/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5917_ _6734_/Q _5656_/X _5672_/X _6699_/Q _5916_/X VGND VGND VPWR VPWR _5917_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4785__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6897_ _6977_/CLK _6897_/D fanout461/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5178__A _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6974__SET_B fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5848_ _6876_/Q _5674_/X _5845_/X _5847_/X VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a211o_1
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5734__A1 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5779_ _6945_/Q _5658_/X _5666_/X _7001_/Q VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold1463_A _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7144__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4021__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold860 hold860/A VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold871 hold871/A VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold882 hold882/A VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold893 hold893/A VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input146_A wb_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2250 hold616/X VGND VGND VPWR VPWR _4142_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2261 _6854_/Q VGND VGND VPWR VPWR hold599/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2272 _6652_/Q VGND VGND VPWR VPWR hold840/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2283 _6732_/Q VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2294 _6688_/Q VGND VGND VPWR VPWR hold578/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1560 hold333/X VGND VGND VPWR VPWR _4060_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1571 hold315/X VGND VGND VPWR VPWR _5369_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1582 _6739_/Q VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1593 _6900_/Q VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4225__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6759__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6437__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5551__A _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6205__A2 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6820_ _7135_/CLK _6820_/D fanout467/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4216__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5964__A1 _6643_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3963_ _3963_/A VGND VGND VPWR VPWR _3963_/Y sky130_fd_sc_hd__inv_2
X_6751_ _6786_/CLK _6751_/D fanout436/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5964__B2 _6633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5702_ _6893_/Q _5662_/X _5672_/X _6949_/Q VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4106__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6682_ _3950_/A1 _6682_/D _4107_/B VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_4
X_3894_ input118/X input119/X _3894_/C _3894_/D VGND VGND VPWR VPWR _3900_/C sky130_fd_sc_hd__and4bb_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5633_ _5633_/A1 _5611_/Y _5634_/B _5632_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__a31o_1
XANTENNA__5716__A1 _6846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5716__B2 _7038_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3945__S _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__B1 _4009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5564_ hold91/X hold43/X _5568_/S VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4515_ _4462_/Y _4464_/Y _4466_/A _4570_/A _4947_/B VGND VGND VPWR VPWR _5151_/D
+ sky130_fd_sc_hd__o32a_1
Xhold101 hold101/A VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold112 hold112/A VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5495_ _5495_/A0 wire371/X _5496_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
Xhold123 hold123/A VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold134 hold134/A VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold145 hold145/A VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4446_ _4498_/B _4663_/D VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__and2b_1
XFILLER_171_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold156 hold156/A VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold167 hold167/A VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold178 hold178/A VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold189 hold189/A VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7165_ _7185_/CLK _7165_/D fanout446/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_1
X_4377_ _4447_/B _4663_/D VGND VGND VPWR VPWR _4717_/A sky130_fd_sc_hd__nor2_8
XANTENNA_fanout396_A _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5461__A _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6116_ _6116_/A0 _6115_/X _6341_/S VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__mux2_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3429_/A hold46/X _3390_/B VGND VGND VPWR VPWR _5222_/A sky130_fd_sc_hd__and3_4
X_7096_ _7140_/CLK _7096_/D fanout473/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6047_ _6926_/Q _5982_/X _6016_/X _7038_/Q _6046_/X VGND VGND VPWR VPWR _6054_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ hold28/X _3259_/B VGND VGND VPWR VPWR _3259_/X sky130_fd_sc_hd__and2_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4207__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5400__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4524__B _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6949_ _7017_/CLK _6949_/D fanout461/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4016__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3718__B1 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold690 hold690/A VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5891__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2080 hold527/X VGND VGND VPWR VPWR _4208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2091 _6450_/Q VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1390 hold160/X VGND VGND VPWR VPWR _5428_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5310__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__A1 _6528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6779__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3709__B1 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput206 _3185_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 _3951_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4300_ _4300_/A0 _5580_/A1 hold65/X VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
Xoutput228 _7223_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput239 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
X_5280_ _5280_/A0 _5577_/A1 _5280_/S VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ _5240_/A0 _5303_/A1 _5236_/C VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5281__A _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ _4162_/A0 hold43/X _4163_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4093_ _4093_/A0 _5543_/A1 _4097_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3660__A2 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6803_ _6803_/CLK _6803_/D fanout442/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_91_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5937__A1 _6572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5937__B2 _6710_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4995_ _4995_/A _4995_/B VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3948__A0 _3239_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6734_ _6736_/CLK _6734_/D _3959_/B VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfstp_4
X_3946_ _6660_/Q input3/X input1/X VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__mux2_8
XANTENNA__3412__A2 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3877_ hold4/A hold1/A _3878_/S VGND VGND VPWR VPWR _6439_/D sky130_fd_sc_hd__mux2_1
X_6665_ _7107_/CLK _6665_/D fanout451/X VGND VGND VPWR VPWR _7210_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5616_ _6491_/Q _5679_/B _5676_/B VGND VGND VPWR VPWR _5620_/S sky130_fd_sc_hd__and3_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _6830_/CLK _6596_/D fanout440/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5175__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5547_ _5547_/A0 _5583_/A1 _5550_/S VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__mux2_1
X_5478_ _5478_/A0 hold71/X _5478_/S VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7217_ _7217_/A VGND VGND VPWR VPWR _7217_/X sky130_fd_sc_hd__clkbuf_2
X_4429_ _4637_/A _4574_/A _4637_/D VGND VGND VPWR VPWR _4808_/B sky130_fd_sc_hd__and3_4
XFILLER_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout400 hold275/X VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout411 _5872_/B VGND VGND VPWR VPWR _5689_/A sky130_fd_sc_hd__buf_8
XANTENNA__5191__A _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5873__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout433 fanout434/X VGND VGND VPWR VPWR fanout433/X sky130_fd_sc_hd__buf_12
X_7148_ _7180_/CLK _7148_/D fanout448/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout444 fanout449/X VGND VGND VPWR VPWR fanout444/X sky130_fd_sc_hd__buf_12
XFILLER_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout455 _6411_/A VGND VGND VPWR VPWR _6430_/A sky130_fd_sc_hd__buf_6
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout466 fanout470/X VGND VGND VPWR VPWR fanout466/X sky130_fd_sc_hd__buf_12
XFILLER_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7079_ _7086_/CLK _7079_/D fanout467/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A wb_adr_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6050__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3939__A0 _6503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input74_A pad_flash_io1_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6105__A1 _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5305__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5864__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4429__B _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5919__A1 _6532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4164__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _6925_/Q _5344_/A _5542_/A _7101_/Q _3799_/X VGND VGND VPWR VPWR _3801_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4780_ _4947_/A _4688_/A _4544_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21a_1
XFILLER_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3731_ _6693_/Q _4256_/A _4262_/A _6698_/Q VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_csclk _6549_/CLK VGND VGND VPWR VPWR _6786_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6450_ _6809_/CLK _6450_/D fanout433/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_4
X_3662_ _6879_/Q _5290_/A _4128_/A _6581_/Q _3661_/X VGND VGND VPWR VPWR _3662_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5401_ _5401_/A0 _5572_/A1 _5406_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
X_6381_ _6380_/X _6381_/A1 _6384_/S VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__mux2_1
X_3593_ _7040_/Q _3325_/Y _5497_/A _7064_/Q VGND VGND VPWR VPWR _3593_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2443_A _6784_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5332_ _5332_/A0 _5575_/A1 _5334_/S VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__mux2_1
X_5263_ _5263_/A _5578_/B VGND VGND VPWR VPWR _5271_/S sky130_fd_sc_hd__and2_4
XFILLER_88_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2805 hold647/X VGND VGND VPWR VPWR _5360_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7002_ _7140_/CLK _7002_/D fanout473/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_4
X_4214_ _4214_/A0 _5238_/A1 _4217_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
Xhold2816 hold953/X VGND VGND VPWR VPWR _5404_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5194_ _5194_/A0 _5194_/A1 _5199_/S VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__mux2_1
Xhold2827 _7050_/Q VGND VGND VPWR VPWR hold966/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2838 _7130_/Q VGND VGND VPWR VPWR hold954/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2849 _6781_/Q VGND VGND VPWR VPWR _3388_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4145_ _4145_/A0 _5189_/A1 _4145_/S VGND VGND VPWR VPWR _4145_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ _4076_/A0 _5189_/A1 _4076_/S VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6280__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4830__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3633__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6032__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4978_ _4491_/Y _4655_/A _4581_/X _4969_/B _4905_/X VGND VGND VPWR VPWR _5103_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6717_ _6835_/CLK _6717_/D fanout435/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3397__B2 _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3929_ _6655_/Q _6658_/Q VGND VGND VPWR VPWR _3929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6648_ _6761_/CLK _6648_/D _6430_/A VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6579_ _6830_/CLK _6579_/D fanout441/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold1543_A _7036_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6099__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5846__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6271__B1 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4821__A1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3624__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6023__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6326__A1 _6643_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap419 _4751_/C VGND VGND VPWR VPWR _4714_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4888__A1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output278_A _6795_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6262__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5950_ _3241_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7081__RESET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4901_ _5149_/A _4901_/B VGND VGND VPWR VPWR _5098_/B sky130_fd_sc_hd__and2_1
X_5881_ _7167_/Q _5880_/X _6341_/S VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4832_ _4831_/X _4832_/B _4832_/C _4832_/D VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__and4b_1
XANTENNA__3379__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3379__B2 _6948_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4477_/C _4765_/B _4972_/A _4955_/D _5150_/C VGND VGND VPWR VPWR _4764_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4114__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6502_ _6936_/CLK _6502_/D fanout463/X VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfrtp_2
X_3714_ _6966_/Q _5389_/A _4158_/A _6605_/Q VGND VGND VPWR VPWR _3714_/X sky130_fd_sc_hd__a22o_1
X_4694_ _4811_/B _4988_/A _4693_/B VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6433_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
X_3645_ _3645_/A _3645_/B _3645_/C _3645_/D VGND VGND VPWR VPWR _3674_/A sky130_fd_sc_hd__nor4_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3953__S _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6364_ _6684_/Q _6364_/A2 _6364_/B1 _4218_/Y VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__a22o_1
X_3576_ _6944_/Q _5362_/A _5202_/A _6807_/Q _3568_/X VGND VGND VPWR VPWR _3580_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5315_ _5315_/A0 _5567_/A1 _5316_/S VGND VGND VPWR VPWR _5315_/X sky130_fd_sc_hd__mux2_1
X_6295_ _6725_/Q _5978_/X _6008_/X _6740_/Q _6294_/X VGND VGND VPWR VPWR _6295_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5828__B1 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2602 _5208_/X VGND VGND VPWR VPWR hold682/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5246_ _5246_/A0 _5534_/A1 _5253_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
Xhold2613 hold502/X VGND VGND VPWR VPWR _5171_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2624 _7051_/Q VGND VGND VPWR VPWR hold738/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2635 _6843_/Q VGND VGND VPWR VPWR hold743/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__clkdlybuf4s15_2
Xhold1901 hold529/X VGND VGND VPWR VPWR _4178_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2646 _5195_/X VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5177_ _5177_/A0 _5238_/A1 _5177_/S VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1912 _5442_/X VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2657 hold859/X VGND VGND VPWR VPWR _4260_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1923 hold669/X VGND VGND VPWR VPWR _3985_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2668 _6743_/Q VGND VGND VPWR VPWR hold559/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1934 hold546/X VGND VGND VPWR VPWR _4130_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2679 _4303_/X VGND VGND VPWR VPWR hold671/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1945 _7122_/Q VGND VGND VPWR VPWR hold612/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1956 hold286/X VGND VGND VPWR VPWR _5387_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4128_ _4128_/A _5533_/B VGND VGND VPWR VPWR _4133_/S sky130_fd_sc_hd__and2_2
Xhold1967 _7088_/Q VGND VGND VPWR VPWR hold780/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1978 hold515/X VGND VGND VPWR VPWR _4312_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1989 _7220_/A VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6253__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4059_ _4059_/A0 _5572_/A1 _4064_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3606__A2 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4024__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6308__A1 _6632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6733__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3542__A1 _7065_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3542__B2 _6534_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6470__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5819__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6861__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5295__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A mgmt_gpio_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6244__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3781__A1 _6957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold508 hold508/A VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold519 hold519/A VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3430_ _3430_/A _3430_/B VGND VGND VPWR VPWR _3523_/B sky130_fd_sc_hd__nand2_8
XFILLER_171_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3361_ _6852_/Q _5254_/A _4241_/A input60/X VGND VGND VPWR VPWR _3361_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5099_/X _5100_/B _5100_/C _5100_/D VGND VGND VPWR VPWR _5101_/C sky130_fd_sc_hd__and4b_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6080_ _7103_/Q _6008_/X _6016_/X _7039_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3292_ _3347_/A _3354_/A VGND VGND VPWR VPWR _5425_/A sky130_fd_sc_hd__nor2_8
XFILLER_183_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5286__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5031_ _4596_/A _4812_/A _4392_/X VGND VGND VPWR VPWR _5032_/C sky130_fd_sc_hd__a21oi_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 hold101/X VGND VGND VPWR VPWR _5250_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1219 _6714_/Q VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6235__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4109__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6982_ _7072_/CLK _6982_/D fanout460/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5933_ _6622_/Q _5686_/X _5929_/X _5932_/X VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5864_ _6644_/Q _5668_/X _5686_/X _6619_/Q _5863_/X VGND VGND VPWR VPWR _5869_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4815_ _4583_/B _4676_/Y _4688_/A _4729_/A VGND VGND VPWR VPWR _4815_/X sky130_fd_sc_hd__o22a_1
X_5795_ _5816_/A1 _5794_/X _6342_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4013__A2 _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4746_ _4746_/A _4746_/B VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_48_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7126_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4071__C _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5761__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4677_ _4677_/A _4677_/B VGND VGND VPWR VPWR _5049_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6416_ _6416_/A _6423_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
XFILLER_135_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3628_ _6694_/Q _4256_/A _4182_/A _6626_/Q VGND VGND VPWR VPWR _3628_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3524__A1 _7089_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3524__B2 _6701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6347_ _3803_/Y hold997/A _6354_/S VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3559_ _3618_/A1 _4112_/A0 _3857_/B VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2410 _6742_/Q VGND VGND VPWR VPWR hold844/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6278_ _6754_/Q _5638_/X _6007_/X _6532_/Q _6277_/X VGND VGND VPWR VPWR _6279_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4343_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6934__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5277__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _3894_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2421 _4287_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4663_/D sky130_fd_sc_hd__clkbuf_16
Xhold2432 _7033_/Q VGND VGND VPWR VPWR hold777/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6362_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2443 _6784_/Q VGND VGND VPWR VPWR hold901/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5229_ hold64/A hold47/X hold9/A VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__and3_2
Xhold2454 _5570_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1720 _4118_/X VGND VGND VPWR VPWR hold197/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5403__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2465 hold802/X VGND VGND VPWR VPWR _5412_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2476 _6997_/Q VGND VGND VPWR VPWR hold877/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1731 hold453/X VGND VGND VPWR VPWR hold1731/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2487 hold803/X VGND VGND VPWR VPWR _5430_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1742 _4157_/X VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2498 hold838/X VGND VGND VPWR VPWR _5574_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1753 hold440/X VGND VGND VPWR VPWR hold1753/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5029__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1764 hold821/X VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1775 _6907_/Q VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6226__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4019__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1786 _4183_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1797 hold403/X VGND VGND VPWR VPWR _4097_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4262__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5752__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3763__A1 _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_90 _6238_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5268__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5313__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output310_A _3966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4779__B1 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3451__B1 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4600_ _4402_/Y _4570_/A _4658_/B _4564_/Y VGND VGND VPWR VPWR _4609_/B sky130_fd_sc_hd__o22a_1
X_5580_ hold200/X _5580_/A1 _5586_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5743__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _5117_/A _4531_/B _5095_/A VGND VGND VPWR VPWR _4533_/C sky130_fd_sc_hd__and3_1
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2356_A _6525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold305 hold305/A VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4462_ _4477_/A _4477_/B _4955_/C VGND VGND VPWR VPWR _4462_/Y sky130_fd_sc_hd__nand3_4
Xhold327 hold327/A VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold338 hold338/A VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6201_ _6980_/Q _5976_/B _5978_/X _7124_/Q _6200_/X VGND VGND VPWR VPWR _6204_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3413_ _7123_/Q _5560_/A _5362_/A _6947_/Q VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__a22o_1
X_4393_ _4720_/C _4649_/B VGND VGND VPWR VPWR _4650_/B sky130_fd_sc_hd__nor2_8
X_7181_ _7184_/CLK _7181_/D fanout443/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6905_/Q _5985_/X _5989_/X _6897_/Q VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__a22o_1
X_3344_ _3563_/A _3764_/A VGND VGND VPWR VPWR _4241_/A sky130_fd_sc_hd__nor2_8
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6056_/X _6058_/X _6063_/C _6339_/B VGND VGND VPWR VPWR _6064_/C sky130_fd_sc_hd__and4bb_1
X_3275_ _3347_/A _3343_/A VGND VGND VPWR VPWR _5452_/A sky130_fd_sc_hd__nor2_8
Xhold1005 _6514_/Q VGND VGND VPWR VPWR _4053_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7141__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1016 hold1/X VGND VGND VPWR VPWR _3982_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1027 _3325_/Y VGND VGND VPWR VPWR _5470_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5014_ _5009_/A _5009_/B _4719_/B VGND VGND VPWR VPWR _5014_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1038 _5541_/S VGND VGND VPWR VPWR _5540_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1049 _5304_/X VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4347__B _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6208__B1 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3251__B _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3690__B1 _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6965_ _6974_/CLK _6965_/D fanout450/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5431__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5916_ _6641_/Q _5655_/X _5663_/X _6631_/Q _5905_/Y VGND VGND VPWR VPWR _5916_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3442__B1 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6896_ _6996_/CLK _6896_/D fanout462/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5178__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3993__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _6956_/Q _5672_/X _5679_/X _6908_/Q _5846_/X VGND VGND VPWR VPWR _5847_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5734__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5778_ _7033_/Q _5655_/X _5668_/X _7057_/Q VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4729_/A _4995_/A VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5498__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold850 hold850/A VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold861 hold861/A VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold872 hold872/A VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold894 hold894/A VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4538__A _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2240 _6791_/Q VGND VGND VPWR VPWR hold566/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2251 _4142_/X VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2262 hold599/X VGND VGND VPWR VPWR _5265_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2273 hold840/X VGND VGND VPWR VPWR _4216_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input139_A wb_dat_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2284 hold781/X VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2295 hold578/X VGND VGND VPWR VPWR _4252_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1550 hold322/X VGND VGND VPWR VPWR _5298_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1992_A _6501_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1561 _6860_/Q VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1572 _5369_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1583 hold512/X VGND VGND VPWR VPWR _4313_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3681__B1 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1594 hold387/X VGND VGND VPWR VPWR _5316_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_60_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3433__B1 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5725__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5489__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output260_A _6803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7164__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6150__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4161__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5551__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3672__B1 _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5413__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _6760_/CLK _6750_/D fanout441/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfrtp_4
X_3962_ _6456_/Q _3962_/B VGND VGND VPWR VPWR _3963_/A sky130_fd_sc_hd__nor2_2
XANTENNA__5964__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5701_ _6981_/Q _5656_/X _5663_/X _7021_/Q _5700_/X VGND VGND VPWR VPWR _5701_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _3950_/A1 _6681_/D _4107_/B VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3893_ input123/X input122/X _3893_/C _3893_/D VGND VGND VPWR VPWR _3900_/B sky130_fd_sc_hd__and4bb_1
XFILLER_176_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5632_ _6491_/Q _6015_/B _6014_/A VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__and3_1
XANTENNA__5716__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__A1 input72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3727__B2 _6488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5563_ _5563_/A0 _5563_/A1 _5568_/S VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4514_ _4729_/A _4514_/B VGND VGND VPWR VPWR _4514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold102 hold102/A VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5494_ _5494_/A0 _5575_/A1 _5496_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
Xhold113 hold113/A VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold124 hold124/A VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold135 hold135/A VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7233_ _7233_/A VGND VGND VPWR VPWR _7233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4445_ _4485_/B _4564_/B VGND VGND VPWR VPWR _4483_/B sky130_fd_sc_hd__and2_4
Xhold146 _4173_/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold157 hold157/A VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7164_ _7185_/CLK _7164_/D fanout446/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
X_4376_ _4649_/B _4560_/A VGND VGND VPWR VPWR _4384_/A sky130_fd_sc_hd__nand2_8
XFILLER_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5461__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6115_ _6840_/Q _6339_/B _6114_/X VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__o21ba_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3327_ _3338_/A _3535_/A VGND VGND VPWR VPWR _5488_/A sky130_fd_sc_hd__nor2_8
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7135_/CLK _7095_/D fanout466/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout389_A _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _7078_/Q _6013_/X _6017_/X _7070_/Q VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4077__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3258_ _3259_/B VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__inv_2
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6681__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3189_ _6680_/D VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3415__B1 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6948_ _6963_/CLK _6948_/D fanout465/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5955__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6879_ _6977_/CLK _6879_/D fanout460/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3718__A1 _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3718__B2 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4032__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6132__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4143__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold680 hold680/A VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold691 hold691/A VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5891__A1 _6570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5371__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5891__B2 _6708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2070 _6956_/Q VGND VGND VPWR VPWR hold357/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2081 _4208_/X VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2092 hold667/X VGND VGND VPWR VPWR _3979_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1380 _6966_/Q VGND VGND VPWR VPWR hold251/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1391 _5428_/X VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6199__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3236_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput218 _7214_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput229 _7224_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6123__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2054_A _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4230_ _4230_/A0 _4229_/X _4240_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5281__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4161_ _4161_/A0 _5581_/A1 _4163_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ _4092_/A _5220_/C VGND VGND VPWR VPWR _4097_/S sky130_fd_sc_hd__and2_2
XFILLER_83_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5501__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6802_ _6821_/CLK _6802_/D fanout442/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_2
X_4994_ _4676_/Y _4812_/Y _4993_/Y _5138_/B VGND VGND VPWR VPWR _5010_/B sky130_fd_sc_hd__o211a_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5937__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6733_ _6733_/CLK _6733_/D _3959_/B VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtp_4
X_3945_ _3944_/X _3966_/B _6456_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_8
XANTENNA__3956__S _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6664_ _7108_/CLK _6664_/D fanout451/X VGND VGND VPWR VPWR _7209_/A sky130_fd_sc_hd__dfrtp_1
X_3876_ hold1/A hold41/A _3878_/S VGND VGND VPWR VPWR _6440_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5615_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5676_/B sky130_fd_sc_hd__nor2_8
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6595_ _6752_/CLK _6595_/D fanout440/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5546_ _5546_/A0 _5582_/A1 _5550_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ _5477_/A0 wire371/X _5478_/S VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4125__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7216_ _7216_/A VGND VGND VPWR VPWR _7216_/X sky130_fd_sc_hd__clkbuf_2
X_4428_ _4637_/B _4637_/A VGND VGND VPWR VPWR _4463_/B sky130_fd_sc_hd__nand2b_4
Xfanout401 hold275/X VGND VGND VPWR VPWR _5561_/A1 sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR net399_2/A
+ sky130_fd_sc_hd__clkbuf_16
Xfanout412 _5872_/B VGND VGND VPWR VPWR _5685_/A sky130_fd_sc_hd__buf_4
XANTENNA__5191__B _5220_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7179_/CLK _7147_/D fanout447/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfstp_4
Xfanout434 _3959_/B VGND VGND VPWR VPWR fanout434/X sky130_fd_sc_hd__buf_12
X_4359_ _4682_/A _4365_/B _4447_/B VGND VGND VPWR VPWR _4360_/B sky130_fd_sc_hd__a21o_1
Xfanout445 fanout449/X VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__buf_6
XFILLER_59_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout456 _6416_/A VGND VGND VPWR VPWR _6413_/A sky130_fd_sc_hd__buf_12
Xfanout467 fanout470/X VGND VGND VPWR VPWR fanout467/X sky130_fd_sc_hd__buf_12
XFILLER_86_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7078_ _7078_/CLK _7078_/D fanout445/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6029_ _7093_/Q _5984_/X _6020_/X _6024_/X _6028_/X VGND VGND VPWR VPWR _6029_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_100_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5411__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1690_A _6689_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4027__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1955_A _6963_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input67_A mgmt_gpio_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6105__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7202__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5321__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5919__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _7094_/Q hold31/A _5178_/A _6785_/Q _3729_/X VGND VGND VPWR VPWR _3735_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3661_ _6550_/Q _4092_/A _4134_/A _6586_/Q VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__a22o_1
X_5400_ _5400_/A0 _5571_/A1 _5406_/S VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__mux2_1
X_6380_ _6686_/Q _6380_/A2 _6380_/B1 _4218_/Y _6379_/X VGND VGND VPWR VPWR _6380_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ _7000_/Q _5425_/A _4304_/A _6735_/Q _3591_/X VGND VGND VPWR VPWR _3595_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5331_/A0 _5529_/A1 _5334_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5262_ _5262_/A0 _5568_/A1 _5262_/S VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7001_ _7001_/CLK _7001_/D fanout466/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2806 _5360_/X VGND VGND VPWR VPWR hold648/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4213_ _4213_/A0 _5543_/A1 _4217_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2817 _6814_/Q VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5193_ _5193_/A0 _5193_/A1 _5199_/S VGND VGND VPWR VPWR _5193_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2828 hold966/X VGND VGND VPWR VPWR _5485_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2839 hold954/X VGND VGND VPWR VPWR _5575_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4144_ _4144_/A0 _5195_/A1 _4145_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _4075_/A0 _5195_/A1 _4076_/S VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5231__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6280__A1 _6631_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6280__B2 _6771_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4830__A2 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6032__A1 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6032__B2 _6869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4977_ _4569_/C _4968_/Y _4971_/Y _4972_/Y VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__o211a_1
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6716_ _7121_/CLK _6716_/D _6399_/A VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3397__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5791__B1 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3928_ _6657_/Q _3904_/A _3904_/Y _3928_/B2 VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__a22o_1
XFILLER_177_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6647_ _6760_/CLK _6647_/D _6433_/A VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6335__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3859_ _6470_/Q _3879_/A _6468_/Q _6654_/Q VGND VGND VPWR VPWR _3860_/S sky130_fd_sc_hd__and4b_1
XFILLER_164_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6578_ _6745_/CLK _6578_/D fanout440/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5529_ _5529_/A0 _5529_/A1 _5532_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5406__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6099__A1 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6099__B2 _6848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5846__B2 _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3609__B1 _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6271__A1 _6586_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input121_A wb_adr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4821__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_csclk_A _3955_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6023__A1 _6877_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6023__B2 _6845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6326__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4337__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap409 _3857_/B VGND VGND VPWR VPWR _3738_/S sky130_fd_sc_hd__buf_4
XFILLER_6_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4888__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output173_A _3973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5316__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6262__A1 _6585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6262__B2 _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4900_ _4947_/B _4570_/D _4616_/A VGND VGND VPWR VPWR _5063_/C sky130_fd_sc_hd__o21a_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5880_ _5869_/Y _5879_/Y _6525_/Q _5678_/Y VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_179_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4831_ _4955_/D _4718_/C _5026_/C _4812_/A VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__a22o_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6390__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3379__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4762_ _4402_/Y _4583_/B _4426_/Y VGND VGND VPWR VPWR _4791_/A sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_6_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6501_ _6936_/CLK _6501_/D fanout463/X VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfrtp_2
X_3713_ _6894_/Q _5308_/A _3539_/Y _6531_/Q _3712_/X VGND VGND VPWR VPWR _3716_/C
+ sky130_fd_sc_hd__a221o_1
X_4693_ _4811_/B _4693_/B VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
X_3644_ _7023_/Q _5452_/A _4237_/S _3879_/B _3643_/X VGND VGND VPWR VPWR _3645_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_162_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6363_ _6362_/X hold273/A _6384_/S VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3575_ _6725_/Q _4292_/A _4164_/A _6612_/Q _3574_/X VGND VGND VPWR VPWR _3580_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5314_ _5314_/A0 _5575_/A1 _5316_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3551__A2 _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6294_ hold67/A _5977_/X _6007_/X _6533_/Q _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5245_ _5245_/A _5569_/B VGND VGND VPWR VPWR _5253_/S sky130_fd_sc_hd__and2_4
Xhold2603 _6692_/Q VGND VGND VPWR VPWR hold692/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2614 _5171_/X VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2625 hold738/X VGND VGND VPWR VPWR _5486_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkbuf_8
Xhold2636 hold743/X VGND VGND VPWR VPWR _5252_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2647 _6801_/Q VGND VGND VPWR VPWR hold805/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1902 _4178_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__buf_2
Xhold1913 _7112_/Q VGND VGND VPWR VPWR hold767/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5176_ _5176_/A0 _5543_/A1 _5177_/S VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__mux2_1
Xhold2658 _4260_/X VGND VGND VPWR VPWR hold860/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1924 _3985_/X VGND VGND VPWR VPWR _6453_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2669 hold559/X VGND VGND VPWR VPWR _4318_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1935 _4130_/X VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1946 hold612/X VGND VGND VPWR VPWR _5566_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4127_ _4127_/A0 _5277_/A1 _4127_/S VGND VGND VPWR VPWR _4127_/X sky130_fd_sc_hd__mux2_1
Xhold1957 _5387_/X VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1968 hold780/X VGND VGND VPWR VPWR _5528_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5056__A2 _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1979 _4312_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4058_ _4058_/A0 _5562_/A1 _4064_/S VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5764__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6308__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4319__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3790__A2 _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4040__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3542__A2 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input169_A wb_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5819__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3781__A2 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold509 hold509/A VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6180__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3360_ _6802_/Q _3319_/Y _3336_/Y input28/X VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a22o_2
XFILLER_124_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3764_/A _3354_/B VGND VGND VPWR VPWR _3291_/Y sky130_fd_sc_hd__nor2_8
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5030_ _4417_/B _4688_/B _4774_/X _4963_/A _4894_/A VGND VGND VPWR VPWR _5149_/B
+ sky130_fd_sc_hd__o2111a_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1209 _5250_/X VGND VGND VPWR VPWR hold102/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2301_A _6608_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6981_ _7001_/CLK _6981_/D fanout466/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfstp_4
X_5932_ _6647_/Q _5668_/X _5684_/X _6607_/Q VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4797__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5863_ _6535_/Q _5651_/X _5658_/X _6692_/Q VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4633__B _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4814_ _4583_/B _4688_/B _4691_/Y _4729_/A VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__o22a_1
XANTENNA__5746__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5794_ _5794_/A0 _5793_/X _6341_/S VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4745_ _5011_/A _4947_/A _4714_/Y VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3964__S _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3772__A2 _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4676_ _4751_/B _4676_/B VGND VGND VPWR VPWR _4676_/Y sky130_fd_sc_hd__nand2_8
XFILLER_147_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6415_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
X_3627_ _3627_/A _3627_/B _3627_/C _3627_/D VGND VGND VPWR VPWR _3675_/A sky130_fd_sc_hd__nor4_2
XANTENNA__6171__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3524__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6346_ _6677_/Q _6346_/B VGND VGND VPWR VPWR _6354_/S sky130_fd_sc_hd__nand2_8
X_3558_ _3558_/A _3558_/B _3558_/C VGND VGND VPWR VPWR _3558_/Y sky130_fd_sc_hd__nand3_2
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6277_ _6626_/Q _6013_/X _6015_/X _6759_/Q VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2400 hold629/X VGND VGND VPWR VPWR _5180_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3489_ _6711_/Q _4274_/A _4256_/A _6696_/Q VGND VGND VPWR VPWR _3489_/X sky130_fd_sc_hd__a22o_1
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4343_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2411 hold844/X VGND VGND VPWR VPWR _4317_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2422 _6643_/Q VGND VGND VPWR VPWR hold865/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5228_ _5228_/A0 _5228_/A1 _5228_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4345_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2433 hold777/X VGND VGND VPWR VPWR _5466_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2444 hold901/X VGND VGND VPWR VPWR _5179_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2455 _7002_/Q VGND VGND VPWR VPWR hold636/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1710 hold976/X VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2466 _5412_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1721 _6543_/Q VGND VGND VPWR VPWR hold969/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2477 hold877/X VGND VGND VPWR VPWR _5426_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1732 _6902_/Q VGND VGND VPWR VPWR hold589/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1743 _6556_/Q VGND VGND VPWR VPWR hold974/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5159_ _5157_/X _5158_/X _5127_/X VGND VGND VPWR VPWR _5159_/Y sky130_fd_sc_hd__a21boi_1
Xhold2488 _5430_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2499 _5574_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1754 _6564_/Q VGND VGND VPWR VPWR hold973/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1765 _4186_/X VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1776 hold306/X VGND VGND VPWR VPWR _5324_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1787 _7131_/Q VGND VGND VPWR VPWR hold247/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1798 _4097_/X VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4788__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4035__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3874__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__A2 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 hold332/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_91 _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6162__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4476__B1 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4779__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6695__RESET_B fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4530_ _4574_/A _4463_/B _4510_/A _4509_/Y _4529_/X VGND VGND VPWR VPWR _4533_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3754__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4461_ _4506_/A _4461_/B VGND VGND VPWR VPWR _4955_/C sky130_fd_sc_hd__nor2_2
XANTENNA__6153__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold317 _5243_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold328 hold328/A VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold339 hold339/A VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6200_ _6932_/Q _5982_/X _5999_/X _6868_/Q VGND VGND VPWR VPWR _6200_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3506__A2 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3412_ _6963_/Q _5380_/A _3407_/X _3409_/X _3411_/X VGND VGND VPWR VPWR _3422_/B
+ sky130_fd_sc_hd__a2111oi_4
X_7180_ _7180_/CLK _7180_/D fanout446/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_1
X_4392_ _4955_/A _5009_/A _4580_/A VGND VGND VPWR VPWR _4392_/X sky130_fd_sc_hd__and3_1
XFILLER_125_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _7113_/Q _5987_/X _6004_/X _6881_/Q _6130_/X VGND VGND VPWR VPWR _6131_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3343_ _3343_/A _3354_/B VGND VGND VPWR VPWR _5380_/A sky130_fd_sc_hd__nor2_8
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5504__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6902_/Q _5985_/X _6059_/X _6061_/X VGND VGND VPWR VPWR _6063_/C sky130_fd_sc_hd__a211oi_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3355_/A hold79/X VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__nand2_8
Xhold1006 hold1210/X VGND VGND VPWR VPWR hold1211/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4628__B _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1017 _3982_/X VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5013_ _4688_/C _4995_/B _5012_/X _4820_/A VGND VGND VPWR VPWR _5023_/C sky130_fd_sc_hd__o211a_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _5470_/X VGND VGND VPWR VPWR _5478_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1039 _5536_/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6208__B2 _6964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3690__A1 _6942_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6964_ _7099_/CLK _6964_/D fanout471/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
X_5915_ _6689_/Q _5659_/X _5687_/X _6601_/Q VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3442__A1 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6895_ _6977_/CLK _6895_/D fanout460/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5719__B1 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5846_ _6940_/Q _5659_/X _5687_/X _6924_/Q VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5195__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _6881_/Q _5667_/X _5673_/X _6865_/Q _5776_/X VGND VGND VPWR VPWR _5782_/B
+ sky130_fd_sc_hd__a221o_2
X_4728_ _5150_/B _4730_/B VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6144__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4659_ _4652_/Y _4677_/B VGND VGND VPWR VPWR _4704_/C sky130_fd_sc_hd__nand2b_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold840 hold840/A VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold851 hold851/A VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 hold862/A VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold873 hold873/A VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold884 _4052_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6329_ _6711_/Q _5992_/X _6012_/X _6751_/Q _6328_/X VGND VGND VPWR VPWR _6329_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold895 hold895/A VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5414__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2230 _4294_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2241 hold566/X VGND VGND VPWR VPWR _5187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2252 _6870_/Q VGND VGND VPWR VPWR hold588/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2263 _5265_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2274 _4216_/X VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2285 _4305_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1540 _6988_/Q VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2296 _4252_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1551 _7060_/Q VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1562 hold365/X VGND VGND VPWR VPWR _5271_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7153__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1573 _6940_/Q VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1584 _4313_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3681__B2 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1595 _5316_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3433__A1 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input97_A usr2_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5186__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6135__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4729__A _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5324__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6969_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3672__A1 _6481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5949__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3961_ _3961_/A VGND VGND VPWR VPWR _3961_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5700_ _7013_/Q _5664_/X _5666_/X _6997_/Q VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6680_ _7203_/CLK _6680_/D _4107_/B VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3892_ _4720_/C _4649_/B _4649_/C _4649_/D VGND VGND VPWR VPWR _4395_/A sky130_fd_sc_hd__a211o_4
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5631_ _5631_/A _6017_/B VGND VGND VPWR VPWR _5634_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5177__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5562_ _5562_/A0 _5562_/A1 _5568_/S VGND VGND VPWR VPWR _5562_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3727__A2 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4513_ _4513_/A _4513_/B _4652_/A VGND VGND VPWR VPWR _4514_/B sky130_fd_sc_hd__nand3_4
XANTENNA__6126__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5493_ _5493_/A0 _5583_/A1 _5496_/S VGND VGND VPWR VPWR _5493_/X sky130_fd_sc_hd__mux2_1
Xhold103 hold103/A VGND VGND VPWR VPWR hold103/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold114 hold114/A VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7232_ _7232_/A VGND VGND VPWR VPWR _7232_/X sky130_fd_sc_hd__clkbuf_2
Xhold125 hold125/A VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4444_ _4506_/A _4469_/B VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__nor2_4
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold147 hold147/A VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold158 _4271_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold169 hold169/A VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7163_ _7185_/CLK _7163_/D fanout443/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_1
X_4375_ _4649_/B _4560_/A VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__and2_4
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5234__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3360__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6114_ _6105_/X _6313_/D _6114_/C _6114_/D VGND VGND VPWR VPWR _6114_/X sky130_fd_sc_hd__and4b_4
XANTENNA__4012__A_N _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3326_ hold30/A hold15/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__nor2_8
X_7094_ _7094_/CLK _7094_/D fanout450/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _7054_/Q _5990_/X _5997_/X _6950_/Q _6044_/X VGND VGND VPWR VPWR _6045_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3257_ hold53/X _5167_/A1 _3998_/S VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3188_ _3188_/A VGND VGND VPWR VPWR _4222_/B sky130_fd_sc_hd__inv_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout451_A fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3415__A1 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6947_ _6992_/CLK _6947_/D fanout465/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6878_ _7063_/CLK _6878_/D fanout460/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5829_ _7067_/Q _5671_/X _5678_/B _6971_/Q _5707_/B VGND VGND VPWR VPWR _5829_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5409__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__A2 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5340__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold670 hold670/A VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4549__A _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 hold681/A VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold692 hold692/A VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input151_A wb_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5891__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4268__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2060 hold919/X VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2071 hold357/X VGND VGND VPWR VPWR _5379_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2082 _6700_/Q VGND VGND VPWR VPWR hold757/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2093 _3979_/X VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3654__A1 _7039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1370 _7009_/Q VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input12_A mask_rev_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1381 hold251/X VGND VGND VPWR VPWR _5391_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _6576_/Q VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5319__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3709__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6108__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput208 _3235_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XANTENNA__3590__B1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput219 _7215_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_max_cap347_A _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5331__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4160_ _4160_/A0 _5580_/A1 _4163_/S VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7075__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ _3385_/Y hold988/A _4091_/S VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6393__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4194__A _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6801_ _6821_/CLK _6801_/D fanout443/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfstp_4
X_4993_ _4993_/A _4993_/B VGND VGND VPWR VPWR _4993_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6732_ _6736_/CLK _6732_/D _3959_/B VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_4
X_3944_ _3943_/X input38/X _6458_/Q VGND VGND VPWR VPWR _3944_/X sky130_fd_sc_hd__mux2_2
XANTENNA__4070__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6347__A0 _3803_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6663_ _6832_/CLK _6663_/D fanout447/X VGND VGND VPWR VPWR _7208_/A sky130_fd_sc_hd__dfrtp_1
X_3875_ hold41/A hold93/A _3878_/S VGND VGND VPWR VPWR _6441_/D sky130_fd_sc_hd__mux2_1
XANTENNA_hold2750_A _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5614_ _5614_/A1 _5613_/B _5611_/Y _5613_/Y VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__a31o_1
XFILLER_176_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6594_ _6752_/CLK _6594_/D fanout440/X VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5570__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5545_ _5545_/A0 _5563_/A1 _5550_/S VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5476_ _5476_/A0 _5584_/A1 _5478_/S VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5858__C1 _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7215_ _7215_/A VGND VGND VPWR VPWR _7215_/X sky130_fd_sc_hd__clkbuf_2
X_4427_ _4637_/B _4637_/A VGND VGND VPWR VPWR _4488_/B sky130_fd_sc_hd__and2b_4
XANTENNA__5322__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout402 hold275/X VGND VGND VPWR VPWR _5579_/A1 sky130_fd_sc_hd__buf_6
Xfanout413 _7150_/Q VGND VGND VPWR VPWR _5872_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold1147_A _7055_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7146_ _7180_/CLK _7146_/D fanout447/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5191__C _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5873__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4358_ _4513_/A _4560_/A VGND VGND VPWR VPWR _4955_/A sky130_fd_sc_hd__and2b_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout435 fanout436/X VGND VGND VPWR VPWR fanout435/X sky130_fd_sc_hd__buf_12
XANTENNA__3884__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout446 fanout448/X VGND VGND VPWR VPWR fanout446/X sky130_fd_sc_hd__buf_12
XFILLER_113_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input4_A mask_rev_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout457 _6411_/A VGND VGND VPWR VPWR _6416_/A sky130_fd_sc_hd__buf_12
Xfanout468 fanout469/X VGND VGND VPWR VPWR fanout468/X sky130_fd_sc_hd__buf_12
XFILLER_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3309_ _3309_/A _3430_/B VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__nand2_8
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7077_ _7078_/CLK _7077_/D fanout447/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfstp_2
X_4289_ hold632/X _5194_/A1 _4291_/S VGND VGND VPWR VPWR _4289_/X sky130_fd_sc_hd__mux2_1
X_6028_ _7101_/Q _6008_/X _6026_/X _6027_/X _5976_/X VGND VGND VPWR VPWR _6028_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_86_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7154__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6050__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4061__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4043__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1948_A _6944_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5561__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5313__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5864__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4824__B1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6041__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6329__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ _6935_/Q _5353_/A _5202_/A _6806_/Q VGND VGND VPWR VPWR _3660_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5552__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3591_ _6647_/Q _4206_/A _4194_/A _6637_/Q VGND VGND VPWR VPWR _3591_/X sky130_fd_sc_hd__a22o_1
X_5330_ _5330_/A0 _5537_/A1 _5334_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5304__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ _5261_/A0 _5567_/A1 _5262_/S VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7000_ _7128_/CLK _7000_/D fanout468/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5855__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4212_ _4212_/A hold9/A VGND VGND VPWR VPWR _4217_/S sky130_fd_sc_hd__and2_2
Xhold2807 _6914_/Q VGND VGND VPWR VPWR hold962/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5192_ hold773/X _5534_/A1 _5199_/S VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__mux2_1
Xhold2818 hold793/X VGND VGND VPWR VPWR _5216_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2829 _6661_/Q VGND VGND VPWR VPWR hold935/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4143_ hold561/X _5194_/A1 _4145_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5512__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4074_ _4074_/A0 _5194_/A1 _4076_/S VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4815__B1 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7177__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6280__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4291__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6032__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4043__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4976_ _4976_/A _4976_/B VGND VGND VPWR VPWR _4985_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6715_ _7121_/CLK hold90/X _6399_/A VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3927_ _3927_/A1 _6437_/Q _3850_/S _3904_/A _3862_/A VGND VGND VPWR VPWR _3927_/Y
+ sky130_fd_sc_hd__o32ai_1
XFILLER_50_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6646_ _6761_/CLK _6646_/D _6430_/A VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfstp_1
X_3858_ _3879_/B _3858_/A1 _3858_/S VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5543__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6577_ _6745_/CLK _6577_/D fanout441/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_4
X_3789_ _6917_/Q _5335_/A _4274_/A _6707_/Q _3788_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_117_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5528_ _5528_/A0 _5582_/A1 _5532_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6099__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5459_ _5459_/A0 _5567_/A1 _5460_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5846__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7129_ _7135_/CLK _7129_/D fanout470/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5422__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3609__A1 _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3609__B2 _6632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6271__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4038__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4282__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input114_A wb_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4821__A3 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3877__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6023__A2 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3793__B1 _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5534__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3545__B1 _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5332__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6262__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4273__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _4417_/B _4633_/B _4384_/A _4658_/A VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__a211o_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4761_ _4625_/A _5033_/A _4976_/A VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6500_ _7125_/CLK _6500_/D fanout468/X VGND VGND VPWR VPWR _7221_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3784__B1 _4009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3712_ _6723_/Q _4292_/A _4146_/A _6595_/Q VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4692_ _4676_/Y _4688_/X _4691_/Y _5011_/B VGND VGND VPWR VPWR _4692_/X sky130_fd_sc_hd__a31o_1
XFILLER_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5525__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6431_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
X_3643_ _6991_/Q _5416_/A _4047_/C input45/X VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5507__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2546_A _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6362_ _6684_/Q _6362_/A2 _6362_/B1 _4218_/Y _6361_/X VGND VGND VPWR VPWR _6362_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3574_ input46/X _4047_/C _5560_/A _7120_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_4
XANTENNA__7090__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5313_ _5313_/A0 _5448_/A1 _5316_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
X_6293_ _6617_/Q _5984_/X _5998_/X _6582_/Q VGND VGND VPWR VPWR _6293_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2713_A _6958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5828__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5244_ _5244_/A0 _5577_/A1 _5244_/S VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2604 hold692/X VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2615 _6588_/Q VGND VGND VPWR VPWR hold931/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2626 _6575_/Q VGND VGND VPWR VPWR hold552/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2637 _5252_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5175_ _5175_/A _5220_/C VGND VGND VPWR VPWR _5177_/S sky130_fd_sc_hd__and2_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__buf_2
Xhold1903 _7214_/A VGND VGND VPWR VPWR hold933/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2648 hold805/X VGND VGND VPWR VPWR _5198_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5242__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1914 hold767/X VGND VGND VPWR VPWR _5555_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2659 _6618_/Q VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1925 _6816_/Q VGND VGND VPWR VPWR hold939/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4126_ _4126_/A0 _5233_/A1 _4127_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
Xhold1936 _6619_/Q VGND VGND VPWR VPWR hold694/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1947 _5566_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1958 _7080_/Q VGND VGND VPWR VPWR hold851/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1969 _5528_/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6253__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4057_ _4057_/A0 _5579_/A1 _4064_/S VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4264__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4016__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5764__A1 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__nor2_1
XFILLER_193_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5516__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6629_ _6794_/CLK _6629_/D fanout434/X VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5417__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5819__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6244__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4255__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__B2 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3766__B1 _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5507__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5327__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3518__B1 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4231__S _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3290_ hold62/X _3290_/B VGND VGND VPWR VPWR _3354_/B sky130_fd_sc_hd__nand2_8
XFILLER_124_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6235__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4246__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6980_ _7107_/CLK _6980_/D fanout452/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5931_ _6533_/Q _5653_/X _5662_/X _6587_/Q _5930_/X VGND VGND VPWR VPWR _5931_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4797__A2 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5862_ _6574_/Q _5667_/X _5688_/X _6579_/Q _5861_/X VGND VGND VPWR VPWR _5869_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _5009_/A _4607_/B _4811_/B VGND VGND VPWR VPWR _5104_/C sky130_fd_sc_hd__o21ai_4
X_5793_ _5782_/Y _5792_/Y _6841_/Q _5678_/Y VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5746__B2 _6959_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3757__B1 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4744_ _4415_/B _4713_/Y _4743_/Y VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__o21ai_1
XFILLER_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4675_ _4675_/A _4683_/A VGND VGND VPWR VPWR _4725_/B sky130_fd_sc_hd__nor2_1
XANTENNA__7200__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5237__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2928_A _6458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3626_ _3971_/A _3431_/Y _4158_/A _6606_/Q _3625_/X VGND VGND VPWR VPWR _3627_/D
+ sky130_fd_sc_hd__a221o_1
X_6414_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
XFILLER_190_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6345_ _6683_/D _3922_/B _6344_/Y _6345_/B2 VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__a22o_1
X_3557_ _3557_/A _3557_/B _3557_/C _3557_/D VGND VGND VPWR VPWR _3558_/C sky130_fd_sc_hd__and4_2
XANTENNA__3980__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6276_ _6729_/Q _5987_/X _6014_/X _6744_/Q _6275_/X VGND VGND VPWR VPWR _6279_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3488_ _3550_/A _3553_/B VGND VGND VPWR VPWR _4256_/A sky130_fd_sc_hd__nor2_8
XFILLER_142_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2401 _5180_/X VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4343_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5227_ _5227_/A0 _5534_/A1 _5228_/S VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__mux2_1
Xhold2412 _4317_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2423 hold865/X VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2434 _5466_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1700 hold198/X VGND VGND VPWR VPWR _4029_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2445 _5179_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1711 hold436/X VGND VGND VPWR VPWR hold1711/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2456 hold636/X VGND VGND VPWR VPWR _5431_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2467 _6534_/Q VGND VGND VPWR VPWR hold878/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1722 hold969/X VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5158_ _4583_/B _4691_/Y _5058_/C _5121_/X VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__o211a_1
Xhold2478 _5426_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1733 _5319_/X VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2489 _6567_/Q VGND VGND VPWR VPWR hold971/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1744 hold974/X VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1755 hold973/X VGND VGND VPWR VPWR hold442/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6226__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4109_ _3737_/Y _4109_/A1 _4115_/S VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1766 _6557_/Q VGND VGND VPWR VPWR hold990/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5089_ _5089_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _5136_/C sky130_fd_sc_hd__and3_1
Xhold1777 _5324_/X VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4237__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1788 hold247/X VGND VGND VPWR VPWR _5576_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1799 _6638_/Q VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5001__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3748__B1 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_70 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_81 hold354/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4051__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A mgmt_gpio_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4476__A1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4226__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3451__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5728__B2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4460_ _4579_/B _4564_/C _4881_/A VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__nand3_4
XFILLER_171_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6153__A1 _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold307 hold307/A VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 hold318/A VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3411_ _6801_/Q _3319_/Y hold16/A _7051_/Q _3410_/X VGND VGND VPWR VPWR _3411_/X
+ sky130_fd_sc_hd__a221o_4
Xhold329 hold329/A VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4391_ _5009_/A _4580_/A VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__5900__A1 _6585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6130_ _6913_/Q _5991_/X _6005_/X _6945_/Q VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3342_ _3343_/A _3346_/A VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__nor2_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6396__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _7134_/Q _5977_/X _5995_/X _6918_/Q _6060_/X VGND VGND VPWR VPWR _6061_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3273_ _3355_/A hold79/X VGND VGND VPWR VPWR _5226_/A sky130_fd_sc_hd__and2_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1007 _7228_/A VGND VGND VPWR VPWR _4248_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_5012_ _5011_/A _4590_/Y _4688_/A VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__a21o_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 hold175/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1029 _5473_/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6208__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5520__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3690__A2 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5967__A1 _6539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6963_ _6963_/CLK _6963_/D fanout464/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3978__A0 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5914_ _6550_/Q _5673_/X _5909_/X _5911_/X _5913_/X VGND VGND VPWR VPWR _5914_/X
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__3442__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6894_ _6967_/CLK _6894_/D fanout465/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5719__A1 _6942_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _6980_/Q _5660_/X _5669_/X _7052_/Q VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5719__B2 _7086_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6351__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _7049_/Q _5669_/X _5687_/X _6921_/Q VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4727_/A _4993_/B VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_hold1177_A _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4658_ _4658_/A _4658_/B VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_2
X_3609_ _7008_/Q _5434_/A _4188_/A _6632_/Q VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__a22o_1
Xhold830 hold830/A VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4589_ _4637_/D _5011_/B VGND VGND VPWR VPWR _5009_/B sky130_fd_sc_hd__nor2_8
Xhold852 hold852/A VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold863 hold863/A VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold874 hold874/A VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6328_ _6701_/Q _5997_/X _6004_/X _6578_/Q VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a22o_1
Xhold885 hold885/A VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold896 hold896/A VGND VGND VPWR VPWR hold896/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2220 _6986_/Q VGND VGND VPWR VPWR hold608/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6259_ _6738_/Q _6008_/X _6016_/X _6451_/Q VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2231 _7034_/Q VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2242 _5187_/X VGND VGND VPWR VPWR hold567/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2253 hold588/X VGND VGND VPWR VPWR _5283_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2264 _6707_/Q VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1530 _5504_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2275 _7068_/Q VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2286 _7100_/Q VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1541 hold364/X VGND VGND VPWR VPWR _5415_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2297 _7037_/Q VGND VGND VPWR VPWR hold751/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1552 hold371/X VGND VGND VPWR VPWR _5496_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1563 _5271_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5430__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1574 hold385/X VGND VGND VPWR VPWR _5361_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1585 _6473_/Q VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3681__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1596 _6892_/Q VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6080__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4046__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3433__A2 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6135__A1 _7065_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5340__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3672__A2 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5949__A1 _6608_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6071__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3960_ _6457_/Q _3960_/B VGND VGND VPWR VPWR _3961_/A sky130_fd_sc_hd__nand2b_2
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3891_ _4649_/C _4649_/D VGND VGND VPWR VPWR _4720_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5630_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6017_/B sky130_fd_sc_hd__and2_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5561_ _5561_/A0 _5561_/A1 _5568_/S VGND VGND VPWR VPWR _5561_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2361_A _7054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4512_ _4719_/A _4638_/B VGND VGND VPWR VPWR _4729_/A sky130_fd_sc_hd__nand2_8
X_5492_ _5492_/A0 _5582_/A1 _5496_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold104 hold104/A VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 hold115/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7231_ _7231_/A VGND VGND VPWR VPWR _7231_/X sky130_fd_sc_hd__clkbuf_2
Xhold126 hold126/A VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4443_ _4486_/A _4485_/B _4598_/B VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__nand3_4
Xhold137 hold137/A VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold148 hold148/A VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold159 hold159/A VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5885__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4374_ _4370_/Y _5011_/A _6686_/Q VGND VGND VPWR VPWR _4374_/Y sky130_fd_sc_hd__o21ai_2
X_7162_ _7185_/CLK _7162_/D fanout443/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6113_/A _6113_/B _6113_/C _6113_/D VGND VGND VPWR VPWR _6114_/D sky130_fd_sc_hd__nor4_1
X_3325_ _3726_/A hold30/X VGND VGND VPWR VPWR _3325_/Y sky130_fd_sc_hd__nor2_8
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/CLK _7093_/D fanout450/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6910_/Q _5991_/X _5993_/X _7006_/Q _6043_/X VGND VGND VPWR VPWR _6044_/X
+ sky130_fd_sc_hd__a221o_1
X_3256_ hold52/X _6657_/Q hold26/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__a21o_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4655__A _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3187_ _3187_/A VGND VGND VPWR VPWR _3187_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3663__A2 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4860__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout444_A fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6946_ _7052_/CLK _6946_/D fanout464/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3415__A2 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6877_ _6977_/CLK _6877_/D fanout461/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfstp_4
X_5828_ _6995_/Q _5929_/B _5681_/X _7091_/Q _5827_/X VGND VGND VPWR VPWR _5835_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5759_ _6888_/Q _5688_/X _5756_/X _5758_/X VGND VGND VPWR VPWR _5760_/C sky130_fd_sc_hd__a211o_1
XFILLER_148_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5876__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _5531_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold671 hold671/A VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold682 hold682/A VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold693 hold693/A VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input144_A wb_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2050 _5309_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2061 _7108_/Q VGND VGND VPWR VPWR hold374/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2072 _5379_/X VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2083 hold757/X VGND VGND VPWR VPWR _4266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2094 _6531_/Q VGND VGND VPWR VPWR hold538/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3654__A2 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1360 _6616_/Q VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1371 hold359/X VGND VGND VPWR VPWR _5439_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1382 _5391_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _4125_/X VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6053__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5800__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6108__B2 _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3590__A1 _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput209 _3234_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XANTENNA__3590__B2 _6811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5867__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4090_ _3422_/Y hold985/A _4091_/S VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6166__S _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4475__A _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4842__A1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2207_A _6845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4194__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6044__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6800_ _6803_/CLK _6800_/D fanout442/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4992_ _4701_/B _4995_/B _4991_/X _5083_/B _5021_/B VGND VGND VPWR VPWR _5000_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6731_ _6731_/CLK _6731_/D _6411_/A VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3943_ _6661_/Q _6781_/Q _6433_/B VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6662_ _6832_/CLK _6662_/D fanout447/X VGND VGND VPWR VPWR _7207_/A sky130_fd_sc_hd__dfrtp_1
X_3874_ hold93/A hold37/A _3878_/S VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5613_ _7148_/Q _5613_/B VGND VGND VPWR VPWR _5613_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6593_ _6817_/CLK _6593_/D fanout436/X VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5544_ hold201/X _5580_/A1 _5550_/S VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3581__A1 _6848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5475_ _5475_/A0 _5583_/A1 _5478_/S VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7214_ _7214_/A VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__clkbuf_2
X_4426_ _4513_/B _5150_/A VGND VGND VPWR VPWR _4426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout403 hold1426/X VGND VGND VPWR VPWR hold1427/A sky130_fd_sc_hd__buf_6
Xfanout414 _6659_/Q VGND VGND VPWR VPWR _3998_/S sky130_fd_sc_hd__buf_12
X_7145_ _7180_/CLK _7145_/D fanout448/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4357_ _4649_/B _4357_/B VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__xor2_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout436 _3959_/B VGND VGND VPWR VPWR fanout436/X sky130_fd_sc_hd__buf_12
XANTENNA_fanout394_A _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout447 fanout448/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__buf_12
XFILLER_100_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3308_ hold87/X hold78/X VGND VGND VPWR VPWR _3430_/B sky130_fd_sc_hd__and2b_4
Xfanout458 _6411_/A VGND VGND VPWR VPWR _6399_/A sky130_fd_sc_hd__clkbuf_16
Xfanout469 fanout470/X VGND VGND VPWR VPWR fanout469/X sky130_fd_sc_hd__buf_12
X_4288_ _4288_/A0 _5193_/A1 _4291_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
X_7076_ _7108_/CLK hold80/X fanout451/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6283__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4385__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3239_ _6840_/Q VGND VGND VPWR VPWR _3239_/Y sky130_fd_sc_hd__clkinv_4
X_6027_ _6901_/Q _5985_/X _6016_/X _7037_/Q VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4833__A1 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1307_A _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6035__B1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6977_/CLK _6929_/D fanout460/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7112_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6767__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6967_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold490 hold490/A VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6274__B1 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 hold1190/A VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6026__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3590_ _7096_/Q hold31/A hold24/A _6811_/Q _3589_/X VGND VGND VPWR VPWR _3595_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4760__B1 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5260_ _5260_/A0 _5584_/A1 _5262_/S VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4211_ _4211_/A0 _5448_/A1 _4211_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _5207_/A _5220_/B _5220_/C VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__and3_4
XFILLER_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2808 hold962/X VGND VGND VPWR VPWR _5332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2819 _6858_/Q VGND VGND VPWR VPWR hold945/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4142_ _4142_/A0 _5193_/A1 _4145_/S VGND VGND VPWR VPWR _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4073_ _4073_/A0 _5193_/A1 _4076_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4815__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4815__B2 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _4564_/B _4934_/B _4881_/B _4572_/Y _4886_/A VGND VGND VPWR VPWR _4976_/B
+ sky130_fd_sc_hd__a311o_2
XANTENNA__5240__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6714_ _6714_/CLK _6714_/D _6399_/A VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3926_ _6437_/Q _6654_/Q _3904_/A _3199_/A VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5791__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6645_ _6826_/CLK _6645_/D _6407_/A VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_4
X_3857_ _6654_/Q _3857_/B VGND VGND VPWR VPWR _3858_/S sky130_fd_sc_hd__nand2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6576_ _6745_/CLK _6576_/D fanout440/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfstp_2
X_3788_ _7037_/Q _3325_/Y _4065_/A _6525_/Q VGND VGND VPWR VPWR _3788_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ _5527_/A0 _5527_/A1 _5532_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5458_ _5458_/A0 _5584_/A1 _5460_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4503__B1 _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4409_ _4574_/A _4637_/D VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__nor2_8
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5389_ _5389_/A _5578_/B VGND VGND VPWR VPWR _5397_/S sky130_fd_sc_hd__and2_4
X_7128_ _7128_/CLK _7128_/D fanout469/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6256__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7059_ _7131_/CLK _7059_/D fanout453/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3609__A2 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6948__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3490__B1 _3389_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A wb_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5231__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4054__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A mgmt_gpio_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4742__B1 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3545__B2 _6588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5298__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6247__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4229__S _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4760_ _4759_/X _4558_/X _5139_/A _4760_/B2 VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ _6846_/Q _5254_/A _5461_/A _7030_/Q _3710_/X VGND VGND VPWR VPWR _3716_/B
+ sky130_fd_sc_hd__a221o_1
X_4691_ _4713_/A _4691_/B VGND VGND VPWR VPWR _4691_/Y sky130_fd_sc_hd__nand2_8
XFILLER_146_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6430_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
X_3642_ _6724_/Q _4292_/A _3539_/Y _6532_/Q _3641_/X VGND VGND VPWR VPWR _3645_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6399__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6361_ _6686_/Q _6361_/A2 _6361_/B1 _6685_/Q VGND VGND VPWR VPWR _6361_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3573_ _6920_/Q _5335_/A _4274_/A _6710_/Q _3572_/X VGND VGND VPWR VPWR _3573_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5312_ _5312_/A0 _5537_/A1 _5316_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
X_6292_ _6292_/A1 _6342_/S _6290_/X _6291_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
XANTENNA__5289__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5243_ _5243_/A0 wire371/X _5244_/S VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5523__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2605 _4257_/X VGND VGND VPWR VPWR hold693/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2616 hold931/X VGND VGND VPWR VPWR _4139_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2627 hold552/X VGND VGND VPWR VPWR _4124_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5174_ _5174_/A0 _5277_/A1 _5174_/S VGND VGND VPWR VPWR _5174_/X sky130_fd_sc_hd__mux2_1
Xhold2638 _7066_/Q VGND VGND VPWR VPWR hold963/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1904 hold933/X VGND VGND VPWR VPWR _4015_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2649 _5198_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1915 _5555_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1926 hold939/X VGND VGND VPWR VPWR _5218_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4125_ hold193/X _5527_/A1 _4127_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1937 hold694/X VGND VGND VPWR VPWR _4177_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1948 _6944_/Q VGND VGND VPWR VPWR hold831/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1959 hold851/X VGND VGND VPWR VPWR _5519_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4056_ _6423_/B _5317_/B _4056_/C VGND VGND VPWR VPWR _4064_/S sky130_fd_sc_hd__and3b_4
XANTENNA__3978__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6354__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5749__C1 _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5213__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4958_ _5044_/A _5044_/B _5032_/B _4958_/D VGND VGND VPWR VPWR _4961_/B sky130_fd_sc_hd__and4_1
XANTENNA__5764__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3775__A1 _6877_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3909_ _6019_/A _6015_/B _6008_/A VGND VGND VPWR VPWR _3909_/X sky130_fd_sc_hd__and3_1
XANTENNA__3775__B2 _6820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4889_ _5138_/A _4889_/B VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__and2_1
XFILLER_192_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6628_ _6830_/CLK _6628_/D _6433_/A VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3527__A1 input16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _7191_/CLK _6559_/D VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5433__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6229__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4049__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6711__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4292__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5204__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3766__A1 _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3518__A1 _6865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3518__B2 _6483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7167__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output276_A _6477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6180__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4191__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5343__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _6577_/Q _5667_/X _5682_/X _6453_/Q VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3454__B1 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ _6687_/Q _5659_/X _5684_/X _6604_/Q VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__a22o_1
X_4812_ _4812_/A _4826_/A VGND VGND VPWR VPWR _4812_/Y sky130_fd_sc_hd__nor2_2
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5792_ _5792_/A _5792_/B _5792_/C _5792_/D VGND VGND VPWR VPWR _5792_/Y sky130_fd_sc_hd__nor4_4
XANTENNA__5746__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _4719_/A _4719_/B _4741_/Y _4742_/Y VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_175_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5518__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4674_ _4682_/A _4691_/B VGND VGND VPWR VPWR _4674_/Y sky130_fd_sc_hd__nand2_4
XFILLER_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6413_ _6413_/A _6423_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
X_3625_ input26/X _3307_/Y _4286_/A _6719_/Q VGND VGND VPWR VPWR _3625_/X sky130_fd_sc_hd__a22o_4
XANTENNA__6171__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6344_ _6344_/A VGND VGND VPWR VPWR _6344_/Y sky130_fd_sc_hd__inv_2
X_3556_ _3556_/A _3556_/B _3556_/C _3556_/D VGND VGND VPWR VPWR _3557_/D sky130_fd_sc_hd__nor4_2
XFILLER_143_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6349__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6275_ _6714_/Q _5973_/X _5988_/X _6571_/Q VGND VGND VPWR VPWR _6275_/X sky130_fd_sc_hd__a22o_1
X_3487_ _3550_/A _3648_/A VGND VGND VPWR VPWR _4274_/A sky130_fd_sc_hd__nor2_8
Xhold2402 _7106_/Q VGND VGND VPWR VPWR hold626/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4343_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5226_ _5226_/A _5226_/B _5569_/B VGND VGND VPWR VPWR _5228_/S sky130_fd_sc_hd__and3_1
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2413 _6604_/Q VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2424 _4205_/X VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2435 _6741_/Q VGND VGND VPWR VPWR hold855/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1701 _4029_/X VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2446 _6946_/Q VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2457 _5431_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1712 _6545_/Q VGND VGND VPWR VPWR hold987/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6684__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2468 hold878/X VGND VGND VPWR VPWR _4076_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5157_ _4570_/C _4523_/Y _4870_/A _4925_/A _5113_/B VGND VGND VPWR VPWR _5157_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold1723 hold422/X VGND VGND VPWR VPWR hold1723/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3693__B1 _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1734 _6547_/Q VGND VGND VPWR VPWR hold988/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout474_A _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2479 _6454_/Q VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_186_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1745 hold424/X VGND VGND VPWR VPWR hold1745/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4108_ _3803_/Y hold991/A _4115_/S VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__mux2_1
Xhold1756 hold442/X VGND VGND VPWR VPWR hold1756/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1767 hold990/X VGND VGND VPWR VPWR hold476/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5088_ _4477_/Y _4938_/X _5027_/X _5087_/X _4791_/B VGND VGND VPWR VPWR _5088_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold1778 _6541_/Q VGND VGND VPWR VPWR hold986/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1789 _5576_/X VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4039_ _4061_/A0 _5529_/A1 _4056_/C VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3445__B1 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3748__A1 _7133_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3748__B2 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5428__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 hold238/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6162__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4173__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5122__B1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input35_A mask_rev_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2980 _6973_/Q VGND VGND VPWR VPWR hold413/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3436__B1 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3987__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5338__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6153__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold319 hold319/A VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3410_ input32/X _3307_/Y _5461_/A _7035_/Q VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4390_ _4717_/A _4712_/A VGND VGND VPWR VPWR _4658_/A sky130_fd_sc_hd__nand2_8
XANTENNA__5900__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3341_ _3550_/A _3686_/A VGND VGND VPWR VPWR _5362_/A sky130_fd_sc_hd__nor2_8
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4478__A _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _7094_/Q _5984_/X _5986_/X _7030_/Q VGND VGND VPWR VPWR _6060_/X sky130_fd_sc_hd__a22o_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold87/A hold78/X VGND VGND VPWR VPWR _3272_/Y sky130_fd_sc_hd__nor2_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6754__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5011_ _5011_/A _5011_/B VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__and2_1
Xhold1008 _6822_/Q VGND VGND VPWR VPWR _5228_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 hold2/X VGND VGND VPWR VPWR _5536_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6962_ _7099_/CLK _6962_/D fanout471/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5967__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5913_ _6611_/Q _5660_/X _5669_/X _6651_/Q _5912_/X VGND VGND VPWR VPWR _5913_/X
+ sky130_fd_sc_hd__a221o_1
X_6893_ _6977_/CLK _6893_/D fanout461/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5844_ _7036_/Q _5655_/X _5656_/X _6988_/Q _5839_/Y VGND VGND VPWR VPWR _5844_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5719__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5775_ _6913_/Q _5670_/X _5671_/X _7065_/Q _5774_/X VGND VGND VPWR VPWR _5782_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4726_ _4726_/A _4726_/B _4738_/B VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__nand3_2
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4657_ _4500_/Y _4640_/Y _5047_/A VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6144__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4155__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_2
Xhold820 hold820/A VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3608_ _6992_/Q _5416_/A _3310_/Y input14/X _3607_/X VGND VGND VPWR VPWR _3614_/B
+ sky130_fd_sc_hd__a221o_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
X_4588_ _4596_/A _4972_/A VGND VGND VPWR VPWR _4986_/C sky130_fd_sc_hd__nand2_4
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold842 hold842/A VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold853 hold853/A VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold864 _5210_/X VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A _6327_/B _6327_/C VGND VGND VPWR VPWR _6339_/C sky130_fd_sc_hd__nor3_4
Xmgmt_gpio_15_buff_inst _3949_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold875 hold875/A VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3539_ _3549_/B _3648_/B VGND VGND VPWR VPWR _3539_/Y sky130_fd_sc_hd__nor2_4
Xhold886 hold886/A VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold897 _5381_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6258_ _6713_/Q _5973_/X _5988_/X _6570_/Q _6257_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2210 hold828/X VGND VGND VPWR VPWR _4096_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2221 hold608/X VGND VGND VPWR VPWR _5413_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2232 hold593/X VGND VGND VPWR VPWR _5467_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2243 _6629_/Q VGND VGND VPWR VPWR hold770/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5209_ _5209_/A0 _5237_/A1 _5209_/S VGND VGND VPWR VPWR _5209_/X sky130_fd_sc_hd__mux2_1
X_6189_ _6170_/X _6189_/B _6189_/C VGND VGND VPWR VPWR _6189_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__3666__B1 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2254 _5283_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1520 hold343/X VGND VGND VPWR VPWR _5370_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2265 hold701/X VGND VGND VPWR VPWR _4275_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2276 hold417/X VGND VGND VPWR VPWR _5505_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1531 _6972_/Q VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2287 hold408/X VGND VGND VPWR VPWR _5541_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1542 _5415_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1553 _5496_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2298 _6597_/Q VGND VGND VPWR VPWR hold891/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1564 _6875_/Q VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 _5361_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1586 hold520/X VGND VGND VPWR VPWR _3991_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1597 hold370/X VGND VGND VPWR VPWR _5307_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3418__B1 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5958__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6080__B2 _7039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4091__A0 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4851__A _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4062__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6135__A2 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4298__A hold64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3657__B1 _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output239_A _3938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4237__S _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3409__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5949__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3890_ _4720_/C _4649_/B VGND VGND VPWR VPWR _3890_/Y sky130_fd_sc_hd__nand2_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A hold9/A VGND VGND VPWR VPWR _5568_/S sky130_fd_sc_hd__and2_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4511_ _4719_/A _4638_/B VGND VGND VPWR VPWR _4955_/D sky130_fd_sc_hd__and2_4
XFILLER_8_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5491_ _5491_/A0 _5581_/A1 _5496_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6126__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7230_ _7230_/A VGND VGND VPWR VPWR _7230_/X sky130_fd_sc_hd__clkbuf_2
Xhold105 hold105/A VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4137__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4442_ _4486_/A _4485_/B _4598_/B VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__and3_2
Xhold116 _4270_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold127 hold127/A VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold138 hold138/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold149 hold149/A VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7161_ _7185_/CLK _7161_/D fanout443/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_1
X_4373_ _4576_/A _4719_/A VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__nand2_8
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6774__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6112_ _7136_/Q _5977_/X _5984_/X _7096_/Q _6111_/X VGND VGND VPWR VPWR _6113_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3360__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3324_ _3764_/A _3535_/A VGND VGND VPWR VPWR _5515_/A sky130_fd_sc_hd__nor2_8
XFILLER_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7108_/CLK _7092_/D fanout451/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _7086_/Q _5638_/X _6012_/X _6998_/Q VGND VGND VPWR VPWR _6043_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3998_/S _3255_/B VGND VGND VPWR VPWR _3255_/Y sky130_fd_sc_hd__nand2b_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5531__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3186_ _6657_/Q VGND VGND VPWR VPWR _3862_/A sky130_fd_sc_hd__inv_2
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4860__A2 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK _6945_/D fanout461/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3986__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6876_ _6963_/CLK _6876_/D fanout463/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout437_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5827_ _6859_/Q _5651_/X _5688_/X _6891_/Q VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5758_ _7032_/Q _5655_/X _5667_/X _6880_/Q _5757_/X VGND VGND VPWR VPWR _5758_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4709_ _4495_/B _4638_/B _4507_/Y _4704_/X _4708_/X VGND VGND VPWR VPWR _4709_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_136_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5689_ _5689_/A _5689_/B _5689_/C VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__and3_4
XFILLER_135_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold650 hold650/A VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold661 hold661/A VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3887__B1 _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold672 hold672/A VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold683 hold683/A VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold694 hold694/A VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2040 hold718/X VGND VGND VPWR VPWR _4057_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__B1 _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2051 _6472_/Q VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5441__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2062 hold374/X VGND VGND VPWR VPWR _5550_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4300__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2073 _6602_/Q VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input137_A wb_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2084 _4266_/X VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4565__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2095 hold538/X VGND VGND VPWR VPWR _4073_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1350 _6581_/Q VGND VGND VPWR VPWR hold170/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 _6621_/Q VGND VGND VPWR VPWR hold166/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1372 _5439_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1383 _7126_/Q VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1394 _6807_/Q VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6053__A1 _7118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3575__C1 _3574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6108__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4119__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3590__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5867__B2 _6707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3878__A0 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5351__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4842__A2 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4668_/Y _4688_/A _4995_/B VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6730_ _6730_/CLK _6730_/D _6411_/A VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfrtp_4
X_3942_ _6666_/Q input77/X _3970_/B VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _6830_/CLK _6661_/D fanout454/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_1
X_3873_ hold37/A hold33/A _3878_/S VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5612_ _5647_/B _5679_/B _5684_/B _5612_/B1 _5605_/Y VGND VGND VPWR VPWR _7147_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6592_ _6817_/CLK _6592_/D fanout436/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5543_ _5543_/A0 _5543_/A1 _5550_/S VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5526__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3581__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5474_ _5474_/A0 _5582_/A1 _5478_/S VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7213_ _7213_/A VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__clkbuf_2
X_4425_ _4513_/B _5150_/A VGND VGND VPWR VPWR _4552_/B sky130_fd_sc_hd__and2_1
XFILLER_133_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7144_ _7179_/CLK _7144_/D fanout448/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout404 _5533_/B VGND VGND VPWR VPWR _5220_/C sky130_fd_sc_hd__buf_8
XANTENNA__4530__A1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4356_ _4492_/B _4356_/B VGND VGND VPWR VPWR _4357_/B sky130_fd_sc_hd__nand2_2
XFILLER_101_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout437 fanout454/X VGND VGND VPWR VPWR _3959_/B sky130_fd_sc_hd__buf_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout448 fanout449/X VGND VGND VPWR VPWR fanout448/X sky130_fd_sc_hd__clkbuf_16
X_3307_ _3764_/B _3553_/B VGND VGND VPWR VPWR _3307_/Y sky130_fd_sc_hd__nor2_8
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7075_ _7131_/CLK _7075_/D fanout453/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout459 input75/X VGND VGND VPWR VPWR _6411_/A sky130_fd_sc_hd__buf_12
XFILLER_101_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4287_ _4287_/A0 _5237_/A1 _4291_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6026_ _6997_/Q _6012_/X _6019_/X _6981_/Q _6025_/X VGND VGND VPWR VPWR _6026_/X
+ sky130_fd_sc_hd__a221o_1
X_3238_ _6848_/Q VGND VGND VPWR VPWR _3238_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4385__B _4751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6035__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5497__A _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6928_ _6936_/CLK _6928_/D fanout463/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6859_ _7131_/CLK _6859_/D fanout452/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5436__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1836_A _6503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3572__A2 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5849__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold480 hold480/A VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold491 hold491/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_2_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _7031_/Q VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1191 _4248_/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6026__A1 _6997_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6026__B2 _6981_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__A _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__C1 _3795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6329__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5346__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4210_ _4210_/A0 _5233_/A1 _4211_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
X_5190_ _5190_/A0 wire375/X _5190_/S VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__mux2_1
Xhold2809 _7083_/Q VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4141_ _4141_/A0 _5237_/A1 _4145_/S VGND VGND VPWR VPWR _4141_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6265__A1 _6526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4072_ _4072_/A0 _5237_/A1 _4076_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4815__A2 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4974_ _5114_/A _4986_/C _5114_/B VGND VGND VPWR VPWR _5061_/B sky130_fd_sc_hd__and3_1
XANTENNA__5776__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6713_ _7121_/CLK _6713_/D _6399_/A VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3925_ _6341_/S _3912_/B _5647_/B VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__o21ai_1
XFILLER_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6644_ _6830_/CLK _6644_/D _6433_/A VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_4
X_3856_ _3807_/B _3904_/A _3855_/X _3856_/B2 _3903_/A VGND VGND VPWR VPWR _6455_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6575_ _6745_/CLK _6575_/D fanout440/X VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfrtp_4
X_3787_ _6965_/Q _5389_/A _5308_/A _6893_/Q _3786_/X VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a221o_1
X_5526_ _5526_/A0 _5562_/A1 _5532_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3554__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5457_ _5457_/A0 _5583_/A1 _5460_/S VGND VGND VPWR VPWR _5457_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4408_ _4391_/Y _4969_/A _4407_/Y VGND VGND VPWR VPWR _4529_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5700__B1 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5388_ _5388_/A0 _5568_/A1 _5388_/S VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7127_ _7133_/CLK _7127_/D fanout468/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3711__C1 _3710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4339_ _4339_/A0 _5448_/A1 _4339_/S VGND VGND VPWR VPWR _4339_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1417_A _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7058_ _7130_/CLK _7058_/D fanout462/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6009_ _5637_/A _6017_/A _6019_/C _5980_/X _5995_/X VGND VGND VPWR VPWR _6010_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5767__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3793__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4742__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3545__A2 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input65_A mgmt_gpio_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6247__A1 _6605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6247__B2 _6728_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__B1 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3710_ _6472_/Q _3988_/A _3977_/A _6451_/Q VGND VGND VPWR VPWR _3710_/X sky130_fd_sc_hd__a22o_2
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3784__A2 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4690_ _4638_/Y _4668_/Y _4688_/X _4990_/B _4689_/Y VGND VGND VPWR VPWR _4703_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3641_ input54/X _4241_/A _3509_/Y _6729_/Q VGND VGND VPWR VPWR _3641_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6183__B1 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6360_ _6684_/Q _6358_/Y _6359_/X _6355_/Y VGND VGND VPWR VPWR _6384_/S sky130_fd_sc_hd__a211o_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5930__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3572_ _6912_/Q _5326_/A _3569_/X _3571_/X VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__a211o_1
X_5311_ _5311_/A0 _5572_/A1 _5316_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6291_ _6490_/Q _6291_/A2 _5649_/Y VGND VGND VPWR VPWR _6291_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5242_ _5242_/A0 wire375/X _5244_/S VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7128_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2606 _6693_/Q VGND VGND VPWR VPWR hold547/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2617 _4139_/X VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5173_ _5173_/A0 _5195_/A1 _5174_/S VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__mux2_1
Xhold2628 _4124_/X VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2639 hold963/X VGND VGND VPWR VPWR _5503_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1905 _4015_/X VGND VGND VPWR VPWR hold934/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1916 _7104_/Q VGND VGND VPWR VPWR hold768/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4124_ _4124_/A0 _5238_/A1 _4127_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1927 _5218_/X VGND VGND VPWR VPWR _5219_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1938 _4177_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1949 hold831/X VGND VGND VPWR VPWR _5366_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_2
X_4055_ _4055_/A0 hold71/X _4055_/S VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7082_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3472__A1 _6985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3472__B2 _6726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ _5067_/A _5023_/A _4957_/C _5034_/C VGND VGND VPWR VPWR _4958_/D sky130_fd_sc_hd__and4_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3994__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6641__SET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3908_ _5637_/A _7156_/Q VGND VGND VPWR VPWR _6008_/A sky130_fd_sc_hd__and2_2
XANTENNA__3775__A2 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4888_ _4574_/A _4463_/B _4568_/Y _4878_/Y _4491_/Y VGND VGND VPWR VPWR _4892_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_177_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6627_ _6760_/CLK _6627_/D fanout441/X VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6174__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3839_ _6460_/Q _6657_/Q _3835_/S _3839_/C1 VGND VGND VPWR VPWR _3841_/A sky130_fd_sc_hd__o211a_1
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3527__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5921__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6558_ _7191_/CLK _6558_/D VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ _5509_/A0 _5527_/A1 _5514_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6489_ _7180_/CLK _6489_/D fanout446/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_133_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1534_A _6486_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4573__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3463__A1 _3462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3766__A2 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3518__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5912__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output269_A _6790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5691__A2 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3454__B2 _6842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ _5860_/A1 _6167_/S _5858_/X _5859_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__o22a_1
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4811_ _4679_/Y _4811_/B VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__nand2b_1
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _6849_/Q _5653_/X _5674_/X _6873_/Q _5790_/X VGND VGND VPWR VPWR _5792_/D
+ sky130_fd_sc_hd__a221o_2
X_4742_ _5011_/A _4947_/A _4713_/Y VGND VGND VPWR VPWR _4742_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3757__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4673_ _4682_/A _4714_/B _4712_/C VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__and3_4
XFILLER_174_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6156__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2551_A _6701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6412_ _6413_/A _6423_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
X_3624_ _7135_/Q _3295_/Y _5434_/A _7007_/Q _3623_/X VGND VGND VPWR VPWR _3627_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6343_ _6676_/Q _6677_/Q _6680_/Q _6683_/Q _3922_/B VGND VGND VPWR VPWR _6344_/A
+ sky130_fd_sc_hd__o41a_1
X_3555_ _7113_/Q _5551_/A _3336_/Y input24/X _3554_/X VGND VGND VPWR VPWR _3556_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5534__S _5540_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6274_ _6704_/Q _5977_/X _5990_/X _6646_/Q _6273_/X VGND VGND VPWR VPWR _6279_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3486_ _3764_/B _3516_/B VGND VGND VPWR VPWR _3486_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5225_ _5225_/A0 _5579_/A1 hold10/X VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2403 hold626/X VGND VGND VPWR VPWR _5548_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2414 hold869/X VGND VGND VPWR VPWR _4159_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2425 _6633_/Q VGND VGND VPWR VPWR hold858/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2436 hold855/X VGND VGND VPWR VPWR _4315_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1702 _6521_/Q VGND VGND VPWR VPWR hold351/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5156_/Y sky130_fd_sc_hd__nand3_1
Xhold2447 hold635/X VGND VGND VPWR VPWR _5368_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2458 _6820_/Q VGND VGND VPWR VPWR hold872/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1713 hold987/X VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2469 _4076_/X VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3693__A1 _7102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1724 _6553_/Q VGND VGND VPWR VPWR hold970/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1735 hold988/X VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1746 _6786_/Q VGND VGND VPWR VPWR hold627/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4107_ _6679_/Q _4107_/B VGND VGND VPWR VPWR _4115_/S sky130_fd_sc_hd__nand2_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1757 _6696_/Q VGND VGND VPWR VPWR hold393/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5087_ _4417_/B _4668_/Y _4777_/X _5117_/B _5117_/A VGND VGND VPWR VPWR _5087_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold1768 hold476/X VGND VGND VPWR VPWR hold1768/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1779 hold986/X VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4038_ _4038_/A0 _4037_/X _4046_/S VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6509__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5198__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _6015_/B _6014_/A _6007_/C VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__and3_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1484_A _7004_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3748__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_50 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_61 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_83 _5377_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1749_A _6719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5370__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5444__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1916_A _7104_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3381__B1 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input167_A wb_sel_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput190 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_95_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5122__B2 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2970 _7144_/Q VGND VGND VPWR VPWR _5600_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input28_A mask_rev_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2981 _6537_/Q VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3436__B2 _7233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5189__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 hold309/A VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5361__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4759__A _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5354__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3340_ _3550_/A _3563_/B VGND VGND VPWR VPWR _5389_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3271_ _3270_/X hold77/X _3998_/S VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_86_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5010_/B VGND VGND VPWR VPWR _5083_/C sky130_fd_sc_hd__and2_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 _6440_/Q VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6961_ _7001_/CLK _6961_/D fanout466/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6673__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5912_ _6571_/Q _5674_/X _5680_/X _6709_/Q VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__a22o_1
X_6892_ _7108_/CLK _6892_/D fanout451/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5843_ _6916_/Q _5670_/X _5685_/X _7076_/Q _5842_/X VGND VGND VPWR VPWR _5843_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5529__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4927__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5774_ _6953_/Q _5672_/X _5682_/X _7041_/Q VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4725_ _5026_/B _4725_/B VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__nand2_2
XFILLER_175_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4656_ _4652_/Y _4656_/B VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__nand2b_1
XFILLER_163_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3607_ _6740_/Q _4310_/A _3539_/Y _6533_/Q VGND VGND VPWR VPWR _3607_/X sky130_fd_sc_hd__a22o_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3973_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold810 _5385_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5352__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold821 hold821/A VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4587_ _4621_/A _4693_/B VGND VGND VPWR VPWR _4901_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__buf_2
Xhold832 hold832/A VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5264__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold843 hold843/A VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3363__B1 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold854 hold854/A VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6326_ _6643_/Q _5986_/X _5998_/X _6583_/Q _6325_/X VGND VGND VPWR VPWR _6327_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3538_ _6937_/Q _5353_/A _4170_/A _6618_/Q _3537_/X VGND VGND VPWR VPWR _3543_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4388__B _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold865 hold865/A VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold876 hold876/A VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold887 hold887/A VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold898 hold898/A VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6257_ _6708_/Q _5992_/X _6012_/X _6748_/Q _6256_/X VGND VGND VPWR VPWR _6257_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2200 hold565/X VGND VGND VPWR VPWR _5454_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6301__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3469_ _3563_/A _3516_/B VGND VGND VPWR VPWR _4292_/A sky130_fd_sc_hd__nor2_4
Xhold2211 _4096_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2222 _5413_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5208_ _5208_/A0 _5543_/A1 _5208_/S VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2233 _5467_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2244 hold770/X VGND VGND VPWR VPWR _4189_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6188_ _6181_/X _6183_/X _6188_/C _6339_/B VGND VGND VPWR VPWR _6189_/C sky130_fd_sc_hd__and4bb_1
Xhold1510 _5277_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2255 _6647_/Q VGND VGND VPWR VPWR hold801/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3666__A1 _7127_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1521 _5370_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2266 _4275_/X VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5139_ _5139_/A _5139_/B _5139_/C VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__and3_1
Xhold2277 _5505_/X VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1532 hold325/X VGND VGND VPWR VPWR _5397_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1543 _7036_/Q VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2288 _7017_/Q VGND VGND VPWR VPWR hold727/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1554 _6452_/Q VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2299 hold891/X VGND VGND VPWR VPWR _4150_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6065__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1565 hold291/X VGND VGND VPWR VPWR _5288_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1576 _7011_/Q VGND VGND VPWR VPWR hold318/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1587 _3991_/X VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1598 _5307_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7157__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6080__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5439__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5343__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4579__A _4751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5894__A2 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4298__B _5184_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4854__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3409__B2 _7011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6071__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output301_A _3745_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4082__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5349__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4909__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5582__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4510_/A _4510_/B VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3593__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5490_ hold598/X _5562_/A1 _5496_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold106 hold106/A VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4441_ _4457_/A _4457_/C _4469_/B VGND VGND VPWR VPWR _4598_/B sky130_fd_sc_hd__a21boi_4
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5334__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold139 hold139/A VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2347_A _6712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5885__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7160_ _7184_/CLK _7160_/D fanout445/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4372_ _4576_/A _4719_/A VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__and2_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6928_/Q _5982_/X _5987_/X _7112_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3323_ _3346_/A _3563_/B VGND VGND VPWR VPWR _5317_/A sky130_fd_sc_hd__nor2_8
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7091_/CLK _7091_/D fanout452/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6066_/A2 _5649_/Y _6041_/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__a21o_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3254_ hold26/X _6657_/Q hold1131/X VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__a21bo_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _6864_/Q VGND VGND VPWR VPWR _3185_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4860__A3 _4683_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6062__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6944_ _7106_/CLK _6944_/D fanout472/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4073__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4671__B _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6875_ _6963_/CLK _6875_/D fanout464/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ _5826_/A _5826_/B _5826_/C VGND VGND VPWR VPWR _5826_/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5573__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ _6856_/Q _5651_/X _5679_/X _6904_/Q VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3584__B1 _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4708_ _4370_/Y _4411_/Y _5067_/A _4707_/X VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__o211a_1
XFILLER_163_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5688_ _5689_/A _5689_/B _5688_/C VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3b_4
XANTENNA__5325__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4639_ _4650_/B _4394_/A _4639_/S VGND VGND VPWR VPWR _4640_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1447_A _6959_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5876__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 hold640/A VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 _5513_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold662 _5549_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold673 hold673/A VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6309_ _6627_/Q _6013_/X _6015_/X _6760_/Q VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold684 hold684/A VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold695 hold695/A VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2030 _4190_/X VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3639__B2 _6631_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2041 _6538_/Q VGND VGND VPWR VPWR hold807/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2052 hold516/X VGND VGND VPWR VPWR _3990_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2063 _6518_/Q VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2074 hold712/X VGND VGND VPWR VPWR _4156_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2085 _6632_/Q VGND VGND VPWR VPWR hold745/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1340 _6694_/Q VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2096 _4073_/X VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1351 _4131_/X VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1362 _4179_/X VGND VGND VPWR VPWR hold167/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1373 _6511_/Q VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1384 hold245/X VGND VGND VPWR VPWR _5571_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 hold412/X VGND VGND VPWR VPWR _5206_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1983_A _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6053__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4064__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5677__B _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5800__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input95_A usr1_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5564__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6780__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5316__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5867__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6044__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4055__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4990_ _5150_/B _4990_/B VGND VGND VPWR VPWR _4990_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_91_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3941_ _6501_/Q _3881_/C _6459_/Q VGND VGND VPWR VPWR _3941_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2297_A _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3872_ hold33/A hold69/A _3878_/S VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__mux2_1
X_6660_ _6835_/CLK _6660_/D _3959_/B VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5004__B1 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5611_ _5611_/A _5647_/B VGND VGND VPWR VPWR _5611_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__5555__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _6817_/CLK _6591_/D fanout435/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_164_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2464_A _6985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5542_ _5542_/A _5578_/B VGND VGND VPWR VPWR _5550_/S sky130_fd_sc_hd__and2_4
XFILLER_129_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5307__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5473_ _7039_/Q _5536_/A1 _5478_/S VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4424_ _4384_/A _4658_/A _4417_/B _4522_/B _4370_/Y VGND VGND VPWR VPWR _4704_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_145_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5858__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7212_ _7212_/A VGND VGND VPWR VPWR _7212_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4355_ _4447_/B _4663_/D _4682_/A _4365_/B VGND VGND VPWR VPWR _4362_/A sky130_fd_sc_hd__nand4_2
X_7143_ _7180_/CLK _7143_/D fanout448/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4947__A _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout405 _5533_/B VGND VGND VPWR VPWR _5569_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__4530__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3306_ _3309_/A _3390_/B VGND VGND VPWR VPWR _3553_/B sky130_fd_sc_hd__nand2_8
Xfanout438 _6407_/A VGND VGND VPWR VPWR _6433_/A sky130_fd_sc_hd__buf_6
XFILLER_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7074_ _7130_/CLK _7074_/D fanout462/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
X_4286_ _4286_/A _5220_/C VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__and2_2
Xfanout449 fanout454/X VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__clkbuf_16
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6283__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6025_ _7085_/Q _5638_/X _6018_/X _6965_/Q VGND VGND VPWR VPWR _6025_/X sky130_fd_sc_hd__a22o_1
X_3237_ _6856_/Q VGND VGND VPWR VPWR _3237_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4294__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6035__A2 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5497__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6927_ _6977_/CLK _6927_/D fanout460/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6858_ _6996_/CLK _6858_/D fanout462/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5546__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5809_ _7034_/Q _5655_/X _5656_/X _6986_/Q _5797_/Y VGND VGND VPWR VPWR _5809_/X
+ sky130_fd_sc_hd__a221o_1
X_6789_ _6793_/CLK _6789_/D fanout434/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1564_A _6875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5849__A2 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold470 hold470/A VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4857__A _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold481 hold481/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7233__A _7233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold492 hold492/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4809__B1 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6274__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4285__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 hold209/X VGND VGND VPWR VPWR _5554_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input10_A mask_rev_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1181 hold220/X VGND VGND VPWR VPWR _5464_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6026__A2 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1192 hold36/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4037__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__B1 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5537__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output299_A _6806_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3548__B1 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4140_ _4140_/A _5220_/C VGND VGND VPWR VPWR _4145_/S sky130_fd_sc_hd__and2_2
XANTENNA__3720__B1 _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4917__D _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6265__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4071_ _5220_/B _5226_/B _5220_/C VGND VGND VPWR VPWR _4076_/S sky130_fd_sc_hd__and3_2
XANTENNA__5473__A0 _7039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4276__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4028__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4973_ _5136_/A _4997_/A _4973_/C VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__and3_2
X_6712_ _6714_/CLK _6712_/D _6399_/A VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3787__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3924_ _6490_/Q _5643_/A VGND VGND VPWR VPWR _3924_/Y sky130_fd_sc_hd__nand2_8
XFILLER_149_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5528__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6643_ _6794_/CLK _6643_/D _3959_/B VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_4
X_3855_ _6657_/Q _6656_/Q _6448_/Q VGND VGND VPWR VPWR _3855_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5537__S _5540_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6574_ _6745_/CLK _6574_/D fanout441/X VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfrtp_4
X_3786_ _6687_/Q _4250_/A _4158_/A _6604_/Q VGND VGND VPWR VPWR _3786_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5525_ _5525_/A0 _5534_/A1 _5532_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
X_5456_ _5456_/A0 _5582_/A1 _5460_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4407_ _4477_/A _4477_/B VGND VGND VPWR VPWR _4407_/Y sky130_fd_sc_hd__nand2_4
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5700__B2 _6997_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5387_ _5387_/A0 _5567_/A1 _5388_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3711__B1 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7126_ _7126_/CLK _7126_/D fanout450/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfstp_1
X_4338_ _4338_/A0 _5233_/A1 _4339_/S VGND VGND VPWR VPWR _4338_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input2_A debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6256__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7057_ _7137_/CLK _7057_/D fanout466/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
X_4269_ _4269_/A0 _5561_/A1 _4273_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4267__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6008_ _6008_/A _6017_/A _6019_/C VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__and3_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3490__A2 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1681_A _6794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5519__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5447__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4742__A2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input58_A mgmt_gpio_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3702__B1 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6247__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4258__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__A1 _7032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5758__B2 _6880_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5357__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _7055_/Q _5488_/A _3977_/A _6452_/Q _3639_/X VGND VGND VPWR VPWR _3645_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4414__A_N _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3571_ input38/X _3293_/Y _3509_/Y _6730_/Q _3570_/X VGND VGND VPWR VPWR _3571_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4733__A2 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5930__B2 _6453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3941__A0 _6501_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5310_ _5310_/A0 _5562_/A1 _5316_/S VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6290_ _6527_/Q _6339_/B _6289_/Y _6341_/S VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4497__A _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5241_ _5241_/A0 hold95/X _5244_/S VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__mux2_1
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5172_ hold504/X _5194_/A1 _5174_/S VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__mux2_1
Xhold2607 hold547/X VGND VGND VPWR VPWR _4258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2618 _6637_/Q VGND VGND VPWR VPWR hold778/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2629 _7035_/Q VGND VGND VPWR VPWR hold737/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1906 hold934/X VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4123_ _4123_/A0 _5543_/A1 _4127_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
Xhold1917 hold768/X VGND VGND VPWR VPWR _5546_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4249__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1928 _6923_/Q VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1939 _6955_/Q VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4054_ _4054_/A0 _5567_/A1 _4055_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4663__C _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3472__A2 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5749__A1 _6839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2963_A _7186_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ _4466_/A _4477_/Y _4934_/Y _4784_/X VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__o31a_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3907_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6015_/B sky130_fd_sc_hd__and2b_4
XFILLER_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ _4947_/B _4570_/A _4986_/C _4885_/X _5023_/A VGND VGND VPWR VPWR _4892_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5267__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout412_A _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6626_ _6761_/CLK _6626_/D _6430_/A VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfstp_2
X_3838_ _3838_/A1 _3835_/S _3837_/X VGND VGND VPWR VPWR _3838_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6557_ _7191_/CLK _6557_/D VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5921__B2 _6581_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3769_ _3769_/A _3769_/B _3769_/C _3769_/D VGND VGND VPWR VPWR _3770_/C sky130_fd_sc_hd__nor4_1
X_5508_ _5508_/A0 _5571_/A1 _5514_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6488_ _6821_/CLK _6488_/D fanout443/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5439_ _5439_/A0 _5529_/A1 _5442_/S VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4200__A _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_2__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6229__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7109_ _7134_/CLK _7109_/D fanout469/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3448__C1 _3434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input112_A wb_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6165__A1 _6842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_63_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4100__A0 _3737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4651__A1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3454__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _4583_/B _4688_/A _4688_/C _4729_/A VGND VGND VPWR VPWR _4820_/A sky130_fd_sc_hd__o22a_1
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _6977_/Q _5660_/X _5662_/X _6897_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
X_4741_ _4415_/B _4712_/Y _4740_/X VGND VGND VPWR VPWR _4741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6156__A1 _7106_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4672_ _4714_/B _4712_/C VGND VGND VPWR VPWR _4672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6156__B2 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6411_ _6411_/A _6423_/B VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__and2_1
X_3623_ _7071_/Q _5506_/A _4328_/A _6754_/Q VGND VGND VPWR VPWR _3623_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6342_ _6342_/A0 _6341_/X _6342_/S VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__mux2_1
X_3554_ _7057_/Q _5488_/A _4176_/A _6623_/Q VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3485_ _6929_/Q _5344_/A _3330_/Y input48/X _3484_/X VGND VGND VPWR VPWR _3499_/A
+ sky130_fd_sc_hd__a221o_1
X_6273_ _6596_/Q _5991_/X _5997_/X _6699_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ _5224_/A0 _5580_/A1 hold10/X VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2404 _6529_/Q VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2415 _4159_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2426 hold858/X VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2437 _4315_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1703 hold351/X VGND VGND VPWR VPWR _4061_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5155_ _5155_/A _5155_/B _5155_/C _5155_/D VGND VGND VPWR VPWR _5156_/C sky130_fd_sc_hd__and4_1
Xhold2448 _5368_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2459 hold872/X VGND VGND VPWR VPWR _5225_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5550__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1714 hold455/X VGND VGND VPWR VPWR hold1714/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3693__A2 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1725 hold970/X VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4106_ _3385_/Y hold981/A _4106_/S VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1736 hold457/X VGND VGND VPWR VPWR hold1736/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5086_ _5086_/A _5086_/B VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__nand2_1
Xhold1747 hold627/X VGND VGND VPWR VPWR _5181_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1758 hold393/X VGND VGND VPWR VPWR _4261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1769 _6566_/Q VGND VGND VPWR VPWR hold978/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4037_ _4060_/A0 _5537_/A1 _4056_/C VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3445__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1108_A _6715_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _6015_/B _6018_/B _6007_/C VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__and3_4
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4939_ _4936_/Y _4938_/X _4776_/Y VGND VGND VPWR VPWR _5117_/B sky130_fd_sc_hd__o21a_1
XANTENNA_40 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_51 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _5244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6756_/CLK _6609_/D fanout441/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_95 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1644_A _6734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3381__B2 _6964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1811_A _6797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5122__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput180 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
XFILLER_121_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput191 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5460__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2960 _7142_/Q VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2971 _7147_/Q VGND VGND VPWR VPWR _5612_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2982 _6766_/Q VGND VGND VPWR VPWR _3187_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6083__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3436__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5830__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6972__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5897__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7052_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3372__A1 _6486_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _3270_/A0 _3879_/B _6657_/Q VGND VGND VPWR VPWR _3270_/X sky130_fd_sc_hd__mux2_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B2 _6720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7073_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5370__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6074__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6960_ _7099_/CLK _6960_/D fanout472/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5821__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5911_ _6754_/Q _5681_/X _5910_/X VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6891_ _7108_/CLK _6891_/D fanout451/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5842_ _6852_/Q _5653_/X _5840_/X _5841_/X VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5773_ _5794_/A0 _5772_/X _6342_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4927__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6642__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2759_A _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4724_ _5001_/A _4724_/B _4724_/C VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__nand3_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5750__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4655_ _4655_/A _4655_/B VGND VGND VPWR VPWR _4656_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5545__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5888__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_2
X_3606_ _6840_/Q _5245_/A _4212_/A _6652_/Q _3605_/X VGND VGND VPWR VPWR _3614_/A
+ sky130_fd_sc_hd__a221o_1
Xhold800 hold800/A VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold811 hold811/A VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_2
X_4586_ _4625_/A _4628_/A VGND VGND VPWR VPWR _4586_/Y sky130_fd_sc_hd__nand2_1
Xhold822 hold822/A VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_6
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3363__A1 _7052_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold844 hold844/A VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6325_ _6613_/Q _5976_/B _5993_/X _6623_/Q VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
Xhold855 hold855/A VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3537_ _7049_/Q hold16/A _3536_/Y _6706_/Q VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__a22o_1
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold877 hold877/A VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1058_A _7081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold888 hold888/A VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold899 hold899/A VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6256_ _6698_/Q _5997_/X _6004_/X _6575_/Q VGND VGND VPWR VPWR _6256_/X sky130_fd_sc_hd__a22o_1
X_3468_ _7073_/Q _5506_/A _4250_/A _6691_/Q _3466_/X VGND VGND VPWR VPWR _3481_/A
+ sky130_fd_sc_hd__a221o_4
XANTENNA__6301__B2 _6735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2201 _5454_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2212 _6612_/Q VGND VGND VPWR VPWR hold824/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5207_ _5207_/A _5222_/A _5533_/B VGND VGND VPWR VPWR _5208_/S sky130_fd_sc_hd__and3_1
Xhold2223 _6758_/Q VGND VGND VPWR VPWR hold580/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2234 _6642_/Q VGND VGND VPWR VPWR hold740/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5280__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6187_ _6923_/Q _5995_/X _6184_/X _6186_/X VGND VGND VPWR VPWR _6188_/C sky130_fd_sc_hd__a211oi_1
XANTENNA__4863__A1 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2245 _4189_/X VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3399_ _6955_/Q _3291_/Y _5326_/A _6915_/Q VGND VGND VPWR VPWR _3399_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3666__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1500 hold111/X VGND VGND VPWR VPWR _4276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1511 _7219_/A VGND VGND VPWR VPWR hold105/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2256 hold801/X VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2267 _6512_/Q VGND VGND VPWR VPWR hold815/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1522 _7123_/Q VGND VGND VPWR VPWR hold282/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1533 _5397_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5138_ _5138_/A _5138_/B _5138_/C VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__and3_1
Xhold2278 _6882_/Q VGND VGND VPWR VPWR hold947/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1544 hold335/X VGND VGND VPWR VPWR _5469_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_11_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2289 hold727/X VGND VGND VPWR VPWR _5448_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1555 hold506/X VGND VGND VPWR VPWR _3983_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1566 _5288_/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1577 hold318/X VGND VGND VPWR VPWR _5441_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1588 _6952_/Q VGND VGND VPWR VPWR hold377/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5069_ _5069_/A _5069_/B VGND VGND VPWR VPWR _5072_/C sky130_fd_sc_hd__and2_1
XANTENNA__3418__A2 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1599 _6703_/Q VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5812__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5455__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4298__C hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input40_A mgmt_gpio_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3657__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4854__B2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7100__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6056__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2790 _7107_/Q VGND VGND VPWR VPWR hold661/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3409__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4909__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3593__A1 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3593__B2 _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5365__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4440_ _4701_/A _4808_/B _4917_/A VGND VGND VPWR VPWR _4457_/C sky130_fd_sc_hd__a21o_1
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold107 hold107/A VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold118 hold118/A VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4489__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold129 hold129/A VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4371_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4719_/A sky130_fd_sc_hd__and2b_4
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7061__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6110_ _6864_/Q _5999_/X _6019_/X _6984_/Q _6109_/X VGND VGND VPWR VPWR _6113_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3355_/A _3322_/B VGND VGND VPWR VPWR _3563_/B sky130_fd_sc_hd__nand2_8
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7090_ _7130_/CLK _7090_/D fanout465/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__B1 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6837_/Q _6339_/B _6029_/X _6040_/Y _5647_/Y VGND VGND VPWR VPWR _6041_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A _3862_/A VGND VGND VPWR VPWR _3253_/Y sky130_fd_sc_hd__nand2_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__B2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3184_ _3921_/A VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6047__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6943_ _7063_/CLK _6943_/D fanout460/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5270__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _6963_/CLK _6874_/D fanout463/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5825_ _6955_/Q _5672_/X _5822_/X _5824_/X VGND VGND VPWR VPWR _5826_/C sky130_fd_sc_hd__a211o_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _6936_/Q _5659_/X _5669_/X _7048_/Q VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3584__A1 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4707_ _4391_/Y _4969_/A _4705_/Y _4832_/D _4640_/Y VGND VGND VPWR VPWR _4707_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3584__B2 _6720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5687_ _5685_/A _5689_/B _5687_/C VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__and3b_4
XANTENNA__5275__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4638_ _4638_/A _4638_/B VGND VGND VPWR VPWR _4638_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__4399__B _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold641 _5333_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4569_ _4569_/A _4569_/B _4569_/C VGND VGND VPWR VPWR _4569_/X sky130_fd_sc_hd__and3_1
Xhold652 hold652/A VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3887__A2 _6434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold663 hold663/A VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6308_ _6632_/Q _5971_/X _5990_/X _6647_/Q _6307_/X VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a221o_1
Xhold674 hold674/A VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold685 hold685/A VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold696 hold696/A VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6286__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6239_ _6233_/X _6339_/B _6239_/C _6239_/D VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__and4b_1
Xhold2020 hold524/X VGND VGND VPWR VPWR _4202_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__A2 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2031 _6771_/Q VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2042 hold807/X VGND VGND VPWR VPWR _4081_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2053 _3990_/X VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2064 hold521/X VGND VGND VPWR VPWR _4058_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 _4156_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1330 _6611_/Q VGND VGND VPWR VPWR _4167_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2086 hold745/X VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6038__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1341 _4259_/X VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2097 _6698_/Q VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1352 _6943_/Q VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1363 _6934_/Q VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1374 hold184/X VGND VGND VPWR VPWR _4050_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1385 _5571_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1396 _5206_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5013__A1 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6210__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input88_A spimemio_flash_io1_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5721__C1 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6277__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5252__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _6502_/Q _3940_/A1 _6458_/Q VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3871_ _3879_/B _3868_/B _3869_/A _3903_/A _3870_/X VGND VGND VPWR VPWR _6445_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6201__B1 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5610_ _5610_/A _6491_/Q VGND VGND VPWR VPWR _5639_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ _6753_/CLK _6590_/D fanout435/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3566__A1 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5541_ _5541_/A0 _5577_/A1 _5541_/S VGND VGND VPWR VPWR _5541_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3566__B2 _6715_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ hold159/X _5580_/A1 _5478_/S VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__mux2_1
X_7211_ _7211_/A VGND VGND VPWR VPWR _7211_/X sky130_fd_sc_hd__clkbuf_2
X_4423_ _4574_/A _4523_/A VGND VGND VPWR VPWR _4522_/B sky130_fd_sc_hd__nand2b_4
XFILLER_133_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4012__B _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7142_ _7180_/CLK _7142_/D fanout448/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
X_4354_ _4447_/B _4663_/D _4682_/A _4365_/B VGND VGND VPWR VPWR _4356_/B sky130_fd_sc_hd__and4_2
Xfanout406 _5317_/B VGND VGND VPWR VPWR _5533_/B sky130_fd_sc_hd__buf_12
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6268__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3305_ hold87/X hold78/X VGND VGND VPWR VPWR _3390_/B sky130_fd_sc_hd__and2_4
X_7073_ _7073_/CLK _7073_/D fanout444/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout439 fanout454/X VGND VGND VPWR VPWR _6407_/A sky130_fd_sc_hd__buf_12
X_4285_ _4285_/A0 _5583_/A1 _4285_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6024_ _7077_/Q _6013_/X _6017_/X _7069_/Q _6023_/X VGND VGND VPWR VPWR _6024_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ _6872_/Q VGND VGND VPWR VPWR _3236_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5491__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5243__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6967_/CLK _6926_/D fanout460/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout442_A fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6857_ _7017_/CLK _6857_/D fanout461/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5808_ _7090_/Q _5681_/X _5803_/X _5804_/X _5807_/X VGND VGND VPWR VPWR _5808_/X
+ sky130_fd_sc_hd__a2111o_2
X_6788_ _6793_/CLK _6788_/D _3959_/B VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ _6871_/Q _5674_/X _5736_/X _5738_/X VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6402__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 hold460/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 hold471/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold482 hold482/A VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6259__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold493 hold493/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4809__A1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4809__B2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input142_A wb_dat_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5482__A1 _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _6596_/Q VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1171 _5554_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1182 _5464_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _7087_/Q VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5234__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4084__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__C _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3796__A1 _6795_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4745__B1 _4714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3428__S _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3547_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3720__A1 _6958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3720__B2 _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4070_ _4070_/A0 _5189_/A1 _4070_/S VGND VGND VPWR VPWR _4070_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5473__A1 _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5225__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4972_ _4972_/A _4972_/B VGND VGND VPWR VPWR _4972_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5776__A2 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6711_ _6746_/CLK _6711_/D _6416_/A VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3923_ _6816_/Q _5610_/A _3197_/Y _3915_/Y VGND VGND VPWR VPWR _3923_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6642_ _6733_/CLK _6642_/D _3959_/B VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3854_ _3903_/A _3199_/A _3807_/B _3854_/B1 VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__a31o_1
XFILLER_177_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _6730_/CLK _6573_/D _6399_/A VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ _6479_/Q _4000_/A _4304_/A _6732_/Q _3784_/X VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a221o_2
X_5524_ _5524_/A _5569_/B VGND VGND VPWR VPWR _5532_/S sky130_fd_sc_hd__and2_4
XFILLER_173_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7203__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5455_ _5455_/A0 _5563_/A1 _5460_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5553__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4406_ _4477_/A _4477_/B VGND VGND VPWR VPWR _5150_/A sky130_fd_sc_hd__and2_2
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5386_ _5386_/A0 _5584_/A1 _5388_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5700__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7125_ _7125_/CLK _7125_/D fanout469/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3711__A1 _6846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4337_ _4337_/A0 _5581_/A1 _4339_/S VGND VGND VPWR VPWR _4337_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout392_A _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7056_ _7112_/CLK _7056_/D fanout468/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4268_ _4268_/A hold9/X VGND VGND VPWR VPWR _4273_/S sky130_fd_sc_hd__and2_2
XANTENNA__5464__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6007_ _6017_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _6007_/X sky130_fd_sc_hd__and3_4
X_3219_ _7000_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4199_ _4199_/A0 _5277_/A1 _4199_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1305_A _6880_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5216__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5767__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6909_ _7094_/CLK _6909_/D fanout450/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5924__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1939_A _6955_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3950__A1 _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5463__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4587__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3702__A1 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3702__B2 _7118_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold290 hold290/A VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5455__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3466__B1 _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5211__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5758__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6183__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3570_ _6597_/Q _4146_/A _4134_/A _6587_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5930__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3941__A1 _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5373__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ _5240_/A0 _5303_/A1 _5244_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4497__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _5171_/A0 _5193_/A1 _5174_/S VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__mux2_1
Xhold2608 _4258_/X VGND VGND VPWR VPWR hold548/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2619 hold778/X VGND VGND VPWR VPWR _4198_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4122_ _4122_/A _5533_/B VGND VGND VPWR VPWR _4127_/S sky130_fd_sc_hd__and2_2
XFILLER_96_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1907 _6622_/Q VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1918 _7217_/A VGND VGND VPWR VPWR hold584/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5446__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1929 hold283/X VGND VGND VPWR VPWR _5342_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4053_ _4053_/A0 hold39/X _4055_/S VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3457__B1 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_4__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5749__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4955_ _4955_/A _4955_/B _4955_/C _4955_/D VGND VGND VPWR VPWR _4957_/C sky130_fd_sc_hd__nand4_1
XANTENNA__5548__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ _7151_/Q _7152_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__and2b_4
XFILLER_177_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4886_ _4886_/A _4976_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6625_ _6826_/CLK _6625_/D _6407_/A VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_4
X_3837_ _6462_/Q _6657_/Q _3830_/Y _3836_/X _3846_/S VGND VGND VPWR VPWR _3837_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6174__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4185__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6556_ _7191_/CLK _6556_/D VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5921__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3768_ _6869_/Q _5281_/A _4334_/A _6757_/Q _3767_/X VGND VGND VPWR VPWR _3769_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout405_A _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__A1 input89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5507_ _5507_/A0 _5534_/A1 _5514_/S VGND VGND VPWR VPWR _5507_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4688__A _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6487_ _6821_/CLK _6487_/D fanout443/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfstp_2
X_3699_ _6822_/Q _5226_/A _5226_/B _5202_/A _6805_/Q VGND VGND VPWR VPWR _3699_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__5283__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1255_A _7038_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5438_ _5438_/A0 _5582_/A1 _5442_/S VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 hold1867/X VGND VGND VPWR VPWR hold479/A sky130_fd_sc_hd__buf_6
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5369_ _5369_/A0 _5567_/A1 _5370_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4200__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7108_ _7108_/CLK _7108_/D fanout451/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5437__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7039_ _7137_/CLK _7039_/D fanout466/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3448__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3999__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A wb_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5458__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7196__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__B1 _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6165__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5912__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A mgmt_gpio_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5193__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5428__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3439__B1 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5222__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6141__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5368__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4740_ _4947_/A _4712_/Y _4728_/Y _4737_/Y _4739_/X VGND VGND VPWR VPWR _4740_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4671_/A _4683_/A VGND VGND VPWR VPWR _4691_/B sky130_fd_sc_hd__nor2_8
XANTENNA__6156__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4167__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6410_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and2_1
XFILLER_174_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3622_ _7015_/Q _5443_/A _5362_/A _6943_/Q _3621_/X VGND VGND VPWR VPWR _3627_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6341_ _6341_/A0 _6340_/X _6341_/S VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__mux2_1
X_3553_ _3553_/A _3553_/B VGND VGND VPWR VPWR _4176_/A sky130_fd_sc_hd__nor2_4
XFILLER_127_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6272_ _6601_/Q _5995_/X _6019_/X _6734_/Q _6271_/X VGND VGND VPWR VPWR _6279_/A
+ sky130_fd_sc_hd__a221o_1
X_3484_ _6633_/Q _4188_/A _4316_/A _6746_/Q VGND VGND VPWR VPWR _3484_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5223_ _6818_/Q _5536_/A1 hold10/X VGND VGND VPWR VPWR _5223_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2405 hold841/X VGND VGND VPWR VPWR _4070_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2416 _6475_/Q VGND VGND VPWR VPWR hold861/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2427 _4193_/X VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5154_ _4402_/Y _4570_/C _4570_/D _4968_/Y _4534_/Y VGND VGND VPWR VPWR _5155_/D
+ sky130_fd_sc_hd__o221a_1
Xhold2438 _6483_/Q VGND VGND VPWR VPWR hold857/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2449 _7025_/Q VGND VGND VPWR VPWR hold835/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1704 _6554_/Q VGND VGND VPWR VPWR hold984/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5419__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1715 _6802_/Q VGND VGND VPWR VPWR hold416/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4890__A2 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1726 hold428/X VGND VGND VPWR VPWR hold1726/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ _3422_/Y hold989/A _4106_/S VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1737 _6546_/Q VGND VGND VPWR VPWR hold985/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5085_ _5143_/A _5139_/C _5165_/B _5006_/Y VGND VGND VPWR VPWR _5085_/X sky130_fd_sc_hd__a31o_1
Xhold1748 _5181_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1759 _4261_/X VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A0 _4035_/X _4046_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5987_ _6019_/A _6008_/A _6019_/C VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__and3_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5278__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4938_ _5011_/A _4601_/A _4466_/A VGND VGND VPWR VPWR _4938_/X sky130_fd_sc_hd__a21o_2
XANTENNA__3602__B1 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4945__A3 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_41 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6147__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4570_/C _4655_/A _4590_/Y _4713_/Y VGND VGND VPWR VPWR _4870_/D sky130_fd_sc_hd__o22a_1
XANTENNA_52 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _6608_/CLK _6608_/D _6413_/A VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_85 _3529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6539_ _6753_/CLK _6539_/D fanout435/X VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6410__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3381__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput181 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3669__B1 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput192 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4330__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2950 _7153_/Q VGND VGND VPWR VPWR _5629_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2961 _7143_/Q VGND VGND VPWR VPWR _5598_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2972 _7156_/Q VGND VGND VPWR VPWR _5640_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2983 _6491_/Q VGND VGND VPWR VPWR _5640_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4149__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3372__A2 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7180__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A2 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4085__A0 _3737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4624__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5910_ _6694_/Q _5658_/X _5664_/X _6759_/Q VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a22o_1
X_6890_ _7108_/CLK _6890_/D fanout451/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5841_ _6860_/Q _5651_/X _5662_/X _6900_/Q VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5772_ _6490_/Q _7162_/Q _5771_/X VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__a21bo_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4723_ _4812_/A _4725_/B VGND VGND VPWR VPWR _4770_/B sky130_fd_sc_hd__nand2_2
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4654_ _4917_/C _4838_/B _4917_/B VGND VGND VPWR VPWR _4655_/B sky130_fd_sc_hd__nand3b_2
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3605_ _7056_/Q _5488_/A _4328_/A _6755_/Q VGND VGND VPWR VPWR _3605_/X sky130_fd_sc_hd__a22o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
X_4585_ _4948_/A _4724_/C VGND VGND VPWR VPWR _4973_/C sky130_fd_sc_hd__nand2_1
Xhold801 hold801/A VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_2
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold812 hold812/A VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold823 hold823/A VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_2
Xhold834 hold834/A VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 uart_enabled VGND VGND VPWR VPWR _3970_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _6633_/Q _5971_/X _6007_/X _6534_/Q _6323_/X VGND VGND VPWR VPWR _6327_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3536_ _3563_/A _3553_/B VGND VGND VPWR VPWR _3536_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__3363__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold856 hold856/A VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold867 hold867/A VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold878 hold878/A VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold889 hold889/A VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6255_ _6255_/A _6255_/B _6255_/C VGND VGND VPWR VPWR _6264_/C sky130_fd_sc_hd__nor3_1
X_3467_ _3550_/A hold88/X VGND VGND VPWR VPWR _4250_/A sky130_fd_sc_hd__nor2_8
XANTENNA__5561__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6301__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2202 _6644_/Q VGND VGND VPWR VPWR hold753/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4312__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5206_ _5206_/A0 _5303_/A1 _5206_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
Xhold2213 hold824/X VGND VGND VPWR VPWR _4168_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2224 hold580/X VGND VGND VPWR VPWR _4336_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6186_ _6851_/Q _6007_/X _6019_/X _6987_/Q _6185_/X VGND VGND VPWR VPWR _6186_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2235 hold740/X VGND VGND VPWR VPWR _4204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3398_ _6891_/Q _5299_/A _3389_/Y _3395_/X _3397_/X VGND VGND VPWR VPWR _3406_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_130_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2246 _7029_/Q VGND VGND VPWR VPWR hold747/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1501 _4276_/X VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1512 hold105/X VGND VGND VPWR VPWR _4025_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5137_ _5086_/Y _5137_/B _5137_/C VGND VGND VPWR VPWR _5137_/X sky130_fd_sc_hd__and3b_1
Xhold2257 _4210_/X VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2268 hold815/X VGND VGND VPWR VPWR _4051_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1523 hold282/X VGND VGND VPWR VPWR _5567_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout472_A fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1534 _6486_/Q VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2279 hold947/X VGND VGND VPWR VPWR _5296_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1545 _5469_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1556 _3983_/X VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1567 _6987_/Q VGND VGND VPWR VPWR hold300/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5068_ _4391_/Y _4580_/Y _4584_/Y _4765_/Y _4438_/Y VGND VGND VPWR VPWR _5069_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1578 _5441_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1589 hold377/X VGND VGND VPWR VPWR _5375_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4019_ _4019_/A0 _4018_/X _4029_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6405__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4206__A _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4579__C _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4551__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5471__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4303__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input33_A mask_rev_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4854__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4087__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6056__A1 _7102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2780 _5351_/X VGND VGND VPWR VPWR hold639/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2791 hold661/X VGND VGND VPWR VPWR _5549_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7140__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4790__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3593__A2 _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold108 hold108/A VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 _7196_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4370_ _4955_/A _4513_/B VGND VGND VPWR VPWR _4370_/Y sky130_fd_sc_hd__nand2_2
XFILLER_153_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3321_ _3563_/A hold15/X VGND VGND VPWR VPWR _5551_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5381__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6040_ _6032_/X _6040_/B _6313_/D VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__6295__B2 _6740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3998_/S hold20/X _3252_/B1 VGND VGND VPWR VPWR _3252_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _6437_/Q VGND VGND VPWR VPWR _3183_/Y sky130_fd_sc_hd__inv_2
XANTENNA_hold2402_A _7106_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6047__B2 _7038_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6942_ _7001_/CLK _6942_/D fanout466/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3805__B1 _3803_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6873_ _7063_/CLK _6873_/D fanout461/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5824_ _6987_/Q _5656_/X _5668_/X _7059_/Q _5823_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5755_ _6992_/Q _5929_/B _5682_/X _7040_/Q _5754_/X VGND VGND VPWR VPWR _5760_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6863__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5556__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4706_ _4826_/A _4735_/B VGND VGND VPWR VPWR _4832_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3584__A2 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5686_ _5689_/A _5686_/B _5688_/C VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__and3_4
XFILLER_175_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4637_ _4637_/A _4637_/B _4637_/C _4637_/D VGND VGND VPWR VPWR _4726_/B sky130_fd_sc_hd__nor4_2
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold620 hold620/A VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4568_ _4568_/A _4881_/B VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__nand2_2
Xhold631 hold631/A VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold642 hold642/A VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap350 _3354_/B VGND VGND VPWR VPWR _3550_/A sky130_fd_sc_hd__buf_12
Xhold653 _4232_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3519_ _6552_/Q _4092_/A _5169_/A _6773_/Q _3518_/X VGND VGND VPWR VPWR _3529_/A
+ sky130_fd_sc_hd__a221o_4
X_6307_ _6592_/Q _5985_/X _5999_/X _6551_/Q VGND VGND VPWR VPWR _6307_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold664 hold664/A VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold675 hold675/A VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4499_ _4682_/A _4693_/B _4447_/B VGND VGND VPWR VPWR _4499_/Y sky130_fd_sc_hd__a21oi_2
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5291__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6286__A1 _6581_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold697 hold697/A VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1335_A _6942_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6238_ _6238_/A _6238_/B _6238_/C _6238_/D VGND VGND VPWR VPWR _6239_/D sky130_fd_sc_hd__nor4_1
XFILLER_104_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2010 _4335_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2021 _4202_/X VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2032 _5172_/X VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2043 _7128_/Q VGND VGND VPWR VPWR hold829/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2054 _7008_/Q VGND VGND VPWR VPWR hold870/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6899_/Q _5989_/X _5994_/X _7067_/Q _6168_/X VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2065 _6846_/Q VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _4215_/X VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1331 _4167_/X VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1502_A _6996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2076 _6932_/Q VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2087 _4192_/X VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1342 _6890_/Q VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2098 hold549/X VGND VGND VPWR VPWR _4264_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1353 hold128/X VGND VGND VPWR VPWR _5365_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1364 hold258/X VGND VGND VPWR VPWR _5355_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1375 _6485_/Q VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _6840_/Q VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _7070_/Q VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5797__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6416__A _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6210__A1 _6996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6821_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5466__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5721__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output237_A _3937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5788__B1 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A _3870_/B VGND VGND VPWR VPWR _3870_/X sky130_fd_sc_hd__and2_1
XFILLER_149_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6201__B2 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5376__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ _5540_/A0 _5567_/A1 _5540_/S VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3566__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5960__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5471_ hold751/X _5579_/A1 _5478_/S VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_54_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4422_ _4574_/A _4495_/B VGND VGND VPWR VPWR _4610_/A sky130_fd_sc_hd__nor2_2
X_7210_ _7210_/A VGND VGND VPWR VPWR _7210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5712__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7141_ _7180_/CLK _7141_/D fanout446/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_2
X_4353_ _4447_/B _4682_/A _4365_/B VGND VGND VPWR VPWR _4360_/A sky130_fd_sc_hd__nand3_2
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout407 hold9/A VGND VGND VPWR VPWR _5578_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__6268__A1 _6591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3304_ hold62/X hold22/X VGND VGND VPWR VPWR _3686_/B sky130_fd_sc_hd__nand2b_4
X_7072_ _7072_/CLK _7072_/D fanout461/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_4
X_4284_ _4284_/A0 hold43/X _4285_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
X_6023_ _6877_/Q _6004_/X _6007_/X _6845_/Q VGND VGND VPWR VPWR _6023_/X sky130_fd_sc_hd__a22o_1
X_3235_ _6880_/Q VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5779__B1 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _7061_/CLK _6925_/D fanout450/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6856_ _7091_/CLK _6856_/D fanout452/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5807_ _6866_/Q _5673_/X _5805_/X _5806_/X VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__a211o_1
X_6787_ _6835_/CLK _6787_/D _3959_/B VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfrtp_4
X_3999_ _3999_/A0 _5577_/A1 _3999_/S VGND VGND VPWR VPWR _3999_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5286__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5951__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5738_ _6951_/Q _5672_/X _5679_/X _6903_/Q _5737_/X VGND VGND VPWR VPWR _5738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5669_ _5689_/A _5689_/B _5687_/C VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__and3_4
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5703__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 hold450/A VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold461 hold461/A VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold483 hold483/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A wb_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1150 _6442_/Q VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3493__A1 _3974_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3493__B2 _6716_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1161 hold202/X VGND VGND VPWR VPWR _4149_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1172 _7119_/Q VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 _6839_/Q VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 hold232/X VGND VGND VPWR VPWR _5527_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6785__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6195__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5196__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4745__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3548__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5942__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5170__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3720__A2 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6489__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3484__A1 _6633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2100_A _6783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4971_ _4971_/A _4981_/B VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__nand2_1
X_6710_ _6731_/CLK hold44/X _6413_/A VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_4
X_3922_ _4222_/B _3922_/B VGND VGND VPWR VPWR _3922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3787__A2 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6641_ _6733_/CLK _6641_/D _3959_/B VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfstp_4
X_3853_ _3853_/A0 _3880_/A0 _3853_/S VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6186__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4304__A _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6572_ _6730_/CLK hold59/X _6399_/A VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfrtp_4
X_3784_ _7029_/Q _5461_/A _4009_/A _6487_/Q VGND VGND VPWR VPWR _3784_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5523_ _5523_/A0 _5577_/A1 _5523_/S VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ _5454_/A0 _5562_/A1 _5460_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4405_ _3890_/Y _4492_/B _4356_/B _4341_/X VGND VGND VPWR VPWR _4477_/B sky130_fd_sc_hd__a31oi_4
XFILLER_117_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5161__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5385_ _5385_/A0 _5583_/A1 _5388_/S VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7124_ _7124_/CLK _7124_/D fanout471/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_4
X_4336_ _4336_/A0 _5238_/A1 _4339_/S VGND VGND VPWR VPWR _4336_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3711__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7133_/CLK _7055_/D fanout469/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_4
X_4267_ _4267_/A0 _5189_/A1 _4267_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6110__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_A _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6006_ _5637_/A _6015_/B _6017_/A _5985_/X _6005_/X VGND VGND VPWR VPWR _6010_/B
+ sky130_fd_sc_hd__a311o_1
X_3218_ _7008_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4693__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4198_ _4198_/A0 _5233_/A1 _4199_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3778__A2 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6908_ _6992_/CLK _6908_/D fanout463/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6839_ _7073_/CLK _6839_/D fanout444/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6177__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6413__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5924__B1 _5914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3702__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold291 hold291/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6101__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6168__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5915__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5391__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5694__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5170_ _5170_/A0 _5237_/A1 _5174_/S VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2609 _6721_/Q VGND VGND VPWR VPWR hold927/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4121_ _4121_/A0 _5583_/A1 hold58/X VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1908 hold818/X VGND VGND VPWR VPWR _4180_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1919 hold584/X VGND VGND VPWR VPWR _4021_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4052_ _4052_/A0 _5583_/A1 _4055_/S VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3457__A1 _7106_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3457__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3203__A _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4954_ _4954_/A _5117_/B _5038_/B _4954_/D VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__and4_1
X_3905_ _6656_/Q _3904_/A _3904_/B _3903_/Y VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__a31o_1
XANTENNA__6159__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4885_ _4391_/Y _4584_/Y _4683_/A VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6624_ _6826_/CLK _6624_/D _6407_/A VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5906__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3836_ _6462_/Q _6461_/Q _6460_/Q hold60/A VGND VGND VPWR VPWR _3836_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5382__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3767_ _6803_/Q _5207_/A hold47/A _5452_/A _7021_/Q VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a32o_1
X_6555_ _7191_/CLK _6555_/D VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5564__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6654__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3393__B1 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5506_ _5506_/A _5533_/B VGND VGND VPWR VPWR _5514_/S sky130_fd_sc_hd__and2_4
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4688__B _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6486_ _6486_/CLK _6486_/D fanout434/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfstp_4
X_3698_ _6743_/Q _4316_/A _4122_/A _6575_/Q _3697_/X VGND VGND VPWR VPWR _3703_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5437_ _5437_/A0 _5572_/A1 _5442_/S VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6331__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput330 hold1849/X VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__buf_6
Xoutput341 hold1771/X VGND VGND VPWR VPWR hold427/A sky130_fd_sc_hd__buf_6
XFILLER_161_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ _5368_/A0 _5584_/A1 _5370_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3696__A1 _6796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7107_ _7107_/CLK _7107_/D fanout451/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4319_ _4319_/A0 _5581_/A1 _4321_/S VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__mux2_1
X_5299_ _5299_/A _5569_/B VGND VGND VPWR VPWR _5307_/S sky130_fd_sc_hd__and2_4
XFILLER_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7038_ _7124_/CLK _7038_/D fanout467/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5373__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5474__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input63_A mgmt_gpio_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3687__A1 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3687__B2 _6783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3439__A1 _7018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3439__B2 _6800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5222__B _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4651__A3 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A1 _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4670_ _4637_/A _4637_/B _4667_/X _4669_/X _4387_/Y VGND VGND VPWR VPWR _4703_/A
+ sky130_fd_sc_hd__o311a_1
X_3621_ _6786_/Q _5178_/A _4206_/A _6646_/Q VGND VGND VPWR VPWR _3621_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5364__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5384__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3375__B1 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6340_ _6529_/Q _6339_/B _6339_/X VGND VGND VPWR VPWR _6340_/X sky130_fd_sc_hd__o21ba_1
X_3552_ _6953_/Q _3291_/Y _3427_/Y _6793_/Q _3551_/X VGND VGND VPWR VPWR _3556_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6271_ _6586_/Q _5989_/X _5999_/X _6550_/Q VGND VGND VPWR VPWR _6271_/X sky130_fd_sc_hd__a22o_1
X_3483_ _3553_/A _3516_/B VGND VGND VPWR VPWR _4316_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2432_A _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5222_ _5222_/A _5226_/B hold9/A VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__and3_1
XFILLER_130_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3678__B2 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2406 _4070_/X VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2417 hold861/X VGND VGND VPWR VPWR _3993_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5153_ _5137_/X _5152_/Y _5147_/X _5146_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__a211o_1
Xhold2428 _7097_/Q VGND VGND VPWR VPWR hold730/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2439 _4005_/X VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1705 hold984/X VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1716 hold416/X VGND VGND VPWR VPWR _5199_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4104_ _3462_/Y hold979/A _4106_/S VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5084_ _4698_/Y _5011_/X _5022_/C _5081_/Y VGND VGND VPWR VPWR _5165_/B sky130_fd_sc_hd__o211a_1
Xhold1727 _6586_/Q VGND VGND VPWR VPWR hold631/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1738 hold985/X VGND VGND VPWR VPWR hold438/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1749 _6719_/Q VGND VGND VPWR VPWR hold632/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4035_ _4059_/A0 _5572_/A1 _4056_/C VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5559__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _6019_/B _6018_/B _6016_/C VGND VGND VPWR VPWR _5986_/X sky130_fd_sc_hd__and3_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _4729_/A _4688_/B _4935_/X _4936_/Y _4539_/Y VGND VGND VPWR VPWR _4954_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_20 _5894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4868_ _4638_/Y _4712_/Y _4922_/C _4867_/X _5063_/B VGND VGND VPWR VPWR _4870_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_42 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5355__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6608_/CLK hold76/X _6399_/A VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_75 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _6654_/Q _3816_/Y _3904_/B _3840_/B VGND VGND VPWR VPWR _3846_/S sky130_fd_sc_hd__o31a_4
XANTENNA__5294__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _3680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4729_/A _4714_/Y _4779_/X _4798_/X _4539_/Y VGND VGND VPWR VPWR _4800_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_97 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3366__B1 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6538_ _6753_/CLK _6538_/D fanout440/X VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6469_ _3958_/A1 _6469_/D _6419_/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3669__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput171 _3972_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
Xoutput182 _5763_/A VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2940 _7172_/Q VGND VGND VPWR VPWR _5970_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2951 _6460_/Q VGND VGND VPWR VPWR _3846_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2962 _6457_/Q VGND VGND VPWR VPWR _3853_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2973 _6491_/Q VGND VGND VPWR VPWR _5622_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6216__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5815__C1 _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6083__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1999_A _7032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4094__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5830__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5469__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5346__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5897__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output267_A _6782_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__B _3960_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6074__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5821__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5379__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _6884_/Q _5667_/X _5682_/X _7044_/Q VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5585__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _3239_/Y _5707_/B _5760_/Y wire346/X _6490_/Q VGND VGND VPWR VPWR _5771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7087__RESET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3596__B1 _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4722_ _5001_/A _4732_/B _4722_/C VGND VGND VPWR VPWR _4722_/X sky130_fd_sc_hd__and3_1
XANTENNA__5337__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4653_ _4682_/A _4693_/B _4504_/X VGND VGND VPWR VPWR _4838_/B sky130_fd_sc_hd__a21o_1
XANTENNA_hold2647_A _6801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3348__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5888__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3604_ _3604_/A _3604_/B _3604_/C _3604_/D VGND VGND VPWR VPWR _3615_/B sky130_fd_sc_hd__nor4_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_2
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_4
X_4584_ _4808_/A _4710_/A VGND VGND VPWR VPWR _4584_/Y sky130_fd_sc_hd__nand2_2
Xhold802 hold802/A VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3965_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold813 hold813/A VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_2
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6323_ _6539_/Q _5983_/X _6005_/X _6696_/Q VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
Xhold824 hold824/A VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold835 hold835/A VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3535_ _3535_/A _3550_/B VGND VGND VPWR VPWR _4170_/A sky130_fd_sc_hd__nor2_8
Xhold846 hold846/A VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold857 hold857/A VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold868 hold868/A VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold879 hold879/A VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3466_ input7/X _3315_/Y _4152_/A _6603_/Q VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__a22o_1
X_6254_ _6610_/Q _5976_/B _5993_/X _6620_/Q _6253_/X VGND VGND VPWR VPWR _6255_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5205_ _5205_/A0 _5527_/A1 _5206_/S VGND VGND VPWR VPWR _5205_/X sky130_fd_sc_hd__mux2_1
Xhold2203 hold753/X VGND VGND VPWR VPWR _4207_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2214 _4168_/X VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3397_ _6995_/Q _5416_/A _4000_/A _6485_/Q _3396_/X VGND VGND VPWR VPWR _3397_/X
+ sky130_fd_sc_hd__a221o_1
X_6185_ _6963_/Q _5992_/X _6012_/X _7003_/Q VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__a22o_1
Xhold2225 _4336_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2236 _4204_/X VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2247 hold747/X VGND VGND VPWR VPWR _5462_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3520__B1 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1502 _6996_/Q VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1513 _4025_/X VGND VGND VPWR VPWR hold106/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5136_ _5136_/A _5136_/B _5136_/C VGND VGND VPWR VPWR _5137_/C sky130_fd_sc_hd__and3_1
Xhold2258 _6790_/Q VGND VGND VPWR VPWR hold579/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2269 _6595_/Q VGND VGND VPWR VPWR hold615/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1524 _5567_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1535 _4008_/X VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6065__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1546 _6615_/Q VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5067_ _5067_/A _5067_/B VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__and2_1
Xhold1557 _6831_/Q VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4076__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1568 hold300/X VGND VGND VPWR VPWR _5414_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1579 _6876_/Q VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout465_A input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1113_A _6983_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4018_ _4050_/A0 _5563_/A1 _4047_/C VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5812__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5289__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5025__B1 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5576__A1 wire371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5969_ _5969_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4206__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5328__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6421__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input165_A wb_sel_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5500__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3511__B1 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input26_A mask_rev_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6056__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2770 _5340_/X VGND VGND VPWR VPWR hold763/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2781 _7091_/Q VGND VGND VPWR VPWR hold659/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2792 _6938_/Q VGND VGND VPWR VPWR hold942/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4067__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5199__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5016__B1 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5567__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4116__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3578__B1 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5319__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4527__C1 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold109 hold109/A VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3971__A _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3320_ _3322_/B hold14/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__nand2_4
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3251_ _5147_/A1 _3998_/S VGND VGND VPWR VPWR _3251_/Y sky130_fd_sc_hd__nand2b_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3502__B1 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3182_ _6460_/Q VGND VGND VPWR VPWR _3182_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6047__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4058__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6941_ _7001_/CLK _6941_/D fanout466/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6872_ _6992_/CLK _6872_/D fanout463/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3211__A _7064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5558__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5823_ _6979_/Q _5660_/X _5669_/X _7051_/Q VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5837__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3569__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5754_ _7016_/Q _5664_/X _5686_/X _7008_/Q VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _5009_/B _5150_/C VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5685_ _5685_/A _5686_/B _5689_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_4
XFILLER_136_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5947__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _4663_/D _4840_/A _4498_/X _3969_/A VGND VGND VPWR VPWR _4636_/X sky130_fd_sc_hd__a31o_2
XFILLER_175_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold610 hold610/A VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold621 hold621/A VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4567_ _4980_/A _4693_/B VGND VGND VPWR VPWR _5100_/C sky130_fd_sc_hd__nand2_1
XANTENNA__5572__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold632 hold632/A VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3741__B1 _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6306_ _6730_/Q _5987_/X _6004_/X _6577_/Q _6305_/X VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a221o_1
Xhold654 hold654/A VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3518_ _6865_/Q _5272_/A _4000_/A _6483_/Q VGND VGND VPWR VPWR _3518_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold665 hold665/A VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold676 hold676/A VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4498_ _4637_/B _4498_/B VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__and2_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold687 hold687/A VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6286__A2 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold698 hold698/A VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6237_ _6584_/Q _5989_/X _6013_/X _6624_/Q _6236_/X VGND VGND VPWR VPWR _6238_/D
+ sky130_fd_sc_hd__a221o_1
Xhold2000 hold827/X VGND VGND VPWR VPWR _5465_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3449_ _3449_/A _3449_/B _3449_/C VGND VGND VPWR VPWR _3461_/A sky130_fd_sc_hd__nor3_1
Xhold2011 _6587_/Q VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4297__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2022 _6614_/Q VGND VGND VPWR VPWR hold688/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2033 _7064_/Q VGND VGND VPWR VPWR hold846/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2044 hold829/X VGND VGND VPWR VPWR _5573_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _7123_/Q _5978_/X _6016_/X _7043_/Q VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__a22o_1
Xhold2055 hold870/X VGND VGND VPWR VPWR _5438_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1310 _7134_/Q VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _6951_/Q VGND VGND VPWR VPWR hold153/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2066 hold534/X VGND VGND VPWR VPWR _5256_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1332 _6476_/Q VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6038__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2077 hold362/X VGND VGND VPWR VPWR _5352_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__nand3_1
Xhold1343 hold259/X VGND VGND VPWR VPWR _5305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2088 _6650_/Q VGND VGND VPWR VPWR hold533/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4049__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1354 _5365_/X VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2099 _4264_/X VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6099_ _7024_/Q _5971_/X _6007_/X _6848_/Q _6098_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1365 _5355_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1376 _4007_/X VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 hold402/X VGND VGND VPWR VPWR _5249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 hold260/X VGND VGND VPWR VPWR _5508_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5549__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7170__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6210__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5048__A _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5482__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3732__B1 _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6277__A2 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4288__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6029__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5788__B2 _7089_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3799__B1 _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6201__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5470_ _5470_/A _5578_/B VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__and2_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4421_ _4955_/A _4955_/B _4477_/C VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__and3_4
XANTENNA__5392__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7140_ _7140_/CLK _7140_/D fanout473/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3723__B1 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4352_ _4682_/A _4365_/B VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout408 _5317_/B VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__buf_12
XANTENNA__6268__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3303_ hold62/X hold22/X VGND VGND VPWR VPWR _5207_/A sky130_fd_sc_hd__and2b_4
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4283_ _4283_/A0 _5581_/A1 _4285_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
X_7071_ _7073_/CLK _7071_/D fanout445/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4279__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3206__A _7104_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6022_ _6853_/Q _5983_/X _5995_/X _6917_/Q _6021_/X VGND VGND VPWR VPWR _6039_/A
+ sky130_fd_sc_hd__a221o_1
X_3234_ _6888_/Q VGND VGND VPWR VPWR _3234_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2979_A _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6924_ _6936_/CLK _6924_/D fanout465/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _6945_/CLK _6855_/D _6416_/A VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5567__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5806_ _6978_/Q _5660_/X _5669_/X _7050_/Q VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6786_ _6786_/CLK _6786_/D fanout435/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4203__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3998_ _3998_/A0 _7202_/Q _3998_/S VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5737_ _6935_/Q _5659_/X _5687_/X _6919_/Q VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1180_A _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1278_A _6888_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5668_ _5689_/A _5684_/B _5687_/C VGND VGND VPWR VPWR _5668_/X sky130_fd_sc_hd__and3_4
XFILLER_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4619_ _4570_/C _4655_/A _4922_/A _4617_/X _4618_/Y VGND VGND VPWR VPWR _4622_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_191_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5703__B2 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5599_ _7142_/Q _7143_/Q _7144_/Q _5599_/D VGND VGND VPWR VPWR _5601_/B sky130_fd_sc_hd__nand4_2
XFILLER_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3714__B1 _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold440 hold440/A VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold451 hold451/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold462 hold462/A VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold473 _4036_/X VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6259__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold484 hold484/A VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold495 _4236_/X VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 hold217/X VGND VGND VPWR VPWR _5572_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 hold37/X VGND VGND VPWR VPWR _3994_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4690__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3493__A2 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _4149_/X VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1173 hold231/X VGND VGND VPWR VPWR _5563_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input128_A wb_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 hold219/X VGND VGND VPWR VPWR _5248_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1195 _5527_/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5477__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__A1 _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input93_A trap VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4745__A2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5942__A1 _6642_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5942__B2 _6632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5506__A _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3705__B1 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3484__A2 _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _4598_/A _5001_/B _4883_/X VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__a21boi_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3921_/A _3921_/B VGND VGND VPWR VPWR _3922_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5387__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6640_ _6794_/CLK _6640_/D _3959_/B VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3852_ _6468_/Q _3852_/B VGND VGND VPWR VPWR _3853_/S sky130_fd_sc_hd__nor2_1
XANTENNA__6186__A1 _6851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6495__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6571_ _6730_/CLK _6571_/D _6413_/A VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4304__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3783_ _3783_/A _3783_/B _3783_/C _3783_/D VGND VGND VPWR VPWR _3802_/B sky130_fd_sc_hd__nor4_1
X_5522_ _5522_/A0 _5549_/A1 _5523_/S VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5453_ hold902/X _5561_/A1 _5460_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5416__A _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4404_ _4492_/B _4356_/B _4650_/B VGND VGND VPWR VPWR _4477_/A sky130_fd_sc_hd__a21o_4
XFILLER_145_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6994_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5384_ _5384_/A0 _5582_/A1 _5388_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7123_ _7124_/CLK _7123_/D fanout471/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_4
X_4335_ _4335_/A0 _5543_/A1 _4339_/S VGND VGND VPWR VPWR _4335_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7054_ _7133_/CLK _7054_/D fanout467/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6110__A1 _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4266_ _4266_/A0 _5195_/A1 _4267_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6110__B2 _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6815_/CLK sky130_fd_sc_hd__clkbuf_16
X_6005_ _6017_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__and3_4
X_3217_ _7016_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
X_4197_ hold177/X _5581_/A1 _4199_/S VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout378_A _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6992_/CLK _6907_/D fanout463/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5297__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6838_ _7078_/CLK _6838_/D fanout444/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_11_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5924__A1 _6527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6769_ _6809_/CLK _6769_/D fanout433/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5326__A _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold270 hold270/A VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold281 _4054_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6101__A1 _7032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6101__B2 _6888_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3466__A2 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A1 _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5915__A1 _6689_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output297_A _6804_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6456__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4140__A _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4351__B1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2043_A _7128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4120_ _4120_/A0 hold43/X hold58/X VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1909 _4180_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4051_ _4051_/A0 _5582_/A1 _4055_/S VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3457__A2 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_2
XANTENNA__5851__B1 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4953_ _4368_/B _4407_/Y _4938_/X _4786_/X VGND VGND VPWR VPWR _4954_/D sky130_fd_sc_hd__o31a_1
XFILLER_33_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3904_ _3904_/A _3904_/B VGND VGND VPWR VPWR _3904_/Y sky130_fd_sc_hd__nand2_1
X_4884_ _4658_/B _4564_/Y _4965_/C _5102_/B _4883_/X VGND VGND VPWR VPWR _4892_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_32_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6623_ _6746_/CLK _6623_/D _6416_/A VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_4
X_3835_ _3831_/B _3834_/X _3835_/S VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ _7191_/CLK _6554_/D VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ _7117_/Q _5560_/A _4322_/A _6747_/Q _3765_/X VGND VGND VPWR VPWR _3769_/C
+ sky130_fd_sc_hd__a221o_1
X_5505_ _5505_/A0 _5577_/A1 _5505_/S VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6485_ _6486_/CLK _6485_/D fanout434/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_4
X_3697_ _7086_/Q _5524_/A _3325_/Y _7038_/Q VGND VGND VPWR VPWR _3697_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4688__C _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5436_ _5436_/A0 _5571_/A1 _5442_/S VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6331__A1 _6741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput320 hold982/X VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__buf_6
XFILLER_133_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput331 hold1887/X VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__buf_6
Xoutput342 hold972/X VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__buf_6
X_5367_ _5367_/A0 _5448_/A1 _5370_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3696__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7106_ _7106_/CLK _7106_/D fanout472/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_4
X_4318_ _4318_/A0 _5238_/A1 _4321_/S VGND VGND VPWR VPWR _4318_/X sky130_fd_sc_hd__mux2_1
X_5298_ _5298_/A0 _5568_/A1 _5298_/S VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6095__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7037_ _7086_/CLK _7037_/D fanout467/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__4196__S _4199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4249_ _4249_/A0 hold71/X _4249_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3448__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1310_A _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3620__A2 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4030__C1 _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input56_A mgmt_gpio_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5490__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3687__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6086__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3439__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5833__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5222__C hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A2 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _6911_/Q _5326_/A _4194_/A _6636_/Q _3619_/X VGND VGND VPWR VPWR _3627_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3551_ _6454_/Q _3977_/A _4286_/A _6721_/Q VGND VGND VPWR VPWR _3551_/X sky130_fd_sc_hd__a22o_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2258_A _6790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _6636_/Q _5994_/X _5996_/X _6651_/Q _6269_/X VGND VGND VPWR VPWR _6270_/X
+ sky130_fd_sc_hd__a221o_1
X_3482_ _3553_/A _3648_/A VGND VGND VPWR VPWR _4188_/A sky130_fd_sc_hd__nor2_8
X_5221_ _5221_/A0 hold275/X _5221_/S VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3678__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2407 _6787_/Q VGND VGND VPWR VPWR hold899/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2425_A _6633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2418 _3993_/X VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5152_ _5152_/A _5152_/B VGND VGND VPWR VPWR _5152_/Y sky130_fd_sc_hd__nand2_1
Xhold2429 hold730/X VGND VGND VPWR VPWR _5538_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6077__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1706 hold450/X VGND VGND VPWR VPWR hold1706/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4103_ _6351_/A0 hold990/A _4106_/S VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__mux2_1
Xhold1717 _5199_/X VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5083_ _5083_/A _5083_/B _5083_/C _5083_/D VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__and4_1
Xhold1728 _4137_/X VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1739 hold438/X VGND VGND VPWR VPWR hold1739/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3214__A _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5824__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4034_ _4034_/A0 _4033_/X _4046_/S VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _6018_/B _6007_/C _6016_/C VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__and3_4
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4936_ _5150_/A _4936_/B VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand2_2
XFILLER_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3602__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _3775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4590_/Y _4712_/Y _4866_/X _4616_/B VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__o211a_1
XANTENNA_32 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5575__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_43 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6608_/CLK _6606_/D _6399_/A VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout410_A _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ _6445_/Q _3863_/A VGND VGND VPWR VPWR _3904_/B sky130_fd_sc_hd__and2_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 hold16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4947_/A _4714_/Y _4797_/X _4536_/Y VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_87 _3769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3366__A1 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_98 _6486_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6745_/CLK _6537_/D fanout440/X VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3366__B2 _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3749_ _6609_/Q _4164_/A _3562_/Y input98/X _3748_/X VGND VGND VPWR VPWR _3750_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6468_ _3958_/A1 _6468_/D _6418_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_4
X_5419_ _5419_/A0 _5572_/A1 _5424_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _6399_/A _6430_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
XFILLER_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput172 _7206_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XANTENNA__3669__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4866__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput183 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput194 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_87_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6068__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2930 _7180_/Q VGND VGND VPWR VPWR _6217_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2941 hold52/A VGND VGND VPWR VPWR _3832_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2952 _3844_/X VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2963 _7186_/Q VGND VGND VPWR VPWR _6345_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2974 _7155_/Q VGND VGND VPWR VPWR _5635_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5291__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input110_A wb_adr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5485__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6059__B1 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5806__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5282__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6231__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5770_ _5770_/A _5770_/B _5770_/C _5770_/D VGND VGND VPWR VPWR _5770_/Y sky130_fd_sc_hd__nor4_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3596__A1 _7032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4721_ _4726_/A _4989_/B _4993_/B VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__nand3_1
XFILLER_148_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__B2 _6642_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5395__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4652_ _4652_/A _4652_/B VGND VGND VPWR VPWR _4652_/Y sky130_fd_sc_hd__nand2_2
XFILLER_147_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__buf_2
X_3603_ _6745_/Q _4316_/A _3977_/A _6453_/Q _3602_/X VGND VGND VPWR VPWR _3604_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_hold64_A hold64/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_2
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
X_4583_ _4658_/A _4583_/B VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__nor2_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3971_/A sky130_fd_sc_hd__buf_8
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3209__A _7080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold803 hold803/A VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold814 hold814/A VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3966_/B sky130_fd_sc_hd__buf_2
X_6322_ _6746_/Q _6014_/X _6320_/X _6321_/X VGND VGND VPWR VPWR _6327_/A sky130_fd_sc_hd__a211o_1
XFILLER_190_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
X_3534_ _6475_/Q _3988_/A _4304_/A _6736_/Q _3532_/X VGND VGND VPWR VPWR _3543_/A
+ sky130_fd_sc_hd__a221o_4
Xhold825 hold825/A VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_2
XFILLER_143_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold836 hold836/A VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6298__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold858 hold858/A VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _6640_/Q _5986_/X _5998_/X _6580_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
Xhold869 hold869/A VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _3550_/A _3533_/B VGND VGND VPWR VPWR _4152_/A sky130_fd_sc_hd__nor2_4
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5204_ _5204_/A0 _5571_/A1 _5206_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
Xhold2204 _4207_/X VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6184_ _6939_/Q _5980_/X _6008_/X _7107_/Q VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a22o_1
Xhold2215 _6471_/Q VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6239__B _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3396_ _7139_/Q _3295_/Y hold31/A _7099_/Q VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__a22o_1
Xhold2226 _6510_/Q VGND VGND VPWR VPWR hold531/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2237 _6755_/Q VGND VGND VPWR VPWR hold820/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1503 hold329/X VGND VGND VPWR VPWR _5424_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5135_ _5135_/A _5135_/B _5135_/C _5135_/D VGND VGND VPWR VPWR _5135_/X sky130_fd_sc_hd__and4_1
Xhold2248 _5462_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1514 hold106/X VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2259 hold579/X VGND VGND VPWR VPWR _5186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1525 _7027_/Q VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1536 _6737_/Q VGND VGND VPWR VPWR _4311_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1547 hold107/X VGND VGND VPWR VPWR _4172_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1558 hold271/X VGND VGND VPWR VPWR _5239_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5066_ _5155_/B _5130_/B _5131_/A VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__and3_1
XANTENNA__5273__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1569 _5414_/X VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4017_ _4017_/A0 _4016_/X _4029_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout458_A _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6222__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5968_ _6529_/Q _5678_/Y _5959_/X _5967_/X _6341_/S VGND VGND VPWR VPWR _5968_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _5115_/B _5047_/C _4919_/C VGND VGND VPWR VPWR _5126_/B sky130_fd_sc_hd__and3_1
X_5899_ _6536_/Q _5651_/X _5653_/X _6531_/Q VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input158_A wb_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2760 hold617/X VGND VGND VPWR VPWR _5377_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2771 _7075_/Q VGND VGND VPWR VPWR hold650/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2782 hold659/X VGND VGND VPWR VPWR _5531_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2793 hold942/X VGND VGND VPWR VPWR _5359_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5264__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A mask_rev_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5016__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4224__C1 _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3578__A1 _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ hold52/A hold19/X _6657_/Q VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__mux2_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3502__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3181_ _6468_/Q VGND VGND VPWR VPWR _3181_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5255__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ _6994_/CLK _6940_/D fanout462/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6871_ _7063_/CLK _6871_/D fanout460/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5822_ _6963_/Q _5680_/X _5685_/X _7075_/Q VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3569__A1 _6952_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5753_ _6960_/Q _5680_/X _5685_/X _7072_/Q _5752_/X VGND VGND VPWR VPWR _5760_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4704_ _4704_/A _5124_/B _4704_/C _4704_/D VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__and4_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5684_ _5689_/A _5684_/B _5687_/C VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__and3b_4
XANTENNA__4781__A3 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4635_ _4986_/C _4880_/B _4632_/X _4965_/B _4561_/X VGND VGND VPWR VPWR _4759_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold600 hold600/A VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold611 hold611/A VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4566_ _4981_/A _4693_/B VGND VGND VPWR VPWR _4616_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3881__B _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3741__A1 _6901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6305_ _6597_/Q _5991_/X _6005_/X _6695_/Q VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__a22o_1
Xhold644 hold644/A VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap352 hold30/X VGND VGND VPWR VPWR _3535_/A sky130_fd_sc_hd__buf_12
XFILLER_116_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3517_ _3553_/B _3535_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__nor2_8
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4497_ _4701_/A _4693_/B VGND VGND VPWR VPWR _4643_/D sky130_fd_sc_hd__nand2_1
XFILLER_143_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold677 hold677/A VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold688 hold688/A VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1056_A _6572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold699 hold699/A VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6236_ _6687_/Q _5980_/X _6017_/X _6769_/Q VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6140__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3448_ _6994_/Q _5416_/A _5308_/A _6898_/Q _3434_/X VGND VGND VPWR VPWR _3449_/C
+ sky130_fd_sc_hd__a221o_1
Xhold2001 _5465_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2012 hold726/X VGND VGND VPWR VPWR _4138_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2023 hold688/X VGND VGND VPWR VPWR _4171_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2034 hold846/X VGND VGND VPWR VPWR _5501_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6191_/A2 _6166_/X _6167_/S VGND VGND VPWR VPWR _6167_/X sky130_fd_sc_hd__mux2_1
Xhold2045 _5573_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1300 _6895_/Q VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3379_ _6876_/Q _5281_/A _5362_/A _6948_/Q VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__a22o_1
Xhold2056 _5438_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1311 _6847_/Q VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 hold153/X VGND VGND VPWR VPWR _5374_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2067 _7000_/Q VGND VGND VPWR VPWR hold808/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _4417_/B _4688_/C _4779_/X _4954_/A VGND VGND VPWR VPWR _5149_/C sky130_fd_sc_hd__o211a_1
Xhold1333 hold250/X VGND VGND VPWR VPWR _3995_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2078 _5352_/X VGND VGND VPWR VPWR hold363/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1344 _5305_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6098_ _6856_/Q _5983_/X _6005_/X _6944_/Q VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__a22o_1
Xhold2089 hold533/X VGND VGND VPWR VPWR _4214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5246__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1355 _6749_/Q VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1366 _7079_/Q VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1377 _6886_/Q VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5049_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__and4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1388 _5249_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1399 _5508_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5797__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5721__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3732__A1 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5237__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2590 _4217_/X VGND VGND VPWR VPWR hold678/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5788__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3966__B _3966_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3420__B1 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4763__A3 _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5960__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4420_ _4420_/A _4461_/B _4420_/C VGND VGND VPWR VPWR _4477_/C sky130_fd_sc_hd__and3_2
XFILLER_172_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5712__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4351_ _4637_/A _4637_/B _4574_/A _4637_/D VGND VGND VPWR VPWR _4365_/B sky130_fd_sc_hd__o211a_4
XFILLER_141_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2240_A _6791_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3302_ hold21/X hold28/A hold55/A VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__and3_1
X_7070_ _7078_/CLK _7070_/D fanout445/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfstp_2
X_4282_ _4282_/A0 _5580_/A1 _4285_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5476__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6021_ _6893_/Q _5989_/X _6015_/X _7013_/Q VGND VGND VPWR VPWR _6021_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3233_ _6896_/Q VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5228__A1 _5228_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5779__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3222__A _6976_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6923_ _6996_/CLK _6923_/D fanout462/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6854_ _7082_/CLK _6854_/D fanout460/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5805_ _6874_/Q _5674_/X _5680_/X _6962_/Q VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__a22o_1
X_6785_ _6835_/CLK _6785_/D _3959_/B VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_4
X_3997_ _3997_/A0 wire371/X _3999_/S VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5400__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _6975_/Q _5660_/X _5669_/X _7047_/Q VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3411__B1 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5951__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5667_ _5689_/A _5686_/B _5688_/C VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3b_4
XFILLER_108_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4618_ _4625_/A _5048_/A _4562_/A VGND VGND VPWR VPWR _4618_/Y sky130_fd_sc_hd__o21ai_1
X_5598_ _5598_/A1 _5591_/Y _5641_/B _5597_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5703__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4199__S _4199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3714__B2 _6605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold441 hold441/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4549_ _4724_/C _4628_/A VGND VGND VPWR VPWR _5138_/A sky130_fd_sc_hd__nand2_1
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold463 hold463/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 hold474/A VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold485 hold485/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
Xhold496 hold496/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5467__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6219_ _6644_/Q _5990_/X _5996_/X _6649_/Q VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7199_ _3950_/A1 _7199_/D _6346_/B VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3478__B1 _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1130 _6467_/Q VGND VGND VPWR VPWR _3253_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _5572_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _3994_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _7023_/Q VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1174 _5563_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _5248_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1196 _6969_/Q VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6195__A2 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5942__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input86_A spimemio_flash_io0_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3953__A1 _6811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5493__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5506__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3705__A1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4130__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3977__A _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3920_ _6435_/Q _3183_/Y _6654_/Q _3904_/A _3920_/B1 VGND VGND VPWR VPWR _3920_/X
+ sky130_fd_sc_hd__a41o_1
X_3851_ _3920_/B1 _3199_/Y _3814_/B _3851_/B1 VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__a31o_1
XANTENNA__6186__A2 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2190_A _6735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4197__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6570_ _7121_/CLK _6570_/D _6399_/A VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3782_ _6949_/Q _3291_/Y _3293_/Y input71/X _3781_/X VGND VGND VPWR VPWR _3783_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5933__A2 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3944__A1 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5521_ _5521_/A0 _5584_/A1 _5523_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2455_A _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4601__A _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5452_ _5452_/A _5578_/B VGND VGND VPWR VPWR _5460_/S sky130_fd_sc_hd__and2_4
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4403_ _4724_/B _4625_/A VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5416__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5383_ _5383_/A0 _5581_/A1 _5388_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3217__A _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7122_ _7139_/CLK _7122_/D fanout471/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4334_ _4334_/A hold9/A VGND VGND VPWR VPWR _4339_/S sky130_fd_sc_hd__and2_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5449__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7053_ _7134_/CLK _7053_/D fanout469/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_87_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4265_ _4265_/A0 _5194_/A1 _4267_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7160__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6110__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6004_ _6015_/B _6017_/A _6007_/C VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__and3_4
XFILLER_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4121__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3216_ _7024_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4196_ _4196_/A0 _5238_/A1 _4199_/S VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout440_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6906_ _6992_/CLK _6906_/D fanout463/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3632__B1 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6837_ _7073_/CLK _6837_/D fanout444/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__6177__A2 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5924__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6768_ _7203_/CLK _6768_/D _6346_/B VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5719_ _6942_/Q _5658_/X _5681_/X _7086_/Q VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__a22o_1
X_6699_ _6736_/CLK _6699_/D fanout436/X VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5326__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3699__B1 _5202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold260 hold260/A VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold282 hold282/A VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold293 _4063_/X VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6101__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input140_A wb_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _4059_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__B1 _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6168__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5915__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5236__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4140__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6340__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7183__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2036_A _6526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ _4050_/A0 _5563_/A1 _4055_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5851__A1 _6964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4952_ _4601_/A _4491_/Y _4514_/B _4947_/A _4802_/B VGND VGND VPWR VPWR _5038_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3903_ _3903_/A _3904_/A VGND VGND VPWR VPWR _3903_/Y sky130_fd_sc_hd__nor2_1
X_4883_ _4438_/Y _4601_/A _4601_/B _4580_/Y _4581_/X VGND VGND VPWR VPWR _4883_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6159__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6622_ _6756_/CLK _6622_/D fanout441/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_4
X_3834_ hold61/A _3247_/Y _3834_/S VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5906__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6553_ _7191_/CLK _6553_/D VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfxtp_1
X_3765_ input11/X _3310_/Y _5209_/S _7206_/A VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a22o_4
XFILLER_192_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3393__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5504_ _5504_/A0 _5567_/A1 _5505_/S VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__mux2_1
X_6484_ _6486_/CLK _6484_/D fanout434/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfstp_4
X_3696_ _6796_/Q _3319_/Y _4164_/A _6610_/Q _3695_/X VGND VGND VPWR VPWR _3703_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpad_flashh_clk_buff_inst _3958_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_133_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5435_ _5435_/A0 _5534_/A1 _5442_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput310 _3966_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6331__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput321 hold1753/X VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__buf_6
Xoutput332 hold1831/X VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__buf_6
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold1783/X VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__buf_6
X_5366_ _5366_/A0 _5582_/A1 _5370_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7105_ _7137_/CLK _7105_/D fanout466/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_4
X_4317_ _4317_/A0 _5543_/A1 _4321_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout390_A _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5297_ _5297_/A0 _5549_/A1 _5298_/S VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6095__A1 _7056_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7036_ _7099_/CLK _7036_/D fanout471/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6095__B2 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4248_ _4248_/A0 hold35/X _4249_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5842__A1 _6852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4179_ hold166/X _5581_/A1 _4181_/S VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__B1 _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4241__A _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4598__D _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6322__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4333__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input49_A mgmt_gpio_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6086__B2 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5833__B2 _7011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6996_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__B _3974_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3375__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3550_ _3550_/A _3550_/B VGND VGND VPWR VPWR _4286_/A sky130_fd_sc_hd__nor2_8
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3481_ _3481_/A _3481_/B _3481_/C _3481_/D VGND VGND VPWR VPWR _3558_/A sky130_fd_sc_hd__nor4_2
XFILLER_115_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4324__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5220_ hold64/X _5220_/B _5220_/C VGND VGND VPWR VPWR _5221_/S sky130_fd_sc_hd__and3_1
XFILLER_142_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5151_ _5150_/X _5151_/B _5151_/C _5151_/D VGND VGND VPWR VPWR _5152_/B sky130_fd_sc_hd__and4b_2
Xhold2408 hold899/X VGND VGND VPWR VPWR _5182_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2419 _6717_/Q VGND VGND VPWR VPWR hold905/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4102_ _3616_/Y hold974/A _4106_/S VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1707 _6901_/Q VGND VGND VPWR VPWR hold620/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5082_ _4578_/A _4990_/B _5108_/A _5023_/A VGND VGND VPWR VPWR _5083_/D sky130_fd_sc_hd__o211a_1
Xhold1718 _6570_/Q VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1729 _6559_/Q VGND VGND VPWR VPWR hold989/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4033_ hold521/X _5562_/A1 _4056_/C VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5984_ _6008_/A _6018_/B _6019_/C VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__and3_4
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4935_ _5011_/A _4601_/A _4663_/D _4465_/B VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2954_A _6434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 _5002_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4638_/Y _4995_/A _4924_/C _4865_/X _5095_/B VGND VGND VPWR VPWR _4866_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_33 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_44 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _6731_/CLK _6605_/D _6413_/A VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_55 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ _6447_/Q _6446_/Q VGND VGND VPWR VPWR _3863_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_66 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4729_/A _4713_/Y _4796_/X _4534_/Y VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__o211a_1
XFILLER_165_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_77 hold31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_88 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3366__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6536_ _6753_/CLK _6536_/D fanout435/X VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_4
X_3748_ _7133_/Q _3295_/Y _3431_/Y input61/X VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__a22o_4
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3679_ _6918_/Q _5335_/A hold89/A _6713_/Q _3678_/X VGND VGND VPWR VPWR _3684_/A
+ sky130_fd_sc_hd__a221o_1
X_6467_ _3547_/A1 _6467_/D _6417_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4315__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5418_ _5418_/A0 _5571_/A1 _5424_/S VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__mux2_1
X_6398_ _6399_/A _6430_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _3973_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
Xoutput184 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
X_5349_ _5349_/A0 _5529_/A1 _5352_/S VGND VGND VPWR VPWR _5349_/X sky130_fd_sc_hd__mux2_1
Xoutput195 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2920 hold86/A VGND VGND VPWR VPWR _4907_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2931 _6659_/Q VGND VGND VPWR VPWR _4223_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2942 _6470_/Q VGND VGND VPWR VPWR _3811_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2953 _6682_/Q VGND VGND VPWR VPWR _3968_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2964 _7154_/Q VGND VGND VPWR VPWR _5633_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5815__A1 _6842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4618__A2 _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2975 _7140_/Q VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6138__D _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7019_ _7131_/CLK _7019_/D fanout452/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6446__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6240__A1 _6525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input103_A wb_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4306__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4146__A _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4649_/B _4720_/B _4720_/C VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__and3b_4
XFILLER_159_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__A2 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4793__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _4590_/Y _4648_/Y _4683_/A _5121_/A VGND VGND VPWR VPWR _4651_/X sky130_fd_sc_hd__o31a_1
XFILLER_159_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_2
X_3602_ input29/X _3307_/Y _3315_/Y input6/X VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__a22o_4
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3348__A2 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4582_ _4724_/B _4724_/C VGND VGND VPWR VPWR _4969_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5742__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_4
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_2
XFILLER_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_12
X_6321_ _6598_/Q _5991_/X _6018_/X _6721_/Q _6318_/X VGND VGND VPWR VPWR _6321_/X
+ sky130_fd_sc_hd__a221o_2
X_3533_ _3553_/A _3533_/B VGND VGND VPWR VPWR _4304_/A sky130_fd_sc_hd__nor2_8
Xhold804 hold804/A VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold815 hold815/A VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3960_/B sky130_fd_sc_hd__buf_4
XANTENNA_hold57_A hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold826 hold826/A VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6636__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_2
Xhold837 hold837/A VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold848 hold848/A VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6298__A1 _6572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6252_ _6630_/Q _5971_/X _6007_/X _6531_/Q _6251_/X VGND VGND VPWR VPWR _6255_/B
+ sky130_fd_sc_hd__a221o_1
Xhold859 hold859/A VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3464_ _3463_/X _3464_/A1 _3739_/S VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5203_ _5203_/A0 _5534_/A1 _5206_/S VGND VGND VPWR VPWR _5203_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7096__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6183_ _7131_/Q _5973_/X _5986_/X _7035_/Q _6182_/X VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2205 _7045_/Q VGND VGND VPWR VPWR hold764/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3395_ _7115_/Q _5551_/A _5263_/A _6859_/Q VGND VGND VPWR VPWR _3395_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3225__A _6960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2216 hold722/X VGND VGND VPWR VPWR _3989_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2227 hold531/X VGND VGND VPWR VPWR _4049_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5134_ _5134_/A _5155_/C VGND VGND VPWR VPWR _5134_/Y sky130_fd_sc_hd__nand2_1
Xhold2238 hold820/X VGND VGND VPWR VPWR _4332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3520__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2249 _6590_/Q VGND VGND VPWR VPWR hold616/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1504 _5424_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1515 _6852_/Q VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1526 hold301/X VGND VGND VPWR VPWR _5459_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6469__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1537 _4311_/X VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5065_ _4570_/C _4968_/Y _4903_/B _4622_/C _4539_/Y VGND VGND VPWR VPWR _5131_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1548 _4172_/X VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1559 _6520_/Q VGND VGND VPWR VPWR hold333/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4016_ hold531/X _5562_/A1 _4047_/C VGND VGND VPWR VPWR _4016_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3879__B _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6222__A1 _6604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6660__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5967_ _6539_/Q _5651_/X _5962_/X _5966_/X VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__a211o_1
X_4918_ _4365_/B _4988_/A _4840_/A _4917_/X VGND VGND VPWR VPWR _4919_/C sky130_fd_sc_hd__a22oi_4
XFILLER_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5898_ _6575_/Q _5667_/X _5682_/X _6451_/Q VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4849_ _5009_/A _4710_/A _4811_/B VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1370_A _7009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5733__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6519_ _6936_/CLK _6519_/D fanout463/X VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1635_A _6904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1802_A _6625_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3511__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2750 _6917_/Q VGND VGND VPWR VPWR hold786/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2761 _7222_/A VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2772 hold650/X VGND VGND VPWR VPWR _5513_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2783 _6957_/Q VGND VGND VPWR VPWR hold896/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2794 _5359_/X VGND VGND VPWR VPWR hold943/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5016__A2 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5496__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3578__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4775__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5724__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output272_A _6473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6709__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3502__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3180_ _6469_/Q VGND VGND VPWR VPWR _3879_/A sky130_fd_sc_hd__inv_2
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _7072_/CLK _6870_/D fanout460/X VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5821_ _6883_/Q _5667_/X _5687_/X _6923_/Q _5820_/X VGND VGND VPWR VPWR _5826_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3569__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5963__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5752_ _7056_/Q _5668_/X _5681_/X _7088_/Q VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4703_ _4703_/A _4703_/B _4703_/C _4703_/D VGND VGND VPWR VPWR _4704_/D sky130_fd_sc_hd__and4_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5683_ _7085_/Q _5681_/X _5682_/X _7037_/Q VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4634_ _5001_/A _4731_/A VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5715__B1 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4565_ _4971_/A _4693_/B VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__nand2_1
Xhold612 hold612/A VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold623 hold623/A VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3881__C _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6304_ _6304_/A _6304_/B _6304_/C _6304_/D VGND VGND VPWR VPWR _6314_/B sky130_fd_sc_hd__nor4_2
Xhold634 hold634/A VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3741__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3516_ _3544_/A _3516_/B VGND VGND VPWR VPWR _4092_/A sky130_fd_sc_hd__nor2_8
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap353 _3686_/B VGND VGND VPWR VPWR _3764_/B sky130_fd_sc_hd__buf_12
X_4496_ _4576_/A _4523_/A VGND VGND VPWR VPWR _4658_/B sky130_fd_sc_hd__nand2_4
Xhold656 hold656/A VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold678 hold678/A VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6140__B1 _6139_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6235_ _6722_/Q _5978_/X _5995_/X _6599_/Q _6234_/X VGND VGND VPWR VPWR _6238_/C
+ sky130_fd_sc_hd__a221o_1
X_3447_ _6890_/Q _5299_/A _5497_/A _7066_/Q _3435_/X VGND VGND VPWR VPWR _3449_/B
+ sky130_fd_sc_hd__a221o_1
Xhold689 hold689/A VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2002 _6579_/Q VGND VGND VPWR VPWR hold766/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2013 _4138_/X VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _4171_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2035 _5501_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6166_ _7177_/Q _6165_/X _6166_/S VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__mux2_1
X_3378_ _7028_/Q _5452_/A _3307_/Y input33/X _3348_/X VGND VGND VPWR VPWR _3383_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 _7136_/Q VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1301 hold139/X VGND VGND VPWR VPWR _5311_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2057 _7215_/A VGND VGND VPWR VPWR hold918/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1312 hold130/X VGND VGND VPWR VPWR _5257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2068 hold808/X VGND VGND VPWR VPWR _5429_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1323 _5374_/X VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A _5117_/B _5117_/C VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__and3_1
Xhold1334 _3995_/X VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2079 _6645_/Q VGND VGND VPWR VPWR hold527/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6097_ _6992_/Q _6014_/X _6095_/X _6096_/X VGND VGND VPWR VPWR _6102_/A sky130_fd_sc_hd__a211o_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout470_A input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1345 _6477_/Q VGND VGND VPWR VPWR hold214/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1216_A _6887_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1356 _4325_/X VGND VGND VPWR VPWR hold169/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5048_ _5048_/A _5048_/B VGND VGND VPWR VPWR _5049_/D sky130_fd_sc_hd__nand2_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1367 hold162/X VGND VGND VPWR VPWR _5518_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1378 hold244/X VGND VGND VPWR VPWR _5301_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1389 _6999_/Q VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _7086_/CLK _6999_/D fanout467/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1585_A _6473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4514__A _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5182__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input170_A wb_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3732__A2 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6131__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input31_A mask_rev_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2580 _6930_/Q VGND VGND VPWR VPWR hold948/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2591 _6793_/Q VGND VGND VPWR VPWR hold904/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1890 _4034_/X VGND VGND VPWR VPWR hold886/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6511__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6198__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3420__B2 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5173__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4350_ _4637_/A _4637_/B VGND VGND VPWR VPWR _4592_/B sky130_fd_sc_hd__nor2_2
XANTENNA__3723__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3301_ _3553_/A _3726_/A VGND VGND VPWR VPWR _5398_/A sky130_fd_sc_hd__nor2_8
XFILLER_99_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4281_ _4281_/A0 _5561_/A1 _4285_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6122__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _6861_/Q _5999_/X _6005_/X _6941_/Q VGND VGND VPWR VPWR _6020_/X sky130_fd_sc_hd__a22o_1
X_3232_ _6904_/Q VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6922_ _7052_/CLK _6922_/D fanout464/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6853_ _6945_/CLK _6853_/D _6416_/A VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4739__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5804_ _6946_/Q _5658_/X _5664_/X _7018_/Q VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5936__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6784_ _6786_/CLK _6784_/D _3959_/B VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_4
X_3996_ _3996_/A0 _7201_/Q _3998_/S VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ _6983_/Q _5656_/X _5663_/X _7023_/Q _5734_/X VGND VGND VPWR VPWR _5735_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3411__A1 _6801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6657__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5666_ _5689_/A _5679_/B _5688_/C VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_3_1_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5164__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4617_ _4522_/B _4570_/D _4614_/X _4616_/X VGND VGND VPWR VPWR _4617_/X sky130_fd_sc_hd__o211a_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5597_ _7142_/Q _7143_/Q _6490_/Q _6492_/Q _3924_/Y VGND VGND VPWR VPWR _5597_/X
+ sky130_fd_sc_hd__o221a_1
Xhold420 hold420/A VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3714__A2 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold431 hold431/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XANTENNA__4911__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4548_ _4574_/A _4463_/B _4569_/B _4546_/X _4770_/A VGND VGND VPWR VPWR _4548_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold442 hold442/A VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold464 hold464/A VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold475 hold475/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4479_ _4486_/A _4485_/B _4881_/A VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__and3_2
Xhold497 _4230_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6218_ _6594_/Q _5991_/X _6018_/X _6717_/Q VGND VGND VPWR VPWR _6218_/X sky130_fd_sc_hd__a22o_1
X_7198_ _3950_/A1 _7198_/D _6346_/B VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3478__B2 _6741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _5217_/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6149_ _7026_/Q _5971_/X _6007_/X _6850_/Q _6148_/X VGND VGND VPWR VPWR _6152_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _3253_/Y VGND VGND VPWR VPWR hold1131/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _6833_/Q VGND VGND VPWR VPWR _4233_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 hold38/X VGND VGND VPWR VPWR hold1153/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 hold208/X VGND VGND VPWR VPWR _5455_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1175 _7135_/Q VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1186 _6443_/Q VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 hold97/X VGND VGND VPWR VPWR _5394_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3650__B2 _6527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1967_A _7088_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5927__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7199__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6352__A0 _3462_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input79_A spi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3705__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6104__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3977__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3641__A1 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5918__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3850_ _3927_/A1 _3850_/A1 _3850_/S VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3781_ _6957_/Q _5380_/A _4152_/A _6599_/Q VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5394__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5520_ _5520_/A0 hold95/X _5523_/S VGND VGND VPWR VPWR _5520_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5451_ _5451_/A0 _5577_/A1 _5451_/S VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4402_ _4523_/A _4590_/B VGND VGND VPWR VPWR _4402_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__5697__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5382_ hold568/X _5562_/A1 _5388_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7121_ _7121_/CLK _7121_/D _6411_/A VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_4
X_4333_ _4333_/A0 _5277_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3932__S _3934_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2615_A _6588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4264_ _4264_/A0 _5193_/A1 _4267_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7052_ _7052_/CLK _7052_/D fanout464/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3215_ _7032_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
X_6003_ _7151_/Q _6007_/C _6016_/C _5989_/X _5997_/X VGND VGND VPWR VPWR _6010_/A
+ sky130_fd_sc_hd__a311o_1
X_4195_ _4195_/A0 _5543_/A1 _4199_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4424__A3 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6905_ _7017_/CLK _6905_/D fanout461/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3632__B2 _6797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6836_ _7091_/CLK _6836_/D fanout452/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5385__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6767_ _7203_/CLK _6767_/D _6346_/B VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_1
X_3979_ _3979_/A0 _5237_/A1 _3987_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3396__B1 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5718_ _5718_/A _5718_/B _5718_/C VGND VGND VPWR VPWR _5718_/Y sky130_fd_sc_hd__nor3_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6698_ _6736_/CLK _6698_/D fanout436/X VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5649_ _6342_/S VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6334__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3699__B2 _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold250 hold250/A VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6775__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold261 hold261/A VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold272 _5239_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold283 hold283/A VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_3_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input133_A wb_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3871__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A1 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6325__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5236__C _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5300__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5851__A2 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3988__A _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4951_ _4368_/A _4462_/Y _4934_/Y _5041_/A _4800_/B VGND VGND VPWR VPWR _5148_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3902_ _6682_/Q _3969_/B _3901_/Y _3921_/A VGND VGND VPWR VPWR _3902_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4882_ _4934_/B _4972_/B VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _6746_/CLK _6621_/D _6416_/A VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5367__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3833_ _3833_/A _3833_/B VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3378__B1 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6552_ _6753_/CLK _6552_/D fanout440/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfrtp_4
X_3764_ _3764_/A _3764_/B VGND VGND VPWR VPWR _5209_/S sky130_fd_sc_hd__nor2_4
XFILLER_146_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5503_ _5503_/A0 _5575_/A1 _5505_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
X_6483_ _6486_/CLK _6483_/D fanout434/X VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfstp_4
X_3695_ _6630_/Q _4188_/A _4322_/A _6748_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 _6807_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5434_ _5434_/A _5569_/B VGND VGND VPWR VPWR _5442_/S sky130_fd_sc_hd__and2_4
Xoutput311 _7232_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput322 hold1780/X VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__buf_6
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput333 hold1846/X VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__buf_6
Xoutput344 hold1726/X VGND VGND VPWR VPWR hold429/A sky130_fd_sc_hd__buf_6
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5365_ _5365_/A0 _5572_/A1 _5370_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5443__A _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7104_ _7112_/CLK _7104_/D fanout473/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4316_ _4316_/A hold9/X VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__and2_4
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5296_ _5296_/A0 _5575_/A1 _5298_/S VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6095__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7035_ _7084_/CLK _7035_/D fanout447/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
X_4247_ _4247_/A0 _5584_/A1 _4249_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout383_A _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1031_A _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5842__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4178_ _4178_/A0 _5238_/A1 _4181_/S VGND VGND VPWR VPWR _4178_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3605__A1 _7056_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6819_ _7086_/CLK _6819_/D fanout467/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5358__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3369__B1 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire427 _4389_/Y VGND VGND VPWR VPWR _4580_/A sky130_fd_sc_hd__buf_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4030__B2 _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4241__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6307__B1 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4869__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5353__A _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3541__B1 _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6086__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4097__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5833__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5499__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7143__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7150__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3780__B1 _5202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ input56/X _4241_/A _4158_/A _6608_/Q _3478_/X VGND VGND VPWR VPWR _3481_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5521__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5263__A _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2146_A _6573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__B1 _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _5150_/A _5150_/B _5150_/C VGND VGND VPWR VPWR _5150_/X sky130_fd_sc_hd__and3_1
XFILLER_69_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2409 _5182_/X VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4101_ _3675_/Y hold977/A _4106_/S VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6077__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5081_ _5081_/A _5081_/B VGND VGND VPWR VPWR _5081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1708 _5318_/X VGND VGND VPWR VPWR hold621/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1719 hold196/X VGND VGND VPWR VPWR _4118_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4032_ _4032_/A0 _4031_/X _4046_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5824__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5983_ _6019_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__and3_4
XFILLER_178_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4934_ _5009_/A _4934_/B VGND VGND VPWR VPWR _4934_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4260__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4865_ _4402_/Y _4570_/A _4651_/X _4856_/X _4864_/X VGND VGND VPWR VPWR _4865_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_20_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_12 _5140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6604_ _6608_/CLK _6604_/D _6413_/A VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3816_ _6656_/Q _3904_/A VGND VGND VPWR VPWR _3816_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_45 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_56 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4796_/A _4796_/B _4796_/C VGND VGND VPWR VPWR _4796_/X sky130_fd_sc_hd__and3_1
XFILLER_192_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_67 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 hold330/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _5880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6753_/CLK _6535_/D fanout440/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_4
X_3747_ _5207_/A _5222_/A _3745_/Y _3746_/X VGND VGND VPWR VPWR _3750_/C sky130_fd_sc_hd__a31o_1
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1079_A _6607_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3771__B1 _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6466_ _3547_/A1 _6466_/D _6416_/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfrtp_1
X_3678_ _6650_/Q _4212_/A _3562_/Y input96/X VGND VGND VPWR VPWR _3678_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5417_ _5417_/A0 hold275/X _5424_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6397_ _6399_/A _6430_/B VGND VGND VPWR VPWR _6397_/X sky130_fd_sc_hd__and2_1
XANTENNA__3392__S _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1246_A _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput174 _3974_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5348_ _5348_/A0 _5537_/A1 _5352_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2910 _3926_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6068__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2921 _7171_/Q VGND VGND VPWR VPWR _5969_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2932 _4223_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2943 _6676_/Q VGND VGND VPWR VPWR _3921_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4079__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5279_ _5279_/A0 _5549_/A1 _5280_/S VGND VGND VPWR VPWR _5279_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2954 _6434_/Q VGND VGND VPWR VPWR _3885_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7018_ _7099_/CLK _7018_/D fanout472/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2965 _7146_/Q VGND VGND VPWR VPWR _5606_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5815__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2976 _6810_/Q VGND VGND VPWR VPWR hold104/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5579__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7173__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6240__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4251__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4003__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input61_A mgmt_gpio_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3514__B1 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6059__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5806__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout390 _5536_/A1 VGND VGND VPWR VPWR _5581_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4146__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6231__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4720_/B _4650_/B VGND VGND VPWR VPWR _4683_/A sky130_fd_sc_hd__nand2_8
XFILLER_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_2
X_3601_ _6984_/Q _5407_/A _4176_/A _6622_/Q _3600_/X VGND VGND VPWR VPWR _3604_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_2
X_4581_ _4560_/B _4560_/C _4652_/A VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__a21bo_4
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5742__B2 _7039_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_2
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3753__B1 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6320_ _6648_/Q _5990_/X _5996_/X _6653_/Q VGND VGND VPWR VPWR _6320_/X sky130_fd_sc_hd__a22o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7232_/A sky130_fd_sc_hd__buf_6
Xhold805 hold805/A VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3532_ _6638_/Q _4194_/A _4322_/A _6751_/Q VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold816 _4051_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3934_/S sky130_fd_sc_hd__buf_8
XFILLER_115_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7231_/A sky130_fd_sc_hd__buf_4
XFILLER_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_2
Xhold827 hold827/A VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold838 hold838/A VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6298__A2 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold849 hold849/A VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6251_ _6536_/Q _5983_/X _6005_/X _6693_/Q VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__a22o_1
X_3463_ _6778_/Q _3462_/Y _3857_/B VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5202_ _5202_/A _5569_/B VGND VGND VPWR VPWR _5206_/S sky130_fd_sc_hd__and2_2
XANTENNA__4101__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6182_ _7091_/Q _5638_/X _5999_/X _6867_/Q VGND VGND VPWR VPWR _6182_/X sky130_fd_sc_hd__a22o_1
X_3394_ _7107_/Q _5542_/A _3336_/Y input27/X VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__a22o_1
Xhold2206 hold764/X VGND VGND VPWR VPWR _5480_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2217 _3989_/X VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2228 _6723_/Q VGND VGND VPWR VPWR hold574/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5133_ _4564_/Y _4968_/Y _5072_/C _5132_/X _4609_/B VGND VGND VPWR VPWR _5155_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold2239 _4332_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3940__S _6458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1505 _7028_/Q VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1516 hold346/X VGND VGND VPWR VPWR _5262_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1527 _5459_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1538 _7099_/Q VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5064_ _4569_/B _4510_/B _4625_/Y _4902_/A _4971_/Y VGND VGND VPWR VPWR _5130_/B
+ sky130_fd_sc_hd__o2111a_1
Xhold1549 _6884_/Q VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4015_ _4015_/A0 _4014_/X _4029_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7196__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4056__B _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6222__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5966_ _6701_/Q _5672_/X _5963_/X _5965_/X VGND VGND VPWR VPWR _5966_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4233__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4917_ _4917_/A _4917_/B _4917_/C _4917_/D VGND VGND VPWR VPWR _4917_/X sky130_fd_sc_hd__and4_1
X_5897_ _6743_/Q _5929_/B _5668_/X _6645_/Q _5884_/X VGND VGND VPWR VPWR _5897_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4848_ _4391_/Y _4580_/Y _4640_/Y VGND VGND VPWR VPWR _5049_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4779_ _4464_/Y _4569_/C _4688_/C _4947_/A VGND VGND VPWR VPWR _4779_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6518_ _6936_/CLK _6518_/D fanout463/X VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6449_ _3940_/A1 _6449_/D _6404_/X VGND VGND VPWR VPWR _6449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6936_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2740 _5282_/X VGND VGND VPWR VPWR hold680/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2751 _5336_/X VGND VGND VPWR VPWR hold787/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2762 hold849/X VGND VGND VPWR VPWR _4242_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2773 _6915_/Q VGND VGND VPWR VPWR hold640/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2784 _6874_/Q VGND VGND VPWR VPWR hold949/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6816_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2795 _6995_/Q VGND VGND VPWR VPWR hold645/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6563__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6788__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4224__B2 _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5724__B2 _6958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output265_A _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2011_A _6587_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2109_A _6782_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _7035_/Q _5655_/X _5679_/X _6907_/Q VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4215__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5751_ _5751_/A1 _6342_/S _5749_/X _5750_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__o22a_1
X_4702_ _5009_/B _4702_/B VGND VGND VPWR VPWR _4702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5682_ _5689_/A _5686_/B _5687_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_4
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4633_ _4658_/A _4633_/B VGND VGND VPWR VPWR _4731_/A sky130_fd_sc_hd__nor2_2
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5715__B2 _6950_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4564_ _4579_/B _4564_/B _4564_/C VGND VGND VPWR VPWR _4564_/Y sky130_fd_sc_hd__nand3_4
Xhold602 hold602/A VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold613 hold613/A VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6303_ _6690_/Q _5980_/X _6016_/X _6453_/Q _6302_/X VGND VGND VPWR VPWR _6304_/D
+ sky130_fd_sc_hd__a221o_1
Xhold624 hold624/A VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3515_ _3515_/A _3515_/B _3515_/C _3515_/D VGND VGND VPWR VPWR _3557_/A sky130_fd_sc_hd__nor4_1
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap354 _3356_/A VGND VGND VPWR VPWR _3563_/A sky130_fd_sc_hd__buf_12
X_4495_ _4718_/A _4495_/B VGND VGND VPWR VPWR _4693_/B sky130_fd_sc_hd__nor2_8
Xhold646 hold646/A VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3236__A _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold657 hold657/A VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold668 hold668/A VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6234_ _6737_/Q _6008_/X _6016_/X _6450_/Q VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a22o_1
Xhold679 hold679/A VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3446_ _6954_/Q _3291_/Y _4237_/S _3970_/A _3445_/X VGND VGND VPWR VPWR _3449_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2003 hold766/X VGND VGND VPWR VPWR _4129_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6842_/Q _6339_/B _6164_/X VGND VGND VPWR VPWR _6165_/X sky130_fd_sc_hd__o21ba_1
Xhold2014 _6535_/Q VGND VGND VPWR VPWR hold717/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _6582_/Q VGND VGND VPWR VPWR hold796/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3377_ _7124_/Q _5560_/A _5353_/A _6940_/Q _3376_/X VGND VGND VPWR VPWR _3383_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2036 _6526_/Q VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2047 hold845/X VGND VGND VPWR VPWR _5582_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1302 _6713_/Q VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5110_/Y _5113_/Y _5115_/X VGND VGND VPWR VPWR _5119_/C sky130_fd_sc_hd__o21ai_1
Xhold1313 _6993_/Q VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2058 hold918/X VGND VGND VPWR VPWR _4017_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _5429_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6096_ _6904_/Q _5985_/X _5994_/X _7064_/Q _6094_/X VGND VGND VPWR VPWR _6096_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1324 _6863_/Q VGND VGND VPWR VPWR hold149/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1335 _6942_/Q VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1346 hold214/X VGND VGND VPWR VPWR _3997_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1357 _6910_/Q VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5047_ _5047_/A _5126_/A _5047_/C VGND VGND VPWR VPWR _5110_/A sky130_fd_sc_hd__and3_1
Xhold1368 _5518_/X VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1379 _5301_/X VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6998_ _7133_/CLK _6998_/D fanout468/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5949_ _6608_/Q _5684_/X _5686_/X _6623_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input163_A wb_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2570 _5408_/X VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input24_A mask_rev_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2581 hold948/X VGND VGND VPWR VPWR _5350_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2592 hold904/X VGND VGND VPWR VPWR _5189_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6969__RESET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1880 hold790/X VGND VGND VPWR VPWR _5492_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1891 hold886/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5300__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3956__A0 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3420__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6459__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3708__B1 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3300_ _3347_/A _3338_/A VGND VGND VPWR VPWR _5416_/A sky130_fd_sc_hd__nor2_8
XFILLER_141_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4280_ hold89/X hold9/A VGND VGND VPWR VPWR _4285_/S sky130_fd_sc_hd__and2_2
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6122__B2 _7073_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3231_ _6912_/Q VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6921_ _6945_/CLK _6921_/D _6416_/A VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6852_ _7099_/CLK _6852_/D fanout471/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ _7066_/Q _5671_/X _5799_/X _5801_/X _5802_/X VGND VGND VPWR VPWR _5803_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4739__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6783_ _6826_/CLK _6783_/D _6407_/A VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__4334__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3995_ _3995_/A0 wire375/X _3999_/S VGND VGND VPWR VPWR _3995_/X sky130_fd_sc_hd__mux2_1
X_5734_ _7031_/Q _5655_/X _5678_/B _6967_/Q _5707_/B VGND VGND VPWR VPWR _5734_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3411__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5665_ _5685_/A _5684_/B _5676_/B VGND VGND VPWR VPWR _5929_/B sky130_fd_sc_hd__and3_4
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4616_ _4616_/A _4616_/B _5063_/B VGND VGND VPWR VPWR _4616_/X sky130_fd_sc_hd__and3_1
XFILLER_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5164__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5596_ _7142_/Q _7143_/Q VGND VGND VPWR VPWR _5641_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4911__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _4625_/B _4607_/B VGND VGND VPWR VPWR _4770_/A sky130_fd_sc_hd__nand2_1
Xhold432 hold432/A VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold443 hold443/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_3_5_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold454 hold454/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
Xhold465 _5240_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold476 hold476/A VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4478_ _4724_/C _4611_/A VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold487 hold487/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6217_ _6217_/A1 _6167_/S _6215_/X _6216_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__o22a_1
X_3429_ _3429_/A hold46/X _3430_/B VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__and3_4
X_7197_ _3950_/A1 _7197_/D _6346_/B VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3478__A2 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6148_ _6858_/Q _5983_/X _6005_/X _6946_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1110 _6744_/Q VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1121 _6855_/Q VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4509__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1132 _3254_/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 hold1143/A VGND VGND VPWR VPWR _5241_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1154 hold1154/A VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6079_ _7127_/Q _5973_/X _5988_/X _6871_/Q _6078_/X VGND VGND VPWR VPWR _6079_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _5455_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1176 hold228/X VGND VGND VPWR VPWR _5581_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1187 hold33/X VGND VGND VPWR VPWR _3996_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _5394_/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4978__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3650__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5927__B2 _6582_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3402__A2 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6104__A1 _6960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6104__B2 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4115__A0 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5863__B1 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3626__C1 _3625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6732__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5091__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3641__A2 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5918__B2 _6452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _6837_/Q _5245_/A _5202_/A _6804_/Q _3779_/X VGND VGND VPWR VPWR _3783_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2176_A _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5450_ _5450_/A0 _5549_/A1 _5451_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4170__A _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4401_ _4495_/B _4454_/A VGND VGND VPWR VPWR _4625_/A sky130_fd_sc_hd__nor2_8
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5381_ hold896/X _5561_/A1 _5388_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7120_ _7121_/CLK _7120_/D _6411_/A VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_4
X_4332_ _4332_/A0 _5233_/A1 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4106__A0 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7051_ _7084_/CLK _7051_/D fanout447/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_4
X_4263_ _4263_/A0 _5237_/A1 _4267_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6002_ _5637_/A _6001_/X _6000_/X _5992_/X _6019_/B VGND VGND VPWR VPWR _6002_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5854__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3214_ _7040_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4194_ _4194_/A _5533_/B VGND VGND VPWR VPWR _4199_/S sky130_fd_sc_hd__and2_4
XFILLER_28_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2977_A _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6904_ _6996_/CLK _6904_/D fanout463/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3632__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6835_ _6835_/CLK _6835_/D _3959_/B VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6031__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6766_ _7203_/CLK _6766_/D _4107_/B VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_2
X_3978_ _3879_/B _3978_/A1 _3998_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3396__A1 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5717_ _6878_/Q _5667_/X _5714_/X _5716_/X VGND VGND VPWR VPWR _5718_/C sky130_fd_sc_hd__a211o_1
XANTENNA__3396__B2 _7099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _6736_/CLK _6697_/D fanout436/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3940_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5648_ _6490_/Q _5643_/A _5647_/Y VGND VGND VPWR VPWR _6167_/S sky130_fd_sc_hd__a21o_4
XANTENNA__6334__A1 _6588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5579_ hold854/X _5579_/A1 _5586_/S VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3699__A2 _5226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold240 hold240/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold251 hold251/A VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold273 hold273/A VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6098__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold284 hold284/A VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold295 hold295/A VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1610_A _6481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5845__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input126_A wb_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6270__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6022__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input91_A spimemio_flash_io3_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3387__A1 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5533__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5836__B1 _6843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6984__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6913__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3988__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6261__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4950_ _4955_/A _4955_/B _4955_/C _4955_/D _4949_/Y VGND VGND VPWR VPWR _4950_/X
+ sky130_fd_sc_hd__a41o_1
X_3901_ _3921_/B VGND VGND VPWR VPWR _3901_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4972_/B sky130_fd_sc_hd__and2_1
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6620_ _6756_/CLK _6620_/D fanout441/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3832_ _3832_/A _3840_/B VGND VGND VPWR VPWR _3833_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6781__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3378__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6551_ _6753_/CLK _6551_/D fanout440/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3378__B2 input33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3763_ _6941_/Q _5362_/A _3509_/Y _6727_/Q _3762_/X VGND VGND VPWR VPWR _3769_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_146_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5502_ _5502_/A0 _5583_/A1 _5505_/S VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6482_ _6486_/CLK _6482_/D fanout434/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3694_ _3694_/A _3694_/B _3694_/C _3694_/D VGND VGND VPWR VPWR _3704_/B sky130_fd_sc_hd__nor4_1
XFILLER_118_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5433_ _5433_/A0 _5568_/A1 _5433_/S VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput301 _3745_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
Xoutput312 _7233_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2725_A _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput323 hold1711/X VGND VGND VPWR VPWR hold437/A sky130_fd_sc_hd__buf_6
Xoutput334 hold1966/X VGND VGND VPWR VPWR hold489/A sky130_fd_sc_hd__buf_6
X_5364_ hold206/X _5580_/A1 _5370_/S VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput345 hold1706/X VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__buf_6
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7135_/CLK _7103_/D fanout470/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_4
X_4315_ _4315_/A0 _5189_/A1 _4315_/S VGND VGND VPWR VPWR _4315_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5443__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5295_ _5295_/A0 _5448_/A1 _5298_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5827__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7034_ _7139_/CLK _7034_/D fanout471/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4246_ _4246_/A0 _5529_/A1 _4249_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4177_ _4177_/A0 _5543_/A1 _4181_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout376_A _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6252__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6818_ _7137_/CLK _6818_/D fanout466/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3369__A1 _7004_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3369__B2 input19/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6749_ _6760_/CLK _6749_/D fanout441/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4030__A2 _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4014__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6307__A1 _6592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4869__B2 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5353__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5818__B1 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5294__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6243__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7183__RESET_B fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7112__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3780__B2 _6804_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5263__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5809__B1 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4100_ _3737_/Y hold984/A _4106_/S VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__mux2_1
X_5080_ _5080_/A _5080_/B _5080_/C VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__and3_1
XANTENNA__5285__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1709 _6542_/Q VGND VGND VPWR VPWR hold976/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4031_ hold718/X _5579_/A1 _4056_/C VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4607__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6234__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5982_ _6014_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__and3_4
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3599__A1 _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4933_ _4374_/Y _5127_/A _4933_/C VGND VGND VPWR VPWR _5044_/C sky130_fd_sc_hd__and3b_1
XANTENNA__3599__B2 _6528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _5049_/B _4913_/A _4928_/C _4864_/D VGND VGND VPWR VPWR _4864_/X sky130_fd_sc_hd__and4_1
XFILLER_178_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _5085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _7045_/CLK _6603_/D fanout444/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_24 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3815_ _6657_/Q _3903_/A VGND VGND VPWR VPWR _3840_/B sky130_fd_sc_hd__nand2_4
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_35 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4464_/Y _4570_/D _4713_/Y _4947_/A VGND VGND VPWR VPWR _4796_/C sky130_fd_sc_hd__o22a_1
XANTENNA_57 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3239__A _6840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_68 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _6817_/CLK _6534_/D fanout435/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfstp_4
X_3746_ _6981_/Q _5407_/A hold89/A _6712_/Q VGND VGND VPWR VPWR _3746_/X sky130_fd_sc_hd__a22o_1
XANTENNA_79 hold191/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6465_ _3547_/A1 _6465_/D _6415_/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_2
XFILLER_173_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3677_ _3676_/X _3677_/A1 _3739_/S VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__mux2_1
X_5416_ _5416_/A _5578_/B VGND VGND VPWR VPWR _5424_/S sky130_fd_sc_hd__and2_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6396_ _6399_/A _6430_/B VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__and2_1
XANTENNA__6835__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5347_ _5347_/A0 _5572_/A1 _5352_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
Xoutput175 _3948_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _3947_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
XFILLER_142_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2900 _6680_/Q VGND VGND VPWR VPWR _3188_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xoutput197 _3237_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
Xhold2911 _7179_/Q VGND VGND VPWR VPWR _6216_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2922 _6435_/Q VGND VGND VPWR VPWR _3927_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5278_ _5278_/A0 _5575_/A1 _5280_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
Xhold2933 _7141_/Q VGND VGND VPWR VPWR _5588_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5276__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2944 _3902_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2955 _6468_/Q VGND VGND VPWR VPWR _3814_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7017_ _7017_/CLK _7017_/D fanout461/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
X_4229_ _5239_/A0 _5527_/A1 _5236_/C VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
Xhold2966 _5606_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2977 _7116_/Q VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5028__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1775_A _6907_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3762__A1 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A mgmt_gpio_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5267__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout380 hold95/X VGND VGND VPWR VPWR _5529_/A1 sky130_fd_sc_hd__buf_12
Xfanout391 _5536_/A1 VGND VGND VPWR VPWR _5572_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5303__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5019__B2 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4778__B1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__B1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3600_ _6798_/Q _3319_/Y _4000_/A _6482_/Q VGND VGND VPWR VPWR _3600_/X sky130_fd_sc_hd__a22o_4
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_2
X_4580_ _4580_/A _4607_/B VGND VGND VPWR VPWR _4580_/Y sky130_fd_sc_hd__nand2_2
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5742__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_4
X_3531_ _3553_/A hold88/X VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__nor2_4
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7233_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_171_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold806 hold806/A VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3962_/B sky130_fd_sc_hd__buf_4
Xhold828 hold828/A VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4637_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_170_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold839 hold839/A VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6250_ _6743_/Q _6014_/X _6244_/X _6249_/X VGND VGND VPWR VPWR _6255_/A sky130_fd_sc_hd__a211o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3462_ _3462_/A _3462_/B VGND VGND VPWR VPWR _3462_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__6089__B _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5201_ _5201_/A0 _5237_/A1 _5201_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6181_ _6979_/Q _5976_/B _5977_/X _7139_/Q _6180_/X VGND VGND VPWR VPWR _6181_/X
+ sky130_fd_sc_hd__a221o_1
X_3393_ _7131_/Q _5569_/A _5236_/C input69/X VGND VGND VPWR VPWR _3393_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2207 _6845_/Q VGND VGND VPWR VPWR hold739/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5132_ _4947_/B _4510_/B _4570_/A VGND VGND VPWR VPWR _5132_/X sky130_fd_sc_hd__a21o_1
Xhold2218 _7042_/Q VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2229 hold574/X VGND VGND VPWR VPWR _4294_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5258__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1506 hold342/X VGND VGND VPWR VPWR _5460_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1517 _6851_/Q VGND VGND VPWR VPWR hold299/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5063_ _5063_/A _5063_/B _5063_/C _5063_/D VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__and4_1
Xhold1528 _7067_/Q VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1539 hold288/X VGND VGND VPWR VPWR _5540_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4014_ hold754/X _5579_/A1 _4047_/C VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6207__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4056__C _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5965_ _6736_/Q _5656_/X _5679_/X _6593_/Q _5964_/X VGND VGND VPWR VPWR _5965_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5430__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4916_ _4969_/A _4652_/Y _4676_/Y _4633_/B VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__o22a_1
XFILLER_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5896_ _6698_/Q _5672_/X _5679_/X _6590_/Q _5883_/X VGND VGND VPWR VPWR _5896_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3441__B1 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3992__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _4638_/Y _4688_/B _5098_/A VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__o21a_1
XFILLER_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5733__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4778_ _4569_/B _4510_/B _4729_/A _4688_/A VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__o22a_1
XFILLER_181_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3729_ _6998_/Q _5425_/A _3536_/Y _6703_/Q VGND VGND VPWR VPWR _3729_/X sky130_fd_sc_hd__a22o_4
X_6517_ _6936_/CLK _6517_/D fanout472/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5184__A _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6448_ _3940_/A1 _6448_/D _6403_/X VGND VGND VPWR VPWR _6448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6379_ _6684_/Q _6379_/A2 _6379_/B1 _6685_/Q VGND VGND VPWR VPWR _6379_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5249__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2730 _5231_/X VGND VGND VPWR VPWR hold542/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2741 _7211_/A VGND VGND VPWR VPWR hold572/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2752 _6829_/Q VGND VGND VPWR VPWR hold908/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2763 _4242_/X VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2774 hold640/X VGND VGND VPWR VPWR _5333_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2785 hold949/X VGND VGND VPWR VPWR _5287_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2796 hold645/X VGND VGND VPWR VPWR _5423_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3680__B1 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4224__A2 _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3432__B1 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3983__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5724__A2 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output258_A _6793_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4160__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3671__B1 _4140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5412__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5750_ _5750_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5963__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4701_ _4701_/A _4701_/B VGND VGND VPWR VPWR _4826_/B sky130_fd_sc_hd__nor2_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5689_/A _5684_/B _5689_/C VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__and3_4
X_4632_ _4594_/A _4463_/B _4568_/Y _4837_/B _4631_/X VGND VGND VPWR VPWR _4632_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5715__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4563_ _4615_/B _4693_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 _4062_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2540_A _6788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6302_ _6607_/Q _5982_/X _5992_/X _6710_/Q VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4112__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3514_ _6913_/Q _5326_/A _5335_/A _6921_/Q _3513_/X VGND VGND VPWR VPWR _3515_/D
+ sky130_fd_sc_hd__a221o_1
Xhold614 hold614/A VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4494_ _4652_/B _4560_/A VGND VGND VPWR VPWR _4840_/A sky130_fd_sc_hd__and2b_2
Xhold636 hold636/A VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold647 hold647/A VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap355 hold56/X VGND VGND VPWR VPWR _3544_/A sky130_fd_sc_hd__buf_12
Xhold658 hold658/A VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6233_ _6712_/Q _5973_/X _5988_/X _6569_/Q _6232_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
Xhold669 hold669/A VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3445_ _7130_/Q _5569_/A _5353_/A _6938_/Q VGND VGND VPWR VPWR _3445_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6140__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7163__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3951__S _6820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4151__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _4129_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6164_ _6155_/X _6339_/B _6164_/C _6164_/D VGND VGND VPWR VPWR _6164_/X sky130_fd_sc_hd__and4b_4
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 hold717/X VGND VGND VPWR VPWR _4078_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3376_ _7116_/Q _5551_/A _3988_/A _6478_/Q VGND VGND VPWR VPWR _3376_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2026 hold796/X VGND VGND VPWR VPWR _4132_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5115_ _5115_/A _5115_/B _5124_/C _5126_/C VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__and4_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 hold511/X VGND VGND VPWR VPWR _4067_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1303 hold183/X VGND VGND VPWR VPWR _4282_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2048 _6893_/Q VGND VGND VPWR VPWR hold676/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2059 _4017_/X VGND VGND VPWR VPWR hold919/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _7056_/Q _5990_/X _5996_/X _7048_/Q VGND VGND VPWR VPWR _6095_/X sky130_fd_sc_hd__a22o_1
Xhold1314 hold303/X VGND VGND VPWR VPWR _5421_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4348__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 hold149/X VGND VGND VPWR VPWR _5275_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1336 _5364_/X VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1347 _3997_/X VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5046_ _5046_/A _5046_/B _5046_/C VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__and3_1
Xhold1358 hold236/X VGND VGND VPWR VPWR _5328_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1369 _6571_/Q VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3662__B1 _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6997_ _7137_/CLK _6997_/D fanout466/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5403__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5948_ _5969_/A1 _6342_/S _5946_/X _5947_/X VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__o22a_1
XANTENNA__3414__B1 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5954__A2 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5879_ _5879_/A _5879_/B _5879_/C _5879_/D VGND VGND VPWR VPWR _5879_/Y sky130_fd_sc_hd__nor4_1
XANTENNA_hold1473_A _6728_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5706__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3717__A1 _6728_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3717__B2 _6526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4022__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6131__A2 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4142__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input156_A wb_dat_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2560 hold663/X VGND VGND VPWR VPWR _5306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2571 _6804_/Q VGND VGND VPWR VPWR hold923/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2582 _5350_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2593 _5189_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1870 _6507_/Q VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1881 _5492_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input17_A mask_rev_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1892 _6634_/Q VGND VGND VPWR VPWR hold782/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6198__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5945__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A1 _3881_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6122__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4133__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3230_ _6920_/Q VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6920_ _6996_/CLK _6920_/D fanout462/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3644__B1 _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4987__A3 _4683_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6851_ _7082_/CLK _6851_/D fanout464/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _7002_/Q _5666_/X _5689_/X _7082_/Q VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__a22o_1
X_3994_ _3994_/A0 _7200_/Q _3998_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
X_6782_ _6826_/CLK _6782_/D _6407_/A VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5936__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3947__A1 _6436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5733_ _6999_/Q _5666_/X _5689_/X _7079_/Q _5732_/X VGND VGND VPWR VPWR _5733_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5664_ _5689_/A _5689_/B _5688_/C VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__and3_4
XFILLER_163_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6832_/CLK sky130_fd_sc_hd__clkbuf_16
X_4615_ _4625_/A _4615_/B VGND VGND VPWR VPWR _5063_/B sky130_fd_sc_hd__nand2_1
XFILLER_190_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5595_ _5595_/A0 _5593_/Y _5599_/D VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
Xhold400 hold400/A VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold411 hold411/A VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4546_ _4569_/A _4601_/A _4543_/X _4544_/Y _4898_/A VGND VGND VPWR VPWR _4546_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_191_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold422 hold422/A VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold433 hold433/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
Xhold444 hold444/A VGND VGND VPWR VPWR hold972/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4477_ _4477_/A _4477_/B _4477_/C VGND VGND VPWR VPWR _4477_/Y sky130_fd_sc_hd__nand3_4
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold477 hold477/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_116_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4124__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold488 hold488/A VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold499 hold499/A VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6216_ _6216_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_69_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6803_/CLK sky130_fd_sc_hd__clkbuf_16
X_3428_ _7172_/Q _6813_/Q _6815_/Q VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__mux2_8
X_7196_ _3950_/A1 _7196_/D _6346_/B VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A mask_rev_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6147_ _6994_/Q _6014_/X _6145_/X _6146_/X VGND VGND VPWR VPWR _6152_/A sky130_fd_sc_hd__a211o_1
Xhold1100 _4209_/X VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3359_ _6908_/Q _5317_/A _5461_/A _7036_/Q VGND VGND VPWR VPWR _3359_/X sky130_fd_sc_hd__a22o_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 hold189/X VGND VGND VPWR VPWR _4319_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 hold181/X VGND VGND VPWR VPWR _5266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_58_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1133 hold27/X VGND VGND VPWR VPWR _3255_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _6606_/Q VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6078_ _6959_/Q _5992_/X _6012_/X _6999_/Q _6077_/X VGND VGND VPWR VPWR _6078_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _4053_/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1166 _6911_/Q VGND VGND VPWR VPWR hold246/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5029_ _4417_/B _4648_/Y _4584_/Y VGND VGND VPWR VPWR _5029_/X sky130_fd_sc_hd__o21a_1
Xhold1177 _7071_/Q VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1188 _3996_/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _7007_/Q VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3635__B1 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5401__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4017__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5927__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6104__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2390 _6584_/Q VGND VGND VPWR VPWR hold898/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3626__B1 _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5311__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5091__A2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5918__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4170__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4400_ _4574_/A _4594_/A VGND VGND VPWR VPWR _4454_/A sky130_fd_sc_hd__nand2_8
X_5380_ _5380_/A _5578_/B VGND VGND VPWR VPWR _5388_/S sky130_fd_sc_hd__and2_4
XFILLER_160_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4331_ _4331_/A0 _5581_/A1 _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7050_ _7052_/CLK _7050_/D fanout464/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A _5220_/C VGND VGND VPWR VPWR _4267_/S sky130_fd_sc_hd__and2_2
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6001_ _6015_/B _6018_/B _6019_/C _6019_/A VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5854__A1 _7004_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3213_ _7048_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4193_ _4193_/A0 _5189_/A1 _4193_/S VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7201__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6903_ _7063_/CLK _6903_/D fanout460/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6834_ _7107_/CLK _6834_/D fanout451/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5909__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6031__A1 _7021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6765_ _7203_/CLK _6765_/D _4107_/B VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfrtp_1
X_3977_ _3977_/A _5220_/C VGND VGND VPWR VPWR _3987_/S sky130_fd_sc_hd__and2_2
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5716_ _6846_/Q _5653_/X _5682_/X _7038_/Q _5715_/X VGND VGND VPWR VPWR _5716_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3396__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5790__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6696_ _6760_/CLK _6696_/D _6407_/A VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _6490_/Q _5647_/B VGND VGND VPWR VPWR _5647_/Y sky130_fd_sc_hd__nor2_8
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6334__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ _5578_/A _5578_/B VGND VGND VPWR VPWR _5578_/X sky130_fd_sc_hd__and2_4
XANTENNA__7062__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3699__A3 _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 hold230/A VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold241 hold241/A VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4529_ _4396_/X _4529_/B _5151_/D _4529_/D VGND VGND VPWR VPWR _4529_/X sky130_fd_sc_hd__and4b_1
Xhold252 hold252/A VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold263 hold263/A VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__A1 _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6098__B2 _6944_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold274 hold274/A VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold285 hold285/A VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5845__B2 _7052_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7179_ _7179_/CLK _7179_/D fanout447/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6449__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__A _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3608__B1 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A wb_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1972_A _6877_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6022__A1 _6853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6022__B2 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input84_A spimemio_flash_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6325__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4336__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5306__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5836__B2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output240_A _3932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_2
XFILLER_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3900_ _4395_/A _3900_/B _3900_/C _3900_/D VGND VGND VPWR VPWR _3921_/B sky130_fd_sc_hd__nand4b_4
XFILLER_189_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _5127_/A _4880_/B VGND VGND VPWR VPWR _4965_/C sky130_fd_sc_hd__and2_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3831_ _3830_/Y _3831_/B _3835_/S VGND VGND VPWR VPWR _3833_/A sky130_fd_sc_hd__and3b_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3378__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6550_ _6753_/CLK _6550_/D fanout440/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_4
X_3762_ _7125_/Q _5569_/A _3536_/Y _6702_/Q VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5501_/A0 _5582_/A1 _5505_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
X_6481_ _6486_/CLK _6481_/D fanout434/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfstp_4
X_3693_ _7102_/Q _5542_/A _4140_/A _6590_/Q _3692_/X VGND VGND VPWR VPWR _3694_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4327__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5432_ _5432_/A0 _5567_/A1 _5433_/S VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput302 _3970_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_133_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput313 _7186_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
Xoutput324 hold1723/X VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__buf_6
X_5363_ hold900/X _5561_/A1 _5370_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
Xoutput335 hold1792/X VGND VGND VPWR VPWR hold481/A sky130_fd_sc_hd__buf_6
XFILLER_160_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7059__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _7134_/CLK _7102_/D fanout469/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfstp_4
X_4314_ _4314_/A0 _5195_/A1 _4315_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5294_ _5294_/A0 _5303_/A1 _5298_/S VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4245_ _4245_/A0 _5582_/A1 _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
X_7033_ _7134_/CLK _7033_/D fanout469/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4176_ _4176_/A hold9/A VGND VGND VPWR VPWR _4181_/S sky130_fd_sc_hd__and2_2
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5055__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6252__B2 _6531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6623__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6817_ _6817_/CLK _6817_/D fanout436/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1386_A _6840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3369__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6748_ _6753_/CLK _6748_/D fanout440/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfrtp_4
Xwire429 _4592_/B VGND VGND VPWR VPWR _4638_/A sky130_fd_sc_hd__buf_12
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6679_ _7203_/CLK _6679_/D _4107_/B VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6307__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4318__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4869__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3541__A2 _3319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5818__A1 _7003_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5818__B2 _6875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmgmt_gpio_14_buff_inst _3950_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
XFILLER_19_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5754__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output288_A _6488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4309__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3780__A2 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3532__A2 _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5809__A1 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5809__B2 _6986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5560__A _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4030_ _3343_/A _6430_/B _4012_/X _4056_/C _5317_/B VGND VGND VPWR VPWR _4046_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_23_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5981_ _7153_/Q _7154_/Q VGND VGND VPWR VPWR _6016_/C sky130_fd_sc_hd__and2b_4
XFILLER_52_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3599__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4932_ _4925_/X _4931_/X _5115_/A VGND VGND VPWR VPWR _4932_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4655_/A _4640_/Y _4655_/B _4704_/C VGND VGND VPWR VPWR _4864_/D sky130_fd_sc_hd__o31a_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6602_ _7045_/CLK _6602_/D fanout444/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_14 _5760_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4115__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4548__A1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _6114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _3814_/A _3814_/B VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__5745__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4729_/A _4712_/Y _4789_/X _4793_/X _5095_/A VGND VGND VPWR VPWR _4796_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_47 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_58 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _6736_/CLK _6533_/D fanout436/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_69 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _3745_/A VGND VGND VPWR VPWR _3745_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3771__A2 _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6464_ _3547_/A1 _6464_/D _6414_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfrtp_1
X_3676_ _3739_/A1 _3675_/Y _3738_/S VGND VGND VPWR VPWR _3676_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ _5415_/A0 _5568_/A1 _5415_/S VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6170__B1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6395_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__and2_1
X_5346_ _5346_/A0 _5562_/A1 _5352_/S VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput176 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
Xhold2901 _3922_/Y VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2912 _7185_/Q VGND VGND VPWR VPWR _6342_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5277_ _5277_/A0 _5277_/A1 _5280_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
Xhold2923 _3927_/Y VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2934 _5588_/X VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2945 _6459_/Q VGND VGND VPWR VPWR _3850_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7016_ _7128_/CLK _7016_/D fanout468/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_4
X_4228_ _4228_/A0 _4227_/X _4240_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
Xhold2956 _6448_/Q VGND VGND VPWR VPWR _3860_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2967 _6455_/Q VGND VGND VPWR VPWR _3856_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2978 _7073_/Q VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4159_ _4159_/A0 _5561_/A1 _4163_/S VGND VGND VPWR VPWR _4159_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5028__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4593__A_N _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4025__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5736__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3762__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6161__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3514__A2 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A mgmt_gpio_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5380__A _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout370 hold1189/X VGND VGND VPWR VPWR hold1190/A sky130_fd_sc_hd__clkbuf_2
Xfanout381 hold1044/X VGND VGND VPWR VPWR hold1045/A sky130_fd_sc_hd__buf_6
XFILLER_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout392 _5536_/A1 VGND VGND VPWR VPWR _5563_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output203_A _3935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4724__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4778__B2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__A_N _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__B2 _3428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3753__A2 _5226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3530_ hold88/X _3535_/A VGND VGND VPWR VPWR _4194_/A sky130_fd_sc_hd__nor2_8
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3881_/C sky130_fd_sc_hd__buf_8
Xhold807 hold807/A VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_2
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_2
Xhold818 hold818/A VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _3461_/A _3461_/B _3461_/C VGND VGND VPWR VPWR _3462_/B sky130_fd_sc_hd__and3_2
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5200_ _5207_/A hold47/X _5569_/B VGND VGND VPWR VPWR _5201_/S sky130_fd_sc_hd__and3_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3392_ _7185_/Q _6814_/Q _6815_/Q VGND VGND VPWR VPWR _3392_/X sky130_fd_sc_hd__mux2_8
X_6180_ _6931_/Q _5982_/X _6004_/X _6883_/Q VGND VGND VPWR VPWR _6180_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5131_ _5131_/A _5131_/B _5131_/C VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__and3_1
Xhold2208 hold739/X VGND VGND VPWR VPWR _5255_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2219 hold601/X VGND VGND VPWR VPWR _5476_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5290__A _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1507 _5460_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5062_ _5062_/A VGND VGND VPWR VPWR _5135_/B sky130_fd_sc_hd__inv_2
Xhold1518 hold299/X VGND VGND VPWR VPWR _5261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1529 hold310/X VGND VGND VPWR VPWR _5504_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4013_ _3648_/A _6430_/B _4012_/X _3330_/Y _5317_/B VGND VGND VPWR VPWR _4029_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3949__S _6819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4634__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4769__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5964_ _6643_/Q _5655_/X _5663_/X _6633_/Q _5950_/Y VGND VGND VPWR VPWR _5964_/X
+ sky130_fd_sc_hd__a221o_1
X_4915_ _5048_/A _4915_/B VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__nand2_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5895_ _6640_/Q _5655_/X _5656_/X _6733_/Q _5885_/Y VGND VGND VPWR VPWR _5895_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3441__B2 _6794_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ _4570_/C _4655_/A _4590_/Y _4691_/Y VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5194__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4777_ _4947_/A _4668_/Y _4531_/B VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6516_ _7125_/CLK hold85/X fanout468/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4941__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3728_ _6886_/Q _5299_/A _5497_/A _7062_/Q _3727_/X VGND VGND VPWR VPWR _3735_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5184__B _5184_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6143__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6447_ _3940_/A1 _6447_/D _6402_/X VGND VGND VPWR VPWR _6447_/Q sky130_fd_sc_hd__dfrtp_1
X_3659_ _7079_/Q _5515_/A _5560_/A _7119_/Q _3658_/X VGND VGND VPWR VPWR _3664_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6378_ _6377_/X _6378_/A1 _6384_/S VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5329_ _5329_/A0 _5572_/A1 _5334_/S VGND VGND VPWR VPWR _5329_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5404__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2720 _5386_/X VGND VGND VPWR VPWR hold624/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2731 _6789_/Q VGND VGND VPWR VPWR hold842/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2742 hold572/X VGND VGND VPWR VPWR _4240_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2753 hold908/X VGND VGND VPWR VPWR _5237_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2764 _6961_/Q VGND VGND VPWR VPWR hold809/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2775 _7019_/Q VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2786 _5287_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2797 _5423_/X VGND VGND VPWR VPWR hold646/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5957__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input101_A wb_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5185__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6134__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5314__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3671__A1 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3671__B2 _6591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3423__A1 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4700_ _4718_/C _4700_/B VGND VGND VPWR VPWR _4701_/B sky130_fd_sc_hd__nand2_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2199_A _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5689_/A _5684_/B _5689_/C VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__and3b_4
XFILLER_148_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4757_/A _4997_/A _4973_/C _4631_/D VGND VGND VPWR VPWR _4631_/X sky130_fd_sc_hd__and4_1
XFILLER_147_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5176__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6744__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4923__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4562_ _4562_/A _4693_/B VGND VGND VPWR VPWR _4894_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold604 hold604/A VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6301_ _6755_/Q _5638_/X _6019_/X _6735_/Q _6300_/X VGND VGND VPWR VPWR _6304_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold615 hold615/A VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3513_ _7017_/Q _5443_/A _4212_/A _6653_/Q VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold626 hold626/A VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6125__B1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4493_ _4649_/B _4639_/S VGND VGND VPWR VPWR _4652_/B sky130_fd_sc_hd__xnor2_1
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold648 hold648/A VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap356 hold56/X VGND VGND VPWR VPWR _3346_/A sky130_fd_sc_hd__buf_12
X_6232_ _6707_/Q _5992_/X _6012_/X _6747_/Q _6231_/X VGND VGND VPWR VPWR _6232_/X
+ sky130_fd_sc_hd__a221o_1
Xhold659 hold659/A VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3444_ _3444_/A _3444_/B _3444_/C _3444_/D VGND VGND VPWR VPWR _3462_/A sky130_fd_sc_hd__nor4_4
XFILLER_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _6892_/Q _5299_/A hold31/A _7100_/Q _3374_/X VGND VGND VPWR VPWR _3384_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6163_ _6163_/A _6163_/B _6163_/C _6163_/D VGND VGND VPWR VPWR _6164_/D sky130_fd_sc_hd__nor4_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _6740_/Q VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _6609_/Q VGND VGND VPWR VPWR hold830/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2027 _4132_/X VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5114_ _5114_/A _5114_/B _5114_/C VGND VGND VPWR VPWR _5126_/C sky130_fd_sc_hd__and3_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _4067_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1304 _4282_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6912_/Q _5991_/X _6018_/X _6968_/Q VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__a22o_1
Xhold2049 hold676/X VGND VGND VPWR VPWR _5309_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1315 _5421_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _5275_/X VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1337 _6871_/Q VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1348 _6636_/Q VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5045_ _4569_/B _4523_/Y _4583_/B _4688_/A VGND VGND VPWR VPWR _5046_/C sky130_fd_sc_hd__o22a_1
Xhold1359 _5328_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3662__B2 _6581_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6996_ _6996_/CLK _6996_/D fanout462/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout449_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5947_ _5947_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__o21ba_1
XFILLER_41_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3414__A1 _6875_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5878_ _6732_/Q _5656_/X _5663_/X _6629_/Q _5877_/X VGND VGND VPWR VPWR _5879_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4829_ _4454_/A _4719_/Y _4821_/X _4828_/X _4922_/B VGND VGND VPWR VPWR _4834_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4914__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4678__B1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5890__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input149_A wb_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2550 _4324_/X VGND VGND VPWR VPWR hold555/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2561 _5306_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2572 hold923/X VGND VGND VPWR VPWR _5203_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2583 _6558_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2594 _7085_/Q VGND VGND VPWR VPWR hold928/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1860 _6508_/Q VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1871 hold500/X VGND VGND VPWR VPWR _4044_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1882 _6984_/Q VGND VGND VPWR VPWR hold806/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1893 hold782/X VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3653__A1 input13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3653__B2 input97/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4850__B1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4274__A _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3405__A1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5158__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5309__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4905__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3708__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output270_A _6791_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6107__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5330__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3644__A1 _7023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3644__B2 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6850_ _7124_/CLK _6850_/D fanout471/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ _7010_/Q _5686_/X _5796_/X _5800_/X VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5397__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6781_ _3958_/A1 _6781_/D _6433_/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtn_1
X_3993_ _3993_/A0 _5189_/A1 _3999_/S VGND VGND VPWR VPWR _3993_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5732_ _6991_/Q _5929_/B _5668_/X _7055_/Q _5731_/X VGND VGND VPWR VPWR _5732_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5663_ _5685_/A _5684_/B _5688_/C VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__and3_4
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2650_A _6772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4614_ _5073_/B _4614_/B _4614_/C _4614_/D VGND VGND VPWR VPWR _4614_/X sky130_fd_sc_hd__and4_1
X_5594_ _5599_/D _5594_/B VGND VGND VPWR VPWR _5601_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4545_ _4625_/B _4724_/C VGND VGND VPWR VPWR _4898_/A sky130_fd_sc_hd__nand2_1
Xhold412 hold412/A VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold423 hold423/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_144_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold434 hold434/A VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold445 hold445/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4476_ _4574_/A _4594_/A _4463_/B VGND VGND VPWR VPWR _4476_/X sky130_fd_sc_hd__a21o_2
Xhold456 hold456/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xhold467 hold467/A VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold478 hold478/A VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6215_ _6844_/Q _6339_/B _6214_/Y _6341_/S VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__o211a_1
Xhold489 hold489/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
X_3427_ _3648_/B _3533_/B VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__5321__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7195_ _3950_/A1 _7195_/D _4107_/B VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout399_A hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1047_A _6889_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6146_ _6906_/Q _5985_/X _5994_/X _7066_/Q _6144_/X VGND VGND VPWR VPWR _6146_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _7020_/Q _5443_/A _5506_/A _7076_/Q VGND VGND VPWR VPWR _3358_/X sky130_fd_sc_hd__a22o_1
Xhold1101 _6438_/Q VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6090__B1_N _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1112 _4319_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1123 _5266_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6077_ _6951_/Q _5997_/X _6004_/X _6879_/Q VGND VGND VPWR VPWR _6077_/X sky130_fd_sc_hd__a22o_1
Xhold1134 _3255_/Y VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 hold216/X VGND VGND VPWR VPWR _4161_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3289_ _3322_/B _3430_/A VGND VGND VPWR VPWR _3764_/A sky130_fd_sc_hd__nand2_8
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 hold40/X VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1167 hold246/X VGND VGND VPWR VPWR _5329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1178 hold218/X VGND VGND VPWR VPWR _5509_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5028_ _4417_/B _4688_/A _4800_/C _4898_/A VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__o211a_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 hold34/X VGND VGND VPWR VPWR hold1189/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7085__SET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5388__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _7107_/CLK _6979_/D fanout452/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3399__B1 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4060__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6337__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4541__B _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4033__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3872__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5312__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold990 hold990/A VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5863__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2380 _6509_/Q VGND VGND VPWR VPWR hold754/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2391 hold898/X VGND VGND VPWR VPWR _4135_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3626__A1 _3971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1690 _6689_/Q VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5379__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7153__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4051__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6328__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4330_ _4330_/A0 _5238_/A1 _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5303__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4261_ _4261_/A0 _5277_/A1 _4261_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2231_A _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6000_ _5637_/A _6014_/A _6019_/C _5984_/X _5998_/X VGND VGND VPWR VPWR _6000_/X
+ sky130_fd_sc_hd__a311o_1
X_3212_ _7056_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5854__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4192_ _4192_/A0 _5195_/A1 _4193_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5502__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3617__A1 _3616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4814__B1 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6902_ _7072_/CLK _6902_/D fanout460/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4290__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6833_ _7108_/CLK hold96/X fanout451/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6031__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6764_ _7203_/CLK _6764_/D _6346_/B VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfrtp_1
X_3976_ _6434_/Q _3976_/A1 _3998_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6829__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5715_ _6934_/Q _5659_/X _5672_/X _6950_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6319__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6695_ _6830_/CLK _6695_/D fanout454/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_4
X_5646_ _5646_/A1 _5643_/B _5645_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__a21o_1
XFILLER_163_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A0 _5577_/A1 _5577_/S VGND VGND VPWR VPWR _5577_/X sky130_fd_sc_hd__mux2_1
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4528_ _4947_/A _4426_/Y _4527_/X _4574_/A VGND VGND VPWR VPWR _4529_/D sky130_fd_sc_hd__o22a_1
Xhold231 hold231/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold242 hold242/A VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold253 hold253/A VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold264 hold264/A VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6098__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold275 hold275/A VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__buf_12
X_4459_ _4485_/B _4564_/C _4881_/A VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__and3_1
Xhold286 hold286/A VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold297 hold297/A VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5845__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7178_ _7179_/CLK _7178_/D fanout447/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6129_/A _6129_/B _6129_/C _6129_/D VGND VGND VPWR VPWR _6139_/B sky130_fd_sc_hd__nor4_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5412__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3608__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__B2 input14/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4028__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6270__A2 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4281__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6022__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input77_A ser_tx VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5322__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6261__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4272__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _6657_/Q _3834_/S VGND VGND VPWR VPWR _3830_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_68_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6735_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ _7085_/Q _5524_/A hold24/A _7141_/Q _3760_/X VGND VGND VPWR VPWR _3769_/A
+ sky130_fd_sc_hd__a221o_2
X_5500_ _5500_/A0 _5572_/A1 _5505_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6480_ _6486_/CLK _6480_/D fanout434/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3692_ _6645_/Q _4206_/A _4194_/A _6635_/Q VGND VGND VPWR VPWR _3692_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ _5431_/A0 _5584_/A1 _5433_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput303 _5643_/A VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold1822/X VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__buf_6
X_5362_ _5362_/A _5578_/B VGND VGND VPWR VPWR _5370_/S sky130_fd_sc_hd__and2_4
Xoutput325 hold1878/X VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__buf_6
Xoutput336 hold1864/X VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__buf_6
X_7101_ _7101_/CLK _7101_/D fanout450/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_1
X_4313_ _4313_/A0 _5194_/A1 _4315_/S VGND VGND VPWR VPWR _4313_/X sky130_fd_sc_hd__mux2_1
X_5293_ _5293_/A0 _5572_/A1 _5298_/S VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7032_ _7128_/CLK _7032_/D fanout468/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5827__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4244_ _4244_/A0 _5563_/A1 _4249_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7199__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4175_ _4175_/A0 _5448_/A1 _4175_/S VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5232__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6252__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4263__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _6816_/CLK _6816_/D fanout446/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout431_A _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6747_ _6753_/CLK _6747_/D fanout440/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_4
X_3959_ _6456_/Q _3959_/B VGND VGND VPWR VPWR _3959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6678_ _3950_/A1 _6678_/D _4107_/B VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5629_ _5629_/A1 _5631_/A _5628_/Y VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5818__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input131_A wb_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6243__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5754__A1 _7016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5754__B2 _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3765__B1 _5209_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5809__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5560__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7121__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5690__B1 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4176__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6234__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5980_ _6017_/B _6018_/B _6007_/C VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__and3_4
XANTENNA__4245__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _5123_/A _4931_/B _4931_/C _4931_/D VGND VGND VPWR VPWR _4931_/X sky130_fd_sc_hd__and4_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2396_A _7065_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4862_ _4638_/Y _4713_/Y _4622_/C VGND VGND VPWR VPWR _4870_/B sky130_fd_sc_hd__o21a_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6601_ _6701_/CLK _6601_/D fanout436/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3813_ _3811_/B _3813_/B VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__and2b_1
XANTENNA_15 _5792_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4548__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _6114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5745__B2 _7015_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4947_/A _4712_/Y _4776_/Y _4792_/X _4531_/B VGND VGND VPWR VPWR _4793_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _6817_/CLK _6532_/D fanout435/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3756__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_59 _3970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ _6457_/Q _6437_/Q _6808_/Q VGND VGND VPWR VPWR _3745_/A sky130_fd_sc_hd__nor3_2
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6463_ _3547_/A1 _6463_/D _6413_/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfrtp_1
X_3675_ _3675_/A _3675_/B _3675_/C VGND VGND VPWR VPWR _3675_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__3508__B1 _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5414_ _5414_/A0 _5567_/A1 _5415_/S VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6170__A1 _7099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6394_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__and2_1
XANTENNA__6170__B2 _6955_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5345_ _5345_/A0 _5534_/A1 _5352_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput177 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
Xhold2902 _6447_/Q VGND VGND VPWR VPWR _3867_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput199 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
Xhold2913 _7165_/Q VGND VGND VPWR VPWR _5817_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5276_ _5276_/A0 _5303_/A1 _5280_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2924 hold60/A VGND VGND VPWR VPWR _3838_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7015_ _7133_/CLK _7015_/D fanout468/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5470__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2935 _7145_/Q VGND VGND VPWR VPWR _3914_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_4227_ _5238_/A0 _5238_/A1 _4237_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
Xhold2946 _6446_/Q VGND VGND VPWR VPWR _3868_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2957 _6492_/Q VGND VGND VPWR VPWR _3916_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2968 _7148_/Q VGND VGND VPWR VPWR _5614_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2979 _7120_/Q VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4158_ _4158_/A hold9/X VGND VGND VPWR VPWR _4163_/S sky130_fd_sc_hd__and2_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6694__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6225__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4089_ _3462_/Y hold987/A _4091_/S VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4787__A2 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1496_A _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5736__B2 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1663_A _6724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4041__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6161__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5380__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout382 _5303_/A1 VGND VGND VPWR VPWR _5195_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout393 _5571_/A1 VGND VGND VPWR VPWR _5193_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4227__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3450__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_4
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3753__A3 _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3970_/A sky130_fd_sc_hd__buf_6
Xhold808 hold808/A VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold819 hold819/A VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 spi_enabled VGND VGND VPWR VPWR _3971_/B sky130_fd_sc_hd__buf_4
X_3460_ _3460_/A _3460_/B _3460_/C _3460_/D VGND VGND VPWR VPWR _3461_/C sky130_fd_sc_hd__nor4_1
X_3391_ hold23/X _3516_/B VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__nor2_8
XFILLER_170_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5130_ _5130_/A _5130_/B _5130_/C VGND VGND VPWR VPWR _5131_/C sky130_fd_sc_hd__and3_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2209 _6551_/Q VGND VGND VPWR VPWR hold828/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5290__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5061_ _5061_/A _5061_/B VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__nand2_2
Xhold1508 _6865_/Q VGND VGND VPWR VPWR hold461/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1519 _6948_/Q VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4012_ _6430_/B _4241_/A VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__and2b_2
XFILLER_77_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6207__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4915__A _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5510__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4769__A2 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5963_ _6691_/Q _5659_/X _5687_/X _6603_/Q VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5966__A1 _6701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4914_ _4633_/B _4688_/C _4871_/B _4898_/B VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__o211a_1
X_5894_ _6580_/Q _5688_/X _5887_/X _5888_/X _5893_/X VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3441__A2 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4845_ _4569_/C _4655_/A _4590_/Y _4688_/B VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2945_A _6459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6341__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _4776_/A _5081_/A VGND VGND VPWR VPWR _4776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6515_ _7125_/CLK _6515_/D fanout469/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_1
X_3727_ input72/X _3293_/Y _4009_/A _6488_/Q VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4941__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5184__C _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6446_ _3940_/A1 _6446_/D _6401_/X VGND VGND VPWR VPWR _6446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3658_ _6596_/Q _4146_/A _3536_/Y _6704_/Q VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6143__B2 _7018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6377_ _6686_/Q _6377_/A2 _6377_/B1 _6685_/Q _6376_/X VGND VGND VPWR VPWR _6377_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3589_ _6792_/Q _3427_/Y _3562_/Y input95/X VGND VGND VPWR VPWR _3589_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1244_A _6848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5328_ _5328_/A0 _5571_/A1 _5334_/S VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__mux2_1
Xhold2710 _6823_/Q VGND VGND VPWR VPWR hold708/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2721 _6830_/Q VGND VGND VPWR VPWR hold586/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2732 hold842/X VGND VGND VPWR VPWR _5185_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5259_ _5259_/A0 _5448_/A1 _5262_/S VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2743 _6706_/Q VGND VGND VPWR VPWR hold775/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2754 _6795_/Q VGND VGND VPWR VPWR hold773/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2765 hold809/X VGND VGND VPWR VPWR _5385_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2776 hold643/X VGND VGND VPWR VPWR _5450_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2787 _6827_/Q VGND VGND VPWR VPWR hold873/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2798 _6898_/Q VGND VGND VPWR VPWR hold944/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5420__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4209__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3680__A2 _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4544__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4036__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3432__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3875__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1153_ clkbuf_0__1153_/X VGND VGND VPWR VPWR _6351_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6134__A1 _7097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6134__B2 _7081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output313_A _7186_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5330__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3671__A2 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4454__B _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6070__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4976_/A _5067_/B _4754_/D _4630_/D VGND VGND VPWR VPWR _4631_/D sky130_fd_sc_hd__and4b_1
XANTENNA_hold2094_A _6531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4561_ _4598_/B _4607_/B _4881_/B _3967_/A VGND VGND VPWR VPWR _4561_/X sky130_fd_sc_hd__a31o_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4923__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6300_ _6700_/Q _5997_/X _6017_/X _6772_/Q VGND VGND VPWR VPWR _6300_/X sky130_fd_sc_hd__a22o_1
X_3512_ _3535_/A _3533_/B VGND VGND VPWR VPWR _4212_/A sky130_fd_sc_hd__nor2_8
Xhold605 hold605/A VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4492_ _4637_/B _4492_/B _4500_/B VGND VGND VPWR VPWR _4639_/S sky130_fd_sc_hd__and3_1
XFILLER_183_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold616 hold616/A VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold627 hold627/A VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold638 hold638/A VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _6697_/Q _5997_/X _6004_/X _6574_/Q VGND VGND VPWR VPWR _6231_/X sky130_fd_sc_hd__a22o_1
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3443_ _6874_/Q _5281_/A _5461_/A _7034_/Q _3438_/X VGND VGND VPWR VPWR _3444_/D
+ sky130_fd_sc_hd__a221o_2
XANTENNA__5505__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5884__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7138_/Q _5977_/X _5984_/X _7098_/Q _6161_/X VGND VGND VPWR VPWR _6163_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _7108_/Q _5542_/A _5515_/A _7084_/Q _3360_/X VGND VGND VPWR VPWR _3374_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 hold706/X VGND VGND VPWR VPWR _4314_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 hold830/X VGND VGND VPWR VPWR _4165_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5113_ _5123_/C _5113_/B VGND VGND VPWR VPWR _5113_/Y sky130_fd_sc_hd__nand2_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _6630_/Q VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2039 _6517_/Q VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6896_/Q _5989_/X _6013_/X _7080_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__a22o_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1305 _6880_/Q VGND VGND VPWR VPWR hold348/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1316 _6975_/Q VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1327 _6519_/Q VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5044_ _5044_/A _5044_/B _5044_/C VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__and3_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1338 hold122/X VGND VGND VPWR VPWR _5284_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1349 _4197_/X VGND VGND VPWR VPWR hold178/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5240__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3662__A2 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6995_ _7131_/CLK _6995_/D fanout452/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6061__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5946_ _6528_/Q _5678_/Y _5940_/X _5945_/X _6341_/S VGND VGND VPWR VPWR _5946_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3414__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6757_/Q _5664_/X _5679_/X _6589_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4828_ _4384_/A _4675_/A _4633_/B _4825_/X _4827_/X VGND VGND VPWR VPWR _4828_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4759_ _5139_/A _4759_/B _4759_/C _4759_/D VGND VGND VPWR VPWR _4759_/X sky130_fd_sc_hd__and4_1
XANTENNA__4914__A2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6429_ _6433_/A _6430_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_108_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4678__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5415__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4678__B2 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5875__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4539__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2540 _6788_/Q VGND VGND VPWR VPWR hold895/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2551 _6701_/Q VGND VGND VPWR VPWR hold893/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2562 _6613_/Q VGND VGND VPWR VPWR hold683/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2573 _5203_/X VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2584 hold979/X VGND VGND VPWR VPWR hold446/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2595 hold928/X VGND VGND VPWR VPWR _5525_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1850 _7194_/Q VGND VGND VPWR VPWR hold999/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1861 hold576/X VGND VGND VPWR VPWR _4046_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1872 _4044_/X VGND VGND VPWR VPWR hold501/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1883 hold806/X VGND VGND VPWR VPWR _5411_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3653__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1894 _4195_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4274__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6052__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3405__A2 _3392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5158__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4905__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6107__A1 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output263_A _6785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4669__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5325__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4669__B2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5866__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6947__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_8
XFILLER_94_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3644__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6043__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5800_ _7058_/Q _5668_/X _5684_/X _6930_/Q VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _3958_/A1 _6780_/D _6432_/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtn_1
X_3992_ _3992_/A0 _5195_/A1 _3999_/S VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__mux2_1
X_5731_ _6927_/Q _5684_/X _5686_/X _7007_/Q VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2476_A _6997_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5662_ _5685_/A _5684_/B _5688_/C VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__and3b_4
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4613_ _4570_/B _4523_/Y _4924_/A _5095_/B VGND VGND VPWR VPWR _4614_/D sky130_fd_sc_hd__o211a_1
X_5593_ _7142_/Q _5594_/B VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4544_ _4971_/A _4607_/B VGND VGND VPWR VPWR _4544_/Y sky130_fd_sc_hd__nand2_1
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4109__A0 _3737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold413 hold413/A VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold424 hold424/A VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold435 hold435/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold446 hold446/A VGND VGND VPWR VPWR hold980/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4475_ _4724_/C _4981_/A VGND VGND VPWR VPWR _5117_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5235__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold468 hold468/A VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6214_ _6195_/X _6214_/B _6214_/C VGND VGND VPWR VPWR _6214_/Y sky130_fd_sc_hd__nand3b_2
Xhold479 hold479/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
X_3426_ _3533_/B VGND VGND VPWR VPWR _5184_/B sky130_fd_sc_hd__inv_2
X_7194_ _7194_/CLK _7194_/D VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6145_ _7058_/Q _5990_/X _5996_/X _7050_/Q VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3764_/B _3550_/B VGND VGND VPWR VPWR _4000_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 hold4/X VGND VGND VPWR VPWR _3980_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1113 _6983_/Q VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _6550_/Q VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6076_ _6076_/A _6076_/B _6076_/C VGND VGND VPWR VPWR _6089_/C sky130_fd_sc_hd__nor3_1
X_3288_ _3429_/A hold46/X VGND VGND VPWR VPWR _3430_/A sky130_fd_sc_hd__and2_4
Xhold1135 hold28/X VGND VGND VPWR VPWR _3276_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 _4161_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6282__B1 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1157 _7015_/Q VGND VGND VPWR VPWR hold221/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5027_ _4947_/A _4995_/A _5034_/D _5034_/A _4509_/Y VGND VGND VPWR VPWR _5027_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1168 _5329_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout461_A fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1179 _5509_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3635__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6034__B1 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ _6994_/CLK _6978_/D fanout462/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3399__A1 _6955_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5929_ _6745_/Q _5929_/B VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__and2_1
XFILLER_167_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1576_A _7011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6337__A1 _6608_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3571__A1 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input161_A wb_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold980 hold980/A VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold991 hold991/A VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2370 hold729/X VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2381 hold754/X VGND VGND VPWR VPWR _4048_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input22_A mask_rev_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6273__B1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2392 _4135_/X VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3626__A2 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1680 _5322_/X VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1691 hold592/X VGND VGND VPWR VPWR _4253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6025__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6328__A1 _6701_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5839__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4260_ _4260_/A0 _5233_/A1 _4261_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3211_ _7064_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__6165__B1_N _6164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4191_ _4191_/A0 _5194_/A1 _4193_/S VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6394__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4814__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4814__B2 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6901_ _7017_/CLK _6901_/D fanout461/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfstp_4
X_6832_ _6832_/CLK _6832_/D fanout447/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6763_ _3950_/A1 _6763_/D _4107_/B VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dfrtp_1
X_3975_ _6686_/Q _3975_/B VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__and2_1
XFILLER_149_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5714_ _7030_/Q _5655_/X _5687_/X _6918_/Q VGND VGND VPWR VPWR _5714_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6694_ _6760_/CLK _6694_/D _6416_/A VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5790__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5645_ _7143_/Q _6492_/Q _5645_/C _7142_/Q VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__and4b_1
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5576_ _5576_/A0 wire371/X _5577_/S VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__mux2_1
Xhold210 hold210/A VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 hold221/A VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4527_ _4462_/Y _4477_/Y _4466_/A _4463_/B VGND VGND VPWR VPWR _4527_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold232 hold232/A VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold243 hold243/A VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold254 hold254/A VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1157_A _7015_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold276 hold276/A VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4458_ _4485_/B _4881_/A VGND VGND VPWR VPWR _4491_/B sky130_fd_sc_hd__and2_2
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold287 hold287/A VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold298 _5215_/X VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3409_ _7091_/Q _5524_/A _5434_/A _7011_/Q _3408_/X VGND VGND VPWR VPWR _3409_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7177_ _7185_/CLK _7177_/D fanout447/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_1
X_4389_ _4447_/B _4663_/D _4917_/A _4701_/A VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__nor4_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _6961_/Q _5992_/X _5999_/X _6865_/Q _6127_/X VGND VGND VPWR VPWR _6129_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6974_/Q _5976_/B _5980_/X _6934_/Q VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__a22o_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3608__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4044__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1958_A _7080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5781__A2 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5297__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7101__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6246__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3480__B1 _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5221__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3760_ _7077_/Q _5515_/A _3336_/Y input20/X VGND VGND VPWR VPWR _3760_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _6790_/Q _3427_/Y _4170_/A _6615_/Q _3690_/X VGND VGND VPWR VPWR _3694_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5430_ _5430_/A0 _5583_/A1 _5433_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput304 _3428_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
X_5361_ _5361_/A0 _5568_/A1 _5361_/S VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__mux2_1
Xoutput315 hold1762/X VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__buf_6
XFILLER_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput326 hold1840/X VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__buf_6
Xoutput337 hold1807/X VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__buf_6
X_4312_ _4312_/A0 _5193_/A1 _4315_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7126_/CLK _7100_/D fanout453/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5292_ _5292_/A0 _5562_/A1 _5298_/S VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5288__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7031_ _7073_/CLK _7031_/D fanout445/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_4
X_4243_ _4243_/A0 _5580_/A1 _4249_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5513__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4174_ _4174_/A0 hold43/X _4175_/S VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6237__B1 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5460__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2975_A _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3471__B1 _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _6815_/CLK hold25/X fanout446/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5212__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6746_ _6746_/CLK _6746_/D _6416_/A VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_4
X_3958_ input83/X _3958_/A1 _6456_/Q VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3774__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _4720_/C _4649_/B VGND VGND VPWR VPWR _4394_/A sky130_fd_sc_hd__and2_1
XFILLER_167_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6677_ _7203_/CLK _6677_/D _4107_/B VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5628_ _7153_/Q _5611_/Y _5631_/A VGND VGND VPWR VPWR _5628_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5559_ hold81/X hold71/X _5559_/S VGND VGND VPWR VPWR _5559_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5279__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7229_ _7229_/A VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__7143__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5423__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4547__B _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6228__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4039__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4047__A_N _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input124_A wb_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3878__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5451__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5203__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4557__A3 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5754__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3765__A1 input11/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4190__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5333__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6219__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5442__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5569__A _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _4930_/A _5049_/C _4930_/C _4930_/D VGND VGND VPWR VPWR _4931_/D sky130_fd_sc_hd__and4_1
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3453__B1 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ _4569_/C _4655_/A _4590_/Y _4714_/Y VGND VGND VPWR VPWR _4871_/C sky130_fd_sc_hd__o22a_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6600_ _7045_/CLK _6600_/D fanout444/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_4
X_3812_ _3181_/Y _3814_/B _3879_/A VGND VGND VPWR VPWR _3813_/B sky130_fd_sc_hd__o21ai_1
X_4792_ _4462_/Y _4464_/Y _4466_/A _4790_/X _4791_/X VGND VGND VPWR VPWR _4792_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA_16 _5808_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5745__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _6189_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_49 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6531_ _6817_/CLK _6531_/D fanout435/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_4
X_3743_ _6997_/Q _5425_/A _4092_/A _6548_/Q _3742_/X VGND VGND VPWR VPWR _3750_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5508__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3674_ _3674_/A _3674_/B _3674_/C _3674_/D VGND VGND VPWR VPWR _3675_/C sky130_fd_sc_hd__and4_1
X_6462_ _3547_/A1 _6462_/D _6412_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3508__A1 _7097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5413_ _5413_/A0 _5584_/A1 _5415_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6393_ _6399_/A _6423_/B VGND VGND VPWR VPWR _6393_/X sky130_fd_sc_hd__and2_1
XANTENNA__5902__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7166__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6170__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5344_ _5344_/A _5533_/B VGND VGND VPWR VPWR _5352_/S sky130_fd_sc_hd__and2_4
XANTENNA__4181__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput178 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5275_/A0 _5572_/A1 _5280_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2903 _3867_/X VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2914 _7183_/Q VGND VGND VPWR VPWR _6292_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5243__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2925 _3838_/X VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7014_ _7086_/CLK _7014_/D fanout467/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfstp_4
X_4226_ _4226_/A0 _4225_/X _4240_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
Xhold2936 _5603_/Y VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2947 _3869_/Y VGND VGND VPWR VPWR _6446_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2958 _6445_/Q VGND VGND VPWR VPWR _3870_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2969 _6461_/Q VGND VGND VPWR VPWR _3839_/C1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4157_ _4157_/A0 _5277_/A1 _4157_/S VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3692__B1 _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4088_ _6351_/A0 _4088_/A1 _4091_/S VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5433__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3995__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5736__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3747__A1 _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6729_ _6730_/CLK _6729_/D _6411_/A VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_183_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5418__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7108_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6161__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1823_A _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4172__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7045_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout372 _5584_/A1 VGND VGND VPWR VPWR _5575_/A1 sky130_fd_sc_hd__buf_8
Xfanout383 _5303_/A1 VGND VGND VPWR VPWR _5233_/A1 sky130_fd_sc_hd__buf_6
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout394 _5571_/A1 VGND VGND VPWR VPWR _5238_/A1 sky130_fd_sc_hd__buf_8
XFILLER_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3683__B1 _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5424__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5389__A _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_62_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__B1 _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4724__C _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3738__A1 _3737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output293_A _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5328__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_2
XFILLER_167_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4232__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3972_/A sky130_fd_sc_hd__clkbuf_8
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _3879_/B sky130_fd_sc_hd__buf_12
XFILLER_182_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold809 hold809/A VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4163__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3390_ hold14/X _3390_/B VGND VGND VPWR VPWR _3516_/B sky130_fd_sc_hd__nand2_8
XFILLER_170_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5060_ _5059_/X _5115_/A VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__and2b_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 hold461/X VGND VGND VPWR VPWR _5277_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4011_ hold270/X _5571_/A1 _4011_/S VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5415__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5299__A _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5962_ _6638_/Q _5671_/X _5960_/X _5961_/X VGND VGND VPWR VPWR _5962_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5966__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4913_ _4913_/A _4913_/B VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__and2_2
XFILLER_33_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5893_ _6549_/Q _5673_/X _5890_/X _5892_/X VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4844_ _4569_/B _4655_/A _4590_/Y _4688_/A VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__o22a_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3729__A1 _6998_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _4729_/A _4674_/Y _5063_/A VGND VGND VPWR VPWR _4796_/A sky130_fd_sc_hd__o21a_1
XANTENNA__5238__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6514_ _7134_/CLK _6514_/D fanout469/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3726_ _3726_/A _3726_/B VGND VGND VPWR VPWR _4009_/A sky130_fd_sc_hd__nor2_8
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6445_ _3940_/A1 _6445_/D _6400_/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_1
X_3657_ _7095_/Q hold31/A _4274_/A _6709_/Q _3656_/X VGND VGND VPWR VPWR _3664_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6143__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4154__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6376_ _6684_/Q _6376_/A2 _6376_/B1 _4218_/Y VGND VGND VPWR VPWR _6376_/X sky130_fd_sc_hd__a22o_1
X_3588_ _7016_/Q _5443_/A _3336_/Y input23/X _3564_/X VGND VGND VPWR VPWR _3595_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5327_ _5327_/A0 hold275/X _5334_/S VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2700 hold686/X VGND VGND VPWR VPWR _4321_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2711 hold708/X VGND VGND VPWR VPWR _5230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2722 hold586/X VGND VGND VPWR VPWR _5238_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2733 _5185_/X VGND VGND VPWR VPWR hold843/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5258_ _5258_/A0 _5537_/A1 _5262_/S VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__mux2_1
Xhold2744 _6950_/Q VGND VGND VPWR VPWR hold596/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2755 _5192_/X VGND VGND VPWR VPWR hold774/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7083__RESET_B fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2766 _6953_/Q VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4209_ _4209_/A0 _5581_/A1 _4211_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
X_5189_ _5189_/A0 _5189_/A1 _5190_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
Xhold2777 _5450_/X VGND VGND VPWR VPWR hold644/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2788 hold873/X VGND VGND VPWR VPWR _5234_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3665__B1 _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2799 hold944/X VGND VGND VPWR VPWR _5314_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5406__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3417__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5957__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4090__A0 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4841__A _4917_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4052__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6134__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4145__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input52_A mgmt_gpio_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4696__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4227__S _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3408__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6070__A1 _7055_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6070__B2 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4560_ _4560_/A _4560_/B _4560_/C _4598_/C VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__and4_2
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3511_ _7129_/Q _5569_/A _5380_/A _6961_/Q _3510_/X VGND VGND VPWR VPWR _3515_/C
+ sky130_fd_sc_hd__a221o_1
Xhold606 hold606/A VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4491_ _4598_/C _4491_/B VGND VGND VPWR VPWR _4491_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__6125__A2 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold617 hold617/A VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4136__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold628 hold628/A VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6230_ _6230_/A _6230_/B _6230_/C VGND VGND VPWR VPWR _6239_/C sky130_fd_sc_hd__nor3_1
Xhold639 hold639/A VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3442_ _7002_/Q _5425_/A _5380_/A _6962_/Q _3441_/X VGND VGND VPWR VPWR _3444_/C
+ sky130_fd_sc_hd__a221o_1
Xmax_cap347 _4237_/S VGND VGND VPWR VPWR _5236_/C sky130_fd_sc_hd__buf_12
Xmax_cap358 _3349_/A VGND VGND VPWR VPWR _3347_/A sky130_fd_sc_hd__buf_12
XANTENNA__6397__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5884__A1 _6605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _6844_/Q _5245_/A _5236_/C _3973_/B _3372_/X VGND VGND VPWR VPWR _3384_/A
+ sky130_fd_sc_hd__a221o_1
X_6161_ _6930_/Q _5982_/X _5987_/X _7114_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _4314_/X VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 _4165_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VGND VPWR VPWR _5113_/B sky130_fd_sc_hd__and4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6116_/A0 _6091_/X _6342_/S VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__mux2_1
Xhold2029 hold525/X VGND VGND VPWR VPWR _4190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7204__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 hold348/X VGND VGND VPWR VPWR _5294_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1317 hold143/X VGND VGND VPWR VPWR _5401_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5043_ _5043_/A _5043_/B VGND VGND VPWR VPWR _5043_/Y sky130_fd_sc_hd__nand2_1
Xhold1328 hold191/X VGND VGND VPWR VPWR _4059_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3647__B1 _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1339 _5284_/X VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5521__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_wbbd_sck _7203_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5939__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6994_ _6994_/CLK _6994_/D fanout462/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__6061__A1 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6061__B2 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5945_ _6700_/Q _5672_/X _5941_/X _5943_/X _5944_/X VGND VGND VPWR VPWR _5945_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_53_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3976__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6352__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6548_/Q _5673_/X _5682_/X _6450_/Q _5875_/X VGND VGND VPWR VPWR _5879_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4411_/Y _4701_/B _4812_/Y _4698_/Y _4928_/B VGND VGND VPWR VPWR _4827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4758_ _4986_/C _4837_/B _4965_/B _4757_/X _4716_/Y VGND VGND VPWR VPWR _4759_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3709_ _7070_/Q _5506_/A _5515_/A _7078_/Q _3708_/X VGND VGND VPWR VPWR _3716_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_10_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4689_ _4710_/A _4719_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__nand2_2
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4127__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6428_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_134_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6359_ _6685_/Q _6356_/Y _6357_/Y _6686_/Q _4836_/A VGND VGND VPWR VPWR _6359_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2530 _6528_/Q VGND VGND VPWR VPWR hold924/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2541 hold895/X VGND VGND VPWR VPWR _5183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2552 hold893/X VGND VGND VPWR VPWR _4267_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2563 hold683/X VGND VGND VPWR VPWR _4169_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5431__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3638__B1 _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2574 _6560_/Q VGND VGND VPWR VPWR hold981/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1840 hold474/X VGND VGND VPWR VPWR hold1840/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2585 _6979_/Q VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2596 _5525_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1851 hold999/X VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1862 _6563_/Q VGND VGND VPWR VPWR hold998/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1873 hold501/X VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1884 _5411_/X VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1895 _6539_/Q VGND VGND VPWR VPWR hold916/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6052__A1 _6894_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6052__B2 _7014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3886__S _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4366__A1 _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6107__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4118__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5341__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5094__A2 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6043__A1 _7086_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6043__B2 _6998_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ _3991_/A0 _5194_/A1 _3999_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5730_ _5750_/A1 _5729_/X _6342_/S VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4481__A _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5661_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5688_/C sky130_fd_sc_hd__and2b_4
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4612_ _4625_/A _4981_/A VGND VGND VPWR VPWR _5095_/B sky130_fd_sc_hd__nand2_1
X_5592_ _6341_/S _3911_/B _3197_/Y VGND VGND VPWR VPWR _5594_/B sky130_fd_sc_hd__o21a_1
X_4543_ _4464_/Y _4569_/C _4540_/X _5149_/A _4542_/Y VGND VGND VPWR VPWR _4543_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5516__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold403 hold403/A VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold414 hold414/A VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold425 hold425/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4474_ _4981_/A VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__clkinv_2
Xhold447 hold447/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xhold458 hold458/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_132_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6213_ _6206_/X _6208_/X _6213_/C _6313_/D VGND VGND VPWR VPWR _6214_/C sky130_fd_sc_hd__and4bb_1
Xhold469 hold469/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
X_3425_ hold14/X _3430_/B VGND VGND VPWR VPWR _3533_/B sky130_fd_sc_hd__nand2_8
X_7193_ _7194_/CLK _7193_/D VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6914_/Q _5991_/X _6018_/X _6970_/Q VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__a22o_1
X_3356_ _3356_/A _3550_/B VGND VGND VPWR VPWR _4237_/S sky130_fd_sc_hd__nor2_8
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1103 _3980_/X VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1114 hold179/X VGND VGND VPWR VPWR _5410_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6347__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _7031_/Q _5986_/X _5998_/X _6887_/Q _6074_/X VGND VGND VPWR VPWR _6076_/C
+ sky130_fd_sc_hd__a221o_1
X_3287_ _3563_/A _3354_/A VGND VGND VPWR VPWR _5569_/A sky130_fd_sc_hd__nor2_8
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 hold186/X VGND VGND VPWR VPWR _4095_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1136 _3279_/Y VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 _7055_/Q VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1158 hold221/X VGND VGND VPWR VPWR _5446_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5026_ _5150_/A _5026_/B _5026_/C VGND VGND VPWR VPWR _5034_/D sky130_fd_sc_hd__nand3_1
XANTENNA__6282__B2 _6641_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1169 _7111_/Q VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout454_A input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6034__A1 _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6034__B2 _6957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _6977_/CLK _6977_/D fanout461/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3399__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5928_ _3224_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5859_ _5859_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__6337__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5426__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3571__A2 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5848__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold970 hold970/A VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold981 hold981/A VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold992 hold992/A VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input154_A wb_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2360 hold728/X VGND VGND VPWR VPWR _5547_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2371 _6718_/Q VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6273__A1 _6596_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4423__A_N _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2382 _6687_/Q VGND VGND VPWR VPWR hold847/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6273__B2 _6699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2393 _7113_/Q VGND VGND VPWR VPWR hold724/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1670 hold308/X VGND VGND VPWR VPWR _5174_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input15_A mask_rev_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1681 _6794_/Q VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1692 _4253_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4036__A0 _4036_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5784__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6328__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4339__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5336__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4240__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3210_ _7072_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4190_ _4190_/A0 _5193_/A1 _4193_/S VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4814__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6900_ _6994_/CLK _6900_/D fanout462/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6831_ _6832_/CLK _6831_/D fanout447/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6762_ _3950_/A1 _6762_/D _4107_/B VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__dfrtp_1
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5775__B1 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3974_ _6822_/Q _3974_/B VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__and2_2
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5713_ _6894_/Q _5662_/X _5674_/X _6870_/Q _5712_/X VGND VGND VPWR VPWR _5718_/B
+ sky130_fd_sc_hd__a221o_1
X_6693_ _6826_/CLK _6693_/D _6407_/A VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6319__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5644_ _5644_/A1 _5643_/B _5643_/Y _6490_/Q VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ _5575_/A0 _5575_/A1 _5577_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
Xhold200 hold200/A VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold211 hold211/A VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4526_ _5009_/A _5001_/A _4751_/B VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__and3_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold244 hold244/A VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6288__D _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4457_ _4457_/A _4469_/B _4457_/C VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__and3_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold266 hold266/A VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold299 hold299/A VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3408_ _7083_/Q _5515_/A _5497_/A _7067_/Q VGND VGND VPWR VPWR _3408_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7176_ _7179_/CLK _7176_/D fanout446/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_1
X_4388_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4712_/A sky130_fd_sc_hd__nor2_8
XFILLER_58_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A mask_rev_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6127_ _6937_/Q _5980_/X _5982_/X _6929_/Q VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4386__A _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3764_/B _3563_/B VGND VGND VPWR VPWR _3988_/A sky130_fd_sc_hd__nor2_8
XFILLER_105_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6058_ _7062_/Q _5994_/X _5996_/X _7046_/Q _6057_/X VGND VGND VPWR VPWR _6058_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5009_/A _5009_/B VGND VGND VPWR VPWR _5009_/Y sky130_fd_sc_hd__nor2_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5929__B _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__B1 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4060__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5793__A1_N _5782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6965__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2190 _6735_/Q VGND VGND VPWR VPWR hold826/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3480__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3480__B2 _6608_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__S _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5757__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3690_ _6942_/Q _5362_/A _4286_/A _6718_/Q VGND VGND VPWR VPWR _3690_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6182__B1 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput305 _3392_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
X_5360_ _5360_/A0 _5549_/A1 _5361_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput316 hold1745/X VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_57_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput327 hold1714/X VGND VGND VPWR VPWR hold456/A sky130_fd_sc_hd__buf_6
Xoutput338 hold1852/X VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__buf_6
X_4311_ _4311_/A0 hold275/X _4315_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ hold668/X _5579_/A1 _5298_/S VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7030_ _7078_/CLK _7030_/D fanout445/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfstp_2
X_4242_ _4242_/A0 _5579_/A1 _4249_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4173_ hold145/X _5581_/A1 _4175_/S VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4799__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3471__B2 _6788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6814_ _6815_/CLK _6814_/D fanout446/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6745_ _6745_/CLK _6745_/D fanout441/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_2
X_3957_ _6457_/Q _3959_/B VGND VGND VPWR VPWR _3957_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3984__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3774__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6676_ _7203_/CLK _6676_/D _4107_/B VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3888_ _6455_/Q _6434_/Q _6423_/B VGND VGND VPWR VPWR _3975_/B sky130_fd_sc_hd__o21ai_1
X_5627_ _5647_/B _6019_/A _6017_/A _5605_/Y _5627_/B2 VGND VGND VPWR VPWR _7152_/D
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6173__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5558_ _5558_/A0 _5567_/A1 _5559_/S VGND VGND VPWR VPWR _5558_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5920__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4509_ _4980_/A _4607_/B VGND VGND VPWR VPWR _4509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5489_ hold892/X _5561_/A1 _5496_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7228_ _7228_/A VGND VGND VPWR VPWR _7228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7159_ _7180_/CLK _7159_/D fanout446/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1601_A _6527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A wb_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4055__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3765__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input82_A spi_sdoenb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5690__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5569__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4860_ _4638_/Y _4683_/A _4683_/B _4586_/Y VGND VGND VPWR VPWR _4872_/C sky130_fd_sc_hd__o31a_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3811_ _3811_/A _3811_/B VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__xor2_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4791_ _4791_/A _4791_/B _4791_/C _5034_/B VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__and4_1
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_17 _5836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_28 _6239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7130__RESET_B fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6817_/CLK _6530_/D fanout436/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3756__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3742_ _7053_/Q _5488_/A hold57/A _6569_/Q VGND VGND VPWR VPWR _3742_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6155__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6461_ _3547_/A1 _6461_/D _6411_/X VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_4
X_3673_ _3673_/A _3673_/B _3673_/C _3673_/D VGND VGND VPWR VPWR _3674_/D sky130_fd_sc_hd__nor4_1
X_5412_ _5412_/A0 _5583_/A1 _5415_/S VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3508__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6392_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__and2_1
X_5343_ _5343_/A0 _5568_/A1 _5343_/S VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _5274_/A0 _5571_/A1 _5280_/S VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2904 _7162_/Q VGND VGND VPWR VPWR _5751_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2915 _7198_/Q VGND VGND VPWR VPWR _6372_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7013_ _7101_/CLK _7013_/D fanout450/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_1
Xhold2926 hold77/A VGND VGND VPWR VPWR _4760_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4225_ _5237_/A0 _5237_/A1 _4237_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
Xhold2937 _7152_/Q VGND VGND VPWR VPWR _5627_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2948 _6437_/Q VGND VGND VPWR VPWR _3880_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2959 _6460_/Q VGND VGND VPWR VPWR _3270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4156_ _4156_/A0 _5195_/A1 _4157_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4087_ _3616_/Y hold969/A _4091_/S VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5479__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5197__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4989_ _5150_/B _4989_/B VGND VGND VPWR VPWR _4995_/B sky130_fd_sc_hd__nor2_4
XFILLER_51_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3747__A2 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6728_ _6731_/CLK _6728_/D _6411_/A VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4944__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4944__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6146__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6659_ _7203_/CLK _6659_/D _4107_/B VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3380__B1 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout351 _6313_/D VGND VGND VPWR VPWR _6339_/B sky130_fd_sc_hd__buf_12
Xfanout373 wire375/X VGND VGND VPWR VPWR _5584_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout384 hold43/X VGND VGND VPWR VPWR _5303_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_101_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3683__A1 input12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout395 _5228_/A1 VGND VGND VPWR VPWR _5571_/A1 sky130_fd_sc_hd__buf_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4574__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__B2 _6484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4935__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_4
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5360__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3371__B1 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4010_ _4010_/A0 _5534_/A1 _4011_/S VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4484__A _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5299__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ _6751_/Q _5666_/X _5689_/X _6628_/Q VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4912_ _4640_/Y _4648_/Y _4679_/Y _4564_/Y _4658_/B VGND VGND VPWR VPWR _4913_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5892_ _6610_/Q _5660_/X _5669_/X _6650_/Q _5891_/X VGND VGND VPWR VPWR _5892_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5179__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4843_ _4500_/Y _4652_/Y _4930_/A VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__o21a_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5519__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3729__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4926__A1 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4774_ _4947_/A _4688_/B _4536_/Y VGND VGND VPWR VPWR _4774_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _6828_/CLK _6513_/D fanout469/X VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3725_ _3725_/A _3725_/B _3725_/C _3725_/D VGND VGND VPWR VPWR _3736_/C sky130_fd_sc_hd__nor4_1
XANTENNA__6128__B1 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6444_ net399_2/A _6444_/D _6399_/X VGND VGND VPWR VPWR _6444_/Q sky130_fd_sc_hd__dfrtp_1
X_3656_ _7047_/Q hold16/A _3521_/Y _6537_/Q VGND VGND VPWR VPWR _3656_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5351__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6375_ _6374_/X _6375_/A1 _6384_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3616_/C sky130_fd_sc_hd__nor4_2
XANTENNA__3362__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5326_ _5326_/A _5569_/B VGND VGND VPWR VPWR _5334_/S sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_3_6__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4378__B _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2701 _4321_/X VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2712 _5230_/X VGND VGND VPWR VPWR hold709/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2723 _7098_/Q VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6300__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5257_ _5257_/A0 _5572_/A1 _5262_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
Xhold2734 _6767_/Q VGND VGND VPWR VPWR _5147_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2745 _6702_/Q VGND VGND VPWR VPWR hold759/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2756 _6691_/Q VGND VGND VPWR VPWR hold852/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4208_ _4208_/A0 _5238_/A1 _4211_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2767 hold791/X VGND VGND VPWR VPWR _5376_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5188_ _5188_/A0 _5195_/A1 _5190_/S VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__mux2_1
Xhold2778 _6931_/Q VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3665__B2 _6689_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2789 _5234_/X VGND VGND VPWR VPWR hold874/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4139_ _4139_/A0 _5189_/A1 _4139_/S VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5429__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6119__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5342__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5893__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A mgmt_gpio_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3656__A1 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4853__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7156__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6070__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4081__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4751__B _4751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5339__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5581__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3592__B1 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3510_ _7105_/Q _5542_/A _3509_/Y _6731_/Q VGND VGND VPWR VPWR _3510_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4490_ _4598_/C _4491_/B VGND VGND VPWR VPWR _4628_/A sky130_fd_sc_hd__and2_2
XFILLER_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold607 hold607/A VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold618 _5377_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5333__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3441_ _6914_/Q _5326_/A _3427_/Y _6794_/Q VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap348 _3330_/Y VGND VGND VPWR VPWR _4047_/C sky130_fd_sc_hd__buf_12
XFILLER_143_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5884__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ _6866_/Q _5999_/X _6019_/X _6986_/Q _6143_/X VGND VGND VPWR VPWR _6163_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _6486_/Q _4000_/A _3369_/X _3371_/X VGND VGND VPWR VPWR _3372_/X sky130_fd_sc_hd__a211o_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5111_ _4990_/B _4995_/A _4699_/Y _4924_/C _4924_/A VGND VGND VPWR VPWR _5112_/D
+ sky130_fd_sc_hd__o2111a_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _6757_/Q VGND VGND VPWR VPWR hold691/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _7174_/Q _6090_/X _6341_/S VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__mux2_1
Xhold2019 _6640_/Q VGND VGND VPWR VPWR hold524/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _6864_/Q VGND VGND VPWR VPWR hold381/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5042_ _5042_/A _5149_/B _5086_/A _5042_/D VGND VGND VPWR VPWR _5043_/B sky130_fd_sc_hd__and4_1
Xhold1318 _5401_/X VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 _7102_/Q VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3647__A1 input5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3647__B2 _6739_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4844__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6993_ _7063_/CLK _6993_/D fanout461/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_51_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7107_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold2783_A _6957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6061__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5944_ _6597_/Q _5670_/X _5685_/X _6772_/Q _5927_/X VGND VGND VPWR VPWR _5944_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4072__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6349__A0 _3675_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5875_ _6747_/Q _5666_/X _5685_/X _6769_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4826_ _4826_/A _4826_/B VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_66_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6701_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5572__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4757_ _4757_/A _4920_/B _4757_/C _4757_/D VGND VGND VPWR VPWR _4757_/X sky130_fd_sc_hd__and4_1
XFILLER_135_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3583__B1 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3708_ _7046_/Q hold16/A _5236_/C input47/X VGND VGND VPWR VPWR _3708_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4688_ _4688_/A _4688_/B _4688_/C VGND VGND VPWR VPWR _4688_/X sky130_fd_sc_hd__and3_1
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5324__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6427_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
X_3639_ input22/X _3336_/Y _4188_/A _6631_/Q VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a22o_4
XFILLER_161_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5875__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6358_ _6358_/A _6358_/B VGND VGND VPWR VPWR _6358_/Y sky130_fd_sc_hd__nand2_2
XFILLER_108_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ _5309_/A0 _5579_/A1 _5316_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6289_ _6270_/X _6289_/B _6289_/C VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__nand3b_4
Xhold2520 _5396_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2531 hold924/X VGND VGND VPWR VPWR _4069_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2542 _5183_/X VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2553 _4267_/X VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__A1 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2564 _4169_/X VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__B2 _6771_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2575 hold981/X VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1830 hold994/X VGND VGND VPWR VPWR hold486/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1841 _7216_/A VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2586 hold658/X VGND VGND VPWR VPWR _5405_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1852 hold470/X VGND VGND VPWR VPWR hold1852/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2597 _6635_/Q VGND VGND VPWR VPWR hold518/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1863 hold998/X VGND VGND VPWR VPWR hold492/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1874 _7213_/A VGND VGND VPWR VPWR hold582/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1885 _7188_/Q VGND VGND VPWR VPWR hold996/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1896 hold916/X VGND VGND VPWR VPWR _4082_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6730_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6052__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4063__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4063__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5012__B1 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5563__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3574__B1 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5315__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5866__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4238__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6043__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xnet399_2 net399_2/A VGND VGND VPWR VPWR _3954_/B sky130_fd_sc_hd__inv_2
XANTENNA__4054__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3990_ _3990_/A0 _5193_/A1 _3999_/S VGND VGND VPWR VPWR _3990_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5660_ _5689_/A _5676_/B _5686_/B VGND VGND VPWR VPWR _5660_/X sky130_fd_sc_hd__and3_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4611_/A _4693_/B VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5554__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5591_ _5599_/D VGND VGND VPWR VPWR _5591_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4542_ _4971_/A _4972_/A VGND VGND VPWR VPWR _4542_/Y sky130_fd_sc_hd__nand2_1
Xhold404 hold404/A VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5306__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4473_ _4485_/B _4598_/B _4564_/C VGND VGND VPWR VPWR _4981_/A sky130_fd_sc_hd__and3_4
Xhold437 hold437/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
Xhold448 hold448/A VGND VGND VPWR VPWR hold982/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5857__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6212_ _7044_/Q _6016_/X _6209_/X _6211_/X VGND VGND VPWR VPWR _6213_/C sky130_fd_sc_hd__a211oi_2
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3424_ _3423_/X _3424_/A1 _3739_/S VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7192_ _7194_/CLK _7192_/D VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _7090_/Q _5638_/X _6015_/X _7018_/Q VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3355_/A _3430_/B VGND VGND VPWR VPWR _3550_/B sky130_fd_sc_hd__nand2_8
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5532__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__1153_ _3558_/Y VGND VGND VPWR VPWR clkbuf_0__1153_/X sky130_fd_sc_hd__clkbuf_16
X_6074_ _6975_/Q _5976_/B _5993_/X _7007_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__a22o_1
Xhold1104 hold120/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1115 _5410_/X VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3309_/A _3322_/B VGND VGND VPWR VPWR _3354_/A sky130_fd_sc_hd__nand2_8
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _4095_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1137 _3521_/Y VGND VGND VPWR VPWR _4077_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5025_ _5015_/X _5024_/Y _5139_/A _5140_/A VGND VGND VPWR VPWR _5025_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6282__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1148 hold207/X VGND VGND VPWR VPWR _5491_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1159 _5446_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4293__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6034__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4045__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout447_A fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6976_ _6996_/CLK _6976_/D fanout463/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ _6538_/Q _5651_/X _5688_/X _6582_/Q VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5793__B2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1297_A _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5858_ _6844_/Q _5678_/Y _5849_/X _5857_/X _6166_/S VGND VGND VPWR VPWR _5858_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5545__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4809_ _4574_/A _4637_/D _4719_/Y _4691_/Y _4583_/B VGND VGND VPWR VPWR _4818_/A
+ sky130_fd_sc_hd__o32a_1
X_5789_ _6937_/Q _5659_/X _5663_/X _7025_/Q _5788_/X VGND VGND VPWR VPWR _5792_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_181_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5848__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold960 _5530_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold971 hold971/A VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold982 hold982/A VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold993 hold993/A VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5442__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input147_A wb_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2350 _6752_/Q VGND VGND VPWR VPWR hold862/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4566__B _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2361 _7054_/Q VGND VGND VPWR VPWR hold598/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2372 hold625/X VGND VGND VPWR VPWR _4288_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6273__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4058__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2383 hold847/X VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4284__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2394 hold724/X VGND VGND VPWR VPWR _5556_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1660 _7223_/A VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1671 _5174_/X VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1682 hold222/X VGND VGND VPWR VPWR _5190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1693 _6977_/Q VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6025__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5784__B2 _7073_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3795__B1 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6925__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5536__A1 _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3547__B1 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5839__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5352__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4275__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6830_ _6830_/CLK _6830_/D _6407_/A VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6761_ _6761_/CLK _6761_/D _6430_/A VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_4
X_3973_ _6821_/Q _3973_/B VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__and2_4
XANTENNA__5775__B2 _7065_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5712_ _7062_/Q _5671_/X _5689_/X _7078_/Q VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3786__B1 _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6692_ _6826_/CLK _6692_/D _6407_/A VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _5643_/A _5643_/B VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5527__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5527__S _5532_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3538__B1 _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ _5574_/A0 _5583_/A1 _5577_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold201 hold201/A VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4525_ _4625_/A _5033_/A VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__nand2_2
XFILLER_116_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold212 hold212/A VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold223 hold223/A VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold234 hold234/A VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold245 hold245/A VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4456_ _4450_/A _4450_/B _4451_/A VGND VGND VPWR VPWR _4564_/C sky130_fd_sc_hd__o21a_4
Xhold256 hold256/A VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold267 hold267/A VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold278 hold278/A VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3407_ _6867_/Q _5272_/A _5344_/A _6931_/Q VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__a22o_1
Xhold289 hold289/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7175_ _7179_/CLK _7175_/D fanout443/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4387_ _4921_/A _4886_/A VGND VGND VPWR VPWR _4387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout397_A _5228_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3710__B1 _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6126_ _7121_/Q _5978_/X _6015_/X _7017_/Q _6125_/X VGND VGND VPWR VPWR _6129_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3338_/A _3563_/A VGND VGND VPWR VPWR _5560_/A sky130_fd_sc_hd__nor2_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6057_ _6854_/Q _5983_/X _5998_/X _6886_/Q VGND VGND VPWR VPWR _6057_/X sky130_fd_sc_hd__a22o_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4266__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3269_ _3269_/A0 hold86/X _3998_/S VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__mux2_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _4683_/A _5007_/Y _4999_/D VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__o21a_1
XFILLER_100_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4018__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__A1 _6848_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6959_ _7001_/CLK _6959_/D fanout466/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5766__B2 _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3777__B1 _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5518__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5437__S _5442_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4741__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold790 hold790/A VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3701__B1 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6246__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2180 hold819/X VGND VGND VPWR VPWR _4254_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4257__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2191 hold826/X VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1490 _6478_/Q VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3480__A2 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5757__A1 _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5757__B2 _6904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3958_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5509__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5347__S _5352_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput306 _3953_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold1768/X VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__buf_6
X_4310_ _4310_/A _5569_/B VGND VGND VPWR VPWR _4315_/S sky130_fd_sc_hd__and2_2
XANTENNA__3940__A0 _6502_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput328 hold1739/X VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__buf_6
XFILLER_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput339 hold1756/X VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__buf_6
X_5290_ _5290_/A hold9/A VGND VGND VPWR VPWR _5298_/S sky130_fd_sc_hd__and2_4
X_4241_ _4241_/A _5578_/B VGND VGND VPWR VPWR _4249_/S sky130_fd_sc_hd__and2_4
XANTENNA__5693__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4172_ _4172_/A0 _5580_/A1 _4175_/S VGND VGND VPWR VPWR _4172_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6237__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold16_A hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4799__A2 _4714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3471__A2 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _6815_/CLK _6813_/D fanout446/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5748__A1 _6887_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3956_ input84/X _3881_/C _6457_/Q VGND VGND VPWR VPWR _3956_/X sky130_fd_sc_hd__mux2_4
X_6744_ _6761_/CLK _6744_/D _6416_/A VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6675_ _7112_/CLK hold74/X fanout473/X VGND VGND VPWR VPWR _7229_/A sky130_fd_sc_hd__dfrtp_1
X_3887_ _6455_/Q _6434_/Q _6423_/B VGND VGND VPWR VPWR _3969_/B sky130_fd_sc_hd__o21a_2
XFILLER_164_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5626_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6017_/A sky130_fd_sc_hd__and2b_4
XANTENNA__6173__A1 _6907_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5557_ _5557_/A0 _5584_/A1 _5559_/S VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5920__A1 _6596_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5920__B2 _6771_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4508_ _4625_/A _4508_/B VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__nand2_2
XFILLER_144_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5488_ _5488_/A _5578_/B VGND VGND VPWR VPWR _5496_/S sky130_fd_sc_hd__and2_4
XFILLER_144_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7227_ _7227_/A VGND VGND VPWR VPWR _7227_/X sky130_fd_sc_hd__clkbuf_2
X_4439_ _4701_/A _4808_/B VGND VGND VPWR VPWR _4469_/B sky130_fd_sc_hd__xnor2_4
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7158_ _7180_/CLK _7158_/D fanout446/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6228__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6109_ _7088_/Q _5638_/X _6015_/X _7016_/Q VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7089_ _7133_/CLK _7089_/D fanout470/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4239__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3447__C1 _3435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input75_A porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6219__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3453__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3810_ _6470_/Q _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3904_/A sky130_fd_sc_hd__and3_4
XFILLER_178_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _4947_/A _4662_/Y _4782_/X VGND VGND VPWR VPWR _4790_/X sky130_fd_sc_hd__o21ba_1
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_18 _5849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _6339_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6901_/Q _5317_/A _4140_/A _6589_/Q _3740_/X VGND VGND VPWR VPWR _3750_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6460_ _3547_/A1 _6460_/D _6410_/X VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_4
X_3672_ _6481_/Q _4000_/A _4170_/A _6616_/Q _3671_/X VGND VGND VPWR VPWR _3673_/D
+ sky130_fd_sc_hd__a221o_1
X_5411_ _5411_/A0 _5582_/A1 _5415_/S VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5902__A1 _6526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6391_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6391_/X sky130_fd_sc_hd__and2_1
X_5342_ _5342_/A0 _5567_/A1 _5343_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5273_ _5273_/A0 _5534_/A1 _5280_/S VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2905 _7184_/Q VGND VGND VPWR VPWR _6341_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7012_ _7131_/CLK _7012_/D fanout452/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4224_ _3550_/B _6430_/B _4012_/X _4237_/S _5578_/B VGND VGND VPWR VPWR _4240_/S
+ sky130_fd_sc_hd__o221a_4
Xhold2916 hold19/A VGND VGND VPWR VPWR _3831_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2927 _6685_/Q VGND VGND VPWR VPWR _3918_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2938 _6489_/Q VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2949 _6686_/Q VGND VGND VPWR VPWR _3919_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4155_ _4155_/A0 _5194_/A1 _4157_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5540__S _5540_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3692__A2 _4206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ _3675_/Y hold976/A _4091_/S VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4988_ _4988_/A _5009_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6727_ _6731_/CLK _6727_/D _6413_/A VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3747__A3 _3745_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3601__C1 _3600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3939_ _6503_/Q _3879_/B _6459_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6658_ _3940_/A1 _6658_/D _6425_/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5684_/B sky130_fd_sc_hd__and2_4
XFILLER_180_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6589_ _6817_/CLK _6589_/D fanout435/X VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3380__B2 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout363 _4411_/Y VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__buf_12
Xfanout374 hold1153/X VGND VGND VPWR VPWR hold1154/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout385 _5537_/A1 VGND VGND VPWR VPWR _5582_/A1 sky130_fd_sc_hd__buf_8
XANTENNA__5450__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout396 _5580_/A1 VGND VGND VPWR VPWR _5562_/A1 sky130_fd_sc_hd__clkbuf_16
XANTENNA__7231__A _7231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3683__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6082__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4935__A2 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output279_A _6796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5896__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6776__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5648__B1 _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5360__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2025_A _6582_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6073__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5960_ _6746_/Q _5929_/B _5668_/X _6648_/Q _5949_/X VGND VGND VPWR VPWR _5960_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5820__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4911_ _4633_/B _4688_/B _4845_/X _4901_/B VGND VGND VPWR VPWR _5107_/A sky130_fd_sc_hd__o211a_1
X_5891_ _6570_/Q _5674_/X _5680_/X _6708_/Q VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4842_ _4590_/Y _4676_/Y _4628_/Y VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__o21a_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4773_ _4729_/A _4688_/C _4542_/Y VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__o21a_1
X_6512_ _6512_/CLK _6512_/D fanout473/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
X_3724_ _6934_/Q _5353_/A _4152_/A _6600_/Q _3723_/X VGND VGND VPWR VPWR _3725_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6128__B2 _6865_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6443_ net399_2/A _6443_/D _6398_/X VGND VGND VPWR VPWR _6443_/Q sky130_fd_sc_hd__dfrtp_1
X_3655_ _3655_/A _3655_/B _3655_/C _3655_/D VGND VGND VPWR VPWR _3674_/B sky130_fd_sc_hd__nor4_1
XANTENNA__5535__S _5540_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6374_ _6686_/Q _6374_/A2 _6374_/B1 _6685_/Q _6373_/X VGND VGND VPWR VPWR _6374_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3586_ _6960_/Q _5380_/A _3431_/Y input64/X _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_4
X_5325_ _5325_/A0 _5568_/A1 _5325_/S VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ _5256_/A0 _5562_/A1 _5262_/S VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__mux2_1
Xhold2702 _6753_/Q VGND VGND VPWR VPWR hold562/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2713 _6958_/Q VGND VGND VPWR VPWR hold568/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2724 hold594/X VGND VGND VPWR VPWR _5539_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6300__B2 _6772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2735 _3251_/Y VGND VGND VPWR VPWR _3252_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4207_ _4207_/A0 _5543_/A1 _4211_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
Xhold2746 hold759/X VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2757 hold852/X VGND VGND VPWR VPWR _4255_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5187_ _5187_/A0 _5194_/A1 _5190_/S VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5270__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2768 _6921_/Q VGND VGND VPWR VPWR hold762/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2779 hold638/X VGND VGND VPWR VPWR _5351_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3665__A2 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4862__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4138_ _4138_/A0 _5195_/A1 _4139_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4069_ _4069_/A0 _5195_/A1 _4070_/S VGND VGND VPWR VPWR _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3417__A2 _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5811__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6114__B _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6119__A1 _7089_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6119__B2 _6889_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5445__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5878__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input38_A mgmt_gpio_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3656__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6055__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3408__A2 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5802__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5030__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3592__A1 _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3592__B2 _6735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold608 hold608/A VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5355__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold619 hold619/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3440_ _7026_/Q _5452_/A _5407_/A _6986_/Q _3437_/X VGND VGND VPWR VPWR _3444_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap349 _3293_/Y VGND VGND VPWR VPWR _4056_/C sky130_fd_sc_hd__buf_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3371_ _7132_/Q _5569_/A _5326_/A _6916_/Q _3370_/X VGND VGND VPWR VPWR _3371_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5110_ _5110_/A _5110_/B VGND VGND VPWR VPWR _5110_/Y sky130_fd_sc_hd__nand2_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6839_/Q _6339_/B _6089_/X VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__o21ba_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2009 hold691/X VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5148_/B _5162_/B VGND VGND VPWR VPWR _5042_/D sky130_fd_sc_hd__and3_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 hold381/X VGND VGND VPWR VPWR _5276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1319 _6651_/Q VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3647__A2 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2407_A _6787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4844__B2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6046__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6992_ _6992_/CLK _6992_/D fanout464/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5943_ _6735_/Q _5656_/X _5679_/X _6592_/Q _5942_/X VGND VGND VPWR VPWR _5943_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5874_ _6594_/Q _5670_/X _5671_/X _6634_/Q _5873_/X VGND VGND VPWR VPWR _5879_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4825_ _4822_/Y _4825_/B _4825_/C _4924_/B VGND VGND VPWR VPWR _4825_/X sky130_fd_sc_hd__and4b_1
XFILLER_178_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4756_ _5009_/B _4732_/B _4811_/B VGND VGND VPWR VPWR _4757_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__3583__A1 _6904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3707_ input15/X _3307_/Y _3389_/Y _3706_/X VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3583__B2 _6880_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4687_ _4712_/A _4691_/B VGND VGND VPWR VPWR _4688_/C sky130_fd_sc_hd__nand2_8
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5265__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6426_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
X_3638_ _7031_/Q _5461_/A _5169_/A _6771_/Q _3637_/X VGND VGND VPWR VPWR _3645_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6357_ _6357_/A _6358_/A VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__nand2_1
X_3569_ _6952_/Q _3291_/Y _5308_/A _6896_/Q _3561_/X VGND VGND VPWR VPWR _3569_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5308_ _5308_/A _5578_/B VGND VGND VPWR VPWR _5316_/S sky130_fd_sc_hd__and2_4
X_6288_ _6281_/X _6283_/X _6288_/C _6313_/D VGND VGND VPWR VPWR _6289_/C sky130_fd_sc_hd__and4bb_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2510 hold921/X VGND VGND VPWR VPWR _5354_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2521 _6736_/Q VGND VGND VPWR VPWR hold875/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2532 _4069_/X VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5239_ _5239_/A0 _5527_/A1 _5244_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
Xhold2543 _6837_/Q VGND VGND VPWR VPWR hold910/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2554 _6750_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1820 _6561_/Q VGND VGND VPWR VPWR hold991/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2565 _6859_/Q VGND VGND VPWR VPWR hold654/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__A2 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1831 hold486/X VGND VGND VPWR VPWR hold1831/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2576 _7210_/A VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1842 hold466/X VGND VGND VPWR VPWR _4019_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2587 _5405_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2598 hold518/X VGND VGND VPWR VPWR _4196_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1853 _6761_/Q VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6037__B1 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1864 hold492/X VGND VGND VPWR VPWR hold1864/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1875 hold582/X VGND VGND VPWR VPWR _4040_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1886 hold996/X VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1897 _7048_/Q VGND VGND VPWR VPWR hold814/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5260__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7202__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5012__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3574__A1 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3574__B2 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5079__A1 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5079__B2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3629__A2 _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__buf_8
XFILLER_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5251__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6200__B1 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _4610_/A _4611_/A VGND VGND VPWR VPWR _4614_/C sky130_fd_sc_hd__nand2_1
X_5590_ _6490_/Q _6492_/Q _6491_/Q _3924_/Y VGND VGND VPWR VPWR _5599_/D sky130_fd_sc_hd__o31a_4
XANTENNA__3565__A1 _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4541_ _4971_/A _4724_/C VGND VGND VPWR VPWR _5149_/A sky130_fd_sc_hd__nand2_2
XFILLER_128_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold416 hold416/A VGND VGND VPWR VPWR hold416/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4472_ _4564_/C _4486_/B VGND VGND VPWR VPWR _4510_/A sky130_fd_sc_hd__nand2_4
XFILLER_144_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold427 hold427/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold438 hold438/A VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3423_ _6779_/Q _3422_/Y _3738_/S VGND VGND VPWR VPWR _3423_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6211_ _7140_/Q _5977_/X _5985_/X _6908_/Q _6210_/X VGND VGND VPWR VPWR _6211_/X
+ sky130_fd_sc_hd__a221o_1
Xhold449 hold449/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7191_ _7191_/CLK _7191_/D VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6142_ _6142_/A1 _6167_/S _6140_/X _6141_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__o22a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3354_/A _3354_/B VGND VGND VPWR VPWR _5353_/A sky130_fd_sc_hd__nor2_8
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7023_/Q _5971_/X _6007_/X _6847_/Q _6068_/X VGND VGND VPWR VPWR _6076_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1105 hold5/X VGND VGND VPWR VPWR _5228_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3285_ hold78/X hold87/X VGND VGND VPWR VPWR _3322_/B sky130_fd_sc_hd__and2b_4
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1116 _6729_/Q VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5024_ _5139_/B _5024_/B VGND VGND VPWR VPWR _5024_/Y sky130_fd_sc_hd__nand2_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _6759_/Q VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1138 _4080_/X VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_100_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1149 _5491_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5490__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6975_ _6977_/CLK _6975_/D fanout460/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5242__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _5947_/A1 _6342_/S _5924_/X _5925_/X VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__o22a_1
XFILLER_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5857_ _6868_/Q _5673_/X _5850_/X _5851_/X _5856_/X VGND VGND VPWR VPWR _5857_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _4808_/A _4808_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6666__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5788_ _7017_/Q _5664_/X _5681_/X _7089_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4739_ _5011_/A _4712_/Y _4727_/Y _4823_/C _4738_/Y VGND VGND VPWR VPWR _4739_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6409_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and2_1
XFILLER_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold950 hold950/A VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7146__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold961 hold961/A VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold972 hold972/A VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold983 hold983/A VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold994 hold994/A VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6258__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2340 _4211_/X VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2351 hold862/X VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2362 _5490_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2373 _4288_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2384 _4251_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5481__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1650 hold354/X VGND VGND VPWR VPWR _5339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2395 _5556_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1661 hold172/X VGND VGND VPWR VPWR _4243_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1672 _6601_/Q VGND VGND VPWR VPWR hold581/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1683 _5190_/X VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1694 hold311/X VGND VGND VPWR VPWR _5403_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5678__B _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4582__B _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5233__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5784__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3547__B2 _7232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output261_A _6783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7091_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6249__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7101_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5472__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5224__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6760_ _6760_/CLK _6760_/D _6407_/A VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_4
X_3972_ _3972_/A input1/X VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__and2_1
XANTENNA__5775__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5711_ _6982_/Q _5656_/X _5663_/X _7022_/Q _5710_/X VGND VGND VPWR VPWR _5718_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3786__B2 _6604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6691_ _7045_/CLK _6691_/D fanout444/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5642_ _5589_/Y _5604_/Y _5641_/Y _6492_/Q VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__a22o_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5573_ _5573_/A0 _5582_/A1 _5577_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7169__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2739_A _6869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4524_ _4596_/A _5048_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__nand2_2
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold213 hold213/A VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7121_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold235 hold235/A VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold246 hold246/A VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4455_ _4590_/B _4488_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__nand2_4
Xhold257 hold257/A VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5543__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold268 hold268/A VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold279 hold279/A VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3406_ _3406_/A _3406_/B VGND VGND VPWR VPWR _3422_/A sky130_fd_sc_hd__nor2_1
X_4386_ _5011_/A _4578_/A VGND VGND VPWR VPWR _4886_/A sky130_fd_sc_hd__nor2_2
X_7174_ _7179_/CLK _7174_/D fanout445/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _6921_/Q _5995_/X _5997_/X _6953_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
X_3337_ hold30/X _3563_/B VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__nor2_8
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1038_A _5541_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _7102_/Q _6008_/X _6018_/X _6966_/Q _6055_/X VGND VGND VPWR VPWR _6056_/X
+ sky130_fd_sc_hd__a221o_1
X_3268_ _3842_/C1 _6460_/Q _6657_/Q VGND VGND VPWR VPWR _3268_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3998__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5463__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5007_ _5009_/B _4735_/B _4677_/B _4733_/X VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4683__A _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3199_ _3199_/A VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3474__B1 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5766__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6958_ _7124_/CLK _6958_/D fanout467/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3777__A1 _6784_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5909_ _6636_/Q _5671_/X _5906_/X _5907_/X _5908_/X VGND VGND VPWR VPWR _5909_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6889_ _7073_/CLK _6889_/D fanout444/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5453__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold780 hold780/A VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3701__A1 input44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6686__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5454__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2170 _6592_/Q VGND VGND VPWR VPWR hold758/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2181 _4254_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input20_A mask_rev_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2192 _4308_/X VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1480 _4187_/X VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1491 hold296/X VGND VGND VPWR VPWR _3999_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5206__A1 _5303_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5757__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3768__A1 _6869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6182__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4193__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _3952_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
XANTENNA__3940__A1 _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput318 hold980/X VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__buf_6
Xoutput329 hold1736/X VGND VGND VPWR VPWR hold458/A sky130_fd_sc_hd__buf_6
XANTENNA__5363__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4240_ _4240_/A0 _4239_/X _4240_/S VGND VGND VPWR VPWR _4240_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5693__A1 _6877_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4171_ _4171_/A0 _5561_/A1 _4175_/S VGND VGND VPWR VPWR _4171_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5445__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3456__B1 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2591_A _6793_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6812_ _6816_/CLK _6812_/D fanout446/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5748__A2 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _6745_/CLK _6743_/D fanout440/X VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfrtp_2
X_3955_ _3998_/S _3955_/A2 _6423_/B _3954_/Y VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5538__S _5540_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6674_ _7112_/CLK _6674_/D fanout473/X VGND VGND VPWR VPWR _7228_/A sky130_fd_sc_hd__dfrtp_1
X_3886_ _7158_/Q _6810_/Q _6815_/Q VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__mux2_8
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5625_ _7152_/Q _7151_/Q _6491_/Q VGND VGND VPWR VPWR _5631_/A sky130_fd_sc_hd__and3_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6173__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4184__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5556_ _5556_/A0 _5583_/A1 _5559_/S VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5920__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3931__A1 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4507_ _4508_/B VGND VGND VPWR VPWR _4507_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5273__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5487_ _5487_/A0 _5568_/A1 hold17/A VGND VGND VPWR VPWR _5487_/X sky130_fd_sc_hd__mux2_1
X_7226_ _7226_/A VGND VGND VPWR VPWR _7226_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ _4598_/A VGND VGND VPWR VPWR _4438_/Y sky130_fd_sc_hd__inv_2
X_7157_ _7180_/CLK _7157_/D fanout446/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4369_ _4955_/A _4513_/B VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__and2_4
XANTENNA__3695__B1 _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6108_ _6936_/Q _5980_/X _6017_/X _7072_/Q _6093_/X VGND VGND VPWR VPWR _6113_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7088_ _7112_/CLK _7088_/D fanout473/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5436__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6039_ _6039_/A _6039_/B _6039_/C _6039_/D VGND VGND VPWR VPWR _6040_/B sky130_fd_sc_hd__nor4_1
XANTENNA__3447__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5448__S _5451_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4175__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5911__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input68_A mgmt_gpio_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5427__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3438__B1 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3989__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5358__S _5361_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_19 _5869_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3740_ _6853_/Q _5263_/A _4122_/A _6574_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3610__B1 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3671_ input37/X _3293_/Y _4140_/A _6591_/Q VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6155__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5410_ _5410_/A0 _5572_/A1 _5415_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4166__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6390_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__and2_1
XANTENNA__5902__A2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3374__C1 _3360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _5341_/A0 _5575_/A1 _5343_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _5272_/A _5533_/B VGND VGND VPWR VPWR _5280_/S sky130_fd_sc_hd__and2_4
XFILLER_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7011_ _7052_/CLK _7011_/D fanout464/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_4
X_4223_ _3184_/Y _4223_/A2 _6680_/D _5139_/A _4222_/Y VGND VGND VPWR VPWR _4223_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold2906 _6317_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2917 _7170_/Q VGND VGND VPWR VPWR _5947_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2928 _6458_/Q VGND VGND VPWR VPWR _3851_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2939 _3923_/Y VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4154_ _4154_/A0 _5193_/A1 _4157_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5418__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4085_ _3737_/Y hold986/A _4091_/S VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4987_ _4384_/A _4990_/B _4683_/B _4823_/A VGND VGND VPWR VPWR _5083_/B sky130_fd_sc_hd__o31a_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5268__S _5271_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6726_ _7045_/CLK _6726_/D fanout444/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_4
X_3938_ _6826_/Q input81/X _3971_/B VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6657_ _3940_/A1 _6657_/D _6424_/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6146__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3869_ _3869_/A _3869_/B VGND VGND VPWR VPWR _3869_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4157__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5608_ _6491_/Q _5679_/B VGND VGND VPWR VPWR _5613_/B sky130_fd_sc_hd__nand2_1
X_6588_ _6786_/CLK _6588_/D fanout435/X VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ _5539_/A0 _5584_/A1 _5541_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5106__B1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3380__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7209_ _7209_/A VGND VGND VPWR VPWR _7209_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3668__B1 _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5409__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout386 hold43/X VGND VGND VPWR VPWR _5537_/A1 sky130_fd_sc_hd__buf_12
Xfanout397 _5228_/A1 VGND VGND VPWR VPWR _5580_/A1 sky130_fd_sc_hd__buf_8
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6862__RESET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input122_A wb_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6082__B2 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4632__A2 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__A2 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4148__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3974_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_171_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output174_A _3974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5207__A _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3371__A2 _5569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3659__B1 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4320__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6073__A1 _7023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4084__A0 _3803_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4910_ _4655_/A _4640_/Y _4655_/B _4704_/C _4791_/A VGND VGND VPWR VPWR _5049_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5820__B2 _6907_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5890_ _6753_/Q _5681_/X _5889_/X VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__a21o_1
X_4841_ _4917_/D _4915_/B VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__nand2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4772_ _5136_/A _4973_/C VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _6512_/CLK _6511_/D fanout473/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3723_ _6990_/Q _5416_/A _5326_/A _6910_/Q VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6128__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4139__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6442_ net399_2/A _6442_/D _6397_/X VGND VGND VPWR VPWR _6442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3654_ _7039_/Q _3325_/Y _4122_/A _6576_/Q _3653_/X VGND VGND VPWR VPWR _3655_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6373_ _6684_/Q _6373_/A2 _6373_/B1 _4218_/Y VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3585_ _6572_/Q hold57/A _4158_/A _6607_/Q VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5324_ _5324_/A0 _5567_/A1 _5325_/S VGND VGND VPWR VPWR _5324_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3362__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2703 hold562/X VGND VGND VPWR VPWR _4330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5255_ _5255_/A0 _5579_/A1 _5262_/S VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__mux2_1
Xhold2714 _5382_/X VGND VGND VPWR VPWR hold569/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6300__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2725 _7114_/Q VGND VGND VPWR VPWR hold604/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4311__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4206_ _4206_/A hold9/X VGND VGND VPWR VPWR _4211_/S sky130_fd_sc_hd__and2_4
Xhold2736 _3252_/Y VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2747 _7227_/A VGND VGND VPWR VPWR hold610/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4675__B _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2758 _4255_/X VGND VGND VPWR VPWR hold853/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5186_ _5186_/A0 _5193_/A1 _5190_/S VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2769 hold762/X VGND VGND VPWR VPWR _5340_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4862__A2 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4137_ hold631/X _5194_/A1 _4139_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout372_A _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4068_ _4068_/A0 _5194_/A1 _4070_/S VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5811__A1 _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1487_A _6605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ _6746_/CLK _6709_/D _6416_/A VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6119__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1654_A _6699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6411__A _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4302__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4585__B _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4853__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6055__B2 _6846_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5802__A1 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5030__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7149__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output291_A _6483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3592__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3370_ input42/X _3293_/Y _5524_/A _7092_/Q VGND VGND VPWR VPWR _3370_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6784__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6294__B2 _6533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5040_ _4454_/A _4463_/B _4570_/D _4954_/D _5039_/Y VGND VGND VPWR VPWR _5162_/B
+ sky130_fd_sc_hd__o311a_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 _5276_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4844__A2 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6991_ _7063_/CLK _6991_/D fanout460/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5942_ _6642_/Q _5655_/X _5663_/X _6632_/Q _5928_/Y VGND VGND VPWR VPWR _5942_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6742_/Q _5929_/B _5678_/B _5872_/Y VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
X_4824_ _4995_/A _4698_/Y _4583_/B VGND VGND VPWR VPWR _4825_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4755_ _4976_/A _4755_/B _4755_/C _4997_/A VGND VGND VPWR VPWR _4757_/C sky130_fd_sc_hd__and4b_1
XFILLER_193_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5546__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3706_ _6974_/Q _5398_/A hold57/A _6570_/Q _3705_/X VGND VGND VPWR VPWR _3706_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3583__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4780__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4686_ _4712_/A _4714_/B _4714_/C VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__and3_1
XFILLER_146_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6425_ _6430_/A _6433_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
X_3637_ _6967_/Q _5389_/A _5497_/A _7063_/Q VGND VGND VPWR VPWR _3637_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4532__A1 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6356_ _6358_/A _6356_/B VGND VGND VPWR VPWR _6356_/Y sky130_fd_sc_hd__nand2_2
XFILLER_1_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3568_ _6602_/Q _4152_/A _4256_/A _6695_/Q VGND VGND VPWR VPWR _3568_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5307_/A0 _5577_/A1 _5307_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6287_ _6452_/Q _6016_/X _6284_/X _6286_/X VGND VGND VPWR VPWR _6288_/C sky130_fd_sc_hd__a211oi_1
Xhold2500 _6885_/Q VGND VGND VPWR VPWR hold906/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3499_ _3499_/A _3499_/B _3499_/C _3499_/D VGND VGND VPWR VPWR _3558_/B sky130_fd_sc_hd__nor4_2
Xhold2511 _5354_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2522 hold875/X VGND VGND VPWR VPWR _4309_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2533 _7093_/Q VGND VGND VPWR VPWR hold926/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5238_ _5238_/A0 _5238_/A1 _5244_/S VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2544 hold910/X VGND VGND VPWR VPWR _5246_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2555 hold799/X VGND VGND VPWR VPWR _4326_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1810 _5495_/X VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1821 hold991/X VGND VGND VPWR VPWR hold482/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2566 hold654/X VGND VGND VPWR VPWR _5270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1832 _6506_/Q VGND VGND VPWR VPWR hold879/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2577 hold494/X VGND VGND VPWR VPWR _4236_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1843 _4019_/X VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5169_ _5169_/A _5220_/C VGND VGND VPWR VPWR _5174_/S sky130_fd_sc_hd__and2_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2588 _6653_/Q VGND VGND VPWR VPWR hold677/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1854 hold725/X VGND VGND VPWR VPWR _4339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2599 _4196_/X VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6037__B2 _7053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1865 _6565_/Q VGND VGND VPWR VPWR _4112_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1876 _6562_/Q VGND VGND VPWR VPWR _4109_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1887 hold462/X VGND VGND VPWR VPWR hold1887/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1898 hold814/X VGND VGND VPWR VPWR _5483_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5012__A2 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5456__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3574__A2 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4771__B2 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5720__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input50_A mgmt_gpio_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3966__A_N _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output304_A _3428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5787__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5220__A hold64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5366__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2085_A _6632_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3565__A2 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4540_ _4601_/A _4569_/C _4537_/X _4894_/A _4539_/Y VGND VGND VPWR VPWR _4540_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4471_ _4485_/B _4564_/C _4568_/A VGND VGND VPWR VPWR _4611_/A sky130_fd_sc_hd__and3_4
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold428 hold428/A VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6210_ _6996_/Q _6014_/X _6017_/X _7076_/Q VGND VGND VPWR VPWR _6210_/X sky130_fd_sc_hd__a22o_1
Xhold439 hold439/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
X_3422_ _3422_/A _3422_/B _3422_/C VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__5711__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7190_ _7194_/CLK _7190_/D VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6141_ _6141_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6141_/X sky130_fd_sc_hd__o21ba_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3563_/B _3726_/B VGND VGND VPWR VPWR _5245_/A sky130_fd_sc_hd__nor2_8
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6072_ _6991_/Q _6014_/X _6070_/X _6071_/X VGND VGND VPWR VPWR _6076_/A sky130_fd_sc_hd__a211o_1
XFILLER_112_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3284_/A hold63/X VGND VGND VPWR VPWR _3295_/A sky130_fd_sc_hd__nand2_8
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _5228_/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 hold187/X VGND VGND VPWR VPWR _4301_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5023_ _5023_/A _5083_/C _5023_/C _5023_/D VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__and4_1
Xhold1128 hold195/X VGND VGND VPWR VPWR _4337_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1139 _7127_/Q VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_66_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6974_ _6974_/CLK _6974_/D fanout454/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5778__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5925_ _6490_/Q _5925_/A2 _5649_/Y VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _6892_/Q _5688_/X _5852_/X _5853_/X _5855_/X VGND VGND VPWR VPWR _5856_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4807_ _4411_/Y _4590_/Y _4370_/Y VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__a21o_2
X_5787_ _6929_/Q _5684_/X _5689_/X _7081_/Q _5786_/X VGND VGND VPWR VPWR _5792_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5276__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4738_ _5009_/A _4738_/B _5150_/C VGND VGND VPWR VPWR _4738_/Y sky130_fd_sc_hd__nand3_1
XFILLER_175_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5950__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _4638_/Y _4995_/A _4668_/Y _4583_/B VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6408_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__and2_1
Xhold940 hold940/A VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5702__B1 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold951 hold951/A VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold962 hold962/A VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold973 hold973/A VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6339_ _6330_/X _6339_/B _6339_/C _6339_/D VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__and4b_2
Xhold984 hold984/A VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6258__A1 _6713_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6258__B2 _6570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2330 _6594_/Q VGND VGND VPWR VPWR hold856/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2341 _7057_/Q VGND VGND VPWR VPWR hold721/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2352 _4329_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2363 _7018_/Q VGND VGND VPWR VPWR hold619/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2374 _7026_/Q VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2385 _6726_/Q VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1640 _4293_/X VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2396 _7065_/Q VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1651 _5339_/X VGND VGND VPWR VPWR hold355/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1662 _4243_/X VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1673 hold581/X VGND VGND VPWR VPWR _4155_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1684 _6862_/Q VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1695 _5403_/X VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5769__B1 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3795__A2 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5969__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input98_A usr2_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__B1 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4090__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3547__A2 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5941__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6739__SET_B fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold9_A hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ _3971_/A _3971_/B VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__and2_1
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5710_ _6998_/Q _5666_/X _5673_/X _6862_/Q VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3786__A2 _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6690_ _6735_/CLK _6690_/D fanout444/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5641_ _5645_/C _5641_/B VGND VGND VPWR VPWR _5641_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6185__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2467_A _6534_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3538__A2 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5572_ _5572_/A0 _5572_/A1 _5577_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5932__B1 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4523_ _4523_/A _4595_/B VGND VGND VPWR VPWR _4523_/Y sky130_fd_sc_hd__nand2_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold214 hold214/A VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold225 hold225/A VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4454_ _4454_/A _4463_/B VGND VGND VPWR VPWR _4724_/C sky130_fd_sc_hd__nor2_8
Xhold247 hold247/A VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold258 hold258/A VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3405_ hold24/A _3392_/X _3402_/X _3403_/X _3404_/X VGND VGND VPWR VPWR _3406_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5160__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7173_ _7185_/CLK _7173_/D fanout445/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_1
X_4385_ _5001_/A _4751_/B VGND VGND VPWR VPWR _4578_/A sky130_fd_sc_hd__nand2_2
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6857_/Q _5983_/X _5993_/X _7009_/Q _6123_/X VGND VGND VPWR VPWR _6129_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3710__A2 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3338_/A _3686_/B VGND VGND VPWR VPWR _3336_/Y sky130_fd_sc_hd__nor2_8
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6862_/Q _5999_/X _6007_/X _6846_/Q VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a22o_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3267_ hold13/X hold46/X VGND VGND VPWR VPWR _3355_/A sky130_fd_sc_hd__and2_4
XFILLER_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5139_/A _5140_/A VGND VGND VPWR VPWR _5006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4683__B _4683_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3198_ _6491_/Q VGND VGND VPWR VPWR _5647_/B sky130_fd_sc_hd__clkinv_4
XFILLER_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3474__B2 _6573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout452_A fanout453/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6957_ _7001_/CLK _6957_/D fanout466/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3777__A2 _5178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5908_ _6749_/Q _5666_/X _5689_/X _6626_/Q VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6888_ _7107_/CLK _6888_/D fanout451/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6176__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5839_ _3243_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6403__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold770 hold770/A VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold792 _5376_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input152_A wb_dat_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3701__A2 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6100__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2160 _6725_/Q VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2171 hold758/X VGND VGND VPWR VPWR _4144_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2182 _7020_/Q VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2193 _6599_/Q VGND VGND VPWR VPWR hold735/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1470 _6989_/Q VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1481 _7115_/Q VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input13_A mask_rev_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1492 _3999_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_55_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4085__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3768__A2 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5390__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _3971_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_126_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput319 hold1731/X VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__buf_6
XFILLER_114_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5142__A1 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5693__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4170_ _4170_/A hold9/X VGND VGND VPWR VPWR _4175_/S sky130_fd_sc_hd__and2_2
XFILLER_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ _6816_/CLK _6811_/D fanout446/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6742_ _6752_/CLK _6742_/D fanout440/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_4
X_3954_ _3998_/S _3954_/B VGND VGND VPWR VPWR _3954_/Y sky130_fd_sc_hd__nor2_2
X_6673_ _7112_/CLK _6673_/D fanout473/X VGND VGND VPWR VPWR _7227_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6158__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3885_ _6449_/Q _3885_/A2 _6656_/Q _3904_/A VGND VGND VPWR VPWR _6434_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5624_ _7152_/Q _7151_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__and2_4
XFILLER_176_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5905__B1 _5677_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5555_ _5555_/A0 _5582_/A1 _5559_/S VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5381__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5554__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4506_ _4506_/A _4840_/A _4917_/B _4917_/C VGND VGND VPWR VPWR _4508_/B sky130_fd_sc_hd__and4_2
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5486_ _5486_/A0 _5549_/A1 hold17/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7225_ _7225_/A VGND VGND VPWR VPWR _7225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4437_ _4560_/B _4560_/C _4341_/X _4394_/Y VGND VGND VPWR VPWR _4598_/A sky130_fd_sc_hd__a211oi_4
XANTENNA__6330__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7156_ _7180_/CLK _7156_/D fanout451/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4368_ _4368_/A _4368_/B VGND VGND VPWR VPWR _4513_/B sky130_fd_sc_hd__nor2_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A mask_rev_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6107_ _7120_/Q _5978_/X _5995_/X _6920_/Q _6106_/X VGND VGND VPWR VPWR _6113_/A
+ sky130_fd_sc_hd__a221o_1
X_3319_ _3686_/B _3549_/B VGND VGND VPWR VPWR _3319_/Y sky130_fd_sc_hd__nor2_8
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7087_ _7093_/CLK _7087_/D fanout450/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4299_ _4299_/A0 _5561_/A1 hold65/X VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6038_ _6909_/Q _5991_/X _5993_/X _7005_/Q _6037_/X VGND VGND VPWR VPWR _6039_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5729__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6149__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3249__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6974_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5372__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5464__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4588__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6321__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3438__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7159__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7001_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4938__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6738__RESET_B fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3610__A1 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3610__B2 _6976_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _6847_/Q _5254_/A _5245_/A _6839_/Q _3669_/X VGND VGND VPWR VPWR _3673_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5363__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5374__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3374__B1 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5340_ _5340_/A0 _5448_/A1 _5343_/S VGND VGND VPWR VPWR _5340_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5271_ _5271_/A0 _5577_/A1 _5271_/S VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7010_ _7130_/CLK _7010_/D fanout463/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_4
X_4222_ _6677_/Q _4222_/B _4222_/C VGND VGND VPWR VPWR _4222_/Y sky130_fd_sc_hd__nand3b_1
Xhold2907 _7177_/Q VGND VGND VPWR VPWR _6142_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2918 _7167_/Q VGND VGND VPWR VPWR _5860_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2929 _6456_/Q VGND VGND VPWR VPWR _3854_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4153_ _4153_/A0 _5237_/A1 _4157_/S VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4084_ _3803_/Y hold975/A _4091_/S VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5549__S _5550_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4986_ _4716_/Y _5127_/B _4986_/C VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__and3b_1
XFILLER_168_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5051__B1 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6725_ _6735_/CLK _6725_/D fanout442/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3937_ _6824_/Q input78/X _3971_/B VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_8
XANTENNA__3601__A1 _6984_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6656_ _3940_/A1 _6656_/D _6423_/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3868_ _3868_/A _3868_/B VGND VGND VPWR VPWR _3869_/B sky130_fd_sc_hd__nor2_1
XANTENNA__6000__C1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ _7147_/Q _7146_/Q VGND VGND VPWR VPWR _5679_/B sky130_fd_sc_hd__nor2_8
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5354__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6587_ _6794_/CLK _6587_/D fanout435/X VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfrtp_4
X_3799_ _6722_/Q _4292_/A _4310_/A _6737_/Q VGND VGND VPWR VPWR _3799_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5284__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3365__B1 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5538_ _5538_/A0 _5583_/A1 _5540_/S VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5469_ _5469_/A0 _5568_/A1 _5469_/S VGND VGND VPWR VPWR _5469_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6303__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5106__B2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1432_A _6842_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7208_ _7208_/A VGND VGND VPWR VPWR _7208_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3668__A1 _6473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__B2 _6699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7139_ _7139_/CLK _7139_/D fanout472/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout365 hold71/X VGND VGND VPWR VPWR _5577_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_143_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout376 _5277_/A1 VGND VGND VPWR VPWR _5189_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout387 hold1012/X VGND VGND VPWR VPWR hold1013/A sky130_fd_sc_hd__buf_6
Xfanout398 hold275/X VGND VGND VPWR VPWR _5237_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6082__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A wb_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5459__S _5460_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input80_A spi_sck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5345__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5194__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5896__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5207__B _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4765__C _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6549__CLK _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4608__B1 _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6073__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5820__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5369__S _5370_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A _4917_/B _4857_/C VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__and3_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5584__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4719_/A _4590_/B _4719_/B _4981_/A _4607_/B VGND VGND VPWR VPWR _4771_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6510_ _6512_/CLK _6510_/D fanout473/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_186_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3722_ _7014_/Q _5443_/A _3648_/Y _6819_/Q _3721_/X VGND VGND VPWR VPWR _3725_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ net399_2/A _6441_/D _6396_/X VGND VGND VPWR VPWR _6441_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5336__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3653_ input13/X _3310_/Y _3562_/Y input97/X VGND VGND VPWR VPWR _3653_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5887__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6372_ _6371_/X _6372_/A1 _6384_/S VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__mux2_1
X_3584_ input55/X _4241_/A _4286_/A _6720_/Q _3566_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_1
X_5323_ _5323_/A0 _5575_/A1 _5325_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5254_ _5254_/A _5578_/B VGND VGND VPWR VPWR _5262_/S sky130_fd_sc_hd__and2_4
Xhold2704 _4330_/X VGND VGND VPWR VPWR hold563/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2715 _6826_/Q VGND VGND VPWR VPWR hold784/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2726 hold604/X VGND VGND VPWR VPWR _5557_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4205_ _4205_/A0 _5189_/A1 _4205_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
Xhold2737 _3291_/Y VGND VGND VPWR VPWR _5371_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5185_ _5185_/A0 _5237_/A1 _5190_/S VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__mux2_1
Xhold2748 hold610/X VGND VGND VPWR VPWR _4247_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X sky130_fd_sc_hd__clkbuf_8
Xhold2759 _6954_/Q VGND VGND VPWR VPWR hold617/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A0 _5193_/A1 _4139_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4972__A _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4067_ _4067_/A0 _5193_/A1 _4070_/S VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4075__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5811__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5279__S _5280_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ _4969_/A _4969_/B VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3586__B1 _3431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6708_ _6731_/CLK _6708_/D _6413_/A VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5327__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6639_ _6733_/CLK _6639_/D fanout433/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6411__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5308__A _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1647_A _6591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5878__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4212__A _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_0_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6055__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4066__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5802__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5566__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3577__B1 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5318__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output284_A _6800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6040__C _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6046__A2 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6753__RESET_B fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6990_ _7107_/CLK _6990_/D fanout451/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5941_ _6690_/Q _5659_/X _5687_/X _6602_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5872_ _6717_/Q _5872_/B VGND VGND VPWR VPWR _5872_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3201__A _6719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4823_ _4823_/A _5083_/A _4823_/C VGND VGND VPWR VPWR _4825_/B sky130_fd_sc_hd__and3_1
XFILLER_34_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5557__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3568__B1 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4754_ _4722_/X _4754_/B _5083_/A _4754_/D VGND VGND VPWR VPWR _4755_/B sky130_fd_sc_hd__and4b_1
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3705_ _7110_/Q _5551_/A _5407_/A _6982_/Q VGND VGND VPWR VPWR _3705_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5309__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4685_ _4717_/B _4691_/B VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__nand2_8
XANTENNA__4780__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2929_A _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6424_ _6430_/A _6433_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
X_3636_ _3636_/A _3636_/B _3636_/C _3636_/D VGND VGND VPWR VPWR _3675_/B sky130_fd_sc_hd__nor4_2
XFILLER_134_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4389__D _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6355_ _6358_/A _6355_/A2 _6682_/Q VGND VGND VPWR VPWR _6355_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_162_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3567_ _6888_/Q _5299_/A _4128_/A _6582_/Q VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5562__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5306_ _5306_/A0 _5549_/A1 _5307_/S VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6286_ _6581_/Q _5998_/X _6004_/X _6576_/Q _6285_/X VGND VGND VPWR VPWR _6286_/X
+ sky130_fd_sc_hd__a221o_1
X_3498_ _6613_/Q _4164_/A _4328_/A _6756_/Q _3495_/X VGND VGND VPWR VPWR _3499_/D
+ sky130_fd_sc_hd__a221o_1
Xhold2501 hold906/X VGND VGND VPWR VPWR _5300_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6285__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5237_ _5237_/A0 _5237_/A1 _5244_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
Xhold2512 _6925_/Q VGND VGND VPWR VPWR hold912/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2523 _4309_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4296__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2534 hold926/X VGND VGND VPWR VPWR _5534_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2545 _5246_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1800 hold399/X VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1811 _6797_/Q VGND VGND VPWR VPWR hold637/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2556 _4326_/X VGND VGND VPWR VPWR hold800/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1822 hold482/X VGND VGND VPWR VPWR hold1822/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2567 _5270_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5168_ _5137_/X _5162_/Y _5167_/X _5159_/Y VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__a211o_1
Xhold2578 _6513_/Q VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1833 hold879/X VGND VGND VPWR VPWR _4042_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2589 hold677/X VGND VGND VPWR VPWR _4217_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1844 _7190_/Q VGND VGND VPWR VPWR hold993/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6037__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1855 _4339_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1866 hold1866/A VGND VGND VPWR VPWR hold478/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4119_ hold164/X _5581_/A1 hold58/X VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__mux2_1
Xhold1877 hold1877/A VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6494__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4048__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5099_ _4611_/A _4981_/B _5095_/Y _4897_/B VGND VGND VPWR VPWR _5099_/X sky130_fd_sc_hd__a211o_1
Xhold1888 _6502_/Q VGND VGND VPWR VPWR hold885/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1899 _5483_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4599__A2 _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5548__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3257__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5472__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3731__B1 _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input43_A mgmt_gpio_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4088__S _4091_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__A2 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4287__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6028__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4039__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5787__B2 _7081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5220__B _5220_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3798__B1 _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5539__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6200__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4211__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4762__A2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire360 _4579_/B VGND VGND VPWR VPWR _4485_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire371 hold35/X VGND VGND VPWR VPWR wire371/X sky130_fd_sc_hd__buf_12
X_4470_ _4485_/B _4568_/A VGND VGND VPWR VPWR _4486_/B sky130_fd_sc_hd__and2_2
Xhold407 hold407/A VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold418 hold418/A VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold429 hold429/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
X_3421_ _3421_/A _3421_/B _3421_/C _3421_/D VGND VGND VPWR VPWR _3422_/C sky130_fd_sc_hd__nor4_2
XANTENNA__5711__B2 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5382__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6140_ _6841_/Q _6339_/B _6139_/Y _6341_/S VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__o211a_1
XFILLER_98_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ hold62/A hold22/X VGND VGND VPWR VPWR _3648_/B sky130_fd_sc_hd__nand2_8
XFILLER_98_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6903_/Q _5985_/X _5994_/X _7063_/Q _6069_/X VGND VGND VPWR VPWR _6071_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3284_/A hold63/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__and2_4
XANTENNA__4278__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5022_ _5022_/A _5080_/B _5022_/C _5140_/B VGND VGND VPWR VPWR _5023_/D sky130_fd_sc_hd__and4_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 hold6/X VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _4301_/X VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1129 _4337_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5778__A1 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6973_ _6974_/CLK _6973_/D fanout450/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3789__B1 _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5924_ _6527_/Q _5678_/Y _5914_/X _5923_/X _6341_/S VGND VGND VPWR VPWR _5924_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_81_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5855_ _7068_/Q _5671_/X _5854_/X VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5557__S _5559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4806_ _4933_/C _5044_/A _4805_/X _4374_/Y VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__a31o_1
XFILLER_22_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4202__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5786_ _6993_/Q _5929_/B _5678_/B _5785_/Y VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4737_ _4718_/X _4733_/X _4734_/Y _4738_/B VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_119_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4668_ _4712_/A _4712_/B _4700_/B VGND VGND VPWR VPWR _4668_/Y sky130_fd_sc_hd__nand3_4
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6407_ _6407_/A _6433_/B VGND VGND VPWR VPWR _6407_/X sky130_fd_sc_hd__and2_1
X_3619_ _6959_/Q _5380_/A hold89/A _6714_/Q VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__a22o_1
Xhold930 hold930/A VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold941 _4094_/X VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5292__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4599_ _4625_/A _5048_/A _4981_/A VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 hold952/A VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1345_A _6477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold963 hold963/A VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6338_ _6338_/A _6338_/B _6338_/C _6338_/D VGND VGND VPWR VPWR _6339_/D sky130_fd_sc_hd__nor4_1
Xhold974 hold974/A VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold985 hold985/A VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold996 hold996/A VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6258__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6269_ _6621_/Q _5993_/X _6018_/X _6719_/Q _6268_/X VGND VGND VPWR VPWR _6269_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2320 hold832/X VGND VGND VPWR VPWR _5543_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4269__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6675__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2331 hold856/X VGND VGND VPWR VPWR _4147_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2342 hold721/X VGND VGND VPWR VPWR _5493_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2353 _6894_/Q VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2364 hold619/X VGND VGND VPWR VPWR _5449_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1630 hold117/X VGND VGND VPWR VPWR _5224_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2375 hold630/X VGND VGND VPWR VPWR _5458_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1641 _6631_/Q VGND VGND VPWR VPWR hold537/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2386 hold848/X VGND VGND VPWR VPWR _4297_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2397 hold732/X VGND VGND VPWR VPWR _5502_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1652 _6800_/Q VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1663 _6724_/Q VGND VGND VPWR VPWR hold575/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1674 _4155_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1685 hold229/X VGND VGND VPWR VPWR _5274_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1696 _6834_/Q VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5769__A1 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5769__B2 _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5467__S _5469_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4744__A2 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4400__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6249__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4680__A1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3970_ _3970_/A _3970_/B VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__and2_1
XFILLER_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5377__S _5379_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5640_ _5640_/A1 _5638_/X _5639_/Y _5640_/B2 VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__a22o_1
XANTENNA__6185__A1 _6963_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6185__B2 _7003_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5571_ _5571_/A0 _5571_/A1 _5577_/S VGND VGND VPWR VPWR _5571_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5932__B2 _6607_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4522_ _4594_/A _4522_/B VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__nor2_8
XFILLER_8_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold204 hold204/A VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold226 hold226/A VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4453_ _4483_/B _4598_/C VGND VGND VPWR VPWR _4569_/B sky130_fd_sc_hd__nand2_4
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5696__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold248 hold248/A VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3404_ input18/X _3310_/Y _4241_/A input59/X _3394_/X VGND VGND VPWR VPWR _3404_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4310__A _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7172_ _7179_/CLK _7172_/D fanout443/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
X_4384_ _4384_/A _4675_/A VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__nor2_8
XANTENNA__5160__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6123_ _7129_/Q _5973_/X _6014_/X _6993_/Q VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__a22o_1
X_3335_ _3354_/B _3726_/A VGND VGND VPWR VPWR _5326_/A sky130_fd_sc_hd__nor2_8
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A _6054_/B _6054_/C _6054_/D VGND VGND VPWR VPWR _6064_/B sky130_fd_sc_hd__nor4_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ _3266_/A0 hold45/X _3998_/S VGND VGND VPWR VPWR _3266_/X sky130_fd_sc_hd__mux2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5114_/B _5005_/B _5124_/C VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__and3_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3197_ _6492_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3474__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6956_ _6963_/CLK _6956_/D fanout464/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_4
X_5907_ _6744_/Q _5929_/B _5686_/X _6621_/Q VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__a22o_1
X_6887_ _7078_/CLK _6887_/D fanout444/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5287__S _5289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6176__A1 _7115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5838_ _5859_/A1 _5837_/X _6342_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__B2 _7011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5923__A1 _6591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5769_ _7024_/Q _5663_/X _5673_/X _6864_/Q _5768_/X VGND VGND VPWR VPWR _5770_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1462_A _6488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1727_A _6586_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold760 _4269_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold771 _6949_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold782 hold782/A VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input145_A wb_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6100__A1 _6976_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2150 _4001_/X VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6100__B2 _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2161 hold817/X VGND VGND VPWR VPWR _4296_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4111__A0 _3616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2172 _4144_/X VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2183 hold379/X VGND VGND VPWR VPWR _5451_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2194 hold735/X VGND VGND VPWR VPWR _4153_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1460 hold401/X VGND VGND VPWR VPWR _4133_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1471 hold421/X VGND VGND VPWR VPWR _5417_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1482 hold269/X VGND VGND VPWR VPWR _5558_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 _6899_/Q VGND VGND VPWR VPWR hold279/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5197__S _5199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput309 _3965_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5226__A _5226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4102__A0 _3616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3456__A2 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5850__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6810_ _6816_/CLK _6810_/D fanout446/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _6803_/CLK _6741_/D fanout442/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3953_ _7159_/Q _6811_/Q _6815_/Q VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6672_ _7128_/CLK _6672_/D fanout468/X VGND VGND VPWR VPWR _7226_/A sky130_fd_sc_hd__dfrtp_1
X_3884_ _3879_/B _3853_/S _3883_/X _3927_/A1 VGND VGND VPWR VPWR _6435_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5623_ _5623_/A VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__inv_2
XFILLER_176_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2744_A _6950_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5554_ _5554_/A0 _5563_/A1 _5559_/S VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3863__B _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4505_ _4643_/D _4643_/C VGND VGND VPWR VPWR _4917_/C sky130_fd_sc_hd__and2_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5485_ _5485_/A0 _5575_/A1 hold17/A VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6455__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7224_ _7224_/A VGND VGND VPWR VPWR _7224_/X sky130_fd_sc_hd__clkbuf_2
X_4436_ _4492_/B _4500_/B _4649_/B VGND VGND VPWR VPWR _4560_/C sky130_fd_sc_hd__a21o_2
XFILLER_132_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6330__A1 _6716_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6330__B2 _6573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4367_ _4420_/A _4420_/C _4461_/B VGND VGND VPWR VPWR _4368_/B sky130_fd_sc_hd__a21bo_4
X_7155_ _7180_/CLK _7155_/D fanout448/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5570__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3695__A2 _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _5228_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3318_ _3355_/A _3390_/B VGND VGND VPWR VPWR _3549_/B sky130_fd_sc_hd__nand2_8
X_6106_ _7104_/Q _6008_/X _6016_/X _7040_/Q VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__a22o_1
X_7086_ _7086_/CLK _7086_/D fanout470/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfstp_2
X_4298_ hold64/X _5184_/B hold9/A VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__and3_1
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6094__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6037_ _6933_/Q _5980_/X _5990_/X _7053_/Q VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a22o_1
X_3249_ hold61/X _3249_/A1 _3998_/S VGND VGND VPWR VPWR _3249_/X sky130_fd_sc_hd__mux2_4
XFILLER_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3447__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5841__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _7131_/CLK _6939_/D fanout452/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6414__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_csclk _3955_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold590 hold590/A VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5480__S hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6085__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3438__A2 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5832__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1290 _6709_/Q VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4938__A2 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3610__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5899__B1 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6707__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5270_ _5270_/A0 _5549_/A1 _5271_/S VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6312__A1 _6587_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4221_ _6678_/Q _6679_/Q _6681_/Q VGND VGND VPWR VPWR _4222_/C sky130_fd_sc_hd__nor3_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2908 _6684_/Q VGND VGND VPWR VPWR _3917_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5390__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2919 _7158_/Q VGND VGND VPWR VPWR _5644_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2325_A _6853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4152_ _4152_/A _5569_/B VGND VGND VPWR VPWR _4157_/S sky130_fd_sc_hd__and2_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4083_ _6681_/Q _4107_/B VGND VGND VPWR VPWR _4091_/S sky130_fd_sc_hd__nand2_8
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3204__A _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5823__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4985_ _5135_/A _5061_/B _4985_/C _4985_/D VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__5051__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5051__B2 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2861_A _6678_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6724_ _6735_/CLK _6724_/D fanout442/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfstp_2
X_3936_ _6823_/Q input80/X _3971_/B VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3601__A2 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_6655_ _3958_/A1 _6655_/D _6422_/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5565__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3867_ _3867_/A1 _3868_/B _3866_/Y _6446_/Q VGND VGND VPWR VPWR _3867_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6000__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5606_ _6491_/Q _5604_/Y _5606_/S VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_A _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6586_ _6786_/CLK _6586_/D fanout435/X VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfstp_4
X_3798_ _6933_/Q _5353_/A _5236_/C _3972_/A _3797_/X VGND VGND VPWR VPWR _3801_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ _5537_/A0 _5537_/A1 _5540_/S VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1160_A _6596_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5106__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5468_ _5468_/A0 _5549_/A1 _5469_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6303__B2 _6453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7207_ _7207_/A VGND VGND VPWR VPWR _7207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4419_ _4955_/A _4955_/B _4936_/B VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__and3_2
XFILLER_87_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5399_ hold413/X hold275/X _5406_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3668__A2 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7138_ _7139_/CLK _7138_/D fanout472/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout366 hold71/X VGND VGND VPWR VPWR _5568_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout377 hold95/X VGND VGND VPWR VPWR _5277_/A1 sky130_fd_sc_hd__buf_8
XFILLER_143_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout388 _5527_/A1 VGND VGND VPWR VPWR _5194_/A1 sky130_fd_sc_hd__buf_12
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7069_ _7073_/CLK _7069_/D fanout445/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout399 hold275/X VGND VGND VPWR VPWR _5543_/A1 sky130_fd_sc_hd__buf_12
XFILLER_101_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A wb_adr_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1961_A _6964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5475__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input73_A pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5207__C _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4856__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__A2 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6058__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5805__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3959__A _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4770_/A _4770_/B VGND VGND VPWR VPWR _5138_/C sky130_fd_sc_hd__and2_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3721_ _6862_/Q _5272_/A _4241_/A input53/X VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5385__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6440_ net399_2/A _6440_/D _6395_/X VGND VGND VPWR VPWR _6440_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3652_ _6641_/Q _4200_/A _4322_/A _6749_/Q _3651_/X VGND VGND VPWR VPWR _3655_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6371_ _6684_/Q _6371_/A2 _6371_/B1 _4218_/Y _6370_/X VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3583_ _6904_/Q _5317_/A _5290_/A _6880_/Q _3567_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_4_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5322_ _5322_/A0 _5448_/A1 _5325_/S VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6297__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5253_ _5253_/A0 _5577_/A1 _5253_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2705 _6792_/Q VGND VGND VPWR VPWR hold811/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4847__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4204_ _4204_/A0 _5195_/A1 _4205_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
Xhold2716 hold784/X VGND VGND VPWR VPWR _5233_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2727 _5557_/X VGND VGND VPWR VPWR hold605/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5184_ _5226_/B _5184_/B _5220_/C VGND VGND VPWR VPWR _5190_/S sky130_fd_sc_hd__and3_4
Xhold2738 _5372_/X VGND VGND VPWR VPWR hold772/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2749 _4247_/X VGND VGND VPWR VPWR hold611/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6049__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4135_ _4135_/A0 _5237_/A1 _4139_/S VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4066_ _4066_/A0 _5534_/A1 _4070_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6221__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4968_ _4981_/B VGND VGND VPWR VPWR _4968_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__3586__A1 _6960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6707_ _6746_/CLK _6707_/D _6416_/A VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3586__B2 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3919_ _3919_/A1 _3969_/B _3919_/B1 VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__a21o_1
XANTENNA__5295__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4899_ _5034_/A _5100_/C VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__and2_1
XANTENNA_hold1375_A _6485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6638_ _6826_/CLK _6638_/D _6407_/A VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5308__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4212__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6569_ _7121_/CLK _6569_/D _6399_/A VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_4_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__C1 _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A1 _7136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__B2 _7104_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4122__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output277_A _6478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _6755_/Q _5681_/X _5935_/X _5936_/X _5939_/X VGND VGND VPWR VPWR _5940_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_93_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5871_ _6639_/Q _5655_/X _5662_/X _6584_/Q _5870_/X VGND VGND VPWR VPWR _5879_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6203__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4822_ _4729_/A _4698_/Y _4689_/Y VGND VGND VPWR VPWR _4822_/Y sky130_fd_sc_hd__o21ai_1
X_4753_ _4752_/X _4753_/B _5138_/B _4770_/B VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__and4b_1
X_3704_ _3704_/A _3704_/B _3704_/C VGND VGND VPWR VPWR _3737_/A sky130_fd_sc_hd__and3_2
X_4684_ _4684_/A _4722_/C VGND VGND VPWR VPWR _4688_/A sky130_fd_sc_hd__nand2_8
X_6423_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3635_ _6951_/Q _3291_/Y _5317_/A _6903_/Q _3634_/X VGND VGND VPWR VPWR _3636_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _3385_/Y hold999/A _6354_/S VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__mux2_1
X_3566_ _7112_/Q _5551_/A hold89/A _6715_/Q VGND VGND VPWR VPWR _3566_/X sky130_fd_sc_hd__a22o_2
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5305_ _5305_/A0 wire375/X _5307_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3740__A1 _6853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3497_ _3535_/A _3648_/A VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__nor2_8
X_6285_ _6606_/Q _5982_/X _6005_/X _6694_/Q VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2502 _5300_/X VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5236_ _6430_/B _5533_/B _5236_/C VGND VGND VPWR VPWR _5244_/S sky130_fd_sc_hd__and3b_4
Xhold2513 hold912/X VGND VGND VPWR VPWR _5345_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2524 _7074_/Q VGND VGND VPWR VPWR hold961/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5493__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2535 _7077_/Q VGND VGND VPWR VPWR hold915/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1801 _4199_/X VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2546 _6941_/Q VGND VGND VPWR VPWR hold900/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2557 _7021_/Q VGND VGND VPWR VPWR hold902/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1812 hold637/X VGND VGND VPWR VPWR _5194_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1823 _6924_/Q VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2568 _6981_/Q VGND VGND VPWR VPWR hold903/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5167_ _5167_/A1 _4836_/A _5135_/X _5156_/Y _5166_/X VGND VGND VPWR VPWR _5167_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2579 hold883/X VGND VGND VPWR VPWR _4052_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1834 _4042_/X VGND VGND VPWR VPWR hold880/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout475_A input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1845 hold993/X VGND VGND VPWR VPWR hold484/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4118_ _4118_/A0 _5580_/A1 hold58/A VGND VGND VPWR VPWR _4118_/X sky130_fd_sc_hd__mux2_1
Xhold1856 _6832_/Q VGND VGND VPWR VPWR hold464/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1867 hold478/X VGND VGND VPWR VPWR hold1867/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5098_ _5098_/A _5098_/B _5098_/C VGND VGND VPWR VPWR _5131_/B sky130_fd_sc_hd__and3_1
Xhold1878 hold490/X VGND VGND VPWR VPWR hold1878/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1889 hold885/X VGND VGND VPWR VPWR _4034_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ _4049_/A0 _5562_/A1 _4055_/S VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5720__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5484__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A mgmt_gpio_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__buf_8
XANTENNA__3495__B1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5787__A2 _5684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5220__C _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3798__B2 _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5229__A hold64/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire361 _4598_/A VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3972__A _3972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold408 hold408/A VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold419 hold419/A VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3420_ _7019_/Q _5443_/A _3315_/Y input9/X _3419_/X VGND VGND VPWR VPWR _3421_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5711__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3722__A1 _7014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3351_ hold62/X hold22/X VGND VGND VPWR VPWR _5226_/B sky130_fd_sc_hd__and2_4
XANTENNA__3722__B2 _6819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3346_/A _3338_/A VGND VGND VPWR VPWR _5272_/A sky130_fd_sc_hd__nor2_8
X_6070_ _7055_/Q _5990_/X _5996_/X _7047_/Q VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__a22o_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5475__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5021_ _5021_/A _5021_/B _5021_/C VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__and3_1
Xhold1108 _6715_/Q VGND VGND VPWR VPWR _4284_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1119 _6815_/Q VGND VGND VPWR VPWR _5217_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5227__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6972_ _7131_/CLK _6972_/D fanout453/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3212__A _7056_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5778__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3789__A1 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _6591_/Q _5679_/X _5915_/X _5917_/X _5922_/X VGND VGND VPWR VPWR _5923_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3789__B2 _6707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5854_ _7004_/Q _5666_/X _5689_/X _7084_/Q VGND VGND VPWR VPWR _5854_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4959_/B _4805_/B _5032_/A _5089_/A VGND VGND VPWR VPWR _4805_/X sky130_fd_sc_hd__and4b_1
X_5785_ _6969_/Q _5872_/B VGND VGND VPWR VPWR _5785_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5139__A _5139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4736_ _4955_/D _5150_/C VGND VGND VPWR VPWR _4736_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3410__B1 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5950__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4667_ _4590_/B _4662_/Y _4995_/A _4638_/B VGND VGND VPWR VPWR _4667_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5573__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6406_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__and2_1
Xhold920 hold920/A VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3618_ _3617_/X _3618_/A1 _3739_/S VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__mux2_1
Xhold931 hold931/A VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5702__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4598_ _4598_/A _4598_/B _4598_/C _4607_/B VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__nand4_2
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold942 hold942/A VGND VGND VPWR VPWR hold942/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3713__A1 _6894_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 hold953/A VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3713__B2 _6531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold964 hold964/A VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6337_ _6608_/Q _5982_/X _5987_/X _6731_/Q _6319_/X VGND VGND VPWR VPWR _6338_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3549_ _3553_/A _3549_/B VGND VGND VPWR VPWR _3977_/A sky130_fd_sc_hd__nor2_8
Xhold975 hold975/A VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold986 hold986/A VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold997 hold997/A VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ _6591_/Q _5985_/X _6012_/X _6749_/Q VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__a22o_1
Xhold2310 _6945_/Q VGND VGND VPWR VPWR hold749/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5466__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2321 _6849_/Q VGND VGND VPWR VPWR hold736/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2332 _4147_/X VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2343 _5493_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5219_ _5569_/B _5219_/B VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__and2_1
XFILLER_29_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ _6940_/Q _5980_/X _6019_/X _6988_/Q _6198_/X VGND VGND VPWR VPWR _6204_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2354 hold609/X VGND VGND VPWR VPWR _5310_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2365 _5449_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1620 _7052_/Q VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1505_A _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1631 _5224_/X VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2376 _5458_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2387 _4297_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1642 hold537/X VGND VGND VPWR VPWR _4191_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2398 _5502_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1653 _5197_/X VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5218__A1 _5534_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1664 hold575/X VGND VGND VPWR VPWR _4295_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6417__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1675 _7084_/Q VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1686 _5274_/X VGND VGND VPWR VPWR hold230/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1697 hold238/X VGND VGND VPWR VPWR _5242_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5769__A2 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6194__A2 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__B1 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5941__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3952__A1 _6812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5483__S hold17/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4099__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5457__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3468__B1 _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5209__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4128__A _4128_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3640__B1 _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6185__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4196__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5570_ _5570_/A0 _5579_/A1 _5577_/S VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5932__A2 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4596_/A _4917_/D VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__nand2_2
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5393__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold205 hold205/A VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4452_ _4483_/B _4598_/C VGND VGND VPWR VPWR _4625_/B sky130_fd_sc_hd__and2_1
Xhold216 hold216/A VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold227 _4006_/X VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold238 hold238/A VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4499__A2 _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold249 hold249/A VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5696__A1 _6869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5696__B2 _6901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3403_ _6979_/Q _5398_/A _3988_/A _6477_/Q _3393_/X VGND VGND VPWR VPWR _3403_/X
+ sky130_fd_sc_hd__a221o_1
X_7171_ _7179_/CLK _7171_/D fanout443/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
X_4383_ _4717_/A _4713_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__nand2_4
XANTENNA__4310__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3207__A _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _7137_/Q _5977_/X _6017_/X _7073_/Q _6121_/X VGND VGND VPWR VPWR _6129_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3347_/A _3563_/B VGND VGND VPWR VPWR _5461_/A sky130_fd_sc_hd__nor2_8
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5448__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _7118_/Q _5978_/X _6014_/X _6990_/Q _6052_/X VGND VGND VPWR VPWR _6054_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3459__B1 _5290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3265_ hold60/X _3840_/A _6657_/Q VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__mux2_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4932_/Y _4964_/X _5003_/X _5139_/A _5004_/B2 VGND VGND VPWR VPWR _6764_/D
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4120__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3196_ _5611_/A VGND VGND VPWR VPWR _5610_/A sky130_fd_sc_hd__inv_2
XFILLER_66_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6963_/CLK _6955_/D fanout464/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5568__S _5568_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5906_ _6646_/Q _5668_/X _5684_/X _6606_/Q VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6886_ _7084_/CLK _6886_/D fanout444/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3631__B1 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ _7165_/Q _5836_/X _6341_/S VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__A2 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4187__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5923__A2 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5768_ _6944_/Q _5658_/X _5687_/X _6920_/Q VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3934__A1 input90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4719_ _4719_/A _4719_/B VGND VGND VPWR VPWR _4719_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ _6853_/Q _5651_/X _5668_/X _7053_/Q _5698_/X VGND VGND VPWR VPWR _5699_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold750 hold750/A VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold761 hold761/A VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold772 hold772/A VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold794 _5216_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5439__A1 _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2140 _5445_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6100__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2151 _6733_/Q VGND VGND VPWR VPWR hold550/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2162 _4296_/X VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2173 _6474_/Q VGND VGND VPWR VPWR hold761/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input138_A wb_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2184 _5451_/X VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2195 _4153_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1450 _7062_/Q VGND VGND VPWR VPWR hold267/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1461 _4133_/X VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1472 _5417_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 _5558_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1494 hold279/X VGND VGND VPWR VPWR _5315_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5478__S _5478_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3622__B1 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6313__D _6313_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4178__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5914__A2 _5673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3925__A1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5226__B _5226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4653__A2 _4693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5850__A1 _6948_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5388__S _5388_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6740_ _6803_/CLK _6740_/D fanout442/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3952_ _7157_/Q _6812_/Q _6815_/Q VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6671_ _7128_/CLK _6671_/D fanout468/X VGND VGND VPWR VPWR _7225_/A sky130_fd_sc_hd__dfrtp_1
X_3883_ _6468_/Q _6437_/Q _3852_/B VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6158__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4169__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5622_ _5604_/Y _5622_/A1 _7151_/Q VGND VGND VPWR VPWR _5623_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5905__A2 _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5553_ _5553_/A0 _5580_/A1 _5559_/S VGND VGND VPWR VPWR _5553_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4504_ _4506_/A _4643_/D VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__and2_1
XANTENNA_hold2737_A _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6315__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5484_ _5484_/A0 _5529_/A1 hold17/A VGND VGND VPWR VPWR _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _7223_/A VGND VGND VPWR VPWR _7223_/X sky130_fd_sc_hd__clkbuf_2
X_4435_ _4649_/B _4492_/B _4500_/B VGND VGND VPWR VPWR _4560_/B sky130_fd_sc_hd__nand3_4
XANTENNA__7182__CLK _7184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6330__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _7180_/CLK _7154_/D fanout448/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_4
X_4366_ _4701_/A _4365_/B _4917_/A VGND VGND VPWR VPWR _4420_/C sky130_fd_sc_hd__a21o_1
XFILLER_116_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6105_ _7128_/Q _5973_/X _5988_/X _6872_/Q _6104_/X VGND VGND VPWR VPWR _6105_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3317_ _3355_/A _3390_/B VGND VGND VPWR VPWR _5220_/B sky130_fd_sc_hd__and2_4
X_7085_ _7094_/CLK _7085_/D fanout453/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfstp_2
X_4297_ _4297_/A0 _5189_/A1 _4297_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout388_A _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _7133_/Q _5977_/X _5998_/X _6885_/Q _6035_/X VGND VGND VPWR VPWR _6039_/C
+ sky130_fd_sc_hd__a221o_1
X_3248_ hold60/X _6657_/Q _3247_/Y VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5298__S _5298_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _6996_/CLK _6938_/D fanout462/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6149__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6869_ _7063_/CLK _6869_/D fanout461/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_168_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6430__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6321__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4332__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold580 hold580/A VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold591 hold591/A VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4883__A2 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6085__B2 _6983_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1280 _5303_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1291 _4277_/X VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5899__B2 _6531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3374__A2 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6312__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4220_ _6682_/Q _4220_/B VGND VGND VPWR VPWR _5139_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__4323__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2909 _6658_/Q VGND VGND VPWR VPWR _3199_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4151_ _4151_/A0 _5189_/A1 _4151_/S VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2220_A _6986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4087__A0 _3616_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4082_ _4082_/A0 _5189_/A1 _4082_/S VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_0_csclk_A _6549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4984_ _5069_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _4985_/D sky130_fd_sc_hd__and3_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3220__A _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5051__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6723_ _6735_/CLK _6723_/D fanout442/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_4
X_3935_ _3204_/Y input82/X _3971_/B VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_8
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6654_ _3940_/A1 _6654_/D _6421_/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3866_ _3868_/B _3869_/A VGND VGND VPWR VPWR _3866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5605_ _5610_/A _5647_/B VGND VGND VPWR VPWR _5605_/Y sky130_fd_sc_hd__nand2_1
X_6585_ _6794_/CLK _6585_/D fanout434/X VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3797_ _6789_/Q _3427_/Y _5169_/A _6769_/Q VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ _7095_/Q _5536_/A1 _5541_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3365__A2 _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5467_ _5467_/A0 _5584_/A1 _5469_/S VGND VGND VPWR VPWR _5467_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6303__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7206_ _7206_/A VGND VGND VPWR VPWR _7206_/X sky130_fd_sc_hd__buf_2
XANTENNA__4314__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4418_ _4917_/A _4461_/B VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5398_ _5398_/A _5569_/B VGND VGND VPWR VPWR _5406_/S sky130_fd_sc_hd__and2_4
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7137_ _7137_/CLK _7137_/D fanout470/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4197__S _4199_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4349_ _4574_/A _4637_/D VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__nand2_8
XFILLER_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout367 hold1053/X VGND VGND VPWR VPWR hold1054/A sky130_fd_sc_hd__clkbuf_2
Xfanout378 _5529_/A1 VGND VGND VPWR VPWR _5583_/A1 sky130_fd_sc_hd__buf_8
XFILLER_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7068_ _7132_/CLK _7068_/D fanout451/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout389 _5536_/A1 VGND VGND VPWR VPWR _5527_/A1 sky130_fd_sc_hd__buf_12
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6019_ _6019_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _6019_/X sky130_fd_sc_hd__and3_4
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input66_A mgmt_gpio_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5491__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4305__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output222_A _3945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3959__B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6445__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _6958_/Q _5380_/A _4182_/A _6625_/Q _3719_/X VGND VGND VPWR VPWR _3725_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _6887_/Q _5299_/A _4316_/A _6744_/Q VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2170_A _6592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6370_ _6686_/Q _6370_/A2 _6370_/B1 _6685_/Q VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5741__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3582_ _6690_/Q _4250_/A _4262_/A _6700_/Q _3581_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5321_ _5321_/A0 _5537_/A1 _5325_/S VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2435_A _6741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5252_ _5252_/A0 _5549_/A1 _5253_/S VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6510__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4847__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2706 hold811/X VGND VGND VPWR VPWR _5188_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4203_ hold540/X _5194_/A1 _4205_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
Xhold2717 _5233_/X VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5183_ _5183_/A0 _5189_/A1 _5183_/S VGND VGND VPWR VPWR _5183_/X sky130_fd_sc_hd__mux2_1
Xhold2728 _6824_/Q VGND VGND VPWR VPWR hold541/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3215__A _7032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6049__A1 _6958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2739 _6869_/Q VGND VGND VPWR VPWR hold679/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4134_ _4134_/A _5220_/C VGND VGND VPWR VPWR _4139_/S sky130_fd_sc_hd__and2_2
XFILLER_95_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4065_ _4065_/A _5569_/B VGND VGND VPWR VPWR _4070_/S sky130_fd_sc_hd__and2_2
XFILLER_37_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4967_ _4595_/B _4476_/X _4522_/B VGND VGND VPWR VPWR _4981_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5576__S _5577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3918_ _3918_/A1 _3969_/B _3918_/B1 VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__a21o_1
X_6706_ _6945_/CLK _6706_/D _6413_/A VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3586__A2 _5380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4898_ _4898_/A _4898_/B VGND VGND VPWR VPWR _4902_/A sky130_fd_sc_hd__and2_1
XFILLER_177_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6637_ _6760_/CLK _6637_/D _6433_/A VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_4
X_3849_ _6654_/Q _3904_/A VGND VGND VPWR VPWR _3850_/S sky130_fd_sc_hd__nand2_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4535__A1 _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6568_ _7191_/CLK _6568_/D VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5732__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5519_ _5519_/A0 _5582_/A1 _5523_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6499_ _7125_/CLK _6499_/D fanout469/X VGND VGND VPWR VPWR _7220_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3510__A2 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6468__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5799__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input120_A wb_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6212__A1 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5486__S hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4774__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__A2 _3295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5723__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5515__A _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7198__RESET_B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _6530_/Q _5653_/X _5689_/X _6624_/Q VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6203__A1 _7036_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6203__B2 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4821_ _4676_/Y _4688_/A _4691_/Y _4812_/Y VGND VGND VPWR VPWR _4821_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5396__S _5397_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2385_A _6726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3568__A2 _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4752_ _4804_/A _4683_/Y _4750_/X _4751_/X VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3703_ _3703_/A _3703_/B _3703_/C _3703_/D VGND VGND VPWR VPWR _3704_/C sky130_fd_sc_hd__nor4_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4683_ _4683_/A _4683_/B VGND VGND VPWR VPWR _4683_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6422_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
XFILLER_162_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5714__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3634_ _6651_/Q _4212_/A _4176_/A _6621_/Q VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5190__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6353_ _3422_/Y hold995/A _6354_/S VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__mux2_1
X_3565_ _6856_/Q _5263_/A _4092_/A _6551_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5425__A _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5304_ _5304_/A0 hold95/X _5307_/S VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3740__A2 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6284_ _6689_/Q _5980_/X _6008_/X _6739_/Q VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3496_ _3550_/A _3549_/B VGND VGND VPWR VPWR _4164_/A sky130_fd_sc_hd__nor2_4
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5235_ _5235_/A0 hold39/X hold48/X VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__mux2_1
Xhold2503 _6965_/Q VGND VGND VPWR VPWR hold922/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2514 _5345_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2525 hold961/X VGND VGND VPWR VPWR _5512_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2536 hold915/X VGND VGND VPWR VPWR _5516_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2547 _5363_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1802 _6625_/Q VGND VGND VPWR VPWR hold530/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1813 _5194_/X VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5166_ _5145_/Y _5165_/Y _5140_/X VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__o21a_1
Xhold2558 _5453_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1824 hold323/X VGND VGND VPWR VPWR _5343_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2569 hold903/X VGND VGND VPWR VPWR _5408_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1835 hold880/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ _4117_/A0 _5561_/A1 hold58/A VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
Xhold1846 hold484/X VGND VGND VPWR VPWR hold1846/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5859__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1857 hold464/X VGND VGND VPWR VPWR _5240_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1868 _7212_/A VGND VGND VPWR VPWR hold570/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5097_ _4569_/C _4968_/Y _4542_/Y VGND VGND VPWR VPWR _5098_/C sky130_fd_sc_hd__o21a_1
Xhold1879 _7056_/Q VGND VGND VPWR VPWR hold790/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4048_ _4048_/A0 _5579_/A1 _4055_/S VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5999_ _6014_/A _6019_/C _6007_/C VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__and3_4
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5953__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1652_A _6800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5181__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5335__A _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3731__A2 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input168_A wb_sel_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6130__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput290 _6482_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3495__A1 _7081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_4
XFILLER_181_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input29_A mask_rev_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3798__A2 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6197__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5944__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5229__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7061_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire362 _3861_/Y VGND VGND VPWR VPWR _3868_/B sky130_fd_sc_hd__clkbuf_2
Xhold409 _5541_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5172__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5245__A _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3722__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3350_ _3354_/A _3535_/A VGND VGND VPWR VPWR _5497_/A sky130_fd_sc_hd__nor2_8
XFILLER_152_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk _6549_/CLK VGND VGND VPWR VPWR _6835_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6121__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3281_ hold79/X _3309_/A VGND VGND VPWR VPWR _3338_/A sky130_fd_sc_hd__nand2_8
XFILLER_140_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _4993_/A _4727_/A _5001_/A VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__o21ai_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _4284_/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6971_ _7131_/CLK _6971_/D fanout452/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5922_ _6586_/Q _5662_/X _5919_/X _5921_/X VGND VGND VPWR VPWR _5922_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3789__A2 _5335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_16
X_5853_ _6996_/Q _5929_/B _5686_/X _7012_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4804_ _4804_/A _4948_/A VGND VGND VPWR VPWR _5032_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5784_ _6857_/Q _5651_/X _5685_/X _7073_/Q _5783_/X VGND VGND VPWR VPWR _5792_/A
+ sky130_fd_sc_hd__a221o_1
X_4735_ _4955_/D _4735_/B VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4666_ _4666_/A _5026_/C VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__nand2_8
XFILLER_190_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6405_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6405_/X sky130_fd_sc_hd__and2_1
XANTENNA__3882__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3617_ _6776_/Q _3616_/Y _3738_/S VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5163__A1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold910 hold910/A VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4597_ _5033_/A _4724_/C VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__nand2_1
Xhold921 hold921/A VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold932 hold932/A VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold943 hold943/A VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4910__A1 _4655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6336_ _6552_/Q _5999_/X _6019_/X _6736_/Q _6335_/X VGND VGND VPWR VPWR _6338_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3713__A2 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold954 hold954/A VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1066_A _6617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3548_ _6905_/Q _5317_/A _3325_/Y _7041_/Q _3547_/X VGND VGND VPWR VPWR _3556_/B
+ sky130_fd_sc_hd__a221o_2
Xhold965 hold965/A VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold976 hold976/A VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold987 hold987/A VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold998 hold998/A VGND VGND VPWR VPWR hold998/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6267_ _6291_/A2 _6266_/X _6342_/S VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6112__B1 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2300 _4150_/X VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3479_ _3550_/A _3516_/B VGND VGND VPWR VPWR _4158_/A sky130_fd_sc_hd__nor2_8
Xhold2311 hold749/X VGND VGND VPWR VPWR _5367_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2322 hold736/X VGND VGND VPWR VPWR _5259_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5218_ _5218_/A0 _5534_/A1 hold24/X VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__mux2_1
Xhold2333 _6720_/Q VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7049__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6198_ _6900_/Q _5989_/X _6013_/X _7084_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
Xhold2344 _7082_/Q VGND VGND VPWR VPWR hold628/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1610 _6481_/Q VGND VGND VPWR VPWR hold513/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2355 _5310_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2366 _6926_/Q VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1621 hold386/X VGND VGND VPWR VPWR _5487_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1632 _6532_/Q VGND VGND VPWR VPWR hold523/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5149_ _5149_/A _5149_/B _5149_/C _5149_/D VGND VGND VPWR VPWR _5152_/A sky130_fd_sc_hd__and4_1
Xhold2377 _6982_/Q VGND VGND VPWR VPWR hold591/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2388 _6850_/Q VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1643 _4191_/X VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1654 _6699_/Q VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2399 _6785_/Q VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1665 _4295_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1676 hold405/X VGND VGND VPWR VPWR _5523_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1687 _6929_/Q VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1698 _6484_/Q VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6613__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__A1 _6907_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6656__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6103__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3468__A1 _7073_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4409__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4128__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3640__A1 _7055_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__B2 _6452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5917__B1 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4520_ _4523_/A _4638_/B VGND VGND VPWR VPWR _4655_/A sky130_fd_sc_hd__nand2_8
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ _4451_/A _4451_/B VGND VGND VPWR VPWR _4598_/C sky130_fd_sc_hd__and2_4
XFILLER_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5145__A1 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold217 hold217/A VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5696__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold239 _5242_/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3402_ _6883_/Q _5290_/A _3399_/X _3401_/X VGND VGND VPWR VPWR _3402_/X sky130_fd_sc_hd__a211o_1
X_7170_ _7184_/CLK _7170_/D fanout443/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4382_ _4717_/A _4713_/A VGND VGND VPWR VPWR _4751_/B sky130_fd_sc_hd__and2_4
XFILLER_171_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6121_ _7033_/Q _5986_/X _5988_/X _6873_/Q VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__a22o_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3346_/A _3354_/A VGND VGND VPWR VPWR _5281_/A sky130_fd_sc_hd__nor2_8
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6894_/Q _5989_/X _6015_/X _7014_/Q VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3264_ hold13/X VGND VGND VPWR VPWR _3429_/A sky130_fd_sc_hd__inv_2
XANTENNA__7142__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5003_ _5061_/A _4985_/Y _5005_/B _5002_/Y _4836_/A VGND VGND VPWR VPWR _5003_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3195_ _6490_/Q VGND VGND VPWR VPWR _6166_/S sky130_fd_sc_hd__inv_4
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _6963_/CLK _6954_/D fanout464/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_4
X_5905_ _3201_/Y _5872_/B _5677_/B VGND VGND VPWR VPWR _5905_/Y sky130_fd_sc_hd__a21oi_1
X_6885_ _7073_/CLK _6885_/D fanout444/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _5826_/Y _5835_/Y _6843_/Q _5678_/Y VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__o2bb2a_2
XANTENNA__5908__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5384__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5767_ _6896_/Q _5662_/X _5684_/X _6928_/Q _5766_/X VGND VGND VPWR VPWR _5770_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1183_A _6839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3395__B1 _5263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4718_ _4718_/A _4719_/A _4718_/C VGND VGND VPWR VPWR _4718_/X sky130_fd_sc_hd__and3_1
X_5698_ _7029_/Q _5655_/X _5678_/B _6965_/Q _5707_/B VGND VGND VPWR VPWR _5698_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4720_/C _4649_/B _4649_/C _4649_/D VGND VGND VPWR VPWR _4677_/A sky130_fd_sc_hd__nor4_4
XFILLER_162_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6333__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1350_A _6581_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold740 hold740/A VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold751 hold751/A VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold762 hold762/A VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold773 hold773/A VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold784 hold784/A VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6319_ _6706_/Q _5977_/X _5984_/X _6618_/Q VGND VGND VPWR VPWR _6319_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold795 hold795/A VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1615_A _6641_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2130 hold750/X VGND VGND VPWR VPWR _5435_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2141 _6522_/Q VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2152 hold550/X VGND VGND VPWR VPWR _4306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2163 _7218_/A VGND VGND VPWR VPWR hold937/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2174 hold761/X VGND VGND VPWR VPWR _3992_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1440 _5247_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2185 _6639_/Q VGND VGND VPWR VPWR hold756/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1451 hold267/X VGND VGND VPWR VPWR _5499_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2196 _6548_/Q VGND VGND VPWR VPWR hold707/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1462 _6488_/Q VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1473 _6728_/Q VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1484 _7004_/Q VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _5315_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6865__RESET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3622__A1 _7015_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input96_A usr1_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5375__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5494__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6324__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5226__C _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5850__A2 _5658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _6506_/Q input93/X _6820_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_4
XFILLER_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3613__A1 _7080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4810__B1 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6670_ _7125_/CLK _6670_/D fanout468/X VGND VGND VPWR VPWR _7224_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3882_ _6413_/A _6423_/B VGND VGND VPWR VPWR _3882_/X sky130_fd_sc_hd__and2_1
XFILLER_188_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5621_ _5621_/A VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__inv_2
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5366__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3377__B1 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5552_ _5552_/A0 _5561_/A1 _5559_/S VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4503_ _4637_/B _4808_/B _4701_/A VGND VGND VPWR VPWR _4643_/C sky130_fd_sc_hd__a21o_1
XANTENNA__5118__A1 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5483_ _5483_/A0 _5582_/A1 hold17/A VGND VGND VPWR VPWR _5483_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6315__B1 _6314_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3218__A _7008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7222_ _7222_/A VGND VGND VPWR VPWR _7222_/X sky130_fd_sc_hd__clkbuf_2
X_4434_ _4447_/B _4663_/D _4682_/A _4808_/B VGND VGND VPWR VPWR _4500_/B sky130_fd_sc_hd__and4_2
XFILLER_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7153_ _7180_/CLK _7153_/D fanout448/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_4
X_4365_ _4701_/A _4365_/B VGND VGND VPWR VPWR _4461_/B sky130_fd_sc_hd__xnor2_4
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6104_ _6960_/Q _5992_/X _6012_/X _7000_/Q _6103_/X VGND VGND VPWR VPWR _6104_/X
+ sky130_fd_sc_hd__a221o_1
X_3316_ _3686_/A hold30/X VGND VGND VPWR VPWR _5506_/A sky130_fd_sc_hd__nor2_8
X_7084_ _7084_/CLK _7084_/D fanout447/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_4
X_4296_ _4296_/A0 _5195_/A1 _4297_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6035_ _7109_/Q _5987_/X _5997_/X _6949_/Q VGND VGND VPWR VPWR _6035_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6094__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3247_ hold19/X _3862_/A VGND VGND VPWR VPWR _3247_/Y sky130_fd_sc_hd__nand2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5841__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3255__A_N _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6937_ _6977_/CLK _6937_/D fanout460/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6868_ _7107_/CLK _6868_/D fanout451/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6003__C1 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5357__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5819_ _6915_/Q _5670_/X _5682_/X _7043_/Q _5818_/X VGND VGND VPWR VPWR _5826_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6799_ _6809_/CLK _6799_/D fanout442/X VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6306__B1 _6004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold570 hold570/A VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold581 hold581/A VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold592 hold592/A VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input150_A wb_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6085__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4096__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5832__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1270 _6912_/Q VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5489__S _5496_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input11_A mask_rev_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1281 _6990_/Q VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1292 _6704_/Q VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5045__B1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5348__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3359__B1 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5899__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4422__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4020__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5520__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2046_A _7136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4150_ _4150_/A0 _5233_/A1 _4151_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6787__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4081_ _4081_/A0 _5233_/A1 _4082_/S VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5823__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5399__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4316__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4983_ _5103_/B _4983_/B _4983_/C VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__and3_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3598__B1 _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6722_ _7045_/CLK _6722_/D fanout444/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_2
X_3934_ _3203_/Y input90/X _3934_/S VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5339__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3865_ _6445_/Q _3870_/B VGND VGND VPWR VPWR _3869_/A sky130_fd_sc_hd__nor2_2
X_6653_ _6746_/CLK _6653_/D _6416_/A VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5604_ _6489_/Q _6491_/Q VGND VGND VPWR VPWR _5604_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4011__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6584_ _6786_/CLK _6584_/D fanout435/X VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfrtp_4
X_3796_ _6795_/Q _3319_/Y _5299_/A _6885_/Q _3795_/X VGND VGND VPWR VPWR _3801_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5535_ _5535_/A0 _5571_/A1 _5540_/S VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5466_ _5466_/A0 _5583_/A1 _5469_/S VGND VGND VPWR VPWR _5466_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4417_ _4947_/A _4417_/B VGND VGND VPWR VPWR _5150_/B sky130_fd_sc_hd__nand2_4
XFILLER_132_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5511__A1 hold95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5397_ _5397_/A0 _5568_/A1 _5397_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7136_ _7136_/CLK _7136_/D fanout468/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_4
X_4348_ _4574_/A _4637_/D VGND VGND VPWR VPWR _4576_/A sky130_fd_sc_hd__and2_4
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A debug_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout368 wire371/X VGND VGND VPWR VPWR _5549_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7067_ _7082_/CLK _7067_/D fanout464/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4078__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4279_ _4279_/A0 _5448_/A1 _4279_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
Xfanout379 _5529_/A1 VGND VGND VPWR VPWR _5448_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_74_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6018_ _6019_/B _6018_/B _6019_/C VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__and3_4
XANTENNA__5814__A2 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4002__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3761__B1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input59_A mgmt_gpio_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5502__A1 _5583_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3513__B1 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6058__A2 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4069__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5805__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4417__A _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6215__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4152__A _4152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3650_ _7087_/Q _5524_/A _4065_/A _6527_/Q _3649_/X VGND VGND VPWR VPWR _3655_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3581_ _6848_/Q _5254_/A _3521_/Y _6538_/Q VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5741__B2 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5320_ _5320_/A0 _5572_/A1 _5325_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5251_ _5251_/A0 wire375/X _5253_/S VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6297__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4202_ _4202_/A0 _5193_/A1 _4205_/S VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2428_A _7097_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5182_ _5182_/A0 _5195_/A1 _5183_/S VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__mux2_1
Xhold2707 _5188_/X VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2718 _6962_/Q VGND VGND VPWR VPWR hold623/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6966__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2729 hold541/X VGND VGND VPWR VPWR _5231_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6049__A2 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4133_ _4133_/A0 _5277_/A1 _4133_/S VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ _4064_/A0 hold71/X _4064_/S VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__mux2_1
XFILLER_110_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6221__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4966_ _4581_/X _4969_/B _4878_/Y _4491_/Y _4628_/Y VGND VGND VPWR VPWR _5074_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6705_ _6730_/CLK hold68/X _6413_/A VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__dfstp_2
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3917_ _3917_/A1 _3969_/B _3917_/B1 VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3440__C1 _3437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4897_ _4921_/B _4897_/B VGND VGND VPWR VPWR _4903_/C sky130_fd_sc_hd__nor2_1
XFILLER_149_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6636_ _6761_/CLK _6636_/D _6416_/A VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_2
X_3848_ _6470_/Q _6468_/Q _6654_/Q VGND VGND VPWR VPWR _3880_/S sky130_fd_sc_hd__and3_1
X_3779_ _6817_/Q hold64/A _5220_/B _4194_/A _6634_/Q VGND VGND VPWR VPWR _3779_/X
+ sky130_fd_sc_hd__a32o_1
X_6567_ _7191_/CLK _6567_/D VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5732__B2 _7055_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5518_ _5518_/A0 _5563_/A1 _5523_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
X_6498_ _7134_/CLK _6498_/D fanout469/X VGND VGND VPWR VPWR _7219_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_145_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5449_ _5449_/A0 _5584_/A1 _5451_/S VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4299__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7119_ _7135_/CLK _7119_/D fanout467/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1897_A _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7195__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input113_A wb_adr_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6385_/A3 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6212__A2 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4774__A2 _4688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5723__A1 _7014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5723__B2 _7054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3734__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5515__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3498__C1 _3495_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6346__B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6562__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6203__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4820_ _4820_/A _4820_/B _4820_/C VGND VGND VPWR VPWR _4834_/A sky130_fd_sc_hd__and3_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4214__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _5009_/A _4751_/B _4751_/C VGND VGND VPWR VPWR _4751_/X sky130_fd_sc_hd__and3_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3702_ _7022_/Q _5452_/A _5560_/A _7118_/Q _3701_/X VGND VGND VPWR VPWR _3703_/D
+ sky130_fd_sc_hd__a221o_4
X_4682_ _4682_/A _4717_/A VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__nand2_4
XFILLER_147_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3633_ _6975_/Q _5398_/A _5281_/A _6871_/Q _3632_/X VGND VGND VPWR VPWR _3636_/C
+ sky130_fd_sc_hd__a221o_1
X_6421_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
XANTENNA__5714__B2 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3564_ _7088_/Q _5524_/A _4170_/A _6617_/Q VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__a22o_1
X_6352_ _3462_/Y hold992/A _6354_/S VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5425__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5303_ _5303_/A0 _5303_/A1 _5307_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6611_/Q _5976_/B _5984_/X _6616_/Q _6282_/X VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3495_ _7081_/Q _5515_/A hold24/A _6810_/Q VGND VGND VPWR VPWR _3495_/X sky130_fd_sc_hd__a22o_4
XANTENNA__3226__A _6952_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6731__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5234_ _5234_/A0 _5583_/A1 hold48/X VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2504 hold922/X VGND VGND VPWR VPWR _5390_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2515 _7069_/Q VGND VGND VPWR VPWR hold907/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2526 _5512_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5165_ _5015_/X _5165_/B _5165_/C VGND VGND VPWR VPWR _5165_/Y sky130_fd_sc_hd__nand3b_1
Xhold2537 _5516_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2548 _6748_/Q VGND VGND VPWR VPWR hold554/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1803 hold530/X VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2559 _6891_/Q VGND VGND VPWR VPWR hold663/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1814 _6756_/Q VGND VGND VPWR VPWR hold396/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1825 _5343_/X VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1836 _6503_/Q VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4116_ hold57/X hold9/A VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__and2_2
XFILLER_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1847 _7187_/Q VGND VGND VPWR VPWR hold997/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5096_ _4611_/A _4981_/B _5095_/Y _4897_/B VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__a211oi_1
Xhold1858 _6813_/Q VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1869 hold570/X VGND VGND VPWR VPWR _4038_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4047_ _6430_/B _5317_/B _4047_/C VGND VGND VPWR VPWR _4055_/S sky130_fd_sc_hd__and3b_4
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4205__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6019_/A _6015_/B _6007_/C VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__and3_4
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5953__A1 _6534_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4949_ _5067_/A _5023_/A VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5953__B2 _6588_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3964__A0 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5705__A1 _6845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6619_ _6756_/CLK _6619_/D fanout441/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5335__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6435__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 _6797_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput291 _6483_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4692__A1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__A2 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4747__A2 _4714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5944__B2 _6772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3955__B1 _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5229__C hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3707__B1 _3389_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5245__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6121__A1 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3280_ _3429_/A hold46/X VGND VGND VPWR VPWR _3309_/A sky130_fd_sc_hd__nor2_8
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5880__B1 _6525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2126_A _7086_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6970_ _6994_/CLK _6970_/D fanout462/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6734__SET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5921_ _6537_/Q _5651_/X _5688_/X _6581_/Q _5920_/X VGND VGND VPWR VPWR _5921_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5852_ _7060_/Q _5668_/X _5684_/X _6932_/Q VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _5108_/B _5138_/C _4803_/C _4803_/D VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__and4_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _7009_/Q _5686_/X _5688_/X _6889_/Q VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2662_A _6960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4734_ _5011_/A _4664_/Y _4584_/Y VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3410__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4738_/B _5026_/C VGND VGND VPWR VPWR _4730_/B sky130_fd_sc_hd__and2_1
XFILLER_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6458__CLK _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5699__B1 _5668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6404_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6404_/X sky130_fd_sc_hd__and2_1
X_3616_ _3573_/X _3616_/B _3616_/C _3616_/D VGND VGND VPWR VPWR _3616_/Y sky130_fd_sc_hd__nand4b_4
Xhold900 hold900/A VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold911 hold911/A VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5163__A2 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4596_ _4596_/A _4934_/B VGND VGND VPWR VPWR _4880_/B sky130_fd_sc_hd__nand2_1
Xhold922 hold922/A VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6335_ _6756_/Q _5638_/X _6015_/X _6761_/Q VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_4
Xhold944 hold944/A VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3547_ _3547_/A1 _5236_/C _3431_/Y _7232_/A VGND VGND VPWR VPWR _3547_/X sky130_fd_sc_hd__a22o_2
Xhold955 hold955/A VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold966 hold966/A VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6112__A1 _7136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold988 hold988/A VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6266_ _6266_/A0 _6265_/X _6341_/S VGND VGND VPWR VPWR _6266_/X sky130_fd_sc_hd__mux2_1
X_3478_ _6857_/Q _5263_/A _4310_/A _6741_/Q VGND VGND VPWR VPWR _3478_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6112__B2 _7096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold999 hold999/A VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2301 _6608_/Q VGND VGND VPWR VPWR hold795/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2312 _5367_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2323 _7041_/Q VGND VGND VPWR VPWR hold720/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5217_ _5217_/A0 _5228_/A1 _5217_/S VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__mux2_1
Xhold2334 hold894/X VGND VGND VPWR VPWR _4290_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6197_ _7132_/Q _5973_/X _5998_/X _6892_/Q _6196_/X VGND VGND VPWR VPWR _6204_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1600 hold115/X VGND VGND VPWR VPWR _4270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_192_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2345 hold628/X VGND VGND VPWR VPWR _5521_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2356 _6525_/Q VGND VGND VPWR VPWR hold839/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1611 _4003_/X VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5871__B1 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2367 hold607/X VGND VGND VPWR VPWR _5346_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1622 _5487_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1633 hold523/X VGND VGND VPWR VPWR _4074_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5148_ _5148_/A _5148_/B _5148_/C VGND VGND VPWR VPWR _5149_/D sky130_fd_sc_hd__and3_1
Xhold2378 hold591/X VGND VGND VPWR VPWR _5409_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1644 _6734_/Q VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2389 hold622/X VGND VGND VPWR VPWR _5260_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1655 hold539/X VGND VGND VPWR VPWR _4265_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1666 _6799_/Q VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1677 _5523_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5079_ _4688_/B _4995_/B _5009_/Y _4688_/C VGND VGND VPWR VPWR _5080_/C sky130_fd_sc_hd__o22a_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1688 hold313/X VGND VGND VPWR VPWR _5349_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1699 _7221_/A VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6653__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4250__A _4250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6103__A1 _6952_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__B2 _6880_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4114__A0 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A mgmt_gpio_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3468__A2 _5506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5862__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2890 hold45/A VGND VGND VPWR VPWR _5078_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6116__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3640__A2 _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5917__A1 _6734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5917__B2 _6699_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4450_ _4450_/A _4450_/B VGND VGND VPWR VPWR _4451_/B sky130_fd_sc_hd__nor2_1
Xhold207 hold207/A VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold218 hold218/A VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold229 hold229/A VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3401_ _6907_/Q _5317_/A _5488_/A _7059_/Q _3400_/X VGND VGND VPWR VPWR _3401_/X
+ sky130_fd_sc_hd__a221o_1
X_4381_ _4701_/A _4917_/A VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__and2b_4
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3332_ _3544_/A _3764_/A VGND VGND VPWR VPWR _5299_/A sky130_fd_sc_hd__nor2_8
X_6120_ _6977_/Q _5976_/B _6008_/X _7105_/Q _6119_/X VGND VGND VPWR VPWR _6120_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4105__A0 _3422_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _7022_/Q _5971_/X _5987_/X _7110_/Q _6050_/X VGND VGND VPWR VPWR _6054_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3263_ _3262_/X hold12/X _3998_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A2 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__B1 _5686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5002_ _5114_/B _5002_/B _5124_/C VGND VGND VPWR VPWR _5002_/Y sky130_fd_sc_hd__nand3_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3194_ _7155_/Q VGND VGND VPWR VPWR _5637_/A sky130_fd_sc_hd__clkinv_4
XFILLER_94_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7182__RESET_B fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6953_ _7121_/CLK _6953_/D _6399_/A VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_4
X_5904_ _5925_/A2 _6342_/S _5902_/X _5903_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__o22a_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ _7091_/CLK _6884_/D fanout452/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3631__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A _5835_/B _5835_/C _5835_/D VGND VGND VPWR VPWR _5835_/Y sky130_fd_sc_hd__nor4_1
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6030__B1 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5766_ _6848_/Q _5653_/X _5656_/X _6984_/Q VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3395__A1 _7115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4717_ _4717_/A _4717_/B _4726_/B VGND VGND VPWR VPWR _4727_/A sky130_fd_sc_hd__and3_2
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5697_ _6925_/Q _5684_/X _5694_/X _5696_/X VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__a211o_1
XFILLER_163_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4648_ _4682_/A _4712_/B VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nand2_4
XFILLER_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold730 hold730/A VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold741 hold741/A VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4579_ _4751_/B _4579_/B _4693_/B VGND VGND VPWR VPWR _4889_/B sky130_fd_sc_hd__nand3_2
Xhold752 hold752/A VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold763 hold763/A VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold774 hold774/A VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6318_ _6593_/Q _5985_/X _5994_/X _6638_/Q VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold785 hold785/A VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold796 hold796/A VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6249_ _6590_/Q _5985_/X _5994_/X _6635_/Q _6243_/X VGND VGND VPWR VPWR _6249_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2120 _5565_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2131 _5435_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2142 hold602/X VGND VGND VPWR VPWR _4062_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5844__B1 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2153 _4306_/X VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2164 hold937/X VGND VGND VPWR VPWR _4023_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1430 hold203/X VGND VGND VPWR VPWR _4244_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2175 _3992_/X VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1441 _7230_/A VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2186 hold756/X VGND VGND VPWR VPWR _4201_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2197 hold707/X VGND VGND VPWR VPWR _4093_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1452 _5499_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1463 _7043_/Q VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1474 hold109/X VGND VGND VPWR VPWR _4300_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 hold319/X VGND VGND VPWR VPWR _5433_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7094_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1496 _7124_/Q VGND VGND VPWR VPWR hold338/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3622__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6021__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input89_A spimemio_flash_io2_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6324__A1 _6633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6324__B2 _6534_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3689__A2 _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output245_A _3942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_29_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7125_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6260__B1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3950_ _6507_/Q _3950_/A1 _6818_/Q VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4810__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3613__A2 _5515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4810__B2 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3881_ _6817_/Q _6864_/Q _3881_/C VGND VGND VPWR VPWR _3881_/Y sky130_fd_sc_hd__nor3_4
XFILLER_189_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5620_ _5619_/Y _5685_/A _5620_/S VGND VGND VPWR VPWR _5621_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3377__A1 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _5551_/A _5578_/B VGND VGND VPWR VPWR _5559_/S sky130_fd_sc_hd__and2_4
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4498_/X _4499_/Y _4500_/Y _4501_/X VGND VGND VPWR VPWR _4917_/B sky130_fd_sc_hd__a2bb2oi_2
XANTENNA_hold2458_A _6820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6315__A1 _6528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5118__A2 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5482_ _5482_/A0 _5536_/A1 hold17/A VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7221_ _7221_/A VGND VGND VPWR VPWR _7221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4433_ _4663_/D _4451_/A VGND VGND VPWR VPWR _4486_/A sky130_fd_sc_hd__nor2_8
XANTENNA__3933__S _3934_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7152_ _7179_/CLK _7152_/D fanout447/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_99_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4364_ _4360_/A _4360_/B _4362_/B _4362_/A VGND VGND VPWR VPWR _4368_/A sky130_fd_sc_hd__a22o_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6079__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6103_ _6952_/Q _5997_/X _6004_/X _6880_/Q VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__a22o_1
X_3315_ _3354_/A _3764_/B VGND VGND VPWR VPWR _3315_/Y sky130_fd_sc_hd__nor2_8
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4295_ _4295_/A0 _5194_/A1 _4297_/S VGND VGND VPWR VPWR _4295_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7083_ _7126_/CLK _7083_/D fanout453/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3234__A _6888_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6034_ _7117_/Q _5978_/X _5992_/X _6957_/Q _6033_/X VGND VGND VPWR VPWR _6039_/B
+ sky130_fd_sc_hd__a221o_1
X_3246_ _6470_/Q _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3857_/B sky130_fd_sc_hd__nor3_4
XFILLER_100_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6264__B _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5054__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _6936_/CLK _6936_/D fanout463/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout443_A fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4801__A1 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6867_ _7091_/CLK _6867_/D fanout452/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6853__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6003__B1 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5818_ _7003_/Q _5666_/X _5674_/X _6875_/Q VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6798_ _6809_/CLK _6798_/D fanout433/X VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_157_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5749_ _6839_/Q _5678_/Y _5740_/X _5748_/X _6166_/S VGND VGND VPWR VPWR _5749_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4868__A1 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold560 hold560/A VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold571 _4038_/X VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 hold582/A VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input143_A wb_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5293__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1260 hold302/X VGND VGND VPWR VPWR _5358_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1271 hold382/X VGND VGND VPWR VPWR _5330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1282 hold205/X VGND VGND VPWR VPWR _5418_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1293 hold157/X VGND VGND VPWR VPWR _4271_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5045__B2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3359__B2 _7036_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4859__A1 _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__1153_ clkbuf_0__1153_/X VGND VGND VPWR VPWR _4112_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_114_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4080_ hold190/X _5527_/A1 _4082_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5284__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6233__B1 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6756__RESET_B fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4982_ _4569_/B _4570_/A _4570_/B _4570_/D _4968_/Y VGND VGND VPWR VPWR _4983_/C
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3598__A1 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6721_ _6786_/CLK _6721_/D fanout435/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_4
X_3933_ _3202_/Y input92/X _3934_/S VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_4
XFILLER_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3598__B2 _6772_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4795__B1 _4713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6652_ _6756_/CLK _6652_/D fanout441/X VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3864_ _3904_/A _3863_/Y _3868_/B VGND VGND VPWR VPWR _3870_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__6989__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5603_ _3193_/Y _5601_/B _5602_/Y VGND VGND VPWR VPWR _5603_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6583_ _6756_/CLK _6583_/D fanout441/X VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfrtp_4
X_3795_ input43/X _4047_/C _4241_/A input52/X VGND VGND VPWR VPWR _3795_/X sky130_fd_sc_hd__a22o_4
XFILLER_191_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5534_ _5534_/A0 _5534_/A1 _5540_/S VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _5465_/A0 _5582_/A1 _5469_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7204_ _3950_/A1 _7204_/D _6346_/B VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4719_/A _4595_/B VGND VGND VPWR VPWR _4417_/B sky130_fd_sc_hd__nand2_8
XFILLER_99_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5396_ _5396_/A0 _5549_/A1 _5397_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
X_7135_ _7135_/CLK _7135_/D fanout470/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3522__B2 _6539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4347_ _4917_/A _4701_/A VGND VGND VPWR VPWR _4682_/A sky130_fd_sc_hd__and2_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout393_A _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1139_A _7127_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout369 hold35/X VGND VGND VPWR VPWR _5567_/A1 sky130_fd_sc_hd__clkbuf_16
X_7066_ _7130_/CLK _7066_/D fanout462/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4278_ _4278_/A0 hold43/X _4279_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5275__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6017_ _6017_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _6017_/X sky130_fd_sc_hd__and3_4
X_3229_ _6928_/Q VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6224__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3955_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A1 _6792_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3589__B2 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6919_ _7063_/CLK _6919_/D fanout460/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold390 hold390/A VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5266__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4417__B _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1090 _3536_/Y VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4152__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ _3580_/A _3580_/B _3580_/C _3580_/D VGND VGND VPWR VPWR _3616_/B sky130_fd_sc_hd__nor4_2
XANTENNA__5741__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6491__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5250_ _5250_/A0 hold95/X _5253_/S VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4201_ _4201_/A0 _5237_/A1 _4205_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2708 _7208_/A VGND VGND VPWR VPWR hold652/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5181_ _5181_/A0 _5194_/A1 _5183_/S VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__mux2_1
Xhold2719 hold623/X VGND VGND VPWR VPWR _5386_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4132_ _4132_/A0 _5233_/A1 _4133_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5257__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4063_ _4063_/A0 _5567_/A1 _4064_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6206__B1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4965_ _4561_/X _4965_/B _4965_/C VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__and3b_1
X_6704_ _6730_/CLK _6704_/D _6413_/A VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_2
X_3916_ _6490_/Q _3909_/X _3912_/B _3915_/Y _3916_/B2 VGND VGND VPWR VPWR _6492_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3440__B1 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4783__A3 _4417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4896_ _5117_/A _4924_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__nand2_2
XFILLER_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3991__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6635_ _6826_/CLK _6635_/D _6407_/A VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _6654_/Q _3847_/B VGND VGND VPWR VPWR _3852_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _7191_/CLK _6566_/D VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout406_A _5317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3778_ _7061_/Q _5497_/A _3539_/Y _6530_/Q _3777_/X VGND VGND VPWR VPWR _3783_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5732__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3743__A1 _6997_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6621__SET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5517_ _5517_/A0 _5571_/A1 _5523_/S VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6497_ _6828_/CLK _6497_/D fanout469/X VGND VGND VPWR VPWR _7218_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1256_A _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ _5448_/A0 _5448_/A1 _5451_/S VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5496__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5379_ _5379_/A0 _5568_/A1 _5379_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7118_ _7124_/CLK _7118_/D fanout467/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5248__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7049_ _7137_/CLK _7049_/D _6411_/A VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5799__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A wb_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5723__A2 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input71_A mgmt_gpio_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5487__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3498__B1 _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5239__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3670__B1 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5411__A1 _5582_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4750_ _4637_/C _4719_/A _4683_/Y _4749_/X VGND VGND VPWR VPWR _4750_/X sky130_fd_sc_hd__a31o_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5962__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3701_ input44/X _4047_/C _5263_/A _6854_/Q VGND VGND VPWR VPWR _3701_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4681_ _4682_/A _4717_/A VGND VGND VPWR VPWR _4722_/C sky130_fd_sc_hd__and2_2
XFILLER_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6420_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
XFILLER_174_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3632_ _6863_/Q _5272_/A _3319_/Y _6797_/Q VGND VGND VPWR VPWR _3632_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5714__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6351_ _6351_/A0 _6351_/A1 _6354_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
X_3563_ _3563_/A _3563_/B VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5302_ _5302_/A0 _5527_/A1 _5307_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4102__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2538_A _7053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6282_ _6537_/Q _5983_/X _5986_/X _6641_/Q VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__a22o_1
X_3494_ input30/X _3307_/Y _4200_/A _6643_/Q _3493_/X VGND VGND VPWR VPWR _3499_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5478__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5233_ _5233_/A0 _5233_/A1 hold48/X VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3489__B1 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3941__S _6459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2505 _5390_/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2705_A _6792_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2516 hold907/X VGND VGND VPWR VPWR _5507_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4150__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2527 _7109_/Q VGND VGND VPWR VPWR hold890/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2538 _7053_/Q VGND VGND VPWR VPWR hold892/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _5011_/A _4691_/Y _4818_/A _5163_/X VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__o211a_1
Xhold1804 _4184_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2549 hold554/X VGND VGND VPWR VPWR _4324_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1815 hold396/X VGND VGND VPWR VPWR _4333_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4115_ _3385_/Y hold983/A _4115_/S VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1826 _6908_/Q VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1837 hold472/X VGND VGND VPWR VPWR _4036_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1848 hold997/X VGND VGND VPWR VPWR hold468/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5095_ _5095_/A _5095_/B VGND VGND VPWR VPWR _5095_/Y sky130_fd_sc_hd__nand2_1
Xhold1859 hold297/X VGND VGND VPWR VPWR _5215_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ _4046_/A0 _4045_/X _4046_/S VGND VGND VPWR VPWR _4046_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3661__B1 _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6019_/A _6017_/B _6007_/C VGND VGND VPWR VPWR _5997_/X sky130_fd_sc_hd__and3_4
XANTENNA__5402__A1 _5537_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5169__A _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _4948_/A _5033_/B VGND VGND VPWR VPWR _5136_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3413__B1 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5953__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3964__A1 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4879_ _4510_/A _4564_/Y _4569_/X _4570_/X _4878_/Y VGND VGND VPWR VPWR _4879_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_137_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6618_ _6731_/CLK _6618_/D _6413_/A VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5705__A2 _5653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6549_ _6549_/CLK _6549_/D fanout440/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5469__A1 _5568_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7162__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput270 _6791_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XANTENNA__6130__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput281 _6798_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput292 _6484_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XANTENNA__4141__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3652__B1 _4322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6197__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_65_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5944__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3404__B1 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3955__A1 _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire364 _4218_/Y VGND VGND VPWR VPWR _4220_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire375 hold39/X VGND VGND VPWR VPWR wire375/X sky130_fd_sc_hd__buf_12
XANTENNA__3707__A1 input15/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6121__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5542__A _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4132__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5880__B2 _5678_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4158__A _4158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _6596_/Q _5670_/X _5685_/X _6771_/Q VGND VGND VPWR VPWR _5920_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3643__B1 _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5851_ _6964_/Q _5680_/X _5681_/X _7092_/Q VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
X_4802_ _5090_/C _4802_/B _4802_/C VGND VGND VPWR VPWR _4803_/D sky130_fd_sc_hd__and3_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4199__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5782_ _5782_/A _5782_/B _5782_/C VGND VGND VPWR VPWR _5782_/Y sky130_fd_sc_hd__nor3_4
XFILLER_15_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5935__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4733_ _4726_/A _4607_/B _4727_/A VGND VGND VPWR VPWR _4733_/X sky130_fd_sc_hd__a21o_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4664_ _5026_/C VGND VGND VPWR VPWR _4664_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5699__A1 _6853_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5699__B2 _7053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6403_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__and2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3615_ _3615_/A _3615_/B _3615_/C VGND VGND VPWR VPWR _3616_/D sky130_fd_sc_hd__and3_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6777__CLK_N _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold901 hold901/A VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7185__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4595_ _4638_/A _4595_/B VGND VGND VPWR VPWR _4633_/B sky130_fd_sc_hd__nand2_8
Xhold912 hold912/A VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3237__A _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold923 hold923/A VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold934 hold934/A VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6334_ _6588_/Q _5989_/X _6013_/X _6628_/Q _6333_/X VGND VGND VPWR VPWR _6338_/B
+ sky130_fd_sc_hd__a221o_1
X_3546_ _6873_/Q _5281_/A _5434_/A _7009_/Q _3545_/X VGND VGND VPWR VPWR _3556_/A
+ sky130_fd_sc_hd__a221o_1
Xhold945 hold945/A VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold956 hold956/A VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold967 hold967/A VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold978 hold978/A VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6265_ _6526_/Q _6339_/B _6264_/X VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__o21ba_1
Xhold989 hold989/A VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3477_ _3535_/A _3549_/B VGND VGND VPWR VPWR _4310_/A sky130_fd_sc_hd__nor2_8
XANTENNA__6112__A2 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5452__A _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4123__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2302 hold795/X VGND VGND VPWR VPWR _4163_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5216_ _5216_/A0 _5549_/A1 _5217_/S VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2313 _7013_/Q VGND VGND VPWR VPWR hold836/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2324 hold720/X VGND VGND VPWR VPWR _5475_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6196_ _6884_/Q _6004_/X _6008_/X _7108_/Q VGND VGND VPWR VPWR _6196_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2335 _4290_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1601 _6527_/Q VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2346 _5521_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2357 hold839/X VGND VGND VPWR VPWR _4066_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1612 _7209_/A VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1623 _6817_/Q VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5147_ _5147_/A1 _4836_/A _5134_/Y _5135_/X _5128_/Y VGND VGND VPWR VPWR _5147_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout473_A input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2368 _5346_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1634 _4074_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2379 _5409_/X VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1645 hold558/X VGND VGND VPWR VPWR _4307_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1656 _4265_/X VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1667 hold320/X VGND VGND VPWR VPWR _5196_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1678 _6905_/Q VGND VGND VPWR VPWR hold613/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5078_ _5078_/A1 _4836_/A _5025_/X _5077_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__a211o_1
Xhold1689 _5349_/X VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4029_ _4029_/A0 _4028_/X _4029_/S VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1490_A _6478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1588_A _6952_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4250__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1922_A _6453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6103__A2 _5997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5362__A _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A mask_rev_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2880 _7196_/Q VGND VGND VPWR VPWR _6366_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2891 _7201_/Q VGND VGND VPWR VPWR _6381_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3625__B1 _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5301__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5917__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold219 hold219/A VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3400_ input50/X _3330_/Y _5245_/A _6843_/Q VGND VGND VPWR VPWR _3400_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4380_ _5009_/A _4811_/B VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__and2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ hold56/X hold15/X VGND VGND VPWR VPWR _5263_/A sky130_fd_sc_hd__nor2_8
XFILLER_124_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5272__A _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7126_/Q _5973_/X _5988_/X _6870_/Q VGND VGND VPWR VPWR _6050_/X sky130_fd_sc_hd__a22o_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3840_/A _3842_/C1 _6657_/Q VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5001_ _5001_/A _5001_/B VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__nand2_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__A1 _6996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4381__A_N _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3193_ _3914_/B VGND VGND VPWR VPWR _3193_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6952_ _7099_/CLK _6952_/D fanout472/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5903_ _5903_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__o21ba_1
XFILLER_81_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6883_ _7091_/CLK _6883_/D fanout452/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5834_ _6947_/Q _5658_/X _5673_/X _6867_/Q _5833_/X VGND VGND VPWR VPWR _5835_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5908__A2 _5666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5765_ _6976_/Q _5660_/X _5689_/X _7080_/Q _5764_/X VGND VGND VPWR VPWR _5770_/B
+ sky130_fd_sc_hd__a221o_1
X_4716_ _4384_/A _4658_/A _4638_/Y _4220_/B VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3395__A2 _5551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5696_ _6869_/Q _5674_/X _5679_/X _6901_/Q _5695_/X VGND VGND VPWR VPWR _5696_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4647_ _4682_/A _4712_/B VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__and2_2
XANTENNA__6333__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5881__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1169_A _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold720 hold720/A VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4578_ _4578_/A _4583_/B VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__nor2_4
XFILLER_150_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold731 hold731/A VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold742 hold742/A VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold753 hold753/A VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold764 hold764/A VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6317_ _6341_/A0 _6342_/S _6315_/X _6316_/X VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3529_ _3529_/A _3529_/B _3529_/C _3529_/D VGND VGND VPWR VPWR _3557_/B sky130_fd_sc_hd__nor4_1
XFILLER_143_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold775 hold775/A VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold786 hold786/A VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold797 hold797/A VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6097__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6248_ _6703_/Q _5977_/X _5984_/X _6615_/Q _6247_/X VGND VGND VPWR VPWR _6263_/B
+ sky130_fd_sc_hd__a221o_2
Xhold2110 hold666/X VGND VGND VPWR VPWR _5176_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2121 _6836_/Q VGND VGND VPWR VPWR hold336/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2132 _7206_/A VGND VGND VPWR VPWR hold863/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5844__A1 _7036_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2143 _7024_/Q VGND VGND VPWR VPWR hold876/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5903__B1_N _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2154 _6533_/Q VGND VGND VPWR VPWR hold765/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6179_ _6179_/A _6179_/B _6179_/C _6179_/D VGND VGND VPWR VPWR _6189_/B sky130_fd_sc_hd__nor4_2
Xhold2165 _4023_/X VGND VGND VPWR VPWR hold938/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1420 _7046_/Q VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 _4244_/X VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2176 _7117_/Q VGND VGND VPWR VPWR hold889/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1442 hold212/X VGND VGND VPWR VPWR _5232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2187 _4201_/X VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7200__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1453 _7089_/Q VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2198 _4093_/X VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1464 hold234/X VGND VGND VPWR VPWR _5477_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1475 _4300_/X VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_176_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1486 _5433_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 hold338/X VGND VGND VPWR VPWR _5568_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5780__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6324__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4335__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4099__A0 _3803_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6338__D _6338_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6448__CLK _3940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4810__A2 _4688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3880_ _3880_/A0 _3879_/X _3880_/S VGND VGND VPWR VPWR _6437_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5550_ _5550_/A0 _5577_/A1 _5550_/S VGND VGND VPWR VPWR _5550_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3377__A2 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ _4637_/B _4498_/B _4663_/D VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ _5481_/A0 _5571_/A1 hold17/A VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6315__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _7220_/A VGND VGND VPWR VPWR _7220_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4326__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2353_A _6894_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4432_ _4447_/B _4457_/A VGND VGND VPWR VPWR _4451_/A sky130_fd_sc_hd__xor2_4
XFILLER_172_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7151_ _7185_/CLK _7151_/D fanout447/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfstp_4
X_4363_ _4465_/B _4363_/B VGND VGND VPWR VPWR _4955_/B sky130_fd_sc_hd__and2_1
XFILLER_113_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6079__A1 _7127_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6102_ _6102_/A _6102_/B _6102_/C VGND VGND VPWR VPWR _6114_/C sky130_fd_sc_hd__nor3_1
XANTENNA__4110__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3314_ _3343_/A hold30/X VGND VGND VPWR VPWR _5524_/A sky130_fd_sc_hd__nor2_8
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7082_ _7082_/CLK _7082_/D fanout464/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_4
X_4294_ _4294_/A0 _5193_/A1 _4297_/S VGND VGND VPWR VPWR _4294_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6033_ _7029_/Q _5986_/X _5996_/X _7045_/Q VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__a22o_1
X_3245_ _4917_/A VGND VGND VPWR VPWR _4506_/A sky130_fd_sc_hd__inv_2
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4065__B _5569_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7078_/CLK _6935_/D fanout445/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4801__A2 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout436_A _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6866_ _6996_/CLK _6866_/D fanout462/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _5817_/A1 _6342_/S _5815_/X _5816_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__o22a_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6797_ _6821_/CLK _6797_/D fanout442/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _6887_/Q _5688_/X _5741_/X _5744_/X _5747_/X VGND VGND VPWR VPWR _5748_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5762__B1 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5679_ _5685_/A _5679_/B _5687_/C VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__and3b_4
XANTENNA__6306__A2 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1453_A _7089_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4317__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4868__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold550 hold550/A VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold561 hold561/A VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold572 hold572/A VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1620_A _7052_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold583 _4040_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4020__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1718_A _6570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input136_A wb_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1250 hold366/X VGND VGND VPWR VPWR _5402_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1261 _5358_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _5330_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4256__A _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1283 _5418_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1294 _6927_/Q VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5045__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7002__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3359__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5753__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4308__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4859__A2 _4638_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR _6358_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5036__A2 _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6233__A1 _6712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6233__B2 _6569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B VGND VGND VPWR VPWR _5063_/D sky130_fd_sc_hd__nand2_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3932_ _6827_/Q input89/X _3934_/S VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_4
X_6720_ _6786_/CLK _6720_/D fanout436/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3598__A2 hold16/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4795__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6651_ _6746_/CLK _6651_/D _6416_/A VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfstp_1
X_3863_ _3863_/A _3878_/S VGND VGND VPWR VPWR _3863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5602_ _3193_/Y _5601_/B _5601_/A VGND VGND VPWR VPWR _5602_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_hold2568_A _6981_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4105__S _4106_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6582_ _6760_/CLK _6582_/D fanout441/X VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3794_ _7069_/Q _5506_/A _4256_/A _6692_/Q _3793_/X VGND VGND VPWR VPWR _3801_/A
+ sky130_fd_sc_hd__a221o_1
X_5533_ hold31/X _5533_/B VGND VGND VPWR VPWR _5541_/S sky130_fd_sc_hd__and2_4
XFILLER_117_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3944__S _6458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5464_ _5464_/A0 _5527_/A1 _5469_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7078_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7203_ _7203_/CLK _7203_/D _6346_/B VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_2
X_4415_ _4594_/A _4415_/B VGND VGND VPWR VPWR _5026_/B sky130_fd_sc_hd__nor2_4
X_5395_ _5395_/A0 _5575_/A1 _5397_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
X_7134_ _7134_/CLK _7134_/D fanout469/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_4
X_4346_ _4346_/A _4346_/B _4346_/C VGND VGND VPWR VPWR _4492_/B sky130_fd_sc_hd__and3_4
XANTENNA__3522__A2 _5362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7065_ _7137_/CLK _7065_/D fanout466/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout359 _6167_/S VGND VGND VPWR VPWR _6342_/S sky130_fd_sc_hd__clkbuf_16
X_4277_ hold141/X _5581_/A1 _4279_/S VGND VGND VPWR VPWR _4277_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout386_A hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6016_ _6017_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__and3_4
X_3228_ _6936_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6763__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A2 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4786__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6918_ _6945_/CLK _6918_/D fanout461/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6714_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6849_ _7017_/CLK _6849_/D fanout461/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1570_A _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4015__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5735__B1 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3761__A2 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6160__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold380 hold380/A VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3513__A2 _5443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold391 hold391/A VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 hold75/X VGND VGND VPWR VPWR _4162_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 _4272_/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4777__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5726__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3752__A2 _5326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6151__B1 _5998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4200_ _4200_/A _5220_/C VGND VGND VPWR VPWR _4205_/S sky130_fd_sc_hd__and2_2
X_5180_ _5180_/A0 _5193_/A1 _5183_/S VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__mux2_1
Xhold2709 hold652/X VGND VGND VPWR VPWR _4232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4131_ hold170/X _5527_/A1 _4133_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2316_A _6998_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4062_ _4062_/A0 _5584_/A1 _4064_/S VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6206__A1 _7052_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6206__B2 _6948_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3939__S _6459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5965__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4964_ _4963_/X _5044_/C VGND VGND VPWR VPWR _4964_/X sky130_fd_sc_hd__and2b_1
X_6703_ _6730_/CLK _6703_/D _6413_/A VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3915_ _7142_/Q _7143_/Q _5645_/C VGND VGND VPWR VPWR _3915_/Y sky130_fd_sc_hd__nand3b_2
X_4895_ _5136_/A _4997_/A VGND VGND VPWR VPWR _4921_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3440__B2 _6986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6634_ _6835_/CLK _6634_/D _3959_/B VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_4
X_3846_ _3845_/X _3846_/A1 _3846_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5193__A1 _5193_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3777_ _6784_/Q _5178_/A _4200_/A _6639_/Q VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6565_ _7191_/CLK _6565_/D VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfxtp_1
X_5516_ _5516_/A0 _5534_/A1 _5523_/S VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3743__A2 _5425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6496_ _6512_/CLK _6496_/D fanout473/X VGND VGND VPWR VPWR _7217_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_161_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5447_ _5447_/A0 _5582_/A1 _5451_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1249_A _6976_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5378_ _5378_/A0 _5567_/A1 _5379_/S VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7121_/CLK _7117_/D _6399_/A VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfstp_2
X_4329_ _4329_/A0 _5543_/A1 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7048_ _7128_/CLK _7048_/D fanout468/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4518__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5956__B1 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5708__B1 _5647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3734__A2 _3315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A mgmt_gpio_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6133__B1 _5990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_61_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5304__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3670__B2 _6839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _7126_/Q _5569_/A _5245_/A _6838_/Q _3699_/X VGND VGND VPWR VPWR _3703_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_159_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4680_ _4590_/Y _4674_/Y _4679_/Y _4668_/Y _4678_/X VGND VGND VPWR VPWR _4703_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3631_ _6999_/Q _5425_/A _5542_/A _7103_/Q _3630_/X VGND VGND VPWR VPWR _3636_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6350_ _3616_/Y hold993/A _6354_/S VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__mux2_1
X_3562_ _3764_/A _3648_/B VGND VGND VPWR VPWR _3562_/Y sky130_fd_sc_hd__nor2_2
XFILLER_143_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5301_ _5301_/A0 _5571_/A1 _5307_/S VGND VGND VPWR VPWR _5301_/X sky130_fd_sc_hd__mux2_1
X_6281_ _6724_/Q _5978_/X _5992_/X _6709_/Q _6280_/X VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6124__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3493_ _3974_/B _3293_/Y hold89/A _6716_/Q VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__a22o_1
X_5232_ _5232_/A0 _5563_/A1 hold48/X VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
Xhold2506 _6751_/Q VGND VGND VPWR VPWR hold929/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2517 _5507_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5163_ _4590_/Y _4691_/Y _4995_/B _4674_/Y VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__o22a_1
Xhold2528 hold890/X VGND VGND VPWR VPWR _5552_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2539 _5489_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1805 _7193_/Q VGND VGND VPWR VPWR hold995/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4114_ _3422_/Y hold971/A _4115_/S VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__mux2_1
Xhold1816 _4333_/X VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1827 hold390/X VGND VGND VPWR VPWR _5325_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5094_ _3187_/Y _5139_/A _5085_/X _5093_/X VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__o211a_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1838 _6544_/Q VGND VGND VPWR VPWR _4088_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1849 hold468/X VGND VGND VPWR VPWR hold1849/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4045_ _4064_/A0 _5568_/A1 _4056_/C VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3661__B2 _6586_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5938__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _6019_/A _6019_/B _6016_/C VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__and3_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5169__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4947_ _4947_/A _4947_/B VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3413__A1 _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3413__B2 _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4878_ _4934_/B _5048_/A VGND VGND VPWR VPWR _4878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _6731_/CLK hold51/X _6413_/A VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3829_ _3829_/A1 _3835_/S _3827_/Y _3828_/X VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__o22a_1
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6548_ _6753_/CLK _6548_/D fanout435/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6479_ _6486_/CLK _6479_/D fanout434/X VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput260 _6803_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 _6479_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6480_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput293 _6485_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4692__A3 _4691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6828__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3652__A1 _6641_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3404__A1 input18/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5794__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3404__B2 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6354__A0 _3385_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3707__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6106__B1 _6016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output268_A _6789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5542__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4439__A _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4158__B hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6290__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3643__B2 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ _6948_/Q _5658_/X _5664_/X _7020_/Q VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__a22o_1
X_4801_ _5011_/A _4729_/A _4514_/B VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5396__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5781_ _6905_/Q _5679_/X _5778_/X _5780_/X VGND VGND VPWR VPWR _5782_/C sky130_fd_sc_hd__a211o_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _4988_/A _4732_/B VGND VGND VPWR VPWR _4755_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4663_ _4447_/B _4917_/A _4701_/A _4663_/D VGND VGND VPWR VPWR _5026_/C sky130_fd_sc_hd__and4bb_4
XFILLER_174_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4621__B _5048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5209__S _5209_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5699__A2 _5651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4113__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3614_ _3614_/A _3614_/B _3614_/C _3614_/D VGND VGND VPWR VPWR _3615_/C sky130_fd_sc_hd__nor4_1
X_6402_ _6430_/A _6423_/B VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__and2_1
XFILLER_174_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4594_ _4594_/A _4990_/B VGND VGND VPWR VPWR _4826_/A sky130_fd_sc_hd__nor2_4
Xhold902 hold902/A VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold913 hold913/A VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold924 hold924/A VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6333_ _6691_/Q _5980_/X _6017_/X _6773_/Q VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a22o_1
X_3545_ _7121_/Q _5560_/A _4134_/A _6588_/Q VGND VGND VPWR VPWR _3545_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold935 hold935/A VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3952__S _6815_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold946 hold946/A VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold957 hold957/A VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold968 _4226_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6264_ _6258_/X _6339_/B _6264_/C _6264_/D VGND VGND VPWR VPWR _6264_/X sky130_fd_sc_hd__and4b_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3476_ _7025_/Q _5452_/A _4206_/A _6648_/Q _3474_/X VGND VGND VPWR VPWR _3481_/C
+ sky130_fd_sc_hd__a221o_1
X_5215_ _5215_/A0 wire375/X _5217_/S VGND VGND VPWR VPWR _5215_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5452__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5320__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2303 _4163_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2314 hold836/X VGND VGND VPWR VPWR _5444_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6195_ _6924_/Q _5995_/X _6018_/X _6972_/Q _6194_/X VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4349__A _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2325 _6853_/Q VGND VGND VPWR VPWR hold825/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2336 _7207_/A VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2347 _6712_/Q VGND VGND VPWR VPWR hold925/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1602 hold510/X VGND VGND VPWR VPWR _4068_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5871__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5146_ _5143_/Y _5145_/Y _5140_/X VGND VGND VPWR VPWR _5146_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2358 _4066_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1613 hold256/X VGND VGND VPWR VPWR _4234_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2369 _7137_/Q VGND VGND VPWR VPWR hold729/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1624 hold304/X VGND VGND VPWR VPWR _5221_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1635 _6904_/Q VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1646 _4307_/X VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6921__RESET_B _6416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1657 _6844_/Q VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5077_ _5043_/Y _5086_/B _5060_/X _5076_/Y VGND VGND VPWR VPWR _5077_/X sky130_fd_sc_hd__a211o_1
Xhold1668 _5196_/X VGND VGND VPWR VPWR hold321/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1679 hold613/X VGND VGND VPWR VPWR _5322_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _4055_/A0 hold71/X _4047_/C VGND VGND VPWR VPWR _4028_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5387__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5979_ _7155_/Q _7156_/Q VGND VGND VPWR VPWR _6007_/C sky130_fd_sc_hd__nor2_8
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3398__B1 _3389_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6336__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4023__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3570__B1 _4134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input166_A wb_sel_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5362__B _5578_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5311__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5862__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2870 _7159_/Q VGND VGND VPWR VPWR _5646_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input27_A mask_rev_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2881 _7164_/Q VGND VGND VPWR VPWR _5816_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2892 _7176_/Q VGND VGND VPWR VPWR _6141_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3625__B2 _6719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5378__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4722__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4050__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5550__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3561__B1 _5353_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3330_ _3563_/A _3648_/A VGND VGND VPWR VPWR _3330_/Y sky130_fd_sc_hd__nor2_4
XFILLER_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5272__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5302__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3261_ hold62/X hold29/X VGND VGND VPWR VPWR _3349_/A sky130_fd_sc_hd__nand2b_4
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A _5000_/B VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__and2_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5853__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3192_ _6654_/Q VGND VGND VPWR VPWR _3903_/A sky130_fd_sc_hd__inv_4
XFILLER_39_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6951_ _7086_/CLK _6951_/D fanout467/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5902_ _6526_/Q _5678_/Y _5894_/X _5901_/X _6341_/S VGND VGND VPWR VPWR _5902_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4108__S _4115_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6882_ _6963_/CLK _6882_/D fanout464/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5369__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5833_ _7019_/Q _5664_/X _5686_/X _7011_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3947__S _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6030__A2 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4041__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5764_ _7000_/Q _5666_/X _5678_/B _5763_/Y VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6909__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4715_ _4651_/X _4709_/X _4636_/X VGND VGND VPWR VPWR _4759_/C sky130_fd_sc_hd__a21o_1
XANTENNA__6318__B1 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3893__D _3893_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5695_ _6941_/Q _5658_/X _5669_/X _7045_/Q VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4056__A_N _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4646_ _4917_/A _4712_/B VGND VGND VPWR VPWR _4718_/C sky130_fd_sc_hd__and2_1
XFILLER_135_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7120__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5541__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4577_ _4811_/B _4710_/A VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__nand2_2
Xhold721 hold721/A VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold732 hold732/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold743 hold743/A VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3552__B1 _3427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold754 hold754/A VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6316_ _7183_/Q _3924_/Y _5647_/Y VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__o21ba_1
Xhold765 hold765/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3528_ _6977_/Q _5398_/A _5299_/A _6889_/Q _3527_/X VGND VGND VPWR VPWR _3529_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold776 _4273_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5829__C1 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold787 hold787/A VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6097__A2 _6014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold798 hold798/A VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2100 _6783_/Q VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3459_ _6946_/Q _5362_/A _5290_/A _6882_/Q _3432_/X VGND VGND VPWR VPWR _3460_/D
+ sky130_fd_sc_hd__a221o_1
X_6247_ _6605_/Q _5982_/X _5987_/X _6728_/Q VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold1231_A _6812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2111 _5176_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2122 hold336/X VGND VGND VPWR VPWR _5244_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1329_A _7102_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2133 hold863/X VGND VGND VPWR VPWR _5209_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5844__A2 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2144 hold876/X VGND VGND VPWR VPWR _5456_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6178_ _6947_/Q _6005_/X _6015_/X _7019_/Q _6177_/X VGND VGND VPWR VPWR _6179_/D
+ sky130_fd_sc_hd__a221o_1
Xhold1410 _5331_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2155 hold765/X VGND VGND VPWR VPWR _4075_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2166 hold938/X VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1421 hold261/X VGND VGND VPWR VPWR _5481_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2177 hold889/X VGND VGND VPWR VPWR _5561_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1432 _6842_/Q VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1443 _5232_/X VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2188 _6883_/Q VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5129_ _4569_/B _4968_/Y _4586_/Y _4550_/Y VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__o211a_1
Xhold1454 hold376/X VGND VGND VPWR VPWR _5529_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2199 _7022_/Q VGND VGND VPWR VPWR hold565/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1465 _6811_/Q VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5402__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1476 _7094_/Q VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1487 _6605_/Q VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4526__B _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 _5568_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3607__A1 _6740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3607__B2 _6533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4018__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1698_A _6484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6006__C1 _6005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6021__A2 _5989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6309__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5780__A1 _6985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3791__B1 _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5532__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5312__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output300_A _6807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6260__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4271__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5771__A1 _3239_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4500_ _4637_/B _4500_/B VGND VGND VPWR VPWR _4500_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3782__B1 _3293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5480_ _5480_/A0 _5534_/A1 hold17/X VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4431_ _4447_/B _4682_/A _4808_/B VGND VGND VPWR VPWR _4498_/B sky130_fd_sc_hd__and3_1
XFILLER_172_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _3383_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5523__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3534__B1 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4362_ _4362_/A _4362_/B VGND VGND VPWR VPWR _4363_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7150_ _7180_/CLK _7150_/D fanout448/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfstp_1
X_6101_ _7032_/Q _5986_/X _5998_/X _6888_/Q _6100_/X VGND VGND VPWR VPWR _6102_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6079__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3313_ hold62/X hold29/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__nand2_4
X_7081_ _7094_/CLK _7081_/D fanout450/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_4
X_4293_ _4293_/A0 hold275/X _4297_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3244_ _4637_/D VGND VGND VPWR VPWR _4594_/A sky130_fd_sc_hd__clkinv_8
X_6032_ _7125_/Q _5973_/X _5988_/X _6869_/Q _6031_/X VGND VGND VPWR VPWR _6032_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6934_ _7061_/CLK _6934_/D fanout450/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfstp_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6865_ _7101_/CLK _6865_/D fanout450/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5816_ _5816_/A1 _3924_/Y _5647_/Y VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4014__A1 _5579_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6796_ _6809_/CLK _6796_/D fanout433/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5747_ _7087_/Q _5681_/X _5745_/X _5746_/X VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5762__B2 _6872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3773__B1 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5678_ _5689_/A _5678_/B VGND VGND VPWR VPWR _5678_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_136_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5514__A1 hold71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4629_ _4522_/B _4491_/Y _5102_/A _4602_/Y _4627_/X VGND VGND VPWR VPWR _4630_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3525__B1 _5308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold540 hold540/A VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold551 hold551/A VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold562 hold562/A VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold573 _4240_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold584 hold584/A VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold595 _5539_/X VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7198__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1240 _5312_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1251 _5402_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1262 _7063_/Q VGND VGND VPWR VPWR hold134/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1273 _7096_/Q VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input129_A wb_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4256__B _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1284 _6919_/Q VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 hold151/X VGND VGND VPWR VPWR _5347_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4005__A1 _5189_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input94_A uart_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5753__A1 _6960_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5753__B2 _7072_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5505__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5307__S _5307_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5808__A2 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6380_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6233__A2 _5973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4244__A1 _5563_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4980_ _4980_/A _4981_/B VGND VGND VPWR VPWR _5100_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3931_ _6828_/Q input91/X _3934_/S VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_4
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_56_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6650_ _6756_/CLK _6650_/D fanout441/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4182__A _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3862_ _3862_/A _6656_/Q _3903_/A VGND VGND VPWR VPWR _3878_/S sky130_fd_sc_hd__nand3_4
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5601_ _5601_/A _5601_/B _5601_/C VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__and3_1
X_6581_ _6760_/CLK _6581_/D fanout441/X VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3793_ _7093_/Q hold31/A _4134_/A _6584_/Q VGND VGND VPWR VPWR _3793_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5532_ _5532_/A0 _5577_/A1 _5532_/S VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5463_ _5463_/A0 _5571_/A1 _5469_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7202_ _3950_/A1 _7202_/D _6346_/B VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4414_ _4574_/A _4637_/D VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__and2b_4
X_5394_ _5394_/A0 hold95/X _5397_/S VGND VGND VPWR VPWR _5394_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7133_ _7133_/CLK _7133_/D fanout469/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfstp_4
X_4345_ _4345_/A _4345_/B _4345_/C _4345_/D VGND VGND VPWR VPWR _4346_/C sky130_fd_sc_hd__and4_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7064_ _7136_/CLK _7064_/D fanout470/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_4
X_4276_ _4276_/A0 _5580_/A1 _4279_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
X_6015_ _6019_/A _6015_/B _6019_/B VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__and3_4
X_3227_ _6944_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout379_A _5529_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1027_A _3325_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6224__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4235__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _6945_/CLK _6917_/D fanout461/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_70_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6848_ _7072_/CLK _6848_/D fanout460/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5735__A1 _6983_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6779_ _3958_/A1 _6779_/D _6431_/X VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__5735__B2 _7023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4031__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6160__B2 _6986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold381 hold381/A VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold392 hold392/A VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 _4278_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _4162_/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6215__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1092 _6626_/Q VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output298_A _6805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6151__A1 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ _4130_/A0 _5238_/A1 _4133_/S VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4061_ _4061_/A0 _5529_/A1 _4064_/S VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6206__A2 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4217__A1 _5448_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5500__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _4963_/A _5148_/A _4963_/C VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__and3_1
XANTENNA__3976__A0 _6434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6702_ _6730_/CLK _6702_/D _6413_/A VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_4
X_3914_ _7144_/Q _3914_/B VGND VGND VPWR VPWR _5645_/C sky130_fd_sc_hd__nor2_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3440__A2 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4894_ _4894_/A _4894_/B VGND VGND VPWR VPWR _4903_/B sky130_fd_sc_hd__and2_1
XFILLER_189_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6633_ _6794_/CLK _6633_/D fanout434/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5717__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3845_ _3182_/Y _3879_/B _6657_/Q VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3728__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6564_ _7191_/CLK _6564_/D VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfxtp_1
X_3776_ _6624_/Q _4182_/A _5175_/A _6782_/Q _3775_/X VGND VGND VPWR VPWR _3783_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5515_ _5515_/A _5569_/B VGND VGND VPWR VPWR _5523_/S sky130_fd_sc_hd__and2_4
X_6495_ _6512_/CLK _6495_/D fanout473/X VGND VGND VPWR VPWR _7216_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_172_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5446_ _5446_/A0 _5572_/A1 _5451_/S VGND VGND VPWR VPWR _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5377_ _5377_/A0 _5584_/A1 _5379_/S VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
X_7116_ _7136_/CLK _7116_/D fanout472/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4328_ _4328_/A hold9/X VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and2_4
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input1_A debug_mode VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7047_ _7134_/CLK _7047_/D fanout469/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4259_ hold147/X _5527_/A1 _4261_/S VGND VGND VPWR VPWR _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4208__A1 _5238_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5410__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A1 _6573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4534__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4026__S _4047_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3719__B1 _5281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6241__S _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4550__A _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input57_A mgmt_gpio_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5892__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4998__A2 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output213_A _3946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5320__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3670__A2 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A0 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6794_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3630_ _5207_/A _5184_/B _3427_/Y _6791_/Q _3389_/Y VGND VGND VPWR VPWR _3630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3561_ _6928_/Q _5344_/A _5353_/A _6936_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _5300_/A0 _5534_/A1 _5307_/S VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6280_ _6631_/Q _5971_/X _6017_/X _6771_/Q VGND VGND VPWR VPWR _6280_/X sky130_fd_sc_hd__a22o_4
X_3492_ _3563_/A hold88/A VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__nor2_4
XFILLER_143_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6124__B2 _7009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5231_ _5231_/A0 _5238_/A1 hold48/X VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3489__A2 _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5883__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2507 hold929/X VGND VGND VPWR VPWR _4327_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2518 _6971_/Q VGND VGND VPWR VPWR hold655/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5162_ _5162_/A _5162_/B _5162_/C VGND VGND VPWR VPWR _5162_/Y sky130_fd_sc_hd__nand3_1
Xhold2529 _5552_/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6608_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4113_ _3462_/Y hold978/A _4115_/S VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__mux2_1
Xhold1806 hold995/X VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1817 _7226_/A VGND VGND VPWR VPWR hold340/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5093_ _5088_/X _5136_/C _5092_/X _5086_/Y VGND VGND VPWR VPWR _5093_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1828 _5325_/X VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1839 hold1839/A VGND VGND VPWR VPWR hold474/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7145__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4044_ _4044_/A0 _4043_/X _4046_/S VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5230__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5995_ _6019_/A _6007_/C _6016_/C VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__and3_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6060__B1 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2962_A _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4946_ _4368_/B _4407_/Y _4935_/X _4800_/A VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__o31a_1
XANTENNA__3413__A2 _5560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _5127_/A _4965_/B _5044_/B _4876_/X _4636_/X VGND VGND VPWR VPWR _4906_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6616_ _6731_/CLK _6616_/D _6413_/A VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout411_A _5872_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3828_ _3832_/A _6657_/Q _3846_/S VGND VGND VPWR VPWR _3828_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6547_ _7194_/CLK _6547_/D VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfxtp_1
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3770_/B sky130_fd_sc_hd__nor4_1
XANTENNA__6115__A1 _6840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6478_ _6809_/CLK _6478_/D fanout433/X VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5429_ _5429_/A0 _5582_/A1 _5433_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput250 _3957_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
XFILLER_133_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput261 _6783_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
XANTENNA__5405__S _5406_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput272 _6473_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XANTENNA__5874__B1 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput283 _6799_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput294 _6486_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1895_A _6539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3652__A2 _4200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input111_A wb_adr_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6051__B1 _5987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3404__A2 _3310_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5157__A2 _4523_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6106__A1 _7104_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6106__B2 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5315__S _5316_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5865__B1 _5687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6290__B1 _6289_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3643__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C _4800_/D VGND VGND VPWR VPWR _4803_/C sky130_fd_sc_hd__and4_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5780_ _6985_/Q _5656_/X _5680_/X _6961_/Q _5779_/X VGND VGND VPWR VPWR _5780_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4731_/A _4993_/B VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4662_ _4666_/A _5150_/C VGND VGND VPWR VPWR _4662_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6401_ _6430_/A _6430_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ _7080_/Q _5515_/A _4334_/A _6760_/Q _3612_/X VGND VGND VPWR VPWR _3614_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4593_ _4574_/A _4638_/A VGND VGND VPWR VPWR _4990_/B sky130_fd_sc_hd__nand2b_4
XFILLER_174_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold903 hold903/A VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold914 hold914/A VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6332_ _6726_/Q _5978_/X _5995_/X _6603_/Q _6331_/X VGND VGND VPWR VPWR _6338_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold925 hold925/A VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3544_ _3544_/A _3648_/A VGND VGND VPWR VPWR _4134_/A sky130_fd_sc_hd__nor2_8
Xhold936 _4228_/X VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4108__A0 _3803_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold947 hold947/A VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold958 hold958/A VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6263_ _6263_/A _6263_/B _6263_/C _6263_/D VGND VGND VPWR VPWR _6264_/D sky130_fd_sc_hd__nor4_1
Xhold969 hold969/A VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3475_ _3535_/A _3516_/B VGND VGND VPWR VPWR _4206_/A sky130_fd_sc_hd__nor2_4
X_5214_ _5214_/A0 _5527_/A1 _5217_/S VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2304 _6697_/Q VGND VGND VPWR VPWR hold769/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6194_ _7060_/Q _5990_/X _5991_/X _6916_/Q _6193_/X VGND VGND VPWR VPWR _6194_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2315 _5444_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2326 hold825/X VGND VGND VPWR VPWR _5264_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2337 hold496/X VGND VGND VPWR VPWR _4230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2348 hold925/X VGND VGND VPWR VPWR _4281_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5145_ _4683_/A _5144_/X _5022_/A VGND VGND VPWR VPWR _5145_/Y sky130_fd_sc_hd__o21ai_2
Xhold1603 _4068_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1614 _4234_/X VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2359 _7105_/Q VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1625 _5221_/X VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1636 hold349/X VGND VGND VPWR VPWR _5321_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1647 _6591_/Q VGND VGND VPWR VPWR hold561/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1658 hold410/X VGND VGND VPWR VPWR _5253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5076_ _5066_/X _5074_/X _5062_/A VGND VGND VPWR VPWR _5076_/Y sky130_fd_sc_hd__a21oi_1
Xhold1669 _6773_/Q VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6281__B1 _5992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4027_ _4027_/A0 _4026_/X _4029_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4365__A _4701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout459_A input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3634__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6033__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5978_ _6008_/A _6014_/A _6019_/C VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__and3_4
X_4929_ _5126_/B _4929_/B _5112_/B VGND VGND VPWR VPWR _4930_/D sky130_fd_sc_hd__and3_1
XFILLER_21_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmgmt_gpio_9_buff_inst _3940_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_134_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3570__B2 _6587_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5847__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input159_A wb_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2860 _6776_/Q VGND VGND VPWR VPWR _3677_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2871 _7178_/Q VGND VGND VPWR VPWR _6191_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2882 _7168_/Q VGND VGND VPWR VPWR _5903_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2893 _7199_/Q VGND VGND VPWR VPWR _6375_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6272__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3625__A2 _3307_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4822__A1 _4729_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6024__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output280_A _6797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ hold21/X _3276_/A hold54/A VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__and3_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _6685_/Q VGND VGND VPWR VPWR _3969_/A sky130_fd_sc_hd__inv_2
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6950_ _7072_/CLK _6950_/D fanout460/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfstp_2
X_5901_ _6630_/Q _5663_/X _5895_/X _5896_/X _5900_/X VGND VGND VPWR VPWR _5901_/X
+ sky130_fd_sc_hd__a2111o_1
X_6881_ _7017_/CLK _6881_/D fanout461/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5832_ _6939_/Q _5659_/X _5663_/X _7027_/Q _5831_/X VGND VGND VPWR VPWR _5835_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5763_ _5763_/A _5872_/B VGND VGND VPWR VPWR _5763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4714_ _4717_/B _4714_/B _4714_/C VGND VGND VPWR VPWR _4714_/Y sky130_fd_sc_hd__nand3_4
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5694_ _6933_/Q _5659_/X _5693_/X VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__a21o_1
XFILLER_190_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4645_ _4447_/B _4663_/D VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__and2b_4
XFILLER_175_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold700 hold700/A VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold711 hold711/A VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4576_ _4576_/A _4638_/A VGND VGND VPWR VPWR _4583_/B sky130_fd_sc_hd__nand2_8
Xhold722 hold722/A VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold733 hold733/A VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6315_ _6528_/Q _6339_/B _6314_/Y _6341_/S VGND VGND VPWR VPWR _6315_/X sky130_fd_sc_hd__o211a_1
Xhold744 hold744/A VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold755 _4048_/X VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3527_ input16/X _3310_/Y _4065_/A _6529_/Q VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__a22o_4
XANTENNA__3552__B2 _6793_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold766 hold766/A VGND VGND VPWR VPWR hold766/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5829__B1 _5678_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold788 hold788/A VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6246_ _6549_/Q _5999_/X _6019_/X _6733_/Q _6245_/X VGND VGND VPWR VPWR _6263_/A
+ sky130_fd_sc_hd__a221o_1
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3458_ input40/X _4056_/C _5317_/A _6906_/Q _3457_/X VGND VGND VPWR VPWR _3460_/C
+ sky130_fd_sc_hd__a221o_1
Xhold2101 hold557/X VGND VGND VPWR VPWR _5177_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2112 _6916_/Q VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2123 _6451_/Q VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2134 _5209_/X VGND VGND VPWR VPWR _5210_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_6177_ _7083_/Q _6013_/X _6017_/X _7075_/Q VGND VGND VPWR VPWR _6177_/X sky130_fd_sc_hd__a22o_1
Xhold2145 _5456_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1400 _6974_/Q VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3389_ _3764_/B hold15/A VGND VGND VPWR VPWR _3389_/Y sky130_fd_sc_hd__nor2_4
Xhold2156 _4075_/X VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1411 _7006_/Q VGND VGND VPWR VPWR hold262/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1422 _5481_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2167 _6530_/Q VGND VGND VPWR VPWR hold748/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1224_A _6806_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1433 hold285/X VGND VGND VPWR VPWR _5251_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5128_ _5121_/X _5123_/X _5127_/X VGND VGND VPWR VPWR _5128_/Y sky130_fd_sc_hd__a21boi_1
Xhold2178 _5561_/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2189 hold642/X VGND VGND VPWR VPWR _5297_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1444 _6967_/Q VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1455 _5529_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__B1 _5993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1466 hold452/X VGND VGND VPWR VPWR _5213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1477 hold277/X VGND VGND VPWR VPWR _5535_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1488 hold113/X VGND VGND VPWR VPWR _4160_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5059_ _5123_/B _5059_/B _5059_/C VGND VGND VPWR VPWR _5059_/X sky130_fd_sc_hd__and3_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3607__A2 _4310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4526__C _4751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1499 _6708_/Q VGND VGND VPWR VPWR hold111/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6006__B1 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4542__B _4972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4034__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5780__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3873__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6190__C1 _6166_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6245__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2690 _4213_/X VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5771__A2 _5707_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3782__B2 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4430_ _4682_/A _4808_/B VGND VGND VPWR VPWR _4457_/A sky130_fd_sc_hd__nand2_4
XANTENNA_2 _3471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4361_ _4447_/B _4682_/A _4365_/B _4663_/D VGND VGND VPWR VPWR _4362_/B sky130_fd_sc_hd__a31o_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ _6976_/Q _5976_/B _5993_/X _7008_/Q VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3312_ _3347_/A _3764_/A VGND VGND VPWR VPWR _5443_/A sky130_fd_sc_hd__nor2_8
X_7080_ _7136_/CLK _7080_/D fanout471/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_4
X_4292_ _4292_/A _5569_/B VGND VGND VPWR VPWR _4297_/S sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_52_csclk_A clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6031_ _7021_/Q _5971_/X _5994_/X _7061_/Q _6030_/X VGND VGND VPWR VPWR _6031_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3243_ _6972_/Q VGND VGND VPWR VPWR _3243_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5503__S _5505_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6236__B1 _6017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6933_ _7078_/CLK _6933_/D fanout445/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfstp_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3958__S _6456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6864_ _7108_/CLK _6864_/D fanout451/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5815_ _6842_/Q _5678_/Y _5808_/X _5814_/X _6166_/S VGND VGND VPWR VPWR _5815_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_179_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6795_ _6803_/CLK _6795_/D fanout442/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_179_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _6863_/Q _5673_/X _5680_/X _6959_/Q VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5762__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3773__B2 _6845_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5677_ _5689_/A _5677_/B VGND VGND VPWR VPWR _5707_/B sky130_fd_sc_hd__nor2_8
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4628_ _4628_/A _4917_/D VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nand2_1
Xhold530 hold530/A VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ _4598_/B _4598_/C VGND VGND VPWR VPWR _4601_/B sky130_fd_sc_hd__nand2_1
Xhold541 hold541/A VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold552 hold552/A VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold563 hold563/A VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold574 hold574/A VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold585 hold585/A VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold596 hold596/A VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ _6639_/Q _5986_/X _5998_/X _6579_/Q _6228_/X VGND VGND VPWR VPWR _6230_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5413__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1230 hold84/X VGND VGND VPWR VPWR _4055_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6227__B1 _6007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1241 _6936_/Q VGND VGND VPWR VPWR hold330/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1252 _7072_/Q VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4029__S _4029_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1263 hold134/X VGND VGND VPWR VPWR _5500_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1274 hold411/X VGND VGND VPWR VPWR _5537_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 hold136/X VGND VGND VPWR VPWR _5338_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _5347_/X VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5450__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1975_A _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5753__A2 _5680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A spimemio_flash_io1_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7142__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5323__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6367_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6383_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6218__B1 _6018_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5441__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3930_ _6656_/Q _3929_/Y _3739_/S VGND VGND VPWR VPWR _6436_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3452__B1 _5389_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ _3879_/A _6468_/Q _3903_/A _3857_/B _3847_/B VGND VGND VPWR VPWR _3861_/Y
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__4182__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5600_ _7142_/Q _7143_/Q _5599_/D _5600_/B1 VGND VGND VPWR VPWR _5601_/C sky130_fd_sc_hd__a31o_1
X_6580_ _6745_/CLK _6580_/D fanout440/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3802_/C sky130_fd_sc_hd__nor4_1
XANTENNA__5744__A2 _5662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5531_ _5531_/A0 _5549_/A1 _5532_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5462_ _5462_/A0 _5534_/A1 _5469_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
X_7201_ _3950_/A1 _7201_/D _6346_/B VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_1
X_4413_ _4804_/A VGND VGND VPWR VPWR _4415_/B sky130_fd_sc_hd__clkinv_2
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5393_ _5393_/A0 _5537_/A1 _5397_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
X_7132_ _7132_/CLK _7132_/D fanout453/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4180__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4344_ _4344_/A _4344_/B _4344_/C _4344_/D VGND VGND VPWR VPWR _4346_/B sky130_fd_sc_hd__and4_1
XFILLER_113_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7063_ _7063_/CLK _7063_/D fanout460/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_4
X_4275_ _4275_/A0 _5561_/A1 _4279_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5233__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _6014_/A _6019_/B _6019_/C VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__and3_4
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3226_ _6952_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6209__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3691__B1 _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5968__C1 _6341_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5432__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _7107_/CLK _6916_/D fanout451/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout441_A fanout454/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3443__B1 _5461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4092__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6847_ _7063_/CLK _6847_/D fanout467/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6778_ _3940_/A1 _6778_/D _6430_/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__5735__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3746__A1 _6981_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5729_ _5729_/A0 _5728_/X _6341_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3746__B2 _6712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5408__S _5415_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5499__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7165__CLK _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6160__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4171__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold360 hold360/A VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold382 hold382/A VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold393 hold393/A VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input141_A wb_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _5520_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3682__B1 _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1071 _6461_/Q VGND VGND VPWR VPWR _3842_/C1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1082 _6730_/Q VGND VGND VPWR VPWR _4302_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1093 hold182/X VGND VGND VPWR VPWR _4185_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5423__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3434__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3985__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5726__A2 _5929_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5318__S _5325_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6151__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4162__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ _4060_/A0 _5537_/A1 _4064_/S VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6682__CLK _3950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5414__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4962_ _5162_/A _4962_/B _4962_/C VGND VGND VPWR VPWR _4963_/C sky130_fd_sc_hd__and3_1
XANTENNA__5965__A2 _5656_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3913_ _6816_/Q _5611_/A _3912_/X _6490_/Q VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__a22o_1
X_6701_ _6701_/CLK _6701_/D fanout436/X VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4893_ _4893_/A _4922_/A VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__and2_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6632_ _6794_/CLK _6632_/D fanout435/X VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfrtp_4
X_3844_ _3846_/A1 _3843_/Y _3842_/X VGND VGND VPWR VPWR _3844_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5717__A2 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _7185_/CLK _6563_/D VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfxtp_1
X_3775_ _6877_/Q _5290_/A _3648_/Y _6820_/Q VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__a22o_2
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5514_ _5514_/A0 hold71/X _5514_/S VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6494_ _6512_/CLK _6494_/D fanout473/X VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__6986__RESET_B fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5445_ _5445_/A0 _5562_/A1 _5451_/S VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4153__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5376_ _5376_/A0 _5583_/A1 _5379_/S VGND VGND VPWR VPWR _5376_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7115_ _7139_/CLK _7115_/D fanout471/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_4
X_4327_ _4327_/A0 _5189_/A1 _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout391_A _5536_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7046_ _7084_/CLK _7046_/D fanout445/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4258_ _4258_/A0 _5238_/A1 _4261_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
X_3209_ _7080_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__clkinv_2
X_4189_ _4189_/A0 _5237_/A1 _4193_/S VGND VGND VPWR VPWR _4189_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5405__A1 _5549_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3416__B1 _5254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5956__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4916__B1 _4676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4042__S _4046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6133__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4144__A1 _5195_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4998__A3 _4683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3407__B1 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A1 _3958_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _3559_/X _6778_/Q _3739_/S VGND VGND VPWR VPWR _6778_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3491_ _3553_/A _3550_/B VGND VGND VPWR VPWR _4200_/A sky130_fd_sc_hd__nor2_8
XANTENNA__6124__A2 _5983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4135__A1 _5237_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2154_A _6533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5230_ _5230_/A0 _5543_/A1 hold48/X VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4188__A _4188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5161_ _4417_/B _4698_/Y _4788_/X _5117_/X _5160_/X VGND VGND VPWR VPWR _5162_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold2508 _4327_/X VGND VGND VPWR VPWR hold930/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2519 hold655/X VGND VGND VPWR VPWR _5396_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4112_/A0 _4112_/A1 _4115_/S VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__mux2_1
Xhold1807 hold459/X VGND VGND VPWR VPWR hold1807/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1818 hold340/X VGND VGND VPWR VPWR _4246_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5092_ _5149_/B _5137_/B _5092_/C VGND VGND VPWR VPWR _5092_/X sky130_fd_sc_hd__and3_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1829 _7189_/Q VGND VGND VPWR VPWR hold994/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4043_ hold292/X _5567_/A1 _4056_/C VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5511__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3646__B1 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5994_ _6017_/B _6019_/B _6018_/B VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__and3_4
XANTENNA__5938__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3949__A1 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4945_ _4368_/A _4477_/Y _4729_/A _4550_/Y _4944_/X VGND VGND VPWR VPWR _5090_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _4522_/B _4507_/Y _5108_/C _5089_/B _4875_/X VGND VGND VPWR VPWR _4876_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3827_ _6657_/Q _3827_/B _3827_/C VGND VGND VPWR VPWR _3827_/Y sky130_fd_sc_hd__nor3_1
XFILLER_119_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6615_ _6731_/CLK _6615_/D _6413_/A VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6546_ _7194_/CLK _6546_/D VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout404_A _5533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3758_ _7013_/Q _5443_/A _4146_/A _6594_/Q _3757_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6115__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6477_ _6809_/CLK _6477_/D fanout433/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_134_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3689_ _6753_/Q _4328_/A _3521_/Y _6536_/Q _3688_/X VGND VGND VPWR VPWR _3694_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4126__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ _5428_/A0 _5563_/A1 _5433_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
Xoutput240 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput251 _3964_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
XFILLER_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput262 _6784_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput273 _6474_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 _6800_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XANTENNA__4098__A _6678_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5359_ _5359_/A0 _5575_/A1 _5361_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
Xoutput295 _6471_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1519_A _6948_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7029_ _7045_/CLK _7029_/D fanout444/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3637__B1 _5497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4545__B _4724_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1888_A _6502_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4037__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6051__A1 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6051__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input104_A wb_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3876__S _3878_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4280__B hold9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6106__A2 _6008_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4117__A1 _5561_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5865__A1 _6569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3628__B1 _4182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5331__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6290__A1 _6527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4730_ _4955_/D _4730_/B VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__nand2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__B1 _5542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4661_ _5150_/C VGND VGND VPWR VPWR _4661_/Y sky130_fd_sc_hd__inv_2
X_6400_ _6430_/A _6433_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3612_ _7128_/Q _5569_/A _4140_/A _6592_/Q _3611_/X VGND VGND VPWR VPWR _3612_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4592_ _4637_/C _4592_/B VGND VGND VPWR VPWR _4989_/B sky130_fd_sc_hd__and2b_2
XFILLER_190_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold904 hold904/A VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6331_ _6741_/Q _6008_/X _6016_/X _6454_/Q VGND VGND VPWR VPWR _6331_/X sky130_fd_sc_hd__a22o_1
X_3543_ _3543_/A _3543_/B _3543_/C VGND VGND VPWR VPWR _3557_/C sky130_fd_sc_hd__nor3_1
Xhold915 hold915/A VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold926 hold926/A VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold937 hold937/A VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 hold948/A VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6262_ _6585_/Q _5989_/X _6013_/X _6625_/Q _6261_/X VGND VGND VPWR VPWR _6263_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold959 hold959/A VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3474_ _6849_/Q _5254_/A hold57/A _6573_/Q VGND VGND VPWR VPWR _3474_/X sky130_fd_sc_hd__a22o_1
X_5213_ _5213_/A0 _5303_/A1 _5217_/S VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6193_ _7028_/Q _5971_/X _5987_/X _7116_/Q VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__a22o_1
Xhold2305 hold769/X VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2316 _6998_/Q VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5144_ _4648_/Y _4995_/B _5011_/X _4661_/Y _4735_/Y VGND VGND VPWR VPWR _5144_/X
+ sky130_fd_sc_hd__o221a_1
Xhold2327 _5264_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2338 _6648_/Q VGND VGND VPWR VPWR hold746/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2349 _4281_/X VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1604 _6928_/Q VGND VGND VPWR VPWR hold331/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1615 _6641_/Q VGND VGND VPWR VPWR hold540/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1626 _6868_/Q VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1637 _5321_/X VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5075_ _4402_/Y _4947_/B _4510_/B _4510_/A VGND VGND VPWR VPWR _5100_/D sky130_fd_sc_hd__a31o_1
Xhold1648 _4143_/X VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5241__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1659 _5253_/X VGND VGND VPWR VPWR _6844_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6281__A1 _6724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4026_ _4054_/A0 _5567_/A1 _4047_/C VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5977_ _6015_/B _6008_/A _6017_/A VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__and3_4
XANTENNA__3398__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4928_ _5100_/C _4928_/B _4928_/C VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__and3_1
XFILLER_178_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4859_ _4701_/A _4638_/Y _4701_/B _5073_/B VGND VGND VPWR VPWR _4859_/X sky130_fd_sc_hd__o31a_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6336__A2 _5999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6529_ _6803_/CLK _6529_/D fanout442/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3570__A2 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3858__A0 _3879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2850 _3388_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6817_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2861 _6678_/Q VGND VGND VPWR VPWR _3917_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2872 _6167_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2883 _5882_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2894 hold12/A VGND VGND VPWR VPWR _5004_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6272__B2 _6734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5783__B1 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4338__A1 _5233_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output273_A _6474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7086_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4230__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3561__A2 _5344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3190_ _6684_/Q VGND VGND VPWR VPWR _3967_/A sky130_fd_sc_hd__inv_2
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4813__A2 _4607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5900_ _6585_/Q _5662_/X _5897_/X _5898_/X _5899_/X VGND VGND VPWR VPWR _5900_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _7091_/CLK _6880_/D fanout452/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_4
X_5831_ _6851_/Q _5653_/X _5662_/X _6899_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5762_ _6912_/Q _5670_/X _5674_/X _6872_/Q _5761_/X VGND VGND VPWR VPWR _5770_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5774__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4713_ _4713_/A _4714_/B _4751_/C VGND VGND VPWR VPWR _4713_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6318__A2 _5985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5693_ _6877_/Q _5667_/X _5688_/X _6885_/Q VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4329__A1 _5543_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4644_ _4732_/B _5048_/B VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__nand2_1
XFILLER_190_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4575_ _4637_/A _4637_/B _4637_/C _4637_/D VGND VGND VPWR VPWR _4710_/A sky130_fd_sc_hd__and4bb_4
Xhold701 hold701/A VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap420 _4666_/A VGND VGND VPWR VPWR _4676_/B sky130_fd_sc_hd__clkbuf_2
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold723 hold723/A VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6314_ _6295_/X _6314_/B _6314_/C VGND VGND VPWR VPWR _6314_/Y sky130_fd_sc_hd__nand3b_4
X_3526_ _3726_/B _3550_/B VGND VGND VPWR VPWR _4065_/A sky130_fd_sc_hd__nor2_8
XANTENNA__3552__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold734 _5295_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold745 hold745/A VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold756 hold756/A VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold767 hold767/A VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold778 hold778/A VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6245_ _6753_/Q _5638_/X _6015_/X _6758_/Q VGND VGND VPWR VPWR _6245_/X sky130_fd_sc_hd__a22o_1
Xhold789 hold789/A VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3457_ _7106_/Q _5542_/A _5551_/A _7114_/Q VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2102 _5177_/X VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2113 hold372/X VGND VGND VPWR VPWR _5334_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2124 hold526/X VGND VGND VPWR VPWR _3981_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6176_ _7115_/Q _5987_/X _5993_/X _7011_/Q _6175_/X VGND VGND VPWR VPWR _6179_/C
+ sky130_fd_sc_hd__a221o_1
X_3388_ _3387_/X _3388_/A1 _3739_/S VGND VGND VPWR VPWR _3388_/X sky130_fd_sc_hd__mux2_1
Xhold2135 _6897_/Q VGND VGND VPWR VPWR hold685/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1401 hold264/X VGND VGND VPWR VPWR _5400_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2146 _6573_/Q VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5127_ _5127_/A _5127_/B _5127_/C _5127_/D VGND VGND VPWR VPWR _5127_/X sky130_fd_sc_hd__and4_1
Xhold1412 hold262/X VGND VGND VPWR VPWR _5436_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2157 _6711_/Q VGND VGND VPWR VPWR hold705/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1423 _7195_/Q VGND VGND VPWR VPWR hold273/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2168 hold748/X VGND VGND VPWR VPWR _4072_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1434 _5251_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2179 _6690_/Q VGND VGND VPWR VPWR hold819/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_183_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1445 hold240/X VGND VGND VPWR VPWR _5392_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1456 _6909_/Q VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1467 _7003_/Q VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5058_ _5108_/B _5110_/A _5058_/C _5058_/D VGND VGND VPWR VPWR _5059_/C sky130_fd_sc_hd__and4_1
Xhold1478 _6628_/Q VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 _4160_/X VGND VGND VPWR VPWR hold114/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4009_/A _5569_/B VGND VGND VPWR VPWR _4011_/S sky130_fd_sc_hd__and2_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5765__B1 _5689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6309__A2 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3791__A2 _3977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3528__C1 _3527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4050__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4740__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6188__D _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A mask_rev_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4286__A _4286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2680 _6666_/Q VGND VGND VPWR VPWR hold543/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2691 _6881_/Q VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1990 hold498/X VGND VGND VPWR VPWR _4027_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4225__S _4237_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5756__B1 _5669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3782__A2 _3291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6181__B1 _5977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4360_ _4360_/A _4360_/B VGND VGND VPWR VPWR _4465_/B sky130_fd_sc_hd__nand2_2
XANTENNA_hold2067_A _7000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3534__A2 _3988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3311_ _3563_/A _3726_/A VGND VGND VPWR VPWR _5542_/A sky130_fd_sc_hd__nor2_8
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4291_ _4291_/A0 _5189_/A1 _4291_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2234_A _6642_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6030_ _6925_/Q _5982_/X _6014_/X _6989_/Q VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3242_ _6970_/Q VGND VGND VPWR VPWR _3242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6395__B _6423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6932_ _7107_/CLK _6932_/D fanout451/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4798__A1 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6863_ _6977_/CLK _6863_/D fanout465/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5814_ _7026_/Q _5663_/X _5809_/X _5811_/X _5813_/X VGND VGND VPWR VPWR _5814_/X
+ sky130_fd_sc_hd__a2111o_4
X_6794_ _6794_/CLK _6794_/D fanout434/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3758__C1 _3757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5745_ _6943_/Q _5658_/X _5664_/X _7015_/Q VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6350__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3773__A2 _5226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5676_ _5679_/B _5676_/B VGND VGND VPWR VPWR _5677_/B sky130_fd_sc_hd__nand2_8
XFILLER_175_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6172__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4627_ _4522_/B _4569_/B _4889_/B _4586_/Y _4626_/X VGND VGND VPWR VPWR _4627_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3525__A2 _5416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold531 hold531/A VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4558_ _4767_/A _5114_/A _4556_/X _4557_/X _4374_/Y VGND VGND VPWR VPWR _4558_/X
+ sky130_fd_sc_hd__a41o_1
Xhold542 hold542/A VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold553 hold553/A VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold564 hold564/A VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold575 hold575/A VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3509_ _3563_/A _3533_/B VGND VGND VPWR VPWR _3509_/Y sky130_fd_sc_hd__nor2_4
XFILLER_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold586 hold586/A VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4489_ _4981_/A _4972_/A VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__nand2_1
Xhold597 _5373_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6228_ _6609_/Q _5976_/B _5993_/X _6619_/Q VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6898_/Q _5989_/X _6013_/X _7082_/Q _6158_/X VGND VGND VPWR VPWR _6163_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1220 hold278/X VGND VGND VPWR VPWR _4283_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _6812_/Q VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1242 hold330/X VGND VGND VPWR VPWR _5357_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1253 hold388/X VGND VGND VPWR VPWR _5510_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1264 _5500_/X VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1275 _6872_/Q VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _5338_/X VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1297 _6856_/Q VGND VGND VPWR VPWR hold347/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4789__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4045__S _4056_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5738__B1 _5679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3185__A _6864_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5910__B1 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6364_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output236_A _3936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6370_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6361_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4463__B _4463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ _3860_/A0 _3879_/B _3860_/S VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3791_ _6450_/Q _3977_/A _4286_/A _6717_/Q _3790_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3755__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5530_ _5530_/A0 _5575_/A1 _5532_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4952__A1 _4601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4952__B2 _4947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5461_ _5461_/A _5569_/B VGND VGND VPWR VPWR _5469_/S sky130_fd_sc_hd__and2_4
XANTENNA__6154__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4412_ _4574_/A _4719_/A VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__and2b_2
X_7200_ _3950_/A1 _7200_/D _6346_/B VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5392_ _5392_/A0 _5572_/A1 _5397_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
X_4343_ _4343_/A _4343_/B _4343_/C _4343_/D VGND VGND VPWR VPWR _4346_/A sky130_fd_sc_hd__and4_1
X_7131_ _7131_/CLK _7131_/D fanout452/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5514__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7062_ _7094_/CLK _7062_/D fanout450/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfstp_1
X_4274_ _4274_/A hold9/X VGND VGND VPWR VPWR _4279_/S sky130_fd_sc_hd__and2_2
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6013_ _6019_/A _6017_/B _6019_/B VGND VGND VPWR VPWR _6013_/X sky130_fd_sc_hd__and3_4
X_3225_ _6960_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6209__B2 _7004_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3691__A1 _6790_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6915_ _7091_/CLK _6915_/D fanout452/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3443__B2 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6846_ _7086_/CLK _6846_/D fanout467/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_50_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5196__A1 _5277_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6777_ _3958_/A1 _6777_/D _6429_/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtn_1
X_3989_ _3989_/A0 _5237_/A1 _3999_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3746__A2 _5407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5728_ _5718_/Y _5727_/Y _6838_/Q _5678_/Y VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6145__B1 _5996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5659_ _5685_/A _5679_/B _5689_/C VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__and3b_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold350 hold350/A VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold361 hold361/A VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5424__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 hold383/A VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold394 hold394/A VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input134_A wb_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _6444_/Q VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3682__B2 _6708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1061 _6766_/Q VGND VGND VPWR VPWR _3249_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1072 _3268_/X VGND VGND VPWR VPWR _3269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1083 _4302_/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1094 _4185_/X VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5187__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6136__B1 _6012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output186_A _3947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5334__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3370__B1 _5524_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4961_ _5151_/C _4961_/B _5042_/A _4961_/D VGND VGND VPWR VPWR _4962_/C sky130_fd_sc_hd__and4_1
XFILLER_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6700_ _6736_/CLK _6700_/D fanout436/X VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2399_A _6785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3912_ _3909_/X _3912_/B VGND VGND VPWR VPWR _3912_/X sky130_fd_sc_hd__and2b_1
X_4892_ _4892_/A _4892_/B _4892_/C _4892_/D VGND VGND VPWR VPWR _4892_/X sky130_fd_sc_hd__and4_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6631_ _6794_/CLK _6631_/D fanout434/X VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3843_ _6461_/Q _3840_/B _3846_/S VGND VGND VPWR VPWR _3843_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5509__S _5514_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3728__A2 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6562_ _7185_/CLK _6562_/D VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfxtp_1
X_3774_ _7109_/Q _5551_/A _3486_/Y _3772_/X _3773_/X VGND VGND VPWR VPWR _3774_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ _5513_/A0 _5549_/A1 _5514_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6127__B1 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6493_ _6512_/CLK _6493_/D fanout473/X VGND VGND VPWR VPWR _7214_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ _5444_/A0 _5543_/A1 _5451_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5375_ _5375_/A0 _5537_/A1 _5379_/S VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5244__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3361__B1 _4241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7114_ _7139_/CLK _7114_/D fanout471/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_4
X_4326_ _4326_/A0 _5233_/A1 _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7045_ _7045_/CLK _7045_/D fanout444/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfstp_2
X_4257_ _4257_/A0 _5543_/A1 _4261_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3703__D _3703_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout384_A hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3208_ _7088_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4188_ _4188_/A _5220_/C VGND VGND VPWR VPWR _4193_/S sky130_fd_sc_hd__and2_2
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4861__B1 _4590_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3416__B2 _6851_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1499_A _6708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6829_ _6835_/CLK _6829_/D _3959_/B VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5419__S _5424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3719__A2 _5317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4916__B2 _4633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6118__B1 _6019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold180 hold180/A VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5892__A2 _5660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold191 hold191/A VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4080__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5329__S _5334_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4233__S _5236_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6109__B1 _6015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5580__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3591__B1 _4194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3490_ _6969_/Q _5389_/A _3389_/Y _3486_/Y _3489_/X VGND VGND VPWR VPWR _3499_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5883__A2 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5160_ _4417_/B _4691_/Y _4785_/X _5152_/B _4893_/A VGND VGND VPWR VPWR _5160_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4188__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2509 _6933_/Q VGND VGND VPWR VPWR hold921/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4111_ _3616_/Y hold973/A _4115_/S VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _4417_/B _4688_/C _4779_/X _4954_/A _5149_/A VGND VGND VPWR VPWR _5092_/C
+ sky130_fd_sc_hd__o2111a_1
Xhold1808 _7059_/Q VGND VGND VPWR VPWR hold252/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1819 _4246_/X VGND VGND VPWR VPWR hold341/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4042_ _4042_/A0 _4041_/X _4046_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3646__A1 _6983_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3646__B2 _6812_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5399__A1 hold275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5993_ _6015_/B _6017_/A _6019_/B VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__and3_4
XANTENNA__7155__CLK _7180_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6060__A2 _5984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4944_ _4601_/A _4491_/Y _4514_/B _4947_/A VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6348__A0 _3737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4875_ _5124_/B _4930_/A _4875_/C _4875_/D VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__and4_1
XANTENNA__5239__S _5244_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7154__RESET_B fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6614_ _6731_/CLK _6614_/D _6413_/A VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_4
X_3826_ hold26/A _3826_/B VGND VGND VPWR VPWR _3827_/C sky130_fd_sc_hd__nor2_1
XANTENNA__5020__B1 _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4374__A2 _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5571__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6545_ _7194_/CLK _6545_/D VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3982__S _3998_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3757_ input4/X _3307_/Y _3988_/A _6471_/Q VGND VGND VPWR VPWR _3757_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5763__A _5763_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3582__B1 _4262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6476_ _6733_/CLK _6476_/D fanout433/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfstp_2
X_3688_ _6688_/Q _4250_/A _4092_/A _6549_/Q VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__a22o_1
Xoutput230 _7225_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
XANTENNA__4379__A _5001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5427_ _5427_/A0 _5562_/A1 _5433_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
Xoutput241 _3931_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
XFILLER_160_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput252 _3961_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _6785_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
XANTENNA__5874__A2 _5670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput274 _6475_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput285 _6801_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XANTENNA__4098__B _6346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5358_ _5358_/A0 _5529_/A1 _5361_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput296 _6472_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4309_ _4309_/A0 _5189_/A1 _4309_/S VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5289_ _5289_/A0 _5568_/A1 _5289_/S VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
X_7028_ _7136_/CLK _7028_/D fanout471/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6051__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4062__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4053__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5562__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire346 _5770_/Y VGND VGND VPWR VPWR wire346/X sky130_fd_sc_hd__clkbuf_2
Xwire357 _3349_/A VGND VGND VPWR VPWR _3553_/A sky130_fd_sc_hd__buf_12
XFILLER_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3573__B1 _4274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A mgmt_gpio_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7093__SET_B fanout450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5865__A2 _5674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6290__A2 _6339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4228__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _4713_/A _4712_/B VGND VGND VPWR VPWR _5150_/C sky130_fd_sc_hd__and2_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ _3881_/C _5236_/C _3536_/Y hold67/A VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5553__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4591_ _4596_/A _5009_/B VGND VGND VPWR VPWR _4837_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3564__B1 _4170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2264_A _6707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6330_ _6716_/Q _5973_/X _5988_/X _6573_/Q _6329_/X VGND VGND VPWR VPWR _6330_/X
+ sky130_fd_sc_hd__a221o_1
Xhold905 hold905/A VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3542_ _7065_/Q _5497_/A _3539_/Y _6534_/Q _3541_/X VGND VGND VPWR VPWR _3543_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6398__B _6430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold916 hold916/A VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold927 hold927/A VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold938 hold938/A VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5305__A1 wire375/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6261_ _6688_/Q _5980_/X _6017_/X _6770_/Q VGND VGND VPWR VPWR _6261_/X sky130_fd_sc_hd__a22o_1
X_3473_ hold56/X hold88/A VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__nor2_8
Xhold949 hold949/A VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5212_ hold104/X hold95/X _5217_/S VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5856__A2 _5688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6192_ _6216_/A1 _6167_/S _6190_/X _6191_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__o22a_1
XFILLER_142_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2306 _4263_/X VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2317 hold606/X VGND VGND VPWR VPWR _5427_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2328 _7138_/Q VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5143_ _5143_/A _5143_/B VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2339 hold746/X VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5522__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1605 hold331/X VGND VGND VPWR VPWR _5348_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1616 _4203_/X VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1627 hold368/X VGND VGND VPWR VPWR _5280_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5074_ _5103_/A _5074_/B _5074_/C _5156_/A VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__and4_1
Xhold1638 _6722_/Q VGND VGND VPWR VPWR hold294/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3619__A1 _6959_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1649 _6920_/Q VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4816__B1 _4688_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4025_ _4025_/A0 _4024_/X _4029_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6281__A2 _5978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6033__A2 _5986_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6353__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5976_ _6973_/Q _5976_/B VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__and2_1
XFILLER_80_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ _4633_/B _4688_/B _4845_/X _5121_/B _4901_/B VGND VGND VPWR VPWR _4931_/C
+ sky130_fd_sc_hd__o2111a_1
X_4858_ _4705_/Y _4857_/Y _4640_/Y VGND VGND VPWR VPWR _4928_/C sky130_fd_sc_hd__a21o_1
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5544__A1 _5580_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3809_ _6470_/Q _6469_/Q VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__and2_1
X_4789_ _4464_/Y _4570_/B _4674_/Y _4947_/A VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3555__B1 _3336_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6528_ _6821_/CLK _6528_/D fanout442/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_csclk _6549_/CLK VGND VGND VPWR VPWR _6745_/CLK sky130_fd_sc_hd__clkbuf_16
X_6459_ _3958_/A1 _6459_/D _6409_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5847__A2 _5672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1629_A _6819_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5432__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2840 _5575_/X VGND VGND VPWR VPWR hold955/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2851 _6780_/Q VGND VGND VPWR VPWR _3424_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2862 _6681_/Q VGND VGND VPWR VPWR _3919_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2873 _7181_/Q VGND VGND VPWR VPWR _6266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2884 _7160_/Q VGND VGND VPWR VPWR _5729_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4048__S _4055_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2895 _7174_/Q VGND VGND VPWR VPWR _6067_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6272__A2 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4283__A1 _5581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6009__C1 _5995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6024__A2 _6013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4035__A1 _5572_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5783__A1 _7009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5783__B2 _6889_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3794__B1 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5535__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__B1 _5434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6640__RESET_B _3959_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output266_A _6788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5342__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ _6931_/Q _5684_/X _5689_/X _7083_/Q _5829_/X VGND VGND VPWR VPWR _5835_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4026__A1 _5567_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5223__A0 _6818_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_mgmt_gpio_in[4]_A mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5761_ _7064_/Q _5671_/X _5672_/X _6952_/Q VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4712_ _4712_/A _4712_/B _4712_/C VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__3785__B1 _4304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5692_ _7061_/Q _5671_/X _5685_/X _7069_/Q _5691_/X VGND VGND VPWR VPWR _5692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4643_ _4506_/A _4642_/Y _4643_/C _4643_/D VGND VGND VPWR VPWR _5048_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__5526__A1 _5562_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6728__RESET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5517__S _5523_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4574_ _4574_/A _4638_/A VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__nand2_4
Xhold702 hold702/A VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap421 _4677_/A VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__clkbuf_4
Xhold713 hold713/A VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6313_ _6306_/X _6308_/X _6313_/C _6313_/D VGND VGND VPWR VPWR _6314_/C sky130_fd_sc_hd__and4bb_2
Xhold735 hold735/A VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3525_ _6993_/Q _5416_/A _5308_/A _6897_/Q _3524_/X VGND VGND VPWR VPWR _3529_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold746 hold746/A VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold757 hold757/A VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold768 hold768/A VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5829__A2 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6244_ _6645_/Q _5990_/X _5996_/X _6650_/Q VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__a22o_1
Xhold779 hold779/A VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3456_ _6858_/Q _5263_/A _5335_/A _6922_/Q _3455_/X VGND VGND VPWR VPWR _3460_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2103 _6760_/Q VGND VGND VPWR VPWR hold804/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2114 _5334_/X VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6348__S _6354_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3387_ _6780_/Q _3385_/Y _3738_/S VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__mux2_1
X_6175_ _6859_/Q _5983_/X _5988_/X _6875_/Q VGND VGND VPWR VPWR _6175_/X sky130_fd_sc_hd__a22o_1
Xhold2125 _3981_/X VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2136 hold685/X VGND VGND VPWR VPWR _5313_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2147 hold649/X VGND VGND VPWR VPWR _4121_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1402 _5400_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5126_ _5126_/A _5126_/B _5126_/C VGND VGND VPWR VPWR _5127_/D sky130_fd_sc_hd__and3_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1413 _5436_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2158 hold705/X VGND VGND VPWR VPWR _4279_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1424 hold273/X VGND VGND VPWR VPWR _3978_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2169 _4072_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1435 _7030_/Q VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6254__A2 _5976_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1446 _5392_/X VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1457 hold414/X VGND VGND VPWR VPWR _5327_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1468 hold266/X VGND VGND VPWR VPWR _5432_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5057_ _4384_/A _4969_/A _5115_/B _4930_/C _5114_/C VGND VGND VPWR VPWR _5058_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_55_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4265__A1 _5194_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1479 hold415/X VGND VGND VPWR VPWR _4187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout464_A fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ hold326/X _5577_/A1 _4008_/S VGND VGND VPWR VPWR _4008_/X sky130_fd_sc_hd__mux2_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5488__A _5488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5765__A1 _6976_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5959_ _6552_/Q _5673_/X _5954_/X _5955_/X _5958_/X VGND VGND VPWR VPWR _5959_/X
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__5765__B2 _7080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1481_A _7115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1579_A _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5517__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5427__S _5433_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1746_A _6786_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__B1 _5299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6190__A1 _6843_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4740__A2 _4712_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1913_A _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input164_A wb_rstn_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3700__B1 _5245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4286__B _5220_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2670 _4318_/X VGND VGND VPWR VPWR hold560/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__buf_4
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input25_A mask_rev_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2681 hold543/X VGND VGND VPWR VPWR _4238_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6245__A2 _5638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2692 hold733/X VGND VGND VPWR VPWR _5295_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__buf_12
Xhold1980 _6585_/Q VGND VGND VPWR VPWR hold528/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1991 _4027_/X VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5398__A _5398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4008__A1 _5577_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5756__B2 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3767__B1 _5452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6729__SET_B _6411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5508__A1 _5571_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6821__RESET_B fanout449/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5337__S _5343_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3519__B1 _5169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6181__B2 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 _3515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3310_ _3764_/B hold88/A VGND VGND VPWR VPWR _3310_/Y sky130_fd_sc_hd__nor2_8
XFILLER_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4290_ _4290_/A0 _5195_/A1 _4291_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3241_ _6721_/Q VGND VGND VPWR VPWR _3241_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5692__B1 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6236__A2 _5980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4247__A1 _5584_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6931_ _7091_/CLK _6931_/D fanout452/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4798__A2 _4714_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6862_ _6969_/CLK _6862_/D fanout450/X VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5813_ _6858_/Q _5651_/X _5688_/X _6890_/Q _5812_/X VGND VGND VPWR VPWR _5813_/X
+ sky130_fd_sc_hd__a221o_1
X_6793_ _6793_/CLK _6793_/D fanout434/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3758__B1 _4146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5744_ _6895_/Q _5662_/X _5742_/X _5743_/X VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__a211o_1
XFILLER_188_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5675_ _5679_/B _5676_/B VGND VGND VPWR VPWR _5678_/B sky130_fd_sc_hd__and2_4
XANTENNA__3773__A3 _5207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6736_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4626_ _4522_/B _4569_/A _4898_/B _4624_/X _4625_/Y VGND VGND VPWR VPWR _4626_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4557_ _4384_/A _4658_/A _4417_/B _5127_/A VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__o31a_1
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold532 _4049_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold543 hold543/A VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold554 hold554/A VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold565 hold565/A VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3508_ _7097_/Q hold31/A _4182_/A _6628_/Q _3506_/X VGND VGND VPWR VPWR _3515_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold576 hold576/A VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4488_ _4595_/B _4488_/B VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__nand2_4
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold587 _5238_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold598 hold598/A VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _6629_/Q _5971_/X _6007_/X _6530_/Q _6226_/X VGND VGND VPWR VPWR _6230_/B
+ sky130_fd_sc_hd__a221o_1
X_3439_ _7018_/Q _5443_/A _3319_/Y _6800_/Q _3433_/X VGND VGND VPWR VPWR _3444_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5683__B1 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6938_/Q _5980_/X _6017_/X _7074_/Q VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__a22o_1
Xhold1210 _6828_/Q VGND VGND VPWR VPWR hold1210/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _4283_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _6746_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1232 hold268/X VGND VGND VPWR VPWR _5214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6227__A2 _5971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5109_ _4500_/Y _4640_/Y _4919_/C _5125_/B _4757_/A VGND VGND VPWR VPWR _5110_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_111_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1243 _5357_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6089_ _6079_/X _6313_/D _6089_/C _6089_/D VGND VGND VPWR VPWR _6089_/X sky130_fd_sc_hd__and4b_4
Xhold1254 _5510_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1265 _6903_/Q VGND VGND VPWR VPWR hold124/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1276 hold398/X VGND VGND VPWR VPWR _5285_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _6991_/Q VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 hold347/X VGND VGND VPWR VPWR _5267_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5011__A _5011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4061__S _4064_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4412__A_N _4574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4345_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6368_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6374_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6365_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6218__A2 _5991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4229__A1 _5527_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4236__S _4240_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3452__A2 _5272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3790_ _6629_/Q _4188_/A _4262_/A _6697_/Q VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _5460_/A0 _5568_/A1 _5460_/S VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6154__B2 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4411_ _4719_/A _4590_/B VGND VGND VPWR VPWR _4411_/Y sky130_fd_sc_hd__nand2_4
X_5391_ _5391_/A0 _5571_/A1 _5397_/S VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7130_ _7130_/CLK _7130_/D fanout465/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4342_ _4720_/C _4395_/A VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__nor2_4
XFILLER_98_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7061_ _7061_/CLK _7061_/D fanout450/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfstp_2
X_4273_ hold775/X _5448_/A1 _4273_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6012_ _6015_/B _6019_/B _6018_/B VGND VGND VPWR VPWR _6012_/X sky130_fd_sc_hd__and3_4
XFILLER_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3224_ _6720_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4000__A _4000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

