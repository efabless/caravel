magic
tech sky130A
magscale 1 2
timestamp 1636495793
<< metal4 >>
rect -1120 140 14840 560
<< metal5 >>
rect 7840 15260 8190 15400
tri 6930 15120 7070 15260 se
rect 7070 15120 8190 15260
tri 6790 14840 6930 14980 se
rect 6930 14840 8190 15120
tri 5670 14700 5810 14840 se
rect 5810 14700 7280 14840
rect 5670 14630 7280 14700
tri 5530 14420 5670 14560 se
rect 5670 14490 7140 14630
tri 7140 14490 7280 14630 nw
rect 5670 14420 5950 14490
tri 5950 14420 6020 14490 nw
rect 5040 14210 5950 14420
rect 7840 14350 8190 14840
rect 7840 14280 9660 14350
rect 5040 14070 5810 14210
tri 5810 14070 5950 14210 nw
tri 7280 14140 7420 14280 se
rect 7420 14140 9660 14280
tri 6510 14070 6580 14140 se
rect 6580 14070 9660 14140
tri 5880 13440 6510 14070 se
rect 6510 14000 9660 14070
rect 6510 13580 9380 14000
tri 9380 13860 9520 14000 nw
rect 6510 13440 9240 13580
tri 9240 13440 9380 13580 nw
tri 5740 12880 5880 13020 se
rect 5880 12880 9240 13440
rect 5740 12600 9240 12880
tri 9240 12600 9380 12740 sw
rect 2800 11620 3150 12320
rect 5740 12040 9380 12600
tri 5740 11900 5880 12040 ne
rect 5880 11900 9380 12040
tri 9380 11900 9660 12180 sw
rect 5880 11760 7280 11900
tri 7280 11760 7420 11900 nw
rect 7840 11760 9660 11900
rect 5880 11620 6650 11760
rect 2380 11200 3500 11620
tri 2380 11060 2520 11200 ne
rect 2520 10780 3360 11200
tri 3360 11060 3500 11200 nw
tri 5880 11107 6393 11620 ne
rect 6393 11107 6650 11620
tri 6650 11480 6930 11760 nw
rect 7840 10990 8260 11760
tri 8960 11480 9240 11760 ne
rect 9240 11480 9660 11760
tri 13580 11620 14000 12040 se
rect 14000 11620 14280 12040
tri 13160 11200 13580 11620 se
rect 7840 10920 10640 10990
tri 7280 10780 7420 10920 se
rect 7420 10780 10640 10920
rect 2800 10430 3150 10780
rect 6160 10640 10640 10780
rect 2800 10360 4340 10430
tri 6020 10360 6160 10500 se
rect 6160 10360 9940 10640
tri 9940 10360 10220 10640 nw
tri 1680 10220 1820 10360 se
rect 1820 10220 4340 10360
rect 840 10080 4340 10220
tri 140 9240 840 9940 se
rect 840 9380 3780 10080
tri 3780 9940 3920 10080 nw
rect 840 9240 3640 9380
tri 3640 9240 3780 9380 nw
tri 4760 9240 5880 10360 se
rect 5880 10080 9940 10360
rect 5880 9240 9520 10080
tri 9520 9660 9940 10080 nw
rect 11410 10010 11760 10500
tri 12180 10220 13160 11200 se
rect 13160 10920 13580 11200
tri 13580 11060 14140 11620 nw
rect 13160 10500 13440 10920
tri 13440 10780 13580 10920 nw
rect 13160 10220 13300 10500
tri 13300 10360 13440 10500 nw
tri 12110 10010 12180 10080 se
rect 12180 10010 13300 10220
rect 11410 9800 13300 10010
tri 0 8680 140 8820 se
rect 140 8680 3640 9240
rect 0 8120 3640 8680
tri 4200 8540 4760 9100 se
rect 4760 8540 9380 9240
tri 9380 9100 9520 9240 nw
tri 11270 9240 11410 9380 se
rect 11410 9240 13160 9800
tri 13160 9660 13300 9800 nw
tri 11200 9100 11270 9170 se
rect 11270 9100 13160 9240
tri 3640 8120 3780 8260 sw
rect 0 7420 3780 8120
tri 0 7280 140 7420 ne
rect 140 6860 3780 7420
rect -980 6580 -560 6650
tri -560 6580 -490 6650 sw
rect -980 6440 -420 6580
tri -420 6440 -280 6580 sw
tri 140 6440 560 6860 ne
rect 560 6720 3780 6860
tri 4130 7910 4200 7980 se
rect 4200 7910 9380 8540
rect 4130 6860 9380 7910
tri 10360 8120 11200 8960 se
rect 11200 8120 13020 9100
tri 13020 8960 13160 9100 nw
tri 10080 7560 10360 7840 se
rect 10360 7560 13020 8120
tri 9870 7280 10080 7490 se
rect 10080 7280 13020 7560
tri 9730 6860 9870 7000 se
rect 9870 6860 13020 7280
rect 4130 6720 13020 6860
tri 13020 6720 13160 6860 sw
rect 560 6580 1820 6720
tri 1820 6580 1960 6720 nw
tri 2380 6580 2520 6720 ne
rect 2520 6580 13160 6720
rect 560 6440 1400 6580
rect -980 6300 -140 6440
tri -700 6160 -560 6300 ne
rect -560 6160 -140 6300
tri -140 6160 140 6440 sw
rect 700 6160 1400 6440
tri 1400 6300 1680 6580 nw
rect 2800 6440 13160 6580
tri -420 5880 -140 6160 ne
rect -140 6090 280 6160
tri 280 6090 350 6160 sw
rect 700 6090 1330 6160
tri 1330 6090 1400 6160 nw
rect -140 5880 1330 6090
tri 0 5740 140 5880 ne
rect 140 5740 1330 5880
tri 280 5600 420 5740 ne
rect 420 5600 2160 5740
tri 560 5460 700 5600 ne
rect 700 5460 2160 5600
tri 2160 5460 2440 5740 sw
rect 2800 5460 3220 6440
tri 3580 6300 3720 6440 ne
rect 3720 6300 13160 6440
tri 3780 6020 4060 6300 ne
rect 4060 6020 13160 6300
rect 700 5180 3220 5460
rect 4060 5880 10500 6020
tri 10500 5880 10640 6020 nw
rect 4060 5740 10080 5880
tri 10080 5740 10220 5880 nw
tri 4060 5180 4620 5740 ne
rect 4620 5320 10080 5740
tri 10080 5320 10360 5600 sw
rect 4620 5180 10360 5320
rect 980 5040 3220 5180
tri 3220 5040 3360 5180 sw
rect 4620 5040 7140 5180
tri 7140 5040 7280 5180 nw
tri 7700 5040 7840 5180 ne
rect 7840 5040 10360 5180
tri 980 4900 1120 5040 ne
rect 1120 4900 3640 5040
tri 3640 4900 3780 5040 sw
tri 1400 4060 2240 4900 ne
rect 2240 3780 4200 4900
rect 4620 4760 6020 5040
tri 6020 4900 6160 5040 nw
tri 4620 4340 5040 4760 ne
rect 5040 4340 5600 4760
tri 5600 4340 6020 4760 nw
rect 7980 4760 10360 5040
tri 4200 3780 4760 4340 sw
tri 5040 4200 5180 4340 ne
rect 5180 3780 5600 4340
tri 2100 3500 2240 3640 se
rect 2240 3500 5600 3780
rect 2100 3360 5600 3500
tri 5600 3360 6020 3780 sw
rect 2100 3220 6300 3360
tri 6300 3220 6440 3360 sw
rect 2100 3080 6860 3220
tri 6860 3080 7000 3220 sw
rect 7980 3080 8540 4760
tri 8960 4620 9100 4760 ne
rect 9100 4620 10360 4760
tri 10360 4620 10780 5040 sw
tri 9660 4340 9940 4620 ne
rect 9940 4480 10780 4620
rect 11340 4480 11760 6020
tri 12180 5880 12320 6020 ne
rect 12320 5880 13160 6020
tri 13160 5880 13440 6160 sw
tri 12600 5320 13160 5880 ne
rect 13160 5320 13440 5880
tri 12460 4620 12740 4900 se
rect 12740 4760 14000 4900
tri 14000 4760 14140 4900 sw
rect 12740 4620 14140 4760
tri 12180 4480 12320 4620 se
rect 12320 4480 14140 4620
rect 9940 4410 14140 4480
rect 9940 4340 14000 4410
tri 10360 4060 10640 4340 ne
rect 10640 4060 14000 4340
rect 10640 3710 14840 4060
rect 10640 3640 14140 3710
tri 9660 3080 10220 3640 se
rect 10220 3500 14140 3640
rect 10220 3080 14000 3500
tri 14000 3360 14140 3500 nw
rect 2100 2800 14000 3080
rect 2100 2660 5950 2800
tri 2100 2520 2240 2660 ne
rect 2240 2380 5950 2660
rect 6300 2660 14000 2800
rect 6300 2380 6790 2660
rect 2240 2240 6790 2380
rect 7140 2520 13720 2660
tri 13720 2520 13860 2660 nw
rect 7140 2240 7700 2520
rect 2240 2100 7700 2240
rect 8050 2100 8540 2520
rect 8890 2100 9380 2520
rect 9730 2100 13720 2520
rect 2240 1960 13720 2100
tri 2240 1820 2380 1960 ne
rect 2380 1540 13580 1960
tri 13580 1820 13720 1960 nw
tri 2380 1400 2520 1540 ne
rect 2520 1260 13160 1540
tri 2520 840 2940 1260 ne
rect 2940 700 13160 1260
tri 13160 1120 13580 1540 nw
tri 2940 560 3080 700 ne
rect 3080 560 13160 700
<< fillblock >>
rect -2520 10640 -2240 10920
rect -1260 10360 15000 15560
rect -1960 9800 15000 10360
rect -1260 0 15000 9800
<< end >>
