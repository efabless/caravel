module caravel (clock,
    flash_clk,
    flash_csb,
    flash_io0,
    flash_io1,
    gpio,
    resetb,
    vccd,
    vccd1,
    vccd2,
    vdda,
    vdda1,
    vdda1_2,
    vdda2,
    vddio,
    vddio_2,
    vssa,
    vssa1,
    vssa1_2,
    vssa2,
    vssd,
    vssd1,
    vssd2,
    vssio,
    vssio_2,
    mprj_io);
 input clock;
 inout flash_clk;
 inout flash_csb;
 inout flash_io0;
 inout flash_io1;
 inout gpio;
 input resetb;
 inout vccd;
 inout vccd1;
 inout vccd2;
 inout vdda;
 inout vdda1;
 inout vdda1_2;
 inout vdda2;
 inout vddio;
 inout vddio_2;
 inout vssa;
 inout vssa1;
 inout vssa1_2;
 inout vssa2;
 inout vssd;
 inout vssd1;
 inout vssd2;
 inout vssio;
 inout vssio_2;
 inout [37:0] mprj_io;

 wire vdda2_core;
 wire vssa2_core;
 wire vdda1_core;
 wire vssa1_core;
 wire \gpio_control_bidir_2[2]/zero ;
 wire \gpio_control_bidir_2[2]/one ;
 wire \gpio_control_bidir_2[1]/resetn ;
 wire \gpio_control_bidir_2[1]/serial_clock ;
 wire \gpio_control_bidir_2[1]/serial_data_in ;
 wire \gpio_control_bidir_2[1]/serial_load ;
 wire \gpio_defaults_block_32/VPWR ;
 wire \gpio_defaults_block_32/VGND ;
 wire \gpio_control_in_1a[5]/zero ;
 wire \gpio_control_in_1a[5]/one ;
 wire \gpio_control_in_1[0]/resetn ;
 wire \gpio_control_in_1[0]/serial_clock ;
 wire \gpio_control_in_1[0]/serial_data_in ;
 wire \gpio_control_in_1[0]/serial_load ;
 wire \gpio_defaults_block_31/VPWR ;
 wire \gpio_defaults_block_31/VGND ;
 wire \gpio_defaults_block_10/VPWR ;
 wire \gpio_defaults_block_10/VGND ;
 wire \gpio_defaults_block_21/VPWR ;
 wire \gpio_defaults_block_21/VGND ;
 wire \gpio_defaults_block_20/VPWR ;
 wire \gpio_defaults_block_20/VGND ;
 wire \por/vss3v3 ;
 wire \por/vdd3v3 ;
 wire \rstb_level/VGND ;
 wire \rstb_level/VPWR ;
 wire vssd1_core;
 wire vccd1_core;
 wire \gpio_defaults_block_30/VPWR ;
 wire \gpio_defaults_block_30/VGND ;
 wire \gpio_control_in_1[8]/zero ;
 wire \gpio_control_in_1[8]/one ;
 wire \gpio_control_in_1[8]/resetn ;
 wire \gpio_control_in_1[8]/serial_clock ;
 wire \gpio_control_in_1[8]/serial_data_in ;
 wire \gpio_control_in_1[8]/serial_load ;
 wire \gpio_control_in_2[2]/zero ;
 wire \gpio_control_in_2[2]/one ;
 wire \gpio_control_in_2[1]/resetn ;
 wire \gpio_control_in_2[1]/serial_clock ;
 wire \gpio_control_in_2[1]/serial_data_in ;
 wire \gpio_control_in_2[1]/serial_load ;
 wire \housekeeping/serial_clock ;
 wire \housekeeping/serial_resetn ;
 wire \housekeeping/serial_load ;
 wire \housekeeping/serial_data_1 ;
 wire \housekeeping/serial_data_2 ;
 wire \soc/flash_clk ;
 wire \soc/flash_io0_di ;
 wire \soc/flash_io0_do ;
 wire \soc/flash_io0_oeb ;
 wire \soc/flash_io1_di ;
 wire \soc/flash_io1_do ;
 wire \soc/flash_io1_oeb ;
 wire \soc/flash_io2_di ;
 wire \soc/flash_io2_do ;
 wire \soc/flash_io2_oeb ;
 wire \soc/flash_io3_di ;
 wire \soc/flash_io3_do ;
 wire \soc/flash_io3_oeb ;
 wire \housekeeping/usr2_vdd_pwrgood ;
 wire \housekeeping/usr1_vdd_pwrgood ;
 wire \housekeeping/usr2_vcc_pwrgood ;
 wire \housekeeping/usr1_vcc_pwrgood ;
 wire \soc/mprj_we_o ;
 wire \gpio_control_bidir_1[1]/zero ;
 wire \gpio_control_bidir_1[1]/one ;
 wire \gpio_control_in_1a[0]/resetn ;
 wire \gpio_control_in_1a[0]/serial_clock ;
 wire \gpio_control_in_1a[0]/serial_data_in ;
 wire \gpio_control_in_1a[0]/serial_load ;
 wire \gpio_control_in_2[4]/zero ;
 wire \gpio_control_in_2[4]/one ;
 wire \gpio_control_in_2[3]/resetn ;
 wire \gpio_control_in_2[3]/serial_clock ;
 wire \gpio_control_in_2[3]/serial_data_in ;
 wire \gpio_control_in_2[3]/serial_load ;
 wire \gpio_control_in_1[1]/zero ;
 wire \gpio_control_in_1[1]/one ;
 wire \gpio_control_in_1[2]/resetn ;
 wire \gpio_control_in_1[2]/serial_clock ;
 wire \gpio_control_in_1[2]/serial_data_in ;
 wire \gpio_control_in_1[2]/serial_load ;
 wire \gpio_control_in_2[6]/zero ;
 wire \gpio_control_in_2[6]/one ;
 wire \gpio_control_in_2[5]/resetn ;
 wire \gpio_control_in_2[5]/serial_clock ;
 wire \gpio_control_in_2[5]/serial_data_in ;
 wire \gpio_control_in_2[5]/serial_load ;
 wire \gpio_control_in_1a[0]/zero ;
 wire \gpio_control_in_1a[0]/one ;
 wire \gpio_control_in_1a[1]/resetn ;
 wire \gpio_control_in_1a[1]/serial_clock ;
 wire \gpio_control_in_1a[1]/serial_data_in ;
 wire \gpio_control_in_1a[1]/serial_load ;
 wire \gpio_control_in_2[11]/zero ;
 wire \gpio_control_in_2[11]/one ;
 wire \gpio_control_in_2[10]/resetn ;
 wire \gpio_control_in_2[10]/serial_clock ;
 wire \gpio_control_in_2[10]/serial_data_in ;
 wire \gpio_control_in_2[10]/serial_load ;
 wire \gpio_control_in_1[3]/zero ;
 wire \gpio_control_in_1[3]/one ;
 wire \gpio_control_in_1[4]/resetn ;
 wire \gpio_control_in_1[4]/serial_clock ;
 wire \gpio_control_in_1[4]/serial_data_in ;
 wire \gpio_control_in_1[4]/serial_load ;
 wire \gpio_control_in_2[8]/zero ;
 wire \gpio_control_in_2[8]/one ;
 wire \gpio_control_in_2[7]/resetn ;
 wire \gpio_control_in_2[7]/serial_clock ;
 wire \gpio_control_in_2[7]/serial_data_in ;
 wire \gpio_control_in_2[7]/serial_load ;
 wire \gpio_control_in_1a[2]/zero ;
 wire \gpio_control_in_1a[2]/one ;
 wire \gpio_control_in_1a[3]/resetn ;
 wire \gpio_control_in_1a[3]/serial_clock ;
 wire \gpio_control_in_1a[3]/serial_data_in ;
 wire \gpio_control_in_1a[3]/serial_load ;
 wire \gpio_control_in_2[13]/zero ;
 wire \gpio_control_in_2[13]/one ;
 wire \gpio_control_in_2[12]/resetn ;
 wire \gpio_control_in_2[12]/serial_clock ;
 wire \gpio_control_in_2[12]/serial_data_in ;
 wire \gpio_control_in_2[12]/serial_load ;
 wire \gpio_control_in_1[5]/zero ;
 wire \gpio_control_in_1[5]/one ;
 wire \gpio_control_in_1[6]/resetn ;
 wire \gpio_control_in_1[6]/serial_clock ;
 wire \gpio_control_in_1[6]/serial_data_in ;
 wire \gpio_control_in_1[6]/serial_load ;
 wire \gpio_control_bidir_2[1]/zero ;
 wire \gpio_control_bidir_2[1]/one ;
 wire \gpio_control_bidir_2[0]/resetn ;
 wire \gpio_control_bidir_2[0]/serial_clock ;
 wire \gpio_control_bidir_2[0]/serial_data_in ;
 wire \gpio_control_bidir_2[0]/serial_load ;
 wire \gpio_control_in_2[15]/zero ;
 wire \gpio_control_in_2[15]/one ;
 wire \gpio_control_in_2[14]/resetn ;
 wire \gpio_control_in_2[14]/serial_clock ;
 wire \gpio_control_in_2[14]/serial_data_in ;
 wire \gpio_control_in_2[14]/serial_load ;
 wire \gpio_defaults_block_9/VPWR ;
 wire \gpio_defaults_block_9/VGND ;
 wire vccd_core;
 wire \pll/resetb ;
 wire vccd2_core;
 wire vssd2_core;
 wire \mprj/user_clock2 ;
 wire \mprj/wbs_we_i ;
 wire \mprj/wbs_stb_i ;
 wire \mprj/wbs_cyc_i ;
 wire \mprj/wbs_ack_o ;
 wire \mprj/wb_rst_i ;
 wire \mprj/wb_clk_i ;
 wire \gpio_control_in_1a[4]/zero ;
 wire \gpio_control_in_1a[4]/one ;
 wire \gpio_control_in_1a[5]/resetn ;
 wire \gpio_control_in_1a[5]/serial_clock ;
 wire \gpio_control_in_1a[5]/serial_data_in ;
 wire \gpio_control_in_1a[5]/serial_load ;
 wire \gpio_defaults_block_8/VPWR ;
 wire \gpio_defaults_block_8/VGND ;
 wire \gpio_control_in_1[7]/zero ;
 wire \gpio_control_in_1[7]/one ;
 wire \gpio_defaults_block_7/VPWR ;
 wire \gpio_defaults_block_7/VGND ;
 wire \gpio_defaults_block_6/VPWR ;
 wire \gpio_defaults_block_6/VGND ;
 wire \gpio_control_in_2[1]/zero ;
 wire \gpio_control_in_2[1]/one ;
 wire \gpio_control_in_2[0]/resetn ;
 wire \gpio_control_in_2[0]/serial_clock ;
 wire \gpio_control_in_2[0]/serial_load ;
 wire \gpio_defaults_block_4/VGND ;
 wire \gpio_defaults_block_4/VPWR ;
 wire \gpio_defaults_block_5/VPWR ;
 wire \gpio_defaults_block_5/VGND ;
 wire \gpio_control_in_1[9]/zero ;
 wire \gpio_control_in_1[9]/one ;
 wire \gpio_control_in_1[9]/resetn ;
 wire \gpio_control_in_1[9]/serial_clock ;
 wire \gpio_control_in_1[9]/serial_data_in ;
 wire \gpio_control_in_1[9]/serial_load ;
 wire \gpio_control_bidir_1[0]/zero ;
 wire \gpio_control_bidir_1[0]/one ;
 wire \gpio_control_bidir_1[1]/resetn ;
 wire \gpio_control_bidir_1[1]/serial_clock ;
 wire \gpio_control_bidir_1[1]/serial_data_in ;
 wire \gpio_control_bidir_1[1]/serial_load ;
 wire \gpio_defaults_block_3/VGND ;
 wire \gpio_defaults_block_3/VPWR ;
 wire \gpio_defaults_block_2/VGND ;
 wire \gpio_defaults_block_2/VPWR ;
 wire \gpio_control_in_2[3]/zero ;
 wire \gpio_control_in_2[3]/one ;
 wire \gpio_control_in_2[2]/resetn ;
 wire \gpio_control_in_2[2]/serial_clock ;
 wire \gpio_control_in_2[2]/serial_data_in ;
 wire \gpio_control_in_2[2]/serial_load ;
 wire \gpio_defaults_block_1/VGND ;
 wire \gpio_defaults_block_1/VPWR ;
 wire \gpio_defaults_block_0/VGND ;
 wire \gpio_defaults_block_0/VPWR ;
 wire \gpio_control_in_1[0]/zero ;
 wire \gpio_control_in_1[0]/one ;
 wire \gpio_control_in_1[1]/resetn ;
 wire \gpio_control_in_1[1]/serial_clock ;
 wire \gpio_control_in_1[1]/serial_data_in ;
 wire \gpio_control_in_1[1]/serial_load ;
 wire \gpio_control_in_2[5]/zero ;
 wire \gpio_control_in_2[5]/one ;
 wire \gpio_control_in_2[4]/resetn ;
 wire \gpio_control_in_2[4]/serial_clock ;
 wire \gpio_control_in_2[4]/serial_data_in ;
 wire \gpio_control_in_2[4]/serial_load ;
 wire \gpio_control_in_1[10]/zero ;
 wire \gpio_control_in_1[10]/one ;
 wire \gpio_control_in_1[10]/resetn ;
 wire \gpio_control_in_1[10]/resetn_out ;
 wire \gpio_control_in_1[10]/serial_clock ;
 wire \gpio_control_in_1[10]/serial_clock_out ;
 wire \gpio_control_in_1[9]/serial_data_out ;
 wire \gpio_control_in_1[10]/serial_data_out ;
 wire \gpio_control_in_1[10]/serial_load ;
 wire \gpio_control_in_1[10]/serial_load_out ;
 wire \gpio_control_in_2[10]/zero ;
 wire \gpio_control_in_2[10]/one ;
 wire \gpio_control_in_2[9]/resetn ;
 wire \gpio_control_in_2[9]/serial_clock ;
 wire \gpio_control_in_2[9]/serial_data_in ;
 wire \gpio_control_in_2[9]/serial_load ;
 wire \gpio_defaults_block_29/VPWR ;
 wire \gpio_defaults_block_29/VGND ;
 wire \gpio_control_in_1[2]/zero ;
 wire \gpio_control_in_1[2]/one ;
 wire \gpio_control_in_1[3]/resetn ;
 wire \gpio_control_in_1[3]/serial_clock ;
 wire \gpio_control_in_1[3]/serial_data_in ;
 wire \gpio_control_in_1[3]/serial_load ;
 wire \gpio_defaults_block_19/VPWR ;
 wire \gpio_defaults_block_19/VGND ;
 wire \gpio_defaults_block_18/VPWR ;
 wire \gpio_defaults_block_18/VGND ;
 wire \clocking/ext_clk_sel ;
 wire \housekeeping/reset ;
 wire \clocking/user_clk ;
 wire \gpio_defaults_block_28/VPWR ;
 wire \gpio_defaults_block_28/VGND ;
 wire \gpio_control_in_2[7]/zero ;
 wire \gpio_control_in_2[7]/one ;
 wire \gpio_control_in_2[6]/resetn ;
 wire \gpio_control_in_2[6]/serial_clock ;
 wire \gpio_control_in_2[6]/serial_data_in ;
 wire \gpio_control_in_2[6]/serial_load ;
 wire \gpio_defaults_block_17/VPWR ;
 wire \gpio_defaults_block_17/VGND ;
 wire \spare_logic_block_3/spare_xib ;
 wire \gpio_control_in_1a[1]/zero ;
 wire \gpio_control_in_1a[1]/one ;
 wire \gpio_control_in_1a[2]/resetn ;
 wire \gpio_control_in_1a[2]/serial_clock ;
 wire \gpio_control_in_1a[2]/serial_data_in ;
 wire \gpio_control_in_1a[2]/serial_load ;
 wire \gpio_control_in_2[12]/zero ;
 wire \gpio_control_in_2[12]/one ;
 wire \gpio_control_in_2[11]/resetn ;
 wire \gpio_control_in_2[11]/serial_clock ;
 wire \gpio_control_in_2[11]/serial_data_in ;
 wire \gpio_control_in_2[11]/serial_load ;
 wire \gpio_defaults_block_27/VPWR ;
 wire \gpio_defaults_block_27/VGND ;
 wire \gpio_defaults_block_16/VPWR ;
 wire \gpio_defaults_block_16/VGND ;
 wire \por/porb_h ;
 wire \por/porb_l ;
 wire vssd_core;
 wire \gpio_defaults_block_37/VPWR ;
 wire \gpio_defaults_block_37/VGND ;
 wire \spare_logic_block_2/spare_xib ;
 wire \gpio_defaults_block_26/VPWR ;
 wire \gpio_defaults_block_26/VGND ;
 wire \gpio_control_in_1[4]/zero ;
 wire \gpio_control_in_1[4]/one ;
 wire \gpio_control_in_1[5]/resetn ;
 wire \gpio_control_in_1[5]/serial_clock ;
 wire \gpio_control_in_1[5]/serial_data_in ;
 wire \gpio_control_in_1[5]/serial_load ;
 wire \gpio_defaults_block_15/VPWR ;
 wire \gpio_defaults_block_15/VGND ;
 wire \spare_logic_block_1/spare_xib ;
 wire \gpio_defaults_block_36/VPWR ;
 wire \gpio_defaults_block_36/VGND ;
 wire \gpio_control_in_2[9]/zero ;
 wire \gpio_control_in_2[9]/one ;
 wire \gpio_control_in_2[8]/resetn ;
 wire \gpio_control_in_2[8]/serial_clock ;
 wire \gpio_control_in_2[8]/serial_data_in ;
 wire \gpio_control_in_2[8]/serial_load ;
 wire \gpio_defaults_block_25/VPWR ;
 wire \gpio_defaults_block_25/VGND ;
 wire \gpio_defaults_block_14/VPWR ;
 wire \gpio_defaults_block_14/VGND ;
 wire \soc/sram_ro_csb ;
 wire \soc/sram_ro_clk ;
 wire \soc/debug_in ;
 wire \soc/debug_mode ;
 wire \soc/debug_oeb ;
 wire \soc/debug_out ;
 wire \soc/trap ;
 wire \soc/spi_sdoenb ;
 wire \soc/spi_sdo ;
 wire \soc/spi_sck ;
 wire \soc/spi_csb ;
 wire \soc/spi_sdi ;
 wire \soc/ser_rx ;
 wire \soc/ser_tx ;
 wire \soc/spi_enabled ;
 wire \soc/uart_enabled ;
 wire \soc/qspi_enabled ;
 wire \soc/hk_ack_i ;
 wire \soc/hk_stb_o ;
 wire \soc/hk_cyc_o ;
 wire \soc/flash_csb ;
 wire \soc/core_clk ;
 wire \soc/core_rstn ;
 wire \soc/mprj_wb_iena ;
 wire \soc/mprj_stb_o ;
 wire \soc/mprj_cyc_o ;
 wire \soc/mprj_ack_i ;
 wire \spare_logic_block_0/spare_xib ;
 wire \gpio_control_bidir_2[0]/zero ;
 wire \gpio_control_bidir_2[0]/one ;
 wire \gpio_control_in_2[15]/resetn ;
 wire \gpio_control_in_2[15]/serial_clock ;
 wire \gpio_control_in_2[15]/serial_data_in ;
 wire \gpio_control_in_2[15]/serial_load ;
 wire \gpio_defaults_block_35/VPWR ;
 wire \gpio_defaults_block_35/VGND ;
 wire \gpio_control_in_2[14]/zero ;
 wire \gpio_control_in_2[14]/one ;
 wire \gpio_control_in_2[13]/resetn ;
 wire \gpio_control_in_2[13]/serial_clock ;
 wire \gpio_control_in_2[13]/serial_data_in ;
 wire \gpio_control_in_2[13]/serial_load ;
 wire \gpio_control_in_1a[3]/zero ;
 wire \gpio_control_in_1a[3]/one ;
 wire \gpio_control_in_1a[4]/resetn ;
 wire \gpio_control_in_1a[4]/serial_clock ;
 wire \gpio_control_in_1a[4]/serial_data_in ;
 wire \gpio_control_in_1a[4]/serial_load ;
 wire \gpio_defaults_block_13/VPWR ;
 wire \gpio_defaults_block_13/VGND ;
 wire \gpio_defaults_block_24/VPWR ;
 wire \gpio_defaults_block_24/VGND ;
 wire \padframe/vssa ;
 wire \padframe/vssd ;
 wire \padframe/vdda ;
 wire \padframe/vssa1 ;
 wire \padframe/vdda1 ;
 wire \padframe/vccd ;
 wire \padframe/vdda2 ;
 wire \padframe/vddio ;
 wire \padframe/vssa2 ;
 wire \padframe/vssio ;
 wire \soc/gpio_outenb_pad ;
 wire \soc/gpio_out_pad ;
 wire \soc/gpio_inenb_pad ;
 wire \soc/gpio_mode0_pad ;
 wire \soc/gpio_in_pad ;
 wire \padframe/flash_io1_do_core ;
 wire \padframe/flash_io1_di_core ;
 wire \padframe/flash_io0_do_core ;
 wire \padframe/flash_io0_di_core ;
 wire \padframe/flash_clk_oeb_core ;
 wire \padframe/flash_clk_core ;
 wire \padframe/flash_clk_ieb_core ;
 wire \padframe/flash_csb_oeb_core ;
 wire \padframe/flash_csb_core ;
 wire \padframe/flash_csb_ieb_core ;
 wire \por/por_l ;
 wire \pll/osc ;
 wire \rstb_level/A ;
 wire \padframe/flash_io1_ieb_core ;
 wire \soc/gpio_mode1_pad ;
 wire \padframe/flash_io0_ieb_core ;
 wire \padframe/flash_io1_oeb_core ;
 wire \padframe/flash_io0_oeb_core ;
 wire \pll/enable ;
 wire \pll/dco ;
 wire \gpio_control_in_2[15]/vccd ;
 wire \gpio_control_in_2[15]/vssd ;
 wire \gpio_defaults_block_12/VPWR ;
 wire \gpio_defaults_block_12/VGND ;
 wire \gpio_control_in_1[6]/zero ;
 wire \gpio_control_in_1[6]/one ;
 wire \gpio_control_in_1[7]/resetn ;
 wire \gpio_control_in_1[7]/serial_clock ;
 wire \gpio_control_in_1[7]/serial_data_in ;
 wire \gpio_control_in_1[7]/serial_load ;
 wire \gpio_defaults_block_23/VPWR ;
 wire \gpio_defaults_block_23/VGND ;
 wire \gpio_defaults_block_33/VPWR ;
 wire \gpio_defaults_block_33/VGND ;
 wire \gpio_defaults_block_11/VPWR ;
 wire \gpio_defaults_block_11/VGND ;
 wire \gpio_defaults_block_22/VPWR ;
 wire \gpio_defaults_block_22/VGND ;
 wire \gpio_control_in_2[0]/zero ;
 wire \gpio_control_in_2[0]/one ;
 wire \gpio_control_in_2[0]/resetn_out ;
 wire \gpio_control_in_2[0]/serial_clock_out ;
 wire \gpio_control_in_2[0]/serial_data_in ;
 wire \gpio_control_in_2[0]/serial_data_out ;
 wire \gpio_control_in_2[0]/serial_load_out ;
 wire [2:0] \clocking/sel ;
 wire [2:0] \clocking/sel2 ;
 wire [12:0] \gpio_control_in_2[15]/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_0/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_1/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_10/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_11/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_12/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_13/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_14/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_15/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_16/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_17/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_18/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_19/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_2/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_20/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_21/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_22/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_23/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_24/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_25/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_26/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_27/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_28/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_29/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_3/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_30/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_31/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_32/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_33/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_35/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_36/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_37/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_4/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_5/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_6/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_7/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_8/gpio_defaults ;
 wire [12:0] \gpio_defaults_block_9/gpio_defaults ;
 wire [37:0] \housekeeping/mgmt_gpio_in ;
 wire [37:0] \housekeeping/mgmt_gpio_oeb ;
 wire [37:0] \housekeeping/mgmt_gpio_out ;
 wire [3:0] \housekeeping/pwr_ctrl_out ;
 wire [28:0] \mprj/analog_io ;
 wire [37:0] \mprj/io_in ;
 wire [37:0] \mprj/io_oeb ;
 wire [37:0] \mprj/io_out ;
 wire [127:0] \mprj/la_data_in ;
 wire [127:0] \mprj/la_data_out ;
 wire [127:0] \mprj/la_oenb ;
 wire [2:0] \mprj/user_irq ;
 wire [31:0] \mprj/wbs_adr_i ;
 wire [31:0] \mprj/wbs_dat_i ;
 wire [31:0] \mprj/wbs_dat_o ;
 wire [3:0] \mprj/wbs_sel_i ;
 wire [37:0] \padframe/mprj_io_analog_en ;
 wire [37:0] \padframe/mprj_io_analog_pol ;
 wire [37:0] \padframe/mprj_io_analog_sel ;
 wire [113:0] \padframe/mprj_io_dm ;
 wire [37:0] \padframe/mprj_io_holdover ;
 wire [37:0] \padframe/mprj_io_ib_mode_sel ;
 wire [37:0] \padframe/mprj_io_in ;
 wire [37:0] \padframe/mprj_io_inp_dis ;
 wire [37:0] \padframe/mprj_io_oeb ;
 wire [37:0] \padframe/mprj_io_out ;
 wire [37:0] \padframe/mprj_io_slow_sel ;
 wire [37:0] \padframe/mprj_io_vtrip_sel ;
 wire [1:0] \pll/clockp ;
 wire [4:0] \pll/div ;
 wire [25:0] \pll/ext_trim ;
 wire [31:0] \soc/hk_dat_i ;
 wire [5:0] \soc/irq ;
 wire [127:0] \soc/la_iena ;
 wire [127:0] \soc/la_input ;
 wire [127:0] \soc/la_oenb ;
 wire [127:0] \soc/la_output ;
 wire [31:0] \soc/mprj_adr_o ;
 wire [31:0] \soc/mprj_dat_i ;
 wire [31:0] \soc/mprj_dat_o ;
 wire [3:0] \soc/mprj_sel_o ;
 wire [7:0] \soc/sram_ro_addr ;
 wire [31:0] \soc/sram_ro_data ;
 wire [2:0] \soc/user_irq_ena ;
 wire [1:0] \spare_logic_block_0/spare_xfq ;
 wire [1:0] \spare_logic_block_0/spare_xfqn ;
 wire [3:0] \spare_logic_block_0/spare_xi ;
 wire [1:0] \spare_logic_block_0/spare_xmx ;
 wire [1:0] \spare_logic_block_0/spare_xna ;
 wire [1:0] \spare_logic_block_0/spare_xno ;
 wire [26:0] \spare_logic_block_0/spare_xz ;
 wire [1:0] \spare_logic_block_1/spare_xfq ;
 wire [1:0] \spare_logic_block_1/spare_xfqn ;
 wire [3:0] \spare_logic_block_1/spare_xi ;
 wire [1:0] \spare_logic_block_1/spare_xmx ;
 wire [1:0] \spare_logic_block_1/spare_xna ;
 wire [1:0] \spare_logic_block_1/spare_xno ;
 wire [26:0] \spare_logic_block_1/spare_xz ;
 wire [1:0] \spare_logic_block_2/spare_xfq ;
 wire [1:0] \spare_logic_block_2/spare_xfqn ;
 wire [3:0] \spare_logic_block_2/spare_xi ;
 wire [1:0] \spare_logic_block_2/spare_xmx ;
 wire [1:0] \spare_logic_block_2/spare_xna ;
 wire [1:0] \spare_logic_block_2/spare_xno ;
 wire [26:0] \spare_logic_block_2/spare_xz ;
 wire [1:0] \spare_logic_block_3/spare_xfq ;
 wire [1:0] \spare_logic_block_3/spare_xfqn ;
 wire [3:0] \spare_logic_block_3/spare_xi ;
 wire [1:0] \spare_logic_block_3/spare_xmx ;
 wire [1:0] \spare_logic_block_3/spare_xna ;
 wire [1:0] \spare_logic_block_3/spare_xno ;
 wire [26:0] \spare_logic_block_3/spare_xz ;
 wire [31:0] \user_id_value/mask_rev ;

 xres_buf rstb_level (.A(\rstb_level/A ),
    .X(\pll/resetb ));
 gpio_defaults_block_1803 gpio_defaults_block_0 (.gpio_defaults({\gpio_defaults_block_0/gpio_defaults [12],
    \gpio_defaults_block_0/gpio_defaults [11],
    \gpio_defaults_block_0/gpio_defaults [10],
    \gpio_defaults_block_0/gpio_defaults [9],
    \gpio_defaults_block_0/gpio_defaults [8],
    \gpio_defaults_block_0/gpio_defaults [7],
    \gpio_defaults_block_0/gpio_defaults [6],
    \gpio_defaults_block_0/gpio_defaults [5],
    \gpio_defaults_block_0/gpio_defaults [4],
    \gpio_defaults_block_0/gpio_defaults [3],
    \gpio_defaults_block_0/gpio_defaults [2],
    \gpio_defaults_block_0/gpio_defaults [1],
    \gpio_defaults_block_0/gpio_defaults [0]}));
 gpio_control_block \gpio_control_bidir_1[0]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [0]),
    .mgmt_gpio_oeb(\housekeeping/mgmt_gpio_oeb [0]),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_out [0]),
    .one(\gpio_control_bidir_1[0]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [0]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [0]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [0]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [0]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [0]),
    .pad_gpio_in(\padframe/mprj_io_in [0]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [0]),
    .pad_gpio_out(\padframe/mprj_io_out [0]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [0]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [0]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [0]),
    .resetn(\housekeeping/serial_resetn ),
    .resetn_out(\gpio_control_bidir_1[1]/resetn ),
    .serial_clock(\housekeeping/serial_clock ),
    .serial_clock_out(\gpio_control_bidir_1[1]/serial_clock ),
    .serial_data_in(\housekeeping/serial_data_1 ),
    .serial_data_out(\gpio_control_bidir_1[1]/serial_data_in ),
    .serial_load(\housekeeping/serial_load ),
    .serial_load_out(\gpio_control_bidir_1[1]/serial_load ),
    .user_gpio_in(\mprj/io_in [0]),
    .user_gpio_oeb(\mprj/io_oeb [0]),
    .user_gpio_out(\mprj/io_out [0]),
    .zero(\gpio_control_bidir_1[0]/zero ),
    .gpio_defaults({\gpio_defaults_block_0/gpio_defaults [12],
    \gpio_defaults_block_0/gpio_defaults [11],
    \gpio_defaults_block_0/gpio_defaults [10],
    \gpio_defaults_block_0/gpio_defaults [9],
    \gpio_defaults_block_0/gpio_defaults [8],
    \gpio_defaults_block_0/gpio_defaults [7],
    \gpio_defaults_block_0/gpio_defaults [6],
    \gpio_defaults_block_0/gpio_defaults [5],
    \gpio_defaults_block_0/gpio_defaults [4],
    \gpio_defaults_block_0/gpio_defaults [3],
    \gpio_defaults_block_0/gpio_defaults [2],
    \gpio_defaults_block_0/gpio_defaults [1],
    \gpio_defaults_block_0/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [2],
    \padframe/mprj_io_dm [1],
    \padframe/mprj_io_dm [0]}));
 simple_por por (.porb_h(\por/porb_h ),
    .por_l(\por/por_l ),
    .porb_l(\por/porb_l ));
 user_id_programming user_id_value (.mask_rev({\user_id_value/mask_rev [31],
    \user_id_value/mask_rev [30],
    \user_id_value/mask_rev [29],
    \user_id_value/mask_rev [28],
    \user_id_value/mask_rev [27],
    \user_id_value/mask_rev [26],
    \user_id_value/mask_rev [25],
    \user_id_value/mask_rev [24],
    \user_id_value/mask_rev [23],
    \user_id_value/mask_rev [22],
    \user_id_value/mask_rev [21],
    \user_id_value/mask_rev [20],
    \user_id_value/mask_rev [19],
    \user_id_value/mask_rev [18],
    \user_id_value/mask_rev [17],
    \user_id_value/mask_rev [16],
    \user_id_value/mask_rev [15],
    \user_id_value/mask_rev [14],
    \user_id_value/mask_rev [13],
    \user_id_value/mask_rev [12],
    \user_id_value/mask_rev [11],
    \user_id_value/mask_rev [10],
    \user_id_value/mask_rev [9],
    \user_id_value/mask_rev [8],
    \user_id_value/mask_rev [7],
    \user_id_value/mask_rev [6],
    \user_id_value/mask_rev [5],
    \user_id_value/mask_rev [4],
    \user_id_value/mask_rev [3],
    \user_id_value/mask_rev [2],
    \user_id_value/mask_rev [1],
    \user_id_value/mask_rev [0]}));
 digital_pll pll (.dco(\pll/dco ),
    .enable(\pll/enable ),
    .osc(\pll/osc ),
    .resetb(\pll/resetb ),
    .clockp({\pll/clockp [1],
    \pll/clockp [0]}),
    .div({\pll/div [4],
    \pll/div [3],
    \pll/div [2],
    \pll/div [1],
    \pll/div [0]}),
    .ext_trim({\pll/ext_trim [25],
    \pll/ext_trim [24],
    \pll/ext_trim [23],
    \pll/ext_trim [22],
    \pll/ext_trim [21],
    \pll/ext_trim [20],
    \pll/ext_trim [19],
    \pll/ext_trim [18],
    \pll/ext_trim [17],
    \pll/ext_trim [16],
    \pll/ext_trim [15],
    \pll/ext_trim [14],
    \pll/ext_trim [13],
    \pll/ext_trim [12],
    \pll/ext_trim [11],
    \pll/ext_trim [10],
    \pll/ext_trim [9],
    \pll/ext_trim [8],
    \pll/ext_trim [7],
    \pll/ext_trim [6],
    \pll/ext_trim [5],
    \pll/ext_trim [4],
    \pll/ext_trim [3],
    \pll/ext_trim [2],
    \pll/ext_trim [1],
    \pll/ext_trim [0]}));
 housekeeping housekeeping (.debug_in(\soc/debug_in ),
    .debug_mode(\soc/debug_mode ),
    .debug_oeb(\soc/debug_oeb ),
    .debug_out(\soc/debug_out ),
    .pad_flash_clk(\padframe/flash_clk_core ),
    .pad_flash_clk_oeb(\padframe/flash_clk_oeb_core ),
    .pad_flash_csb(\padframe/flash_csb_core ),
    .pad_flash_csb_oeb(\padframe/flash_csb_oeb_core ),
    .pad_flash_io0_di(\padframe/flash_io0_di_core ),
    .pad_flash_io0_do(\padframe/flash_io0_do_core ),
    .pad_flash_io0_ieb(\padframe/flash_io0_ieb_core ),
    .pad_flash_io0_oeb(\padframe/flash_io0_oeb_core ),
    .pad_flash_io1_di(\padframe/flash_io1_di_core ),
    .pad_flash_io1_do(\padframe/flash_io1_do_core ),
    .pad_flash_io1_ieb(\padframe/flash_io1_ieb_core ),
    .pad_flash_io1_oeb(\padframe/flash_io1_oeb_core ),
    .pll_bypass(\clocking/ext_clk_sel ),
    .pll_dco_ena(\pll/dco ),
    .pll_ena(\pll/enable ),
    .porb(\por/porb_l ),
    .qspi_enabled(\soc/qspi_enabled ),
    .reset(\housekeeping/reset ),
    .ser_rx(\soc/ser_rx ),
    .ser_tx(\soc/ser_tx ),
    .serial_clock(\housekeeping/serial_clock ),
    .serial_data_1(\housekeeping/serial_data_1 ),
    .serial_data_2(\housekeeping/serial_data_2 ),
    .serial_load(\housekeeping/serial_load ),
    .serial_resetn(\housekeeping/serial_resetn ),
    .spi_csb(\soc/spi_csb ),
    .spi_enabled(\soc/spi_enabled ),
    .spi_sck(\soc/spi_sck ),
    .spi_sdi(\soc/spi_sdi ),
    .spi_sdo(\soc/spi_sdo ),
    .spi_sdoenb(\soc/spi_sdoenb ),
    .spimemio_flash_clk(\soc/flash_clk ),
    .spimemio_flash_csb(\soc/flash_csb ),
    .spimemio_flash_io0_di(\soc/flash_io0_di ),
    .spimemio_flash_io0_do(\soc/flash_io0_do ),
    .spimemio_flash_io0_oeb(\soc/flash_io0_oeb ),
    .spimemio_flash_io1_di(\soc/flash_io1_di ),
    .spimemio_flash_io1_do(\soc/flash_io1_do ),
    .spimemio_flash_io1_oeb(\soc/flash_io1_oeb ),
    .spimemio_flash_io2_di(\soc/flash_io2_di ),
    .spimemio_flash_io2_do(\soc/flash_io2_do ),
    .spimemio_flash_io2_oeb(\soc/flash_io2_oeb ),
    .spimemio_flash_io3_di(\soc/flash_io3_di ),
    .spimemio_flash_io3_do(\soc/flash_io3_do ),
    .spimemio_flash_io3_oeb(\soc/flash_io3_oeb ),
    .sram_ro_clk(\soc/sram_ro_clk ),
    .sram_ro_csb(\soc/sram_ro_csb ),
    .trap(\soc/trap ),
    .uart_enabled(\soc/uart_enabled ),
    .user_clock(\clocking/user_clk ),
    .usr1_vcc_pwrgood(\housekeeping/usr1_vcc_pwrgood ),
    .usr1_vdd_pwrgood(\housekeeping/usr1_vdd_pwrgood ),
    .usr2_vcc_pwrgood(\housekeeping/usr2_vcc_pwrgood ),
    .usr2_vdd_pwrgood(\housekeeping/usr2_vdd_pwrgood ),
    .wb_ack_o(\soc/hk_ack_i ),
    .wb_clk_i(\soc/core_clk ),
    .wb_cyc_i(\soc/hk_cyc_o ),
    .wb_rstn_i(\soc/core_rstn ),
    .wb_stb_i(\soc/hk_stb_o ),
    .wb_we_i(\soc/mprj_we_o ),
    .irq({\soc/irq [5],
    \soc/irq [4],
    \soc/irq [3]}),
    .mask_rev_in({\user_id_value/mask_rev [31],
    \user_id_value/mask_rev [30],
    \user_id_value/mask_rev [29],
    \user_id_value/mask_rev [28],
    \user_id_value/mask_rev [27],
    \user_id_value/mask_rev [26],
    \user_id_value/mask_rev [25],
    \user_id_value/mask_rev [24],
    \user_id_value/mask_rev [23],
    \user_id_value/mask_rev [22],
    \user_id_value/mask_rev [21],
    \user_id_value/mask_rev [20],
    \user_id_value/mask_rev [19],
    \user_id_value/mask_rev [18],
    \user_id_value/mask_rev [17],
    \user_id_value/mask_rev [16],
    \user_id_value/mask_rev [15],
    \user_id_value/mask_rev [14],
    \user_id_value/mask_rev [13],
    \user_id_value/mask_rev [12],
    \user_id_value/mask_rev [11],
    \user_id_value/mask_rev [10],
    \user_id_value/mask_rev [9],
    \user_id_value/mask_rev [8],
    \user_id_value/mask_rev [7],
    \user_id_value/mask_rev [6],
    \user_id_value/mask_rev [5],
    \user_id_value/mask_rev [4],
    \user_id_value/mask_rev [3],
    \user_id_value/mask_rev [2],
    \user_id_value/mask_rev [1],
    \user_id_value/mask_rev [0]}),
    .mgmt_gpio_in({\housekeeping/mgmt_gpio_in [37],
    \housekeeping/mgmt_gpio_in [36],
    \housekeeping/mgmt_gpio_in [35],
    \housekeeping/mgmt_gpio_in [34],
    \housekeeping/mgmt_gpio_in [33],
    \housekeeping/mgmt_gpio_in [32],
    \housekeeping/mgmt_gpio_in [31],
    \housekeeping/mgmt_gpio_in [30],
    \housekeeping/mgmt_gpio_in [29],
    \housekeeping/mgmt_gpio_in [28],
    \housekeeping/mgmt_gpio_in [27],
    \housekeeping/mgmt_gpio_in [26],
    \housekeeping/mgmt_gpio_in [25],
    \housekeeping/mgmt_gpio_in [24],
    \housekeeping/mgmt_gpio_in [23],
    \housekeeping/mgmt_gpio_in [22],
    \housekeeping/mgmt_gpio_in [21],
    \housekeeping/mgmt_gpio_in [20],
    \housekeeping/mgmt_gpio_in [19],
    \housekeeping/mgmt_gpio_in [18],
    \housekeeping/mgmt_gpio_in [17],
    \housekeeping/mgmt_gpio_in [16],
    \housekeeping/mgmt_gpio_in [15],
    \housekeeping/mgmt_gpio_in [14],
    \housekeeping/mgmt_gpio_in [13],
    \housekeeping/mgmt_gpio_in [12],
    \housekeeping/mgmt_gpio_in [11],
    \housekeeping/mgmt_gpio_in [10],
    \housekeeping/mgmt_gpio_in [9],
    \housekeeping/mgmt_gpio_in [8],
    \housekeeping/mgmt_gpio_in [7],
    \housekeeping/mgmt_gpio_in [6],
    \housekeeping/mgmt_gpio_in [5],
    \housekeeping/mgmt_gpio_in [4],
    \housekeeping/mgmt_gpio_in [3],
    \housekeeping/mgmt_gpio_in [2],
    \housekeeping/mgmt_gpio_in [1],
    \housekeeping/mgmt_gpio_in [0]}),
    .mgmt_gpio_oeb({\housekeeping/mgmt_gpio_oeb [37],
    \housekeeping/mgmt_gpio_oeb [36],
    \housekeeping/mgmt_gpio_oeb [35],
    \housekeeping/mgmt_gpio_oeb [34],
    \housekeeping/mgmt_gpio_oeb [33],
    \housekeeping/mgmt_gpio_oeb [32],
    \housekeeping/mgmt_gpio_oeb [31],
    \housekeeping/mgmt_gpio_oeb [30],
    \housekeeping/mgmt_gpio_oeb [29],
    \housekeeping/mgmt_gpio_oeb [28],
    \housekeeping/mgmt_gpio_oeb [27],
    \housekeeping/mgmt_gpio_oeb [26],
    \housekeeping/mgmt_gpio_oeb [25],
    \housekeeping/mgmt_gpio_oeb [24],
    \housekeeping/mgmt_gpio_oeb [23],
    \housekeeping/mgmt_gpio_oeb [22],
    \housekeeping/mgmt_gpio_oeb [21],
    \housekeeping/mgmt_gpio_oeb [20],
    \housekeeping/mgmt_gpio_oeb [19],
    \housekeeping/mgmt_gpio_oeb [18],
    \housekeeping/mgmt_gpio_oeb [17],
    \housekeeping/mgmt_gpio_oeb [16],
    \housekeeping/mgmt_gpio_oeb [15],
    \housekeeping/mgmt_gpio_oeb [14],
    \housekeeping/mgmt_gpio_oeb [13],
    \housekeeping/mgmt_gpio_oeb [12],
    \housekeeping/mgmt_gpio_oeb [11],
    \housekeeping/mgmt_gpio_oeb [10],
    \housekeeping/mgmt_gpio_oeb [9],
    \housekeeping/mgmt_gpio_oeb [8],
    \housekeeping/mgmt_gpio_oeb [7],
    \housekeeping/mgmt_gpio_oeb [6],
    \housekeeping/mgmt_gpio_oeb [5],
    \housekeeping/mgmt_gpio_oeb [4],
    \housekeeping/mgmt_gpio_oeb [3],
    \housekeeping/mgmt_gpio_oeb [2],
    \housekeeping/mgmt_gpio_oeb [1],
    \housekeeping/mgmt_gpio_oeb [0]}),
    .mgmt_gpio_out({\housekeeping/mgmt_gpio_out [37],
    \housekeeping/mgmt_gpio_out [36],
    \housekeeping/mgmt_gpio_out [35],
    \housekeeping/mgmt_gpio_in [34],
    \housekeeping/mgmt_gpio_in [33],
    \housekeeping/mgmt_gpio_in [32],
    \housekeeping/mgmt_gpio_in [31],
    \housekeeping/mgmt_gpio_in [30],
    \housekeeping/mgmt_gpio_in [29],
    \housekeeping/mgmt_gpio_in [28],
    \housekeeping/mgmt_gpio_in [27],
    \housekeeping/mgmt_gpio_in [26],
    \housekeeping/mgmt_gpio_in [25],
    \housekeeping/mgmt_gpio_in [24],
    \housekeeping/mgmt_gpio_in [23],
    \housekeeping/mgmt_gpio_in [22],
    \housekeeping/mgmt_gpio_in [21],
    \housekeeping/mgmt_gpio_in [20],
    \housekeeping/mgmt_gpio_in [19],
    \housekeeping/mgmt_gpio_in [18],
    \housekeeping/mgmt_gpio_in [17],
    \housekeeping/mgmt_gpio_in [16],
    \housekeeping/mgmt_gpio_in [15],
    \housekeeping/mgmt_gpio_in [14],
    \housekeeping/mgmt_gpio_in [13],
    \housekeeping/mgmt_gpio_in [12],
    \housekeeping/mgmt_gpio_in [11],
    \housekeeping/mgmt_gpio_in [10],
    \housekeeping/mgmt_gpio_in [9],
    \housekeeping/mgmt_gpio_in [8],
    \housekeeping/mgmt_gpio_in [7],
    \housekeeping/mgmt_gpio_in [6],
    \housekeeping/mgmt_gpio_in [5],
    \housekeeping/mgmt_gpio_in [4],
    \housekeeping/mgmt_gpio_in [3],
    \housekeeping/mgmt_gpio_in [2],
    \housekeeping/mgmt_gpio_out [1],
    \housekeeping/mgmt_gpio_out [0]}),
    .pll90_sel({\clocking/sel2 [2],
    \clocking/sel2 [1],
    \clocking/sel2 [0]}),
    .pll_div({\pll/div [4],
    \pll/div [3],
    \pll/div [2],
    \pll/div [1],
    \pll/div [0]}),
    .pll_sel({\clocking/sel [2],
    \clocking/sel [1],
    \clocking/sel [0]}),
    .pll_trim({\pll/ext_trim [25],
    \pll/ext_trim [24],
    \pll/ext_trim [23],
    \pll/ext_trim [22],
    \pll/ext_trim [21],
    \pll/ext_trim [20],
    \pll/ext_trim [19],
    \pll/ext_trim [18],
    \pll/ext_trim [17],
    \pll/ext_trim [16],
    \pll/ext_trim [15],
    \pll/ext_trim [14],
    \pll/ext_trim [13],
    \pll/ext_trim [12],
    \pll/ext_trim [11],
    \pll/ext_trim [10],
    \pll/ext_trim [9],
    \pll/ext_trim [8],
    \pll/ext_trim [7],
    \pll/ext_trim [6],
    \pll/ext_trim [5],
    \pll/ext_trim [4],
    \pll/ext_trim [3],
    \pll/ext_trim [2],
    \pll/ext_trim [1],
    \pll/ext_trim [0]}),
    .pwr_ctrl_out({\housekeeping/pwr_ctrl_out [3],
    \housekeeping/pwr_ctrl_out [2],
    \housekeeping/pwr_ctrl_out [1],
    \housekeeping/pwr_ctrl_out [0]}),
    .sram_ro_addr({\soc/sram_ro_addr [7],
    \soc/sram_ro_addr [6],
    \soc/sram_ro_addr [5],
    \soc/sram_ro_addr [4],
    \soc/sram_ro_addr [3],
    \soc/sram_ro_addr [2],
    \soc/sram_ro_addr [1],
    \soc/sram_ro_addr [0]}),
    .sram_ro_data({\soc/sram_ro_data [31],
    \soc/sram_ro_data [30],
    \soc/sram_ro_data [29],
    \soc/sram_ro_data [28],
    \soc/sram_ro_data [27],
    \soc/sram_ro_data [26],
    \soc/sram_ro_data [25],
    \soc/sram_ro_data [24],
    \soc/sram_ro_data [23],
    \soc/sram_ro_data [22],
    \soc/sram_ro_data [21],
    \soc/sram_ro_data [20],
    \soc/sram_ro_data [19],
    \soc/sram_ro_data [18],
    \soc/sram_ro_data [17],
    \soc/sram_ro_data [16],
    \soc/sram_ro_data [15],
    \soc/sram_ro_data [14],
    \soc/sram_ro_data [13],
    \soc/sram_ro_data [12],
    \soc/sram_ro_data [11],
    \soc/sram_ro_data [10],
    \soc/sram_ro_data [9],
    \soc/sram_ro_data [8],
    \soc/sram_ro_data [7],
    \soc/sram_ro_data [6],
    \soc/sram_ro_data [5],
    \soc/sram_ro_data [4],
    \soc/sram_ro_data [3],
    \soc/sram_ro_data [2],
    \soc/sram_ro_data [1],
    \soc/sram_ro_data [0]}),
    .wb_adr_i({\soc/mprj_adr_o [31],
    \soc/mprj_adr_o [30],
    \soc/mprj_adr_o [29],
    \soc/mprj_adr_o [28],
    \soc/mprj_adr_o [27],
    \soc/mprj_adr_o [26],
    \soc/mprj_adr_o [25],
    \soc/mprj_adr_o [24],
    \soc/mprj_adr_o [23],
    \soc/mprj_adr_o [22],
    \soc/mprj_adr_o [21],
    \soc/mprj_adr_o [20],
    \soc/mprj_adr_o [19],
    \soc/mprj_adr_o [18],
    \soc/mprj_adr_o [17],
    \soc/mprj_adr_o [16],
    \soc/mprj_adr_o [15],
    \soc/mprj_adr_o [14],
    \soc/mprj_adr_o [13],
    \soc/mprj_adr_o [12],
    \soc/mprj_adr_o [11],
    \soc/mprj_adr_o [10],
    \soc/mprj_adr_o [9],
    \soc/mprj_adr_o [8],
    \soc/mprj_adr_o [7],
    \soc/mprj_adr_o [6],
    \soc/mprj_adr_o [5],
    \soc/mprj_adr_o [4],
    \soc/mprj_adr_o [3],
    \soc/mprj_adr_o [2],
    \soc/mprj_adr_o [1],
    \soc/mprj_adr_o [0]}),
    .wb_dat_i({\soc/mprj_dat_o [31],
    \soc/mprj_dat_o [30],
    \soc/mprj_dat_o [29],
    \soc/mprj_dat_o [28],
    \soc/mprj_dat_o [27],
    \soc/mprj_dat_o [26],
    \soc/mprj_dat_o [25],
    \soc/mprj_dat_o [24],
    \soc/mprj_dat_o [23],
    \soc/mprj_dat_o [22],
    \soc/mprj_dat_o [21],
    \soc/mprj_dat_o [20],
    \soc/mprj_dat_o [19],
    \soc/mprj_dat_o [18],
    \soc/mprj_dat_o [17],
    \soc/mprj_dat_o [16],
    \soc/mprj_dat_o [15],
    \soc/mprj_dat_o [14],
    \soc/mprj_dat_o [13],
    \soc/mprj_dat_o [12],
    \soc/mprj_dat_o [11],
    \soc/mprj_dat_o [10],
    \soc/mprj_dat_o [9],
    \soc/mprj_dat_o [8],
    \soc/mprj_dat_o [7],
    \soc/mprj_dat_o [6],
    \soc/mprj_dat_o [5],
    \soc/mprj_dat_o [4],
    \soc/mprj_dat_o [3],
    \soc/mprj_dat_o [2],
    \soc/mprj_dat_o [1],
    \soc/mprj_dat_o [0]}),
    .wb_dat_o({\soc/hk_dat_i [31],
    \soc/hk_dat_i [30],
    \soc/hk_dat_i [29],
    \soc/hk_dat_i [28],
    \soc/hk_dat_i [27],
    \soc/hk_dat_i [26],
    \soc/hk_dat_i [25],
    \soc/hk_dat_i [24],
    \soc/hk_dat_i [23],
    \soc/hk_dat_i [22],
    \soc/hk_dat_i [21],
    \soc/hk_dat_i [20],
    \soc/hk_dat_i [19],
    \soc/hk_dat_i [18],
    \soc/hk_dat_i [17],
    \soc/hk_dat_i [16],
    \soc/hk_dat_i [15],
    \soc/hk_dat_i [14],
    \soc/hk_dat_i [13],
    \soc/hk_dat_i [12],
    \soc/hk_dat_i [11],
    \soc/hk_dat_i [10],
    \soc/hk_dat_i [9],
    \soc/hk_dat_i [8],
    \soc/hk_dat_i [7],
    \soc/hk_dat_i [6],
    \soc/hk_dat_i [5],
    \soc/hk_dat_i [4],
    \soc/hk_dat_i [3],
    \soc/hk_dat_i [2],
    \soc/hk_dat_i [1],
    \soc/hk_dat_i [0]}),
    .wb_sel_i({\soc/mprj_sel_o [3],
    \soc/mprj_sel_o [2],
    \soc/mprj_sel_o [1],
    \soc/mprj_sel_o [0]}));
 caravel_clocking clocking (.core_clk(\soc/core_clk ),
    .ext_clk(\pll/osc ),
    .ext_clk_sel(\clocking/ext_clk_sel ),
    .ext_reset(\housekeeping/reset ),
    .pll_clk(\pll/clockp [1]),
    .pll_clk90(\pll/clockp [0]),
    .resetb(\pll/resetb ),
    .resetb_sync(\soc/core_rstn ),
    .user_clk(\clocking/user_clk ),
    .sel({\clocking/sel [2],
    \clocking/sel [1],
    \clocking/sel [0]}),
    .sel2({\clocking/sel2 [2],
    \clocking/sel2 [1],
    \clocking/sel2 [0]}));
 mgmt_core_wrapper soc (.core_clk(\soc/core_clk ),
    .core_rstn(\soc/core_rstn ),
    .debug_in(\soc/debug_in ),
    .debug_mode(\soc/debug_mode ),
    .debug_oeb(\soc/debug_oeb ),
    .debug_out(\soc/debug_out ),
    .flash_clk(\soc/flash_clk ),
    .flash_csb(\soc/flash_csb ),
    .flash_io0_di(\soc/flash_io0_di ),
    .flash_io0_do(\soc/flash_io0_do ),
    .flash_io0_oeb(\soc/flash_io0_oeb ),
    .flash_io1_di(\soc/flash_io1_di ),
    .flash_io1_do(\soc/flash_io1_do ),
    .flash_io1_oeb(\soc/flash_io1_oeb ),
    .flash_io2_di(\soc/flash_io2_di ),
    .flash_io2_do(\soc/flash_io2_do ),
    .flash_io2_oeb(\soc/flash_io2_oeb ),
    .flash_io3_di(\soc/flash_io3_di ),
    .flash_io3_do(\soc/flash_io3_do ),
    .flash_io3_oeb(\soc/flash_io3_oeb ),
    .gpio_in_pad(\soc/gpio_in_pad ),
    .gpio_inenb_pad(\soc/gpio_inenb_pad ),
    .gpio_mode0_pad(\soc/gpio_mode0_pad ),
    .gpio_mode1_pad(\soc/gpio_mode1_pad ),
    .gpio_out_pad(\soc/gpio_out_pad ),
    .gpio_outenb_pad(\soc/gpio_outenb_pad ),
    .hk_ack_i(\soc/hk_ack_i ),
    .hk_cyc_o(\soc/hk_cyc_o ),
    .hk_stb_o(\soc/hk_stb_o ),
    .mprj_ack_i(\soc/mprj_ack_i ),
    .mprj_cyc_o(\soc/mprj_cyc_o ),
    .mprj_stb_o(\soc/mprj_stb_o ),
    .mprj_wb_iena(\soc/mprj_wb_iena ),
    .mprj_we_o(\soc/mprj_we_o ),
    .qspi_enabled(\soc/qspi_enabled ),
    .ser_rx(\soc/ser_rx ),
    .ser_tx(\soc/ser_tx ),
    .spi_csb(\soc/spi_csb ),
    .spi_enabled(\soc/spi_enabled ),
    .spi_sck(\soc/spi_sck ),
    .spi_sdi(\soc/spi_sdi ),
    .spi_sdo(\soc/spi_sdo ),
    .spi_sdoenb(\soc/spi_sdoenb ),
    .sram_ro_clk(\soc/sram_ro_clk ),
    .sram_ro_csb(\soc/sram_ro_csb ),
    .trap(\soc/trap ),
    .uart_enabled(\soc/uart_enabled ),
    .hk_dat_i({\soc/hk_dat_i [31],
    \soc/hk_dat_i [30],
    \soc/hk_dat_i [29],
    \soc/hk_dat_i [28],
    \soc/hk_dat_i [27],
    \soc/hk_dat_i [26],
    \soc/hk_dat_i [25],
    \soc/hk_dat_i [24],
    \soc/hk_dat_i [23],
    \soc/hk_dat_i [22],
    \soc/hk_dat_i [21],
    \soc/hk_dat_i [20],
    \soc/hk_dat_i [19],
    \soc/hk_dat_i [18],
    \soc/hk_dat_i [17],
    \soc/hk_dat_i [16],
    \soc/hk_dat_i [15],
    \soc/hk_dat_i [14],
    \soc/hk_dat_i [13],
    \soc/hk_dat_i [12],
    \soc/hk_dat_i [11],
    \soc/hk_dat_i [10],
    \soc/hk_dat_i [9],
    \soc/hk_dat_i [8],
    \soc/hk_dat_i [7],
    \soc/hk_dat_i [6],
    \soc/hk_dat_i [5],
    \soc/hk_dat_i [4],
    \soc/hk_dat_i [3],
    \soc/hk_dat_i [2],
    \soc/hk_dat_i [1],
    \soc/hk_dat_i [0]}),
    .irq({\soc/irq [5],
    \soc/irq [4],
    \soc/irq [3],
    \soc/irq [2],
    \soc/irq [1],
    \soc/irq [0]}),
    .la_iena({\soc/la_iena [127],
    \soc/la_iena [126],
    \soc/la_iena [125],
    \soc/la_iena [124],
    \soc/la_iena [123],
    \soc/la_iena [122],
    \soc/la_iena [121],
    \soc/la_iena [120],
    \soc/la_iena [119],
    \soc/la_iena [118],
    \soc/la_iena [117],
    \soc/la_iena [116],
    \soc/la_iena [115],
    \soc/la_iena [114],
    \soc/la_iena [113],
    \soc/la_iena [112],
    \soc/la_iena [111],
    \soc/la_iena [110],
    \soc/la_iena [109],
    \soc/la_iena [108],
    \soc/la_iena [107],
    \soc/la_iena [106],
    \soc/la_iena [105],
    \soc/la_iena [104],
    \soc/la_iena [103],
    \soc/la_iena [102],
    \soc/la_iena [101],
    \soc/la_iena [100],
    \soc/la_iena [99],
    \soc/la_iena [98],
    \soc/la_iena [97],
    \soc/la_iena [96],
    \soc/la_iena [95],
    \soc/la_iena [94],
    \soc/la_iena [93],
    \soc/la_iena [92],
    \soc/la_iena [91],
    \soc/la_iena [90],
    \soc/la_iena [89],
    \soc/la_iena [88],
    \soc/la_iena [87],
    \soc/la_iena [86],
    \soc/la_iena [85],
    \soc/la_iena [84],
    \soc/la_iena [83],
    \soc/la_iena [82],
    \soc/la_iena [81],
    \soc/la_iena [80],
    \soc/la_iena [79],
    \soc/la_iena [78],
    \soc/la_iena [77],
    \soc/la_iena [76],
    \soc/la_iena [75],
    \soc/la_iena [74],
    \soc/la_iena [73],
    \soc/la_iena [72],
    \soc/la_iena [71],
    \soc/la_iena [70],
    \soc/la_iena [69],
    \soc/la_iena [68],
    \soc/la_iena [67],
    \soc/la_iena [66],
    \soc/la_iena [65],
    \soc/la_iena [64],
    \soc/la_iena [63],
    \soc/la_iena [62],
    \soc/la_iena [61],
    \soc/la_iena [60],
    \soc/la_iena [59],
    \soc/la_iena [58],
    \soc/la_iena [57],
    \soc/la_iena [56],
    \soc/la_iena [55],
    \soc/la_iena [54],
    \soc/la_iena [53],
    \soc/la_iena [52],
    \soc/la_iena [51],
    \soc/la_iena [50],
    \soc/la_iena [49],
    \soc/la_iena [48],
    \soc/la_iena [47],
    \soc/la_iena [46],
    \soc/la_iena [45],
    \soc/la_iena [44],
    \soc/la_iena [43],
    \soc/la_iena [42],
    \soc/la_iena [41],
    \soc/la_iena [40],
    \soc/la_iena [39],
    \soc/la_iena [38],
    \soc/la_iena [37],
    \soc/la_iena [36],
    \soc/la_iena [35],
    \soc/la_iena [34],
    \soc/la_iena [33],
    \soc/la_iena [32],
    \soc/la_iena [31],
    \soc/la_iena [30],
    \soc/la_iena [29],
    \soc/la_iena [28],
    \soc/la_iena [27],
    \soc/la_iena [26],
    \soc/la_iena [25],
    \soc/la_iena [24],
    \soc/la_iena [23],
    \soc/la_iena [22],
    \soc/la_iena [21],
    \soc/la_iena [20],
    \soc/la_iena [19],
    \soc/la_iena [18],
    \soc/la_iena [17],
    \soc/la_iena [16],
    \soc/la_iena [15],
    \soc/la_iena [14],
    \soc/la_iena [13],
    \soc/la_iena [12],
    \soc/la_iena [11],
    \soc/la_iena [10],
    \soc/la_iena [9],
    \soc/la_iena [8],
    \soc/la_iena [7],
    \soc/la_iena [6],
    \soc/la_iena [5],
    \soc/la_iena [4],
    \soc/la_iena [3],
    \soc/la_iena [2],
    \soc/la_iena [1],
    \soc/la_iena [0]}),
    .la_input({\soc/la_input [127],
    \soc/la_input [126],
    \soc/la_input [125],
    \soc/la_input [124],
    \soc/la_input [123],
    \soc/la_input [122],
    \soc/la_input [121],
    \soc/la_input [120],
    \soc/la_input [119],
    \soc/la_input [118],
    \soc/la_input [117],
    \soc/la_input [116],
    \soc/la_input [115],
    \soc/la_input [114],
    \soc/la_input [113],
    \soc/la_input [112],
    \soc/la_input [111],
    \soc/la_input [110],
    \soc/la_input [109],
    \soc/la_input [108],
    \soc/la_input [107],
    \soc/la_input [106],
    \soc/la_input [105],
    \soc/la_input [104],
    \soc/la_input [103],
    \soc/la_input [102],
    \soc/la_input [101],
    \soc/la_input [100],
    \soc/la_input [99],
    \soc/la_input [98],
    \soc/la_input [97],
    \soc/la_input [96],
    \soc/la_input [95],
    \soc/la_input [94],
    \soc/la_input [93],
    \soc/la_input [92],
    \soc/la_input [91],
    \soc/la_input [90],
    \soc/la_input [89],
    \soc/la_input [88],
    \soc/la_input [87],
    \soc/la_input [86],
    \soc/la_input [85],
    \soc/la_input [84],
    \soc/la_input [83],
    \soc/la_input [82],
    \soc/la_input [81],
    \soc/la_input [80],
    \soc/la_input [79],
    \soc/la_input [78],
    \soc/la_input [77],
    \soc/la_input [76],
    \soc/la_input [75],
    \soc/la_input [74],
    \soc/la_input [73],
    \soc/la_input [72],
    \soc/la_input [71],
    \soc/la_input [70],
    \soc/la_input [69],
    \soc/la_input [68],
    \soc/la_input [67],
    \soc/la_input [66],
    \soc/la_input [65],
    \soc/la_input [64],
    \soc/la_input [63],
    \soc/la_input [62],
    \soc/la_input [61],
    \soc/la_input [60],
    \soc/la_input [59],
    \soc/la_input [58],
    \soc/la_input [57],
    \soc/la_input [56],
    \soc/la_input [55],
    \soc/la_input [54],
    \soc/la_input [53],
    \soc/la_input [52],
    \soc/la_input [51],
    \soc/la_input [50],
    \soc/la_input [49],
    \soc/la_input [48],
    \soc/la_input [47],
    \soc/la_input [46],
    \soc/la_input [45],
    \soc/la_input [44],
    \soc/la_input [43],
    \soc/la_input [42],
    \soc/la_input [41],
    \soc/la_input [40],
    \soc/la_input [39],
    \soc/la_input [38],
    \soc/la_input [37],
    \soc/la_input [36],
    \soc/la_input [35],
    \soc/la_input [34],
    \soc/la_input [33],
    \soc/la_input [32],
    \soc/la_input [31],
    \soc/la_input [30],
    \soc/la_input [29],
    \soc/la_input [28],
    \soc/la_input [27],
    \soc/la_input [26],
    \soc/la_input [25],
    \soc/la_input [24],
    \soc/la_input [23],
    \soc/la_input [22],
    \soc/la_input [21],
    \soc/la_input [20],
    \soc/la_input [19],
    \soc/la_input [18],
    \soc/la_input [17],
    \soc/la_input [16],
    \soc/la_input [15],
    \soc/la_input [14],
    \soc/la_input [13],
    \soc/la_input [12],
    \soc/la_input [11],
    \soc/la_input [10],
    \soc/la_input [9],
    \soc/la_input [8],
    \soc/la_input [7],
    \soc/la_input [6],
    \soc/la_input [5],
    \soc/la_input [4],
    \soc/la_input [3],
    \soc/la_input [2],
    \soc/la_input [1],
    \soc/la_input [0]}),
    .la_oenb({\soc/la_oenb [127],
    \soc/la_oenb [126],
    \soc/la_oenb [125],
    \soc/la_oenb [124],
    \soc/la_oenb [123],
    \soc/la_oenb [122],
    \soc/la_oenb [121],
    \soc/la_oenb [120],
    \soc/la_oenb [119],
    \soc/la_oenb [118],
    \soc/la_oenb [117],
    \soc/la_oenb [116],
    \soc/la_oenb [115],
    \soc/la_oenb [114],
    \soc/la_oenb [113],
    \soc/la_oenb [112],
    \soc/la_oenb [111],
    \soc/la_oenb [110],
    \soc/la_oenb [109],
    \soc/la_oenb [108],
    \soc/la_oenb [107],
    \soc/la_oenb [106],
    \soc/la_oenb [105],
    \soc/la_oenb [104],
    \soc/la_oenb [103],
    \soc/la_oenb [102],
    \soc/la_oenb [101],
    \soc/la_oenb [100],
    \soc/la_oenb [99],
    \soc/la_oenb [98],
    \soc/la_oenb [97],
    \soc/la_oenb [96],
    \soc/la_oenb [95],
    \soc/la_oenb [94],
    \soc/la_oenb [93],
    \soc/la_oenb [92],
    \soc/la_oenb [91],
    \soc/la_oenb [90],
    \soc/la_oenb [89],
    \soc/la_oenb [88],
    \soc/la_oenb [87],
    \soc/la_oenb [86],
    \soc/la_oenb [85],
    \soc/la_oenb [84],
    \soc/la_oenb [83],
    \soc/la_oenb [82],
    \soc/la_oenb [81],
    \soc/la_oenb [80],
    \soc/la_oenb [79],
    \soc/la_oenb [78],
    \soc/la_oenb [77],
    \soc/la_oenb [76],
    \soc/la_oenb [75],
    \soc/la_oenb [74],
    \soc/la_oenb [73],
    \soc/la_oenb [72],
    \soc/la_oenb [71],
    \soc/la_oenb [70],
    \soc/la_oenb [69],
    \soc/la_oenb [68],
    \soc/la_oenb [67],
    \soc/la_oenb [66],
    \soc/la_oenb [65],
    \soc/la_oenb [64],
    \soc/la_oenb [63],
    \soc/la_oenb [62],
    \soc/la_oenb [61],
    \soc/la_oenb [60],
    \soc/la_oenb [59],
    \soc/la_oenb [58],
    \soc/la_oenb [57],
    \soc/la_oenb [56],
    \soc/la_oenb [55],
    \soc/la_oenb [54],
    \soc/la_oenb [53],
    \soc/la_oenb [52],
    \soc/la_oenb [51],
    \soc/la_oenb [50],
    \soc/la_oenb [49],
    \soc/la_oenb [48],
    \soc/la_oenb [47],
    \soc/la_oenb [46],
    \soc/la_oenb [45],
    \soc/la_oenb [44],
    \soc/la_oenb [43],
    \soc/la_oenb [42],
    \soc/la_oenb [41],
    \soc/la_oenb [40],
    \soc/la_oenb [39],
    \soc/la_oenb [38],
    \soc/la_oenb [37],
    \soc/la_oenb [36],
    \soc/la_oenb [35],
    \soc/la_oenb [34],
    \soc/la_oenb [33],
    \soc/la_oenb [32],
    \soc/la_oenb [31],
    \soc/la_oenb [30],
    \soc/la_oenb [29],
    \soc/la_oenb [28],
    \soc/la_oenb [27],
    \soc/la_oenb [26],
    \soc/la_oenb [25],
    \soc/la_oenb [24],
    \soc/la_oenb [23],
    \soc/la_oenb [22],
    \soc/la_oenb [21],
    \soc/la_oenb [20],
    \soc/la_oenb [19],
    \soc/la_oenb [18],
    \soc/la_oenb [17],
    \soc/la_oenb [16],
    \soc/la_oenb [15],
    \soc/la_oenb [14],
    \soc/la_oenb [13],
    \soc/la_oenb [12],
    \soc/la_oenb [11],
    \soc/la_oenb [10],
    \soc/la_oenb [9],
    \soc/la_oenb [8],
    \soc/la_oenb [7],
    \soc/la_oenb [6],
    \soc/la_oenb [5],
    \soc/la_oenb [4],
    \soc/la_oenb [3],
    \soc/la_oenb [2],
    \soc/la_oenb [1],
    \soc/la_oenb [0]}),
    .la_output({\soc/la_output [127],
    \soc/la_output [126],
    \soc/la_output [125],
    \soc/la_output [124],
    \soc/la_output [123],
    \soc/la_output [122],
    \soc/la_output [121],
    \soc/la_output [120],
    \soc/la_output [119],
    \soc/la_output [118],
    \soc/la_output [117],
    \soc/la_output [116],
    \soc/la_output [115],
    \soc/la_output [114],
    \soc/la_output [113],
    \soc/la_output [112],
    \soc/la_output [111],
    \soc/la_output [110],
    \soc/la_output [109],
    \soc/la_output [108],
    \soc/la_output [107],
    \soc/la_output [106],
    \soc/la_output [105],
    \soc/la_output [104],
    \soc/la_output [103],
    \soc/la_output [102],
    \soc/la_output [101],
    \soc/la_output [100],
    \soc/la_output [99],
    \soc/la_output [98],
    \soc/la_output [97],
    \soc/la_output [96],
    \soc/la_output [95],
    \soc/la_output [94],
    \soc/la_output [93],
    \soc/la_output [92],
    \soc/la_output [91],
    \soc/la_output [90],
    \soc/la_output [89],
    \soc/la_output [88],
    \soc/la_output [87],
    \soc/la_output [86],
    \soc/la_output [85],
    \soc/la_output [84],
    \soc/la_output [83],
    \soc/la_output [82],
    \soc/la_output [81],
    \soc/la_output [80],
    \soc/la_output [79],
    \soc/la_output [78],
    \soc/la_output [77],
    \soc/la_output [76],
    \soc/la_output [75],
    \soc/la_output [74],
    \soc/la_output [73],
    \soc/la_output [72],
    \soc/la_output [71],
    \soc/la_output [70],
    \soc/la_output [69],
    \soc/la_output [68],
    \soc/la_output [67],
    \soc/la_output [66],
    \soc/la_output [65],
    \soc/la_output [64],
    \soc/la_output [63],
    \soc/la_output [62],
    \soc/la_output [61],
    \soc/la_output [60],
    \soc/la_output [59],
    \soc/la_output [58],
    \soc/la_output [57],
    \soc/la_output [56],
    \soc/la_output [55],
    \soc/la_output [54],
    \soc/la_output [53],
    \soc/la_output [52],
    \soc/la_output [51],
    \soc/la_output [50],
    \soc/la_output [49],
    \soc/la_output [48],
    \soc/la_output [47],
    \soc/la_output [46],
    \soc/la_output [45],
    \soc/la_output [44],
    \soc/la_output [43],
    \soc/la_output [42],
    \soc/la_output [41],
    \soc/la_output [40],
    \soc/la_output [39],
    \soc/la_output [38],
    \soc/la_output [37],
    \soc/la_output [36],
    \soc/la_output [35],
    \soc/la_output [34],
    \soc/la_output [33],
    \soc/la_output [32],
    \soc/la_output [31],
    \soc/la_output [30],
    \soc/la_output [29],
    \soc/la_output [28],
    \soc/la_output [27],
    \soc/la_output [26],
    \soc/la_output [25],
    \soc/la_output [24],
    \soc/la_output [23],
    \soc/la_output [22],
    \soc/la_output [21],
    \soc/la_output [20],
    \soc/la_output [19],
    \soc/la_output [18],
    \soc/la_output [17],
    \soc/la_output [16],
    \soc/la_output [15],
    \soc/la_output [14],
    \soc/la_output [13],
    \soc/la_output [12],
    \soc/la_output [11],
    \soc/la_output [10],
    \soc/la_output [9],
    \soc/la_output [8],
    \soc/la_output [7],
    \soc/la_output [6],
    \soc/la_output [5],
    \soc/la_output [4],
    \soc/la_output [3],
    \soc/la_output [2],
    \soc/la_output [1],
    \soc/la_output [0]}),
    .mprj_adr_o({\soc/mprj_adr_o [31],
    \soc/mprj_adr_o [30],
    \soc/mprj_adr_o [29],
    \soc/mprj_adr_o [28],
    \soc/mprj_adr_o [27],
    \soc/mprj_adr_o [26],
    \soc/mprj_adr_o [25],
    \soc/mprj_adr_o [24],
    \soc/mprj_adr_o [23],
    \soc/mprj_adr_o [22],
    \soc/mprj_adr_o [21],
    \soc/mprj_adr_o [20],
    \soc/mprj_adr_o [19],
    \soc/mprj_adr_o [18],
    \soc/mprj_adr_o [17],
    \soc/mprj_adr_o [16],
    \soc/mprj_adr_o [15],
    \soc/mprj_adr_o [14],
    \soc/mprj_adr_o [13],
    \soc/mprj_adr_o [12],
    \soc/mprj_adr_o [11],
    \soc/mprj_adr_o [10],
    \soc/mprj_adr_o [9],
    \soc/mprj_adr_o [8],
    \soc/mprj_adr_o [7],
    \soc/mprj_adr_o [6],
    \soc/mprj_adr_o [5],
    \soc/mprj_adr_o [4],
    \soc/mprj_adr_o [3],
    \soc/mprj_adr_o [2],
    \soc/mprj_adr_o [1],
    \soc/mprj_adr_o [0]}),
    .mprj_dat_i({\soc/mprj_dat_i [31],
    \soc/mprj_dat_i [30],
    \soc/mprj_dat_i [29],
    \soc/mprj_dat_i [28],
    \soc/mprj_dat_i [27],
    \soc/mprj_dat_i [26],
    \soc/mprj_dat_i [25],
    \soc/mprj_dat_i [24],
    \soc/mprj_dat_i [23],
    \soc/mprj_dat_i [22],
    \soc/mprj_dat_i [21],
    \soc/mprj_dat_i [20],
    \soc/mprj_dat_i [19],
    \soc/mprj_dat_i [18],
    \soc/mprj_dat_i [17],
    \soc/mprj_dat_i [16],
    \soc/mprj_dat_i [15],
    \soc/mprj_dat_i [14],
    \soc/mprj_dat_i [13],
    \soc/mprj_dat_i [12],
    \soc/mprj_dat_i [11],
    \soc/mprj_dat_i [10],
    \soc/mprj_dat_i [9],
    \soc/mprj_dat_i [8],
    \soc/mprj_dat_i [7],
    \soc/mprj_dat_i [6],
    \soc/mprj_dat_i [5],
    \soc/mprj_dat_i [4],
    \soc/mprj_dat_i [3],
    \soc/mprj_dat_i [2],
    \soc/mprj_dat_i [1],
    \soc/mprj_dat_i [0]}),
    .mprj_dat_o({\soc/mprj_dat_o [31],
    \soc/mprj_dat_o [30],
    \soc/mprj_dat_o [29],
    \soc/mprj_dat_o [28],
    \soc/mprj_dat_o [27],
    \soc/mprj_dat_o [26],
    \soc/mprj_dat_o [25],
    \soc/mprj_dat_o [24],
    \soc/mprj_dat_o [23],
    \soc/mprj_dat_o [22],
    \soc/mprj_dat_o [21],
    \soc/mprj_dat_o [20],
    \soc/mprj_dat_o [19],
    \soc/mprj_dat_o [18],
    \soc/mprj_dat_o [17],
    \soc/mprj_dat_o [16],
    \soc/mprj_dat_o [15],
    \soc/mprj_dat_o [14],
    \soc/mprj_dat_o [13],
    \soc/mprj_dat_o [12],
    \soc/mprj_dat_o [11],
    \soc/mprj_dat_o [10],
    \soc/mprj_dat_o [9],
    \soc/mprj_dat_o [8],
    \soc/mprj_dat_o [7],
    \soc/mprj_dat_o [6],
    \soc/mprj_dat_o [5],
    \soc/mprj_dat_o [4],
    \soc/mprj_dat_o [3],
    \soc/mprj_dat_o [2],
    \soc/mprj_dat_o [1],
    \soc/mprj_dat_o [0]}),
    .mprj_sel_o({\soc/mprj_sel_o [3],
    \soc/mprj_sel_o [2],
    \soc/mprj_sel_o [1],
    \soc/mprj_sel_o [0]}),
    .sram_ro_addr({\soc/sram_ro_addr [7],
    \soc/sram_ro_addr [6],
    \soc/sram_ro_addr [5],
    \soc/sram_ro_addr [4],
    \soc/sram_ro_addr [3],
    \soc/sram_ro_addr [2],
    \soc/sram_ro_addr [1],
    \soc/sram_ro_addr [0]}),
    .sram_ro_data({\soc/sram_ro_data [31],
    \soc/sram_ro_data [30],
    \soc/sram_ro_data [29],
    \soc/sram_ro_data [28],
    \soc/sram_ro_data [27],
    \soc/sram_ro_data [26],
    \soc/sram_ro_data [25],
    \soc/sram_ro_data [24],
    \soc/sram_ro_data [23],
    \soc/sram_ro_data [22],
    \soc/sram_ro_data [21],
    \soc/sram_ro_data [20],
    \soc/sram_ro_data [19],
    \soc/sram_ro_data [18],
    \soc/sram_ro_data [17],
    \soc/sram_ro_data [16],
    \soc/sram_ro_data [15],
    \soc/sram_ro_data [14],
    \soc/sram_ro_data [13],
    \soc/sram_ro_data [12],
    \soc/sram_ro_data [11],
    \soc/sram_ro_data [10],
    \soc/sram_ro_data [9],
    \soc/sram_ro_data [8],
    \soc/sram_ro_data [7],
    \soc/sram_ro_data [6],
    \soc/sram_ro_data [5],
    \soc/sram_ro_data [4],
    \soc/sram_ro_data [3],
    \soc/sram_ro_data [2],
    \soc/sram_ro_data [1],
    \soc/sram_ro_data [0]}),
    .user_irq_ena({\soc/user_irq_ena [2],
    \soc/user_irq_ena [1],
    \soc/user_irq_ena [0]}));
 gpio_control_block \gpio_control_bidir_2[2]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [37]),
    .mgmt_gpio_oeb(\housekeeping/mgmt_gpio_oeb [37]),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_out [37]),
    .one(\gpio_control_bidir_2[2]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [37]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [37]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [37]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [37]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [37]),
    .pad_gpio_in(\padframe/mprj_io_in [37]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [37]),
    .pad_gpio_out(\padframe/mprj_io_out [37]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [37]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [37]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [37]),
    .resetn(\housekeeping/serial_resetn ),
    .resetn_out(\gpio_control_bidir_2[1]/resetn ),
    .serial_clock(\housekeeping/serial_clock ),
    .serial_clock_out(\gpio_control_bidir_2[1]/serial_clock ),
    .serial_data_in(\housekeeping/serial_data_2 ),
    .serial_data_out(\gpio_control_bidir_2[1]/serial_data_in ),
    .serial_load(\housekeeping/serial_load ),
    .serial_load_out(\gpio_control_bidir_2[1]/serial_load ),
    .user_gpio_in(\mprj/io_in [37]),
    .user_gpio_oeb(\mprj/io_oeb [37]),
    .user_gpio_out(\mprj/io_out [37]),
    .zero(\gpio_control_bidir_2[2]/zero ),
    .gpio_defaults({\gpio_defaults_block_37/gpio_defaults [12],
    \gpio_defaults_block_37/gpio_defaults [11],
    \gpio_defaults_block_37/gpio_defaults [10],
    \gpio_defaults_block_37/gpio_defaults [9],
    \gpio_defaults_block_37/gpio_defaults [8],
    \gpio_defaults_block_37/gpio_defaults [7],
    \gpio_defaults_block_37/gpio_defaults [6],
    \gpio_defaults_block_37/gpio_defaults [5],
    \gpio_defaults_block_37/gpio_defaults [4],
    \gpio_defaults_block_37/gpio_defaults [3],
    \gpio_defaults_block_37/gpio_defaults [2],
    \gpio_defaults_block_37/gpio_defaults [1],
    \gpio_defaults_block_37/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [113],
    \padframe/mprj_io_dm [112],
    \padframe/mprj_io_dm [111]}));
 gpio_defaults_block_1803 gpio_defaults_block_1 (.gpio_defaults({\gpio_defaults_block_1/gpio_defaults [12],
    \gpio_defaults_block_1/gpio_defaults [11],
    \gpio_defaults_block_1/gpio_defaults [10],
    \gpio_defaults_block_1/gpio_defaults [9],
    \gpio_defaults_block_1/gpio_defaults [8],
    \gpio_defaults_block_1/gpio_defaults [7],
    \gpio_defaults_block_1/gpio_defaults [6],
    \gpio_defaults_block_1/gpio_defaults [5],
    \gpio_defaults_block_1/gpio_defaults [4],
    \gpio_defaults_block_1/gpio_defaults [3],
    \gpio_defaults_block_1/gpio_defaults [2],
    \gpio_defaults_block_1/gpio_defaults [1],
    \gpio_defaults_block_1/gpio_defaults [0]}));
 gpio_control_block \gpio_control_bidir_1[1]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [1]),
    .mgmt_gpio_oeb(\housekeeping/mgmt_gpio_oeb [1]),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_out [1]),
    .one(\gpio_control_bidir_1[1]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [1]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [1]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [1]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [1]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [1]),
    .pad_gpio_in(\padframe/mprj_io_in [1]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [1]),
    .pad_gpio_out(\padframe/mprj_io_out [1]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [1]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [1]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [1]),
    .resetn(\gpio_control_bidir_1[1]/resetn ),
    .resetn_out(\gpio_control_in_1a[0]/resetn ),
    .serial_clock(\gpio_control_bidir_1[1]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[0]/serial_clock ),
    .serial_data_in(\gpio_control_bidir_1[1]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[0]/serial_data_in ),
    .serial_load(\gpio_control_bidir_1[1]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[0]/serial_load ),
    .user_gpio_in(\mprj/io_in [1]),
    .user_gpio_oeb(\mprj/io_oeb [1]),
    .user_gpio_out(\mprj/io_out [1]),
    .zero(\gpio_control_bidir_1[1]/zero ),
    .gpio_defaults({\gpio_defaults_block_1/gpio_defaults [12],
    \gpio_defaults_block_1/gpio_defaults [11],
    \gpio_defaults_block_1/gpio_defaults [10],
    \gpio_defaults_block_1/gpio_defaults [9],
    \gpio_defaults_block_1/gpio_defaults [8],
    \gpio_defaults_block_1/gpio_defaults [7],
    \gpio_defaults_block_1/gpio_defaults [6],
    \gpio_defaults_block_1/gpio_defaults [5],
    \gpio_defaults_block_1/gpio_defaults [4],
    \gpio_defaults_block_1/gpio_defaults [3],
    \gpio_defaults_block_1/gpio_defaults [2],
    \gpio_defaults_block_1/gpio_defaults [1],
    \gpio_defaults_block_1/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [5],
    \padframe/mprj_io_dm [4],
    \padframe/mprj_io_dm [3]}));
 gpio_control_block \gpio_control_bidir_2[1]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [36]),
    .mgmt_gpio_oeb(\housekeeping/mgmt_gpio_oeb [36]),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_out [36]),
    .one(\gpio_control_bidir_2[1]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [36]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [36]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [36]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [36]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [36]),
    .pad_gpio_in(\padframe/mprj_io_in [36]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [36]),
    .pad_gpio_out(\padframe/mprj_io_out [36]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [36]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [36]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [36]),
    .resetn(\gpio_control_bidir_2[1]/resetn ),
    .resetn_out(\gpio_control_bidir_2[0]/resetn ),
    .serial_clock(\gpio_control_bidir_2[1]/serial_clock ),
    .serial_clock_out(\gpio_control_bidir_2[0]/serial_clock ),
    .serial_data_in(\gpio_control_bidir_2[1]/serial_data_in ),
    .serial_data_out(\gpio_control_bidir_2[0]/serial_data_in ),
    .serial_load(\gpio_control_bidir_2[1]/serial_load ),
    .serial_load_out(\gpio_control_bidir_2[0]/serial_load ),
    .user_gpio_in(\mprj/io_in [36]),
    .user_gpio_oeb(\mprj/io_oeb [36]),
    .user_gpio_out(\mprj/io_out [36]),
    .zero(\gpio_control_bidir_2[1]/zero ),
    .gpio_defaults({\gpio_defaults_block_36/gpio_defaults [12],
    \gpio_defaults_block_36/gpio_defaults [11],
    \gpio_defaults_block_36/gpio_defaults [10],
    \gpio_defaults_block_36/gpio_defaults [9],
    \gpio_defaults_block_36/gpio_defaults [8],
    \gpio_defaults_block_36/gpio_defaults [7],
    \gpio_defaults_block_36/gpio_defaults [6],
    \gpio_defaults_block_36/gpio_defaults [5],
    \gpio_defaults_block_36/gpio_defaults [4],
    \gpio_defaults_block_36/gpio_defaults [3],
    \gpio_defaults_block_36/gpio_defaults [2],
    \gpio_defaults_block_36/gpio_defaults [1],
    \gpio_defaults_block_36/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [110],
    \padframe/mprj_io_dm [109],
    \padframe/mprj_io_dm [108]}));
 gpio_defaults_block gpio_defaults_block_37 (.gpio_defaults({\gpio_defaults_block_37/gpio_defaults [12],
    \gpio_defaults_block_37/gpio_defaults [11],
    \gpio_defaults_block_37/gpio_defaults [10],
    \gpio_defaults_block_37/gpio_defaults [9],
    \gpio_defaults_block_37/gpio_defaults [8],
    \gpio_defaults_block_37/gpio_defaults [7],
    \gpio_defaults_block_37/gpio_defaults [6],
    \gpio_defaults_block_37/gpio_defaults [5],
    \gpio_defaults_block_37/gpio_defaults [4],
    \gpio_defaults_block_37/gpio_defaults [3],
    \gpio_defaults_block_37/gpio_defaults [2],
    \gpio_defaults_block_37/gpio_defaults [1],
    \gpio_defaults_block_37/gpio_defaults [0]}));
 spare_logic_block spare_logic_block_1 (.spare_xib(\spare_logic_block_1/spare_xib ),
    .spare_xfq({\spare_logic_block_1/spare_xfq [1],
    \spare_logic_block_1/spare_xfq [0]}),
    .spare_xfqn({\spare_logic_block_1/spare_xfqn [1],
    \spare_logic_block_1/spare_xfqn [0]}),
    .spare_xi({\spare_logic_block_1/spare_xi [3],
    \spare_logic_block_1/spare_xi [2],
    \spare_logic_block_1/spare_xi [1],
    \spare_logic_block_1/spare_xi [0]}),
    .spare_xmx({\spare_logic_block_1/spare_xmx [1],
    \spare_logic_block_1/spare_xmx [0]}),
    .spare_xna({\spare_logic_block_1/spare_xna [1],
    \spare_logic_block_1/spare_xna [0]}),
    .spare_xno({\spare_logic_block_1/spare_xno [1],
    \spare_logic_block_1/spare_xno [0]}),
    .spare_xz({\spare_logic_block_1/spare_xz [26],
    \spare_logic_block_1/spare_xz [25],
    \spare_logic_block_1/spare_xz [24],
    \spare_logic_block_1/spare_xz [23],
    \spare_logic_block_1/spare_xz [22],
    \spare_logic_block_1/spare_xz [21],
    \spare_logic_block_1/spare_xz [20],
    \spare_logic_block_1/spare_xz [19],
    \spare_logic_block_1/spare_xz [18],
    \spare_logic_block_1/spare_xz [17],
    \spare_logic_block_1/spare_xz [16],
    \spare_logic_block_1/spare_xz [15],
    \spare_logic_block_1/spare_xz [14],
    \spare_logic_block_1/spare_xz [13],
    \spare_logic_block_1/spare_xz [12],
    \spare_logic_block_1/spare_xz [11],
    \spare_logic_block_1/spare_xz [10],
    \spare_logic_block_1/spare_xz [9],
    \spare_logic_block_1/spare_xz [8],
    \spare_logic_block_1/spare_xz [7],
    \spare_logic_block_1/spare_xz [6],
    \spare_logic_block_1/spare_xz [5],
    \spare_logic_block_1/spare_xz [4],
    \spare_logic_block_1/spare_xz [3],
    \spare_logic_block_1/spare_xz [2],
    \spare_logic_block_1/spare_xz [1],
    \spare_logic_block_1/spare_xz [0]}));
 spare_logic_block spare_logic_block_3 (.spare_xib(\spare_logic_block_3/spare_xib ),
    .spare_xfq({\spare_logic_block_3/spare_xfq [1],
    \spare_logic_block_3/spare_xfq [0]}),
    .spare_xfqn({\spare_logic_block_3/spare_xfqn [1],
    \spare_logic_block_3/spare_xfqn [0]}),
    .spare_xi({\spare_logic_block_3/spare_xi [3],
    \spare_logic_block_3/spare_xi [2],
    \spare_logic_block_3/spare_xi [1],
    \spare_logic_block_3/spare_xi [0]}),
    .spare_xmx({\spare_logic_block_3/spare_xmx [1],
    \spare_logic_block_3/spare_xmx [0]}),
    .spare_xna({\spare_logic_block_3/spare_xna [1],
    \spare_logic_block_3/spare_xna [0]}),
    .spare_xno({\spare_logic_block_3/spare_xno [1],
    \spare_logic_block_3/spare_xno [0]}),
    .spare_xz({\spare_logic_block_3/spare_xz [26],
    \spare_logic_block_3/spare_xz [25],
    \spare_logic_block_3/spare_xz [24],
    \spare_logic_block_3/spare_xz [23],
    \spare_logic_block_3/spare_xz [22],
    \spare_logic_block_3/spare_xz [21],
    \spare_logic_block_3/spare_xz [20],
    \spare_logic_block_3/spare_xz [19],
    \spare_logic_block_3/spare_xz [18],
    \spare_logic_block_3/spare_xz [17],
    \spare_logic_block_3/spare_xz [16],
    \spare_logic_block_3/spare_xz [15],
    \spare_logic_block_3/spare_xz [14],
    \spare_logic_block_3/spare_xz [13],
    \spare_logic_block_3/spare_xz [12],
    \spare_logic_block_3/spare_xz [11],
    \spare_logic_block_3/spare_xz [10],
    \spare_logic_block_3/spare_xz [9],
    \spare_logic_block_3/spare_xz [8],
    \spare_logic_block_3/spare_xz [7],
    \spare_logic_block_3/spare_xz [6],
    \spare_logic_block_3/spare_xz [5],
    \spare_logic_block_3/spare_xz [4],
    \spare_logic_block_3/spare_xz [3],
    \spare_logic_block_3/spare_xz [2],
    \spare_logic_block_3/spare_xz [1],
    \spare_logic_block_3/spare_xz [0]}));
 mgmt_protect mgmt_buffers (.caravel_clk(\soc/core_clk ),
    .caravel_clk2(\clocking/user_clk ),
    .caravel_rstn(\soc/core_rstn ),
    .mprj_ack_i_core(\soc/mprj_ack_i ),
    .mprj_ack_i_user(\mprj/wbs_ack_o ),
    .mprj_cyc_o_core(\soc/mprj_cyc_o ),
    .mprj_cyc_o_user(\mprj/wbs_cyc_i ),
    .mprj_iena_wb(\soc/mprj_wb_iena ),
    .mprj_stb_o_core(\soc/mprj_stb_o ),
    .mprj_stb_o_user(\mprj/wbs_stb_i ),
    .mprj_we_o_core(\soc/mprj_we_o ),
    .mprj_we_o_user(\mprj/wbs_we_i ),
    .user1_vcc_powergood(\housekeeping/usr1_vcc_pwrgood ),
    .user1_vdd_powergood(\housekeeping/usr1_vdd_pwrgood ),
    .user2_vcc_powergood(\housekeeping/usr2_vcc_pwrgood ),
    .user2_vdd_powergood(\housekeeping/usr2_vdd_pwrgood ),
    .user_clock(\mprj/wb_clk_i ),
    .user_clock2(\mprj/user_clock2 ),
    .user_reset(\mprj/wb_rst_i ),
    .la_data_in_core({\mprj/la_data_in [127],
    \mprj/la_data_in [126],
    \mprj/la_data_in [125],
    \mprj/la_data_in [124],
    \mprj/la_data_in [123],
    \mprj/la_data_in [122],
    \mprj/la_data_in [121],
    \mprj/la_data_in [120],
    \mprj/la_data_in [119],
    \mprj/la_data_in [118],
    \mprj/la_data_in [117],
    \mprj/la_data_in [116],
    \mprj/la_data_in [115],
    \mprj/la_data_in [114],
    \mprj/la_data_in [113],
    \mprj/la_data_in [112],
    \mprj/la_data_in [111],
    \mprj/la_data_in [110],
    \mprj/la_data_in [109],
    \mprj/la_data_in [108],
    \mprj/la_data_in [107],
    \mprj/la_data_in [106],
    \mprj/la_data_in [105],
    \mprj/la_data_in [104],
    \mprj/la_data_in [103],
    \mprj/la_data_in [102],
    \mprj/la_data_in [101],
    \mprj/la_data_in [100],
    \mprj/la_data_in [99],
    \mprj/la_data_in [98],
    \mprj/la_data_in [97],
    \mprj/la_data_in [96],
    \mprj/la_data_in [95],
    \mprj/la_data_in [94],
    \mprj/la_data_in [93],
    \mprj/la_data_in [92],
    \mprj/la_data_in [91],
    \mprj/la_data_in [90],
    \mprj/la_data_in [89],
    \mprj/la_data_in [88],
    \mprj/la_data_in [87],
    \mprj/la_data_in [86],
    \mprj/la_data_in [85],
    \mprj/la_data_in [84],
    \mprj/la_data_in [83],
    \mprj/la_data_in [82],
    \mprj/la_data_in [81],
    \mprj/la_data_in [80],
    \mprj/la_data_in [79],
    \mprj/la_data_in [78],
    \mprj/la_data_in [77],
    \mprj/la_data_in [76],
    \mprj/la_data_in [75],
    \mprj/la_data_in [74],
    \mprj/la_data_in [73],
    \mprj/la_data_in [72],
    \mprj/la_data_in [71],
    \mprj/la_data_in [70],
    \mprj/la_data_in [69],
    \mprj/la_data_in [68],
    \mprj/la_data_in [67],
    \mprj/la_data_in [66],
    \mprj/la_data_in [65],
    \mprj/la_data_in [64],
    \mprj/la_data_in [63],
    \mprj/la_data_in [62],
    \mprj/la_data_in [61],
    \mprj/la_data_in [60],
    \mprj/la_data_in [59],
    \mprj/la_data_in [58],
    \mprj/la_data_in [57],
    \mprj/la_data_in [56],
    \mprj/la_data_in [55],
    \mprj/la_data_in [54],
    \mprj/la_data_in [53],
    \mprj/la_data_in [52],
    \mprj/la_data_in [51],
    \mprj/la_data_in [50],
    \mprj/la_data_in [49],
    \mprj/la_data_in [48],
    \mprj/la_data_in [47],
    \mprj/la_data_in [46],
    \mprj/la_data_in [45],
    \mprj/la_data_in [44],
    \mprj/la_data_in [43],
    \mprj/la_data_in [42],
    \mprj/la_data_in [41],
    \mprj/la_data_in [40],
    \mprj/la_data_in [39],
    \mprj/la_data_in [38],
    \mprj/la_data_in [37],
    \mprj/la_data_in [36],
    \mprj/la_data_in [35],
    \mprj/la_data_in [34],
    \mprj/la_data_in [33],
    \mprj/la_data_in [32],
    \mprj/la_data_in [31],
    \mprj/la_data_in [30],
    \mprj/la_data_in [29],
    \mprj/la_data_in [28],
    \mprj/la_data_in [27],
    \mprj/la_data_in [26],
    \mprj/la_data_in [25],
    \mprj/la_data_in [24],
    \mprj/la_data_in [23],
    \mprj/la_data_in [22],
    \mprj/la_data_in [21],
    \mprj/la_data_in [20],
    \mprj/la_data_in [19],
    \mprj/la_data_in [18],
    \mprj/la_data_in [17],
    \mprj/la_data_in [16],
    \mprj/la_data_in [15],
    \mprj/la_data_in [14],
    \mprj/la_data_in [13],
    \mprj/la_data_in [12],
    \mprj/la_data_in [11],
    \mprj/la_data_in [10],
    \mprj/la_data_in [9],
    \mprj/la_data_in [8],
    \mprj/la_data_in [7],
    \mprj/la_data_in [6],
    \mprj/la_data_in [5],
    \mprj/la_data_in [4],
    \mprj/la_data_in [3],
    \mprj/la_data_in [2],
    \mprj/la_data_in [1],
    \mprj/la_data_in [0]}),
    .la_data_in_mprj({\soc/la_input [127],
    \soc/la_input [126],
    \soc/la_input [125],
    \soc/la_input [124],
    \soc/la_input [123],
    \soc/la_input [122],
    \soc/la_input [121],
    \soc/la_input [120],
    \soc/la_input [119],
    \soc/la_input [118],
    \soc/la_input [117],
    \soc/la_input [116],
    \soc/la_input [115],
    \soc/la_input [114],
    \soc/la_input [113],
    \soc/la_input [112],
    \soc/la_input [111],
    \soc/la_input [110],
    \soc/la_input [109],
    \soc/la_input [108],
    \soc/la_input [107],
    \soc/la_input [106],
    \soc/la_input [105],
    \soc/la_input [104],
    \soc/la_input [103],
    \soc/la_input [102],
    \soc/la_input [101],
    \soc/la_input [100],
    \soc/la_input [99],
    \soc/la_input [98],
    \soc/la_input [97],
    \soc/la_input [96],
    \soc/la_input [95],
    \soc/la_input [94],
    \soc/la_input [93],
    \soc/la_input [92],
    \soc/la_input [91],
    \soc/la_input [90],
    \soc/la_input [89],
    \soc/la_input [88],
    \soc/la_input [87],
    \soc/la_input [86],
    \soc/la_input [85],
    \soc/la_input [84],
    \soc/la_input [83],
    \soc/la_input [82],
    \soc/la_input [81],
    \soc/la_input [80],
    \soc/la_input [79],
    \soc/la_input [78],
    \soc/la_input [77],
    \soc/la_input [76],
    \soc/la_input [75],
    \soc/la_input [74],
    \soc/la_input [73],
    \soc/la_input [72],
    \soc/la_input [71],
    \soc/la_input [70],
    \soc/la_input [69],
    \soc/la_input [68],
    \soc/la_input [67],
    \soc/la_input [66],
    \soc/la_input [65],
    \soc/la_input [64],
    \soc/la_input [63],
    \soc/la_input [62],
    \soc/la_input [61],
    \soc/la_input [60],
    \soc/la_input [59],
    \soc/la_input [58],
    \soc/la_input [57],
    \soc/la_input [56],
    \soc/la_input [55],
    \soc/la_input [54],
    \soc/la_input [53],
    \soc/la_input [52],
    \soc/la_input [51],
    \soc/la_input [50],
    \soc/la_input [49],
    \soc/la_input [48],
    \soc/la_input [47],
    \soc/la_input [46],
    \soc/la_input [45],
    \soc/la_input [44],
    \soc/la_input [43],
    \soc/la_input [42],
    \soc/la_input [41],
    \soc/la_input [40],
    \soc/la_input [39],
    \soc/la_input [38],
    \soc/la_input [37],
    \soc/la_input [36],
    \soc/la_input [35],
    \soc/la_input [34],
    \soc/la_input [33],
    \soc/la_input [32],
    \soc/la_input [31],
    \soc/la_input [30],
    \soc/la_input [29],
    \soc/la_input [28],
    \soc/la_input [27],
    \soc/la_input [26],
    \soc/la_input [25],
    \soc/la_input [24],
    \soc/la_input [23],
    \soc/la_input [22],
    \soc/la_input [21],
    \soc/la_input [20],
    \soc/la_input [19],
    \soc/la_input [18],
    \soc/la_input [17],
    \soc/la_input [16],
    \soc/la_input [15],
    \soc/la_input [14],
    \soc/la_input [13],
    \soc/la_input [12],
    \soc/la_input [11],
    \soc/la_input [10],
    \soc/la_input [9],
    \soc/la_input [8],
    \soc/la_input [7],
    \soc/la_input [6],
    \soc/la_input [5],
    \soc/la_input [4],
    \soc/la_input [3],
    \soc/la_input [2],
    \soc/la_input [1],
    \soc/la_input [0]}),
    .la_data_out_core({\mprj/la_data_out [127],
    \mprj/la_data_out [126],
    \mprj/la_data_out [125],
    \mprj/la_data_out [124],
    \mprj/la_data_out [123],
    \mprj/la_data_out [122],
    \mprj/la_data_out [121],
    \mprj/la_data_out [120],
    \mprj/la_data_out [119],
    \mprj/la_data_out [118],
    \mprj/la_data_out [117],
    \mprj/la_data_out [116],
    \mprj/la_data_out [115],
    \mprj/la_data_out [114],
    \mprj/la_data_out [113],
    \mprj/la_data_out [112],
    \mprj/la_data_out [111],
    \mprj/la_data_out [110],
    \mprj/la_data_out [109],
    \mprj/la_data_out [108],
    \mprj/la_data_out [107],
    \mprj/la_data_out [106],
    \mprj/la_data_out [105],
    \mprj/la_data_out [104],
    \mprj/la_data_out [103],
    \mprj/la_data_out [102],
    \mprj/la_data_out [101],
    \mprj/la_data_out [100],
    \mprj/la_data_out [99],
    \mprj/la_data_out [98],
    \mprj/la_data_out [97],
    \mprj/la_data_out [96],
    \mprj/la_data_out [95],
    \mprj/la_data_out [94],
    \mprj/la_data_out [93],
    \mprj/la_data_out [92],
    \mprj/la_data_out [91],
    \mprj/la_data_out [90],
    \mprj/la_data_out [89],
    \mprj/la_data_out [88],
    \mprj/la_data_out [87],
    \mprj/la_data_out [86],
    \mprj/la_data_out [85],
    \mprj/la_data_out [84],
    \mprj/la_data_out [83],
    \mprj/la_data_out [82],
    \mprj/la_data_out [81],
    \mprj/la_data_out [80],
    \mprj/la_data_out [79],
    \mprj/la_data_out [78],
    \mprj/la_data_out [77],
    \mprj/la_data_out [76],
    \mprj/la_data_out [75],
    \mprj/la_data_out [74],
    \mprj/la_data_out [73],
    \mprj/la_data_out [72],
    \mprj/la_data_out [71],
    \mprj/la_data_out [70],
    \mprj/la_data_out [69],
    \mprj/la_data_out [68],
    \mprj/la_data_out [67],
    \mprj/la_data_out [66],
    \mprj/la_data_out [65],
    \mprj/la_data_out [64],
    \mprj/la_data_out [63],
    \mprj/la_data_out [62],
    \mprj/la_data_out [61],
    \mprj/la_data_out [60],
    \mprj/la_data_out [59],
    \mprj/la_data_out [58],
    \mprj/la_data_out [57],
    \mprj/la_data_out [56],
    \mprj/la_data_out [55],
    \mprj/la_data_out [54],
    \mprj/la_data_out [53],
    \mprj/la_data_out [52],
    \mprj/la_data_out [51],
    \mprj/la_data_out [50],
    \mprj/la_data_out [49],
    \mprj/la_data_out [48],
    \mprj/la_data_out [47],
    \mprj/la_data_out [46],
    \mprj/la_data_out [45],
    \mprj/la_data_out [44],
    \mprj/la_data_out [43],
    \mprj/la_data_out [42],
    \mprj/la_data_out [41],
    \mprj/la_data_out [40],
    \mprj/la_data_out [39],
    \mprj/la_data_out [38],
    \mprj/la_data_out [37],
    \mprj/la_data_out [36],
    \mprj/la_data_out [35],
    \mprj/la_data_out [34],
    \mprj/la_data_out [33],
    \mprj/la_data_out [32],
    \mprj/la_data_out [31],
    \mprj/la_data_out [30],
    \mprj/la_data_out [29],
    \mprj/la_data_out [28],
    \mprj/la_data_out [27],
    \mprj/la_data_out [26],
    \mprj/la_data_out [25],
    \mprj/la_data_out [24],
    \mprj/la_data_out [23],
    \mprj/la_data_out [22],
    \mprj/la_data_out [21],
    \mprj/la_data_out [20],
    \mprj/la_data_out [19],
    \mprj/la_data_out [18],
    \mprj/la_data_out [17],
    \mprj/la_data_out [16],
    \mprj/la_data_out [15],
    \mprj/la_data_out [14],
    \mprj/la_data_out [13],
    \mprj/la_data_out [12],
    \mprj/la_data_out [11],
    \mprj/la_data_out [10],
    \mprj/la_data_out [9],
    \mprj/la_data_out [8],
    \mprj/la_data_out [7],
    \mprj/la_data_out [6],
    \mprj/la_data_out [5],
    \mprj/la_data_out [4],
    \mprj/la_data_out [3],
    \mprj/la_data_out [2],
    \mprj/la_data_out [1],
    \mprj/la_data_out [0]}),
    .la_data_out_mprj({\soc/la_output [127],
    \soc/la_output [126],
    \soc/la_output [125],
    \soc/la_output [124],
    \soc/la_output [123],
    \soc/la_output [122],
    \soc/la_output [121],
    \soc/la_output [120],
    \soc/la_output [119],
    \soc/la_output [118],
    \soc/la_output [117],
    \soc/la_output [116],
    \soc/la_output [115],
    \soc/la_output [114],
    \soc/la_output [113],
    \soc/la_output [112],
    \soc/la_output [111],
    \soc/la_output [110],
    \soc/la_output [109],
    \soc/la_output [108],
    \soc/la_output [107],
    \soc/la_output [106],
    \soc/la_output [105],
    \soc/la_output [104],
    \soc/la_output [103],
    \soc/la_output [102],
    \soc/la_output [101],
    \soc/la_output [100],
    \soc/la_output [99],
    \soc/la_output [98],
    \soc/la_output [97],
    \soc/la_output [96],
    \soc/la_output [95],
    \soc/la_output [94],
    \soc/la_output [93],
    \soc/la_output [92],
    \soc/la_output [91],
    \soc/la_output [90],
    \soc/la_output [89],
    \soc/la_output [88],
    \soc/la_output [87],
    \soc/la_output [86],
    \soc/la_output [85],
    \soc/la_output [84],
    \soc/la_output [83],
    \soc/la_output [82],
    \soc/la_output [81],
    \soc/la_output [80],
    \soc/la_output [79],
    \soc/la_output [78],
    \soc/la_output [77],
    \soc/la_output [76],
    \soc/la_output [75],
    \soc/la_output [74],
    \soc/la_output [73],
    \soc/la_output [72],
    \soc/la_output [71],
    \soc/la_output [70],
    \soc/la_output [69],
    \soc/la_output [68],
    \soc/la_output [67],
    \soc/la_output [66],
    \soc/la_output [65],
    \soc/la_output [64],
    \soc/la_output [63],
    \soc/la_output [62],
    \soc/la_output [61],
    \soc/la_output [60],
    \soc/la_output [59],
    \soc/la_output [58],
    \soc/la_output [57],
    \soc/la_output [56],
    \soc/la_output [55],
    \soc/la_output [54],
    \soc/la_output [53],
    \soc/la_output [52],
    \soc/la_output [51],
    \soc/la_output [50],
    \soc/la_output [49],
    \soc/la_output [48],
    \soc/la_output [47],
    \soc/la_output [46],
    \soc/la_output [45],
    \soc/la_output [44],
    \soc/la_output [43],
    \soc/la_output [42],
    \soc/la_output [41],
    \soc/la_output [40],
    \soc/la_output [39],
    \soc/la_output [38],
    \soc/la_output [37],
    \soc/la_output [36],
    \soc/la_output [35],
    \soc/la_output [34],
    \soc/la_output [33],
    \soc/la_output [32],
    \soc/la_output [31],
    \soc/la_output [30],
    \soc/la_output [29],
    \soc/la_output [28],
    \soc/la_output [27],
    \soc/la_output [26],
    \soc/la_output [25],
    \soc/la_output [24],
    \soc/la_output [23],
    \soc/la_output [22],
    \soc/la_output [21],
    \soc/la_output [20],
    \soc/la_output [19],
    \soc/la_output [18],
    \soc/la_output [17],
    \soc/la_output [16],
    \soc/la_output [15],
    \soc/la_output [14],
    \soc/la_output [13],
    \soc/la_output [12],
    \soc/la_output [11],
    \soc/la_output [10],
    \soc/la_output [9],
    \soc/la_output [8],
    \soc/la_output [7],
    \soc/la_output [6],
    \soc/la_output [5],
    \soc/la_output [4],
    \soc/la_output [3],
    \soc/la_output [2],
    \soc/la_output [1],
    \soc/la_output [0]}),
    .la_iena_mprj({\soc/la_iena [127],
    \soc/la_iena [126],
    \soc/la_iena [125],
    \soc/la_iena [124],
    \soc/la_iena [123],
    \soc/la_iena [122],
    \soc/la_iena [121],
    \soc/la_iena [120],
    \soc/la_iena [119],
    \soc/la_iena [118],
    \soc/la_iena [117],
    \soc/la_iena [116],
    \soc/la_iena [115],
    \soc/la_iena [114],
    \soc/la_iena [113],
    \soc/la_iena [112],
    \soc/la_iena [111],
    \soc/la_iena [110],
    \soc/la_iena [109],
    \soc/la_iena [108],
    \soc/la_iena [107],
    \soc/la_iena [106],
    \soc/la_iena [105],
    \soc/la_iena [104],
    \soc/la_iena [103],
    \soc/la_iena [102],
    \soc/la_iena [101],
    \soc/la_iena [100],
    \soc/la_iena [99],
    \soc/la_iena [98],
    \soc/la_iena [97],
    \soc/la_iena [96],
    \soc/la_iena [95],
    \soc/la_iena [94],
    \soc/la_iena [93],
    \soc/la_iena [92],
    \soc/la_iena [91],
    \soc/la_iena [90],
    \soc/la_iena [89],
    \soc/la_iena [88],
    \soc/la_iena [87],
    \soc/la_iena [86],
    \soc/la_iena [85],
    \soc/la_iena [84],
    \soc/la_iena [83],
    \soc/la_iena [82],
    \soc/la_iena [81],
    \soc/la_iena [80],
    \soc/la_iena [79],
    \soc/la_iena [78],
    \soc/la_iena [77],
    \soc/la_iena [76],
    \soc/la_iena [75],
    \soc/la_iena [74],
    \soc/la_iena [73],
    \soc/la_iena [72],
    \soc/la_iena [71],
    \soc/la_iena [70],
    \soc/la_iena [69],
    \soc/la_iena [68],
    \soc/la_iena [67],
    \soc/la_iena [66],
    \soc/la_iena [65],
    \soc/la_iena [64],
    \soc/la_iena [63],
    \soc/la_iena [62],
    \soc/la_iena [61],
    \soc/la_iena [60],
    \soc/la_iena [59],
    \soc/la_iena [58],
    \soc/la_iena [57],
    \soc/la_iena [56],
    \soc/la_iena [55],
    \soc/la_iena [54],
    \soc/la_iena [53],
    \soc/la_iena [52],
    \soc/la_iena [51],
    \soc/la_iena [50],
    \soc/la_iena [49],
    \soc/la_iena [48],
    \soc/la_iena [47],
    \soc/la_iena [46],
    \soc/la_iena [45],
    \soc/la_iena [44],
    \soc/la_iena [43],
    \soc/la_iena [42],
    \soc/la_iena [41],
    \soc/la_iena [40],
    \soc/la_iena [39],
    \soc/la_iena [38],
    \soc/la_iena [37],
    \soc/la_iena [36],
    \soc/la_iena [35],
    \soc/la_iena [34],
    \soc/la_iena [33],
    \soc/la_iena [32],
    \soc/la_iena [31],
    \soc/la_iena [30],
    \soc/la_iena [29],
    \soc/la_iena [28],
    \soc/la_iena [27],
    \soc/la_iena [26],
    \soc/la_iena [25],
    \soc/la_iena [24],
    \soc/la_iena [23],
    \soc/la_iena [22],
    \soc/la_iena [21],
    \soc/la_iena [20],
    \soc/la_iena [19],
    \soc/la_iena [18],
    \soc/la_iena [17],
    \soc/la_iena [16],
    \soc/la_iena [15],
    \soc/la_iena [14],
    \soc/la_iena [13],
    \soc/la_iena [12],
    \soc/la_iena [11],
    \soc/la_iena [10],
    \soc/la_iena [9],
    \soc/la_iena [8],
    \soc/la_iena [7],
    \soc/la_iena [6],
    \soc/la_iena [5],
    \soc/la_iena [4],
    \soc/la_iena [3],
    \soc/la_iena [2],
    \soc/la_iena [1],
    \soc/la_iena [0]}),
    .la_oenb_core({\mprj/la_oenb [127],
    \mprj/la_oenb [126],
    \mprj/la_oenb [125],
    \mprj/la_oenb [124],
    \mprj/la_oenb [123],
    \mprj/la_oenb [122],
    \mprj/la_oenb [121],
    \mprj/la_oenb [120],
    \mprj/la_oenb [119],
    \mprj/la_oenb [118],
    \mprj/la_oenb [117],
    \mprj/la_oenb [116],
    \mprj/la_oenb [115],
    \mprj/la_oenb [114],
    \mprj/la_oenb [113],
    \mprj/la_oenb [112],
    \mprj/la_oenb [111],
    \mprj/la_oenb [110],
    \mprj/la_oenb [109],
    \mprj/la_oenb [108],
    \mprj/la_oenb [107],
    \mprj/la_oenb [106],
    \mprj/la_oenb [105],
    \mprj/la_oenb [104],
    \mprj/la_oenb [103],
    \mprj/la_oenb [102],
    \mprj/la_oenb [101],
    \mprj/la_oenb [100],
    \mprj/la_oenb [99],
    \mprj/la_oenb [98],
    \mprj/la_oenb [97],
    \mprj/la_oenb [96],
    \mprj/la_oenb [95],
    \mprj/la_oenb [94],
    \mprj/la_oenb [93],
    \mprj/la_oenb [92],
    \mprj/la_oenb [91],
    \mprj/la_oenb [90],
    \mprj/la_oenb [89],
    \mprj/la_oenb [88],
    \mprj/la_oenb [87],
    \mprj/la_oenb [86],
    \mprj/la_oenb [85],
    \mprj/la_oenb [84],
    \mprj/la_oenb [83],
    \mprj/la_oenb [82],
    \mprj/la_oenb [81],
    \mprj/la_oenb [80],
    \mprj/la_oenb [79],
    \mprj/la_oenb [78],
    \mprj/la_oenb [77],
    \mprj/la_oenb [76],
    \mprj/la_oenb [75],
    \mprj/la_oenb [74],
    \mprj/la_oenb [73],
    \mprj/la_oenb [72],
    \mprj/la_oenb [71],
    \mprj/la_oenb [70],
    \mprj/la_oenb [69],
    \mprj/la_oenb [68],
    \mprj/la_oenb [67],
    \mprj/la_oenb [66],
    \mprj/la_oenb [65],
    \mprj/la_oenb [64],
    \mprj/la_oenb [63],
    \mprj/la_oenb [62],
    \mprj/la_oenb [61],
    \mprj/la_oenb [60],
    \mprj/la_oenb [59],
    \mprj/la_oenb [58],
    \mprj/la_oenb [57],
    \mprj/la_oenb [56],
    \mprj/la_oenb [55],
    \mprj/la_oenb [54],
    \mprj/la_oenb [53],
    \mprj/la_oenb [52],
    \mprj/la_oenb [51],
    \mprj/la_oenb [50],
    \mprj/la_oenb [49],
    \mprj/la_oenb [48],
    \mprj/la_oenb [47],
    \mprj/la_oenb [46],
    \mprj/la_oenb [45],
    \mprj/la_oenb [44],
    \mprj/la_oenb [43],
    \mprj/la_oenb [42],
    \mprj/la_oenb [41],
    \mprj/la_oenb [40],
    \mprj/la_oenb [39],
    \mprj/la_oenb [38],
    \mprj/la_oenb [37],
    \mprj/la_oenb [36],
    \mprj/la_oenb [35],
    \mprj/la_oenb [34],
    \mprj/la_oenb [33],
    \mprj/la_oenb [32],
    \mprj/la_oenb [31],
    \mprj/la_oenb [30],
    \mprj/la_oenb [29],
    \mprj/la_oenb [28],
    \mprj/la_oenb [27],
    \mprj/la_oenb [26],
    \mprj/la_oenb [25],
    \mprj/la_oenb [24],
    \mprj/la_oenb [23],
    \mprj/la_oenb [22],
    \mprj/la_oenb [21],
    \mprj/la_oenb [20],
    \mprj/la_oenb [19],
    \mprj/la_oenb [18],
    \mprj/la_oenb [17],
    \mprj/la_oenb [16],
    \mprj/la_oenb [15],
    \mprj/la_oenb [14],
    \mprj/la_oenb [13],
    \mprj/la_oenb [12],
    \mprj/la_oenb [11],
    \mprj/la_oenb [10],
    \mprj/la_oenb [9],
    \mprj/la_oenb [8],
    \mprj/la_oenb [7],
    \mprj/la_oenb [6],
    \mprj/la_oenb [5],
    \mprj/la_oenb [4],
    \mprj/la_oenb [3],
    \mprj/la_oenb [2],
    \mprj/la_oenb [1],
    \mprj/la_oenb [0]}),
    .la_oenb_mprj({\soc/la_oenb [127],
    \soc/la_oenb [126],
    \soc/la_oenb [125],
    \soc/la_oenb [124],
    \soc/la_oenb [123],
    \soc/la_oenb [122],
    \soc/la_oenb [121],
    \soc/la_oenb [120],
    \soc/la_oenb [119],
    \soc/la_oenb [118],
    \soc/la_oenb [117],
    \soc/la_oenb [116],
    \soc/la_oenb [115],
    \soc/la_oenb [114],
    \soc/la_oenb [113],
    \soc/la_oenb [112],
    \soc/la_oenb [111],
    \soc/la_oenb [110],
    \soc/la_oenb [109],
    \soc/la_oenb [108],
    \soc/la_oenb [107],
    \soc/la_oenb [106],
    \soc/la_oenb [105],
    \soc/la_oenb [104],
    \soc/la_oenb [103],
    \soc/la_oenb [102],
    \soc/la_oenb [101],
    \soc/la_oenb [100],
    \soc/la_oenb [99],
    \soc/la_oenb [98],
    \soc/la_oenb [97],
    \soc/la_oenb [96],
    \soc/la_oenb [95],
    \soc/la_oenb [94],
    \soc/la_oenb [93],
    \soc/la_oenb [92],
    \soc/la_oenb [91],
    \soc/la_oenb [90],
    \soc/la_oenb [89],
    \soc/la_oenb [88],
    \soc/la_oenb [87],
    \soc/la_oenb [86],
    \soc/la_oenb [85],
    \soc/la_oenb [84],
    \soc/la_oenb [83],
    \soc/la_oenb [82],
    \soc/la_oenb [81],
    \soc/la_oenb [80],
    \soc/la_oenb [79],
    \soc/la_oenb [78],
    \soc/la_oenb [77],
    \soc/la_oenb [76],
    \soc/la_oenb [75],
    \soc/la_oenb [74],
    \soc/la_oenb [73],
    \soc/la_oenb [72],
    \soc/la_oenb [71],
    \soc/la_oenb [70],
    \soc/la_oenb [69],
    \soc/la_oenb [68],
    \soc/la_oenb [67],
    \soc/la_oenb [66],
    \soc/la_oenb [65],
    \soc/la_oenb [64],
    \soc/la_oenb [63],
    \soc/la_oenb [62],
    \soc/la_oenb [61],
    \soc/la_oenb [60],
    \soc/la_oenb [59],
    \soc/la_oenb [58],
    \soc/la_oenb [57],
    \soc/la_oenb [56],
    \soc/la_oenb [55],
    \soc/la_oenb [54],
    \soc/la_oenb [53],
    \soc/la_oenb [52],
    \soc/la_oenb [51],
    \soc/la_oenb [50],
    \soc/la_oenb [49],
    \soc/la_oenb [48],
    \soc/la_oenb [47],
    \soc/la_oenb [46],
    \soc/la_oenb [45],
    \soc/la_oenb [44],
    \soc/la_oenb [43],
    \soc/la_oenb [42],
    \soc/la_oenb [41],
    \soc/la_oenb [40],
    \soc/la_oenb [39],
    \soc/la_oenb [38],
    \soc/la_oenb [37],
    \soc/la_oenb [36],
    \soc/la_oenb [35],
    \soc/la_oenb [34],
    \soc/la_oenb [33],
    \soc/la_oenb [32],
    \soc/la_oenb [31],
    \soc/la_oenb [30],
    \soc/la_oenb [29],
    \soc/la_oenb [28],
    \soc/la_oenb [27],
    \soc/la_oenb [26],
    \soc/la_oenb [25],
    \soc/la_oenb [24],
    \soc/la_oenb [23],
    \soc/la_oenb [22],
    \soc/la_oenb [21],
    \soc/la_oenb [20],
    \soc/la_oenb [19],
    \soc/la_oenb [18],
    \soc/la_oenb [17],
    \soc/la_oenb [16],
    \soc/la_oenb [15],
    \soc/la_oenb [14],
    \soc/la_oenb [13],
    \soc/la_oenb [12],
    \soc/la_oenb [11],
    \soc/la_oenb [10],
    \soc/la_oenb [9],
    \soc/la_oenb [8],
    \soc/la_oenb [7],
    \soc/la_oenb [6],
    \soc/la_oenb [5],
    \soc/la_oenb [4],
    \soc/la_oenb [3],
    \soc/la_oenb [2],
    \soc/la_oenb [1],
    \soc/la_oenb [0]}),
    .mprj_adr_o_core({\soc/mprj_adr_o [31],
    \soc/mprj_adr_o [30],
    \soc/mprj_adr_o [29],
    \soc/mprj_adr_o [28],
    \soc/mprj_adr_o [27],
    \soc/mprj_adr_o [26],
    \soc/mprj_adr_o [25],
    \soc/mprj_adr_o [24],
    \soc/mprj_adr_o [23],
    \soc/mprj_adr_o [22],
    \soc/mprj_adr_o [21],
    \soc/mprj_adr_o [20],
    \soc/mprj_adr_o [19],
    \soc/mprj_adr_o [18],
    \soc/mprj_adr_o [17],
    \soc/mprj_adr_o [16],
    \soc/mprj_adr_o [15],
    \soc/mprj_adr_o [14],
    \soc/mprj_adr_o [13],
    \soc/mprj_adr_o [12],
    \soc/mprj_adr_o [11],
    \soc/mprj_adr_o [10],
    \soc/mprj_adr_o [9],
    \soc/mprj_adr_o [8],
    \soc/mprj_adr_o [7],
    \soc/mprj_adr_o [6],
    \soc/mprj_adr_o [5],
    \soc/mprj_adr_o [4],
    \soc/mprj_adr_o [3],
    \soc/mprj_adr_o [2],
    \soc/mprj_adr_o [1],
    \soc/mprj_adr_o [0]}),
    .mprj_adr_o_user({\mprj/wbs_adr_i [31],
    \mprj/wbs_adr_i [30],
    \mprj/wbs_adr_i [29],
    \mprj/wbs_adr_i [28],
    \mprj/wbs_adr_i [27],
    \mprj/wbs_adr_i [26],
    \mprj/wbs_adr_i [25],
    \mprj/wbs_adr_i [24],
    \mprj/wbs_adr_i [23],
    \mprj/wbs_adr_i [22],
    \mprj/wbs_adr_i [21],
    \mprj/wbs_adr_i [20],
    \mprj/wbs_adr_i [19],
    \mprj/wbs_adr_i [18],
    \mprj/wbs_adr_i [17],
    \mprj/wbs_adr_i [16],
    \mprj/wbs_adr_i [15],
    \mprj/wbs_adr_i [14],
    \mprj/wbs_adr_i [13],
    \mprj/wbs_adr_i [12],
    \mprj/wbs_adr_i [11],
    \mprj/wbs_adr_i [10],
    \mprj/wbs_adr_i [9],
    \mprj/wbs_adr_i [8],
    \mprj/wbs_adr_i [7],
    \mprj/wbs_adr_i [6],
    \mprj/wbs_adr_i [5],
    \mprj/wbs_adr_i [4],
    \mprj/wbs_adr_i [3],
    \mprj/wbs_adr_i [2],
    \mprj/wbs_adr_i [1],
    \mprj/wbs_adr_i [0]}),
    .mprj_dat_i_core({\soc/mprj_dat_i [31],
    \soc/mprj_dat_i [30],
    \soc/mprj_dat_i [29],
    \soc/mprj_dat_i [28],
    \soc/mprj_dat_i [27],
    \soc/mprj_dat_i [26],
    \soc/mprj_dat_i [25],
    \soc/mprj_dat_i [24],
    \soc/mprj_dat_i [23],
    \soc/mprj_dat_i [22],
    \soc/mprj_dat_i [21],
    \soc/mprj_dat_i [20],
    \soc/mprj_dat_i [19],
    \soc/mprj_dat_i [18],
    \soc/mprj_dat_i [17],
    \soc/mprj_dat_i [16],
    \soc/mprj_dat_i [15],
    \soc/mprj_dat_i [14],
    \soc/mprj_dat_i [13],
    \soc/mprj_dat_i [12],
    \soc/mprj_dat_i [11],
    \soc/mprj_dat_i [10],
    \soc/mprj_dat_i [9],
    \soc/mprj_dat_i [8],
    \soc/mprj_dat_i [7],
    \soc/mprj_dat_i [6],
    \soc/mprj_dat_i [5],
    \soc/mprj_dat_i [4],
    \soc/mprj_dat_i [3],
    \soc/mprj_dat_i [2],
    \soc/mprj_dat_i [1],
    \soc/mprj_dat_i [0]}),
    .mprj_dat_i_user({\mprj/wbs_dat_o [31],
    \mprj/wbs_dat_o [30],
    \mprj/wbs_dat_o [29],
    \mprj/wbs_dat_o [28],
    \mprj/wbs_dat_o [27],
    \mprj/wbs_dat_o [26],
    \mprj/wbs_dat_o [25],
    \mprj/wbs_dat_o [24],
    \mprj/wbs_dat_o [23],
    \mprj/wbs_dat_o [22],
    \mprj/wbs_dat_o [21],
    \mprj/wbs_dat_o [20],
    \mprj/wbs_dat_o [19],
    \mprj/wbs_dat_o [18],
    \mprj/wbs_dat_o [17],
    \mprj/wbs_dat_o [16],
    \mprj/wbs_dat_o [15],
    \mprj/wbs_dat_o [14],
    \mprj/wbs_dat_o [13],
    \mprj/wbs_dat_o [12],
    \mprj/wbs_dat_o [11],
    \mprj/wbs_dat_o [10],
    \mprj/wbs_dat_o [9],
    \mprj/wbs_dat_o [8],
    \mprj/wbs_dat_o [7],
    \mprj/wbs_dat_o [6],
    \mprj/wbs_dat_o [5],
    \mprj/wbs_dat_o [4],
    \mprj/wbs_dat_o [3],
    \mprj/wbs_dat_o [2],
    \mprj/wbs_dat_o [1],
    \mprj/wbs_dat_o [0]}),
    .mprj_dat_o_core({\soc/mprj_dat_o [31],
    \soc/mprj_dat_o [30],
    \soc/mprj_dat_o [29],
    \soc/mprj_dat_o [28],
    \soc/mprj_dat_o [27],
    \soc/mprj_dat_o [26],
    \soc/mprj_dat_o [25],
    \soc/mprj_dat_o [24],
    \soc/mprj_dat_o [23],
    \soc/mprj_dat_o [22],
    \soc/mprj_dat_o [21],
    \soc/mprj_dat_o [20],
    \soc/mprj_dat_o [19],
    \soc/mprj_dat_o [18],
    \soc/mprj_dat_o [17],
    \soc/mprj_dat_o [16],
    \soc/mprj_dat_o [15],
    \soc/mprj_dat_o [14],
    \soc/mprj_dat_o [13],
    \soc/mprj_dat_o [12],
    \soc/mprj_dat_o [11],
    \soc/mprj_dat_o [10],
    \soc/mprj_dat_o [9],
    \soc/mprj_dat_o [8],
    \soc/mprj_dat_o [7],
    \soc/mprj_dat_o [6],
    \soc/mprj_dat_o [5],
    \soc/mprj_dat_o [4],
    \soc/mprj_dat_o [3],
    \soc/mprj_dat_o [2],
    \soc/mprj_dat_o [1],
    \soc/mprj_dat_o [0]}),
    .mprj_dat_o_user({\mprj/wbs_dat_i [31],
    \mprj/wbs_dat_i [30],
    \mprj/wbs_dat_i [29],
    \mprj/wbs_dat_i [28],
    \mprj/wbs_dat_i [27],
    \mprj/wbs_dat_i [26],
    \mprj/wbs_dat_i [25],
    \mprj/wbs_dat_i [24],
    \mprj/wbs_dat_i [23],
    \mprj/wbs_dat_i [22],
    \mprj/wbs_dat_i [21],
    \mprj/wbs_dat_i [20],
    \mprj/wbs_dat_i [19],
    \mprj/wbs_dat_i [18],
    \mprj/wbs_dat_i [17],
    \mprj/wbs_dat_i [16],
    \mprj/wbs_dat_i [15],
    \mprj/wbs_dat_i [14],
    \mprj/wbs_dat_i [13],
    \mprj/wbs_dat_i [12],
    \mprj/wbs_dat_i [11],
    \mprj/wbs_dat_i [10],
    \mprj/wbs_dat_i [9],
    \mprj/wbs_dat_i [8],
    \mprj/wbs_dat_i [7],
    \mprj/wbs_dat_i [6],
    \mprj/wbs_dat_i [5],
    \mprj/wbs_dat_i [4],
    \mprj/wbs_dat_i [3],
    \mprj/wbs_dat_i [2],
    \mprj/wbs_dat_i [1],
    \mprj/wbs_dat_i [0]}),
    .mprj_sel_o_core({\soc/mprj_sel_o [3],
    \soc/mprj_sel_o [2],
    \soc/mprj_sel_o [1],
    \soc/mprj_sel_o [0]}),
    .mprj_sel_o_user({\mprj/wbs_sel_i [3],
    \mprj/wbs_sel_i [2],
    \mprj/wbs_sel_i [1],
    \mprj/wbs_sel_i [0]}),
    .user_irq({\soc/irq [2],
    \soc/irq [1],
    \soc/irq [0]}),
    .user_irq_core({\mprj/user_irq [2],
    \mprj/user_irq [1],
    \mprj/user_irq [0]}),
    .user_irq_ena({\soc/user_irq_ena [2],
    \soc/user_irq_ena [1],
    \soc/user_irq_ena [0]}));
 spare_logic_block spare_logic_block_2 (.spare_xib(\spare_logic_block_2/spare_xib ),
    .spare_xfq({\spare_logic_block_2/spare_xfq [1],
    \spare_logic_block_2/spare_xfq [0]}),
    .spare_xfqn({\spare_logic_block_2/spare_xfqn [1],
    \spare_logic_block_2/spare_xfqn [0]}),
    .spare_xi({\spare_logic_block_2/spare_xi [3],
    \spare_logic_block_2/spare_xi [2],
    \spare_logic_block_2/spare_xi [1],
    \spare_logic_block_2/spare_xi [0]}),
    .spare_xmx({\spare_logic_block_2/spare_xmx [1],
    \spare_logic_block_2/spare_xmx [0]}),
    .spare_xna({\spare_logic_block_2/spare_xna [1],
    \spare_logic_block_2/spare_xna [0]}),
    .spare_xno({\spare_logic_block_2/spare_xno [1],
    \spare_logic_block_2/spare_xno [0]}),
    .spare_xz({\spare_logic_block_2/spare_xz [26],
    \spare_logic_block_2/spare_xz [25],
    \spare_logic_block_2/spare_xz [24],
    \spare_logic_block_2/spare_xz [23],
    \spare_logic_block_2/spare_xz [22],
    \spare_logic_block_2/spare_xz [21],
    \spare_logic_block_2/spare_xz [20],
    \spare_logic_block_2/spare_xz [19],
    \spare_logic_block_2/spare_xz [18],
    \spare_logic_block_2/spare_xz [17],
    \spare_logic_block_2/spare_xz [16],
    \spare_logic_block_2/spare_xz [15],
    \spare_logic_block_2/spare_xz [14],
    \spare_logic_block_2/spare_xz [13],
    \spare_logic_block_2/spare_xz [12],
    \spare_logic_block_2/spare_xz [11],
    \spare_logic_block_2/spare_xz [10],
    \spare_logic_block_2/spare_xz [9],
    \spare_logic_block_2/spare_xz [8],
    \spare_logic_block_2/spare_xz [7],
    \spare_logic_block_2/spare_xz [6],
    \spare_logic_block_2/spare_xz [5],
    \spare_logic_block_2/spare_xz [4],
    \spare_logic_block_2/spare_xz [3],
    \spare_logic_block_2/spare_xz [2],
    \spare_logic_block_2/spare_xz [1],
    \spare_logic_block_2/spare_xz [0]}));
 spare_logic_block spare_logic_block_0 (.spare_xib(\spare_logic_block_0/spare_xib ),
    .spare_xfq({\spare_logic_block_0/spare_xfq [1],
    \spare_logic_block_0/spare_xfq [0]}),
    .spare_xfqn({\spare_logic_block_0/spare_xfqn [1],
    \spare_logic_block_0/spare_xfqn [0]}),
    .spare_xi({\spare_logic_block_0/spare_xi [3],
    \spare_logic_block_0/spare_xi [2],
    \spare_logic_block_0/spare_xi [1],
    \spare_logic_block_0/spare_xi [0]}),
    .spare_xmx({\spare_logic_block_0/spare_xmx [1],
    \spare_logic_block_0/spare_xmx [0]}),
    .spare_xna({\spare_logic_block_0/spare_xna [1],
    \spare_logic_block_0/spare_xna [0]}),
    .spare_xno({\spare_logic_block_0/spare_xno [1],
    \spare_logic_block_0/spare_xno [0]}),
    .spare_xz({\spare_logic_block_0/spare_xz [26],
    \spare_logic_block_0/spare_xz [25],
    \spare_logic_block_0/spare_xz [24],
    \spare_logic_block_0/spare_xz [23],
    \spare_logic_block_0/spare_xz [22],
    \spare_logic_block_0/spare_xz [21],
    \spare_logic_block_0/spare_xz [20],
    \spare_logic_block_0/spare_xz [19],
    \spare_logic_block_0/spare_xz [18],
    \spare_logic_block_0/spare_xz [17],
    \spare_logic_block_0/spare_xz [16],
    \spare_logic_block_0/spare_xz [15],
    \spare_logic_block_0/spare_xz [14],
    \spare_logic_block_0/spare_xz [13],
    \spare_logic_block_0/spare_xz [12],
    \spare_logic_block_0/spare_xz [11],
    \spare_logic_block_0/spare_xz [10],
    \spare_logic_block_0/spare_xz [9],
    \spare_logic_block_0/spare_xz [8],
    \spare_logic_block_0/spare_xz [7],
    \spare_logic_block_0/spare_xz [6],
    \spare_logic_block_0/spare_xz [5],
    \spare_logic_block_0/spare_xz [4],
    \spare_logic_block_0/spare_xz [3],
    \spare_logic_block_0/spare_xz [2],
    \spare_logic_block_0/spare_xz [1],
    \spare_logic_block_0/spare_xz [0]}));
 gpio_defaults_block_0403 gpio_defaults_block_2 (.gpio_defaults({\gpio_defaults_block_2/gpio_defaults [12],
    \gpio_defaults_block_2/gpio_defaults [11],
    \gpio_defaults_block_2/gpio_defaults [10],
    \gpio_defaults_block_2/gpio_defaults [9],
    \gpio_defaults_block_2/gpio_defaults [8],
    \gpio_defaults_block_2/gpio_defaults [7],
    \gpio_defaults_block_2/gpio_defaults [6],
    \gpio_defaults_block_2/gpio_defaults [5],
    \gpio_defaults_block_2/gpio_defaults [4],
    \gpio_defaults_block_2/gpio_defaults [3],
    \gpio_defaults_block_2/gpio_defaults [2],
    \gpio_defaults_block_2/gpio_defaults [1],
    \gpio_defaults_block_2/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1a[0]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [2]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[0]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [2]),
    .one(\gpio_control_in_1a[0]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [2]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [2]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [2]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [2]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [2]),
    .pad_gpio_in(\padframe/mprj_io_in [2]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [2]),
    .pad_gpio_out(\padframe/mprj_io_out [2]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [2]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [2]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [2]),
    .resetn(\gpio_control_in_1a[0]/resetn ),
    .resetn_out(\gpio_control_in_1a[1]/resetn ),
    .serial_clock(\gpio_control_in_1a[0]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[1]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[0]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[1]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[0]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[1]/serial_load ),
    .user_gpio_in(\mprj/io_in [2]),
    .user_gpio_oeb(\mprj/io_oeb [2]),
    .user_gpio_out(\mprj/io_out [2]),
    .zero(\gpio_control_in_1a[0]/zero ),
    .gpio_defaults({\gpio_defaults_block_2/gpio_defaults [12],
    \gpio_defaults_block_2/gpio_defaults [11],
    \gpio_defaults_block_2/gpio_defaults [10],
    \gpio_defaults_block_2/gpio_defaults [9],
    \gpio_defaults_block_2/gpio_defaults [8],
    \gpio_defaults_block_2/gpio_defaults [7],
    \gpio_defaults_block_2/gpio_defaults [6],
    \gpio_defaults_block_2/gpio_defaults [5],
    \gpio_defaults_block_2/gpio_defaults [4],
    \gpio_defaults_block_2/gpio_defaults [3],
    \gpio_defaults_block_2/gpio_defaults [2],
    \gpio_defaults_block_2/gpio_defaults [1],
    \gpio_defaults_block_2/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [8],
    \padframe/mprj_io_dm [7],
    \padframe/mprj_io_dm [6]}));
 gpio_defaults_block gpio_defaults_block_36 (.gpio_defaults({\gpio_defaults_block_36/gpio_defaults [12],
    \gpio_defaults_block_36/gpio_defaults [11],
    \gpio_defaults_block_36/gpio_defaults [10],
    \gpio_defaults_block_36/gpio_defaults [9],
    \gpio_defaults_block_36/gpio_defaults [8],
    \gpio_defaults_block_36/gpio_defaults [7],
    \gpio_defaults_block_36/gpio_defaults [6],
    \gpio_defaults_block_36/gpio_defaults [5],
    \gpio_defaults_block_36/gpio_defaults [4],
    \gpio_defaults_block_36/gpio_defaults [3],
    \gpio_defaults_block_36/gpio_defaults [2],
    \gpio_defaults_block_36/gpio_defaults [1],
    \gpio_defaults_block_36/gpio_defaults [0]}));
 gpio_defaults_block_0403 gpio_defaults_block_3 (.gpio_defaults({\gpio_defaults_block_3/gpio_defaults [12],
    \gpio_defaults_block_3/gpio_defaults [11],
    \gpio_defaults_block_3/gpio_defaults [10],
    \gpio_defaults_block_3/gpio_defaults [9],
    \gpio_defaults_block_3/gpio_defaults [8],
    \gpio_defaults_block_3/gpio_defaults [7],
    \gpio_defaults_block_3/gpio_defaults [6],
    \gpio_defaults_block_3/gpio_defaults [5],
    \gpio_defaults_block_3/gpio_defaults [4],
    \gpio_defaults_block_3/gpio_defaults [3],
    \gpio_defaults_block_3/gpio_defaults [2],
    \gpio_defaults_block_3/gpio_defaults [1],
    \gpio_defaults_block_3/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1a[1]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [3]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[1]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [3]),
    .one(\gpio_control_in_1a[1]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [3]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [3]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [3]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [3]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [3]),
    .pad_gpio_in(\padframe/mprj_io_in [3]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [3]),
    .pad_gpio_out(\padframe/mprj_io_out [3]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [3]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [3]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [3]),
    .resetn(\gpio_control_in_1a[1]/resetn ),
    .resetn_out(\gpio_control_in_1a[2]/resetn ),
    .serial_clock(\gpio_control_in_1a[1]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[2]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[1]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[2]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[1]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[2]/serial_load ),
    .user_gpio_in(\mprj/io_in [3]),
    .user_gpio_oeb(\mprj/io_oeb [3]),
    .user_gpio_out(\mprj/io_out [3]),
    .zero(\gpio_control_in_1a[1]/zero ),
    .gpio_defaults({\gpio_defaults_block_3/gpio_defaults [12],
    \gpio_defaults_block_3/gpio_defaults [11],
    \gpio_defaults_block_3/gpio_defaults [10],
    \gpio_defaults_block_3/gpio_defaults [9],
    \gpio_defaults_block_3/gpio_defaults [8],
    \gpio_defaults_block_3/gpio_defaults [7],
    \gpio_defaults_block_3/gpio_defaults [6],
    \gpio_defaults_block_3/gpio_defaults [5],
    \gpio_defaults_block_3/gpio_defaults [4],
    \gpio_defaults_block_3/gpio_defaults [3],
    \gpio_defaults_block_3/gpio_defaults [2],
    \gpio_defaults_block_3/gpio_defaults [1],
    \gpio_defaults_block_3/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [11],
    \padframe/mprj_io_dm [10],
    \padframe/mprj_io_dm [9]}));
 gpio_control_block \gpio_control_bidir_2[0]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [35]),
    .mgmt_gpio_oeb(\housekeeping/mgmt_gpio_oeb [35]),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_out [35]),
    .one(\gpio_control_bidir_2[0]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [35]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [35]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [35]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [35]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [35]),
    .pad_gpio_in(\padframe/mprj_io_in [35]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [35]),
    .pad_gpio_out(\padframe/mprj_io_out [35]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [35]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [35]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [35]),
    .resetn(\gpio_control_bidir_2[0]/resetn ),
    .resetn_out(\gpio_control_in_2[15]/resetn ),
    .serial_clock(\gpio_control_bidir_2[0]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[15]/serial_clock ),
    .serial_data_in(\gpio_control_bidir_2[0]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[15]/serial_data_in ),
    .serial_load(\gpio_control_bidir_2[0]/serial_load ),
    .serial_load_out(\gpio_control_in_2[15]/serial_load ),
    .user_gpio_in(\mprj/io_in [35]),
    .user_gpio_oeb(\mprj/io_oeb [35]),
    .user_gpio_out(\mprj/io_out [35]),
    .zero(\gpio_control_bidir_2[0]/zero ),
    .gpio_defaults({\gpio_defaults_block_35/gpio_defaults [12],
    \gpio_defaults_block_35/gpio_defaults [11],
    \gpio_defaults_block_35/gpio_defaults [10],
    \gpio_defaults_block_35/gpio_defaults [9],
    \gpio_defaults_block_35/gpio_defaults [8],
    \gpio_defaults_block_35/gpio_defaults [7],
    \gpio_defaults_block_35/gpio_defaults [6],
    \gpio_defaults_block_35/gpio_defaults [5],
    \gpio_defaults_block_35/gpio_defaults [4],
    \gpio_defaults_block_35/gpio_defaults [3],
    \gpio_defaults_block_35/gpio_defaults [2],
    \gpio_defaults_block_35/gpio_defaults [1],
    \gpio_defaults_block_35/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [107],
    \padframe/mprj_io_dm [106],
    \padframe/mprj_io_dm [105]}));
 gpio_defaults_block gpio_defaults_block_35 (.gpio_defaults({\gpio_defaults_block_35/gpio_defaults [12],
    \gpio_defaults_block_35/gpio_defaults [11],
    \gpio_defaults_block_35/gpio_defaults [10],
    \gpio_defaults_block_35/gpio_defaults [9],
    \gpio_defaults_block_35/gpio_defaults [8],
    \gpio_defaults_block_35/gpio_defaults [7],
    \gpio_defaults_block_35/gpio_defaults [6],
    \gpio_defaults_block_35/gpio_defaults [5],
    \gpio_defaults_block_35/gpio_defaults [4],
    \gpio_defaults_block_35/gpio_defaults [3],
    \gpio_defaults_block_35/gpio_defaults [2],
    \gpio_defaults_block_35/gpio_defaults [1],
    \gpio_defaults_block_35/gpio_defaults [0]}));
 gpio_defaults_block_0403 gpio_defaults_block_4 (.gpio_defaults({\gpio_defaults_block_4/gpio_defaults [12],
    \gpio_defaults_block_4/gpio_defaults [11],
    \gpio_defaults_block_4/gpio_defaults [10],
    \gpio_defaults_block_4/gpio_defaults [9],
    \gpio_defaults_block_4/gpio_defaults [8],
    \gpio_defaults_block_4/gpio_defaults [7],
    \gpio_defaults_block_4/gpio_defaults [6],
    \gpio_defaults_block_4/gpio_defaults [5],
    \gpio_defaults_block_4/gpio_defaults [4],
    \gpio_defaults_block_4/gpio_defaults [3],
    \gpio_defaults_block_4/gpio_defaults [2],
    \gpio_defaults_block_4/gpio_defaults [1],
    \gpio_defaults_block_4/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1a[2]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [4]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[2]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [4]),
    .one(\gpio_control_in_1a[2]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [4]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [4]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [4]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [4]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [4]),
    .pad_gpio_in(\padframe/mprj_io_in [4]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [4]),
    .pad_gpio_out(\padframe/mprj_io_out [4]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [4]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [4]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [4]),
    .resetn(\gpio_control_in_1a[2]/resetn ),
    .resetn_out(\gpio_control_in_1a[3]/resetn ),
    .serial_clock(\gpio_control_in_1a[2]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[3]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[2]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[3]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[2]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[3]/serial_load ),
    .user_gpio_in(\mprj/io_in [4]),
    .user_gpio_oeb(\mprj/io_oeb [4]),
    .user_gpio_out(\mprj/io_out [4]),
    .zero(\gpio_control_in_1a[2]/zero ),
    .gpio_defaults({\gpio_defaults_block_4/gpio_defaults [12],
    \gpio_defaults_block_4/gpio_defaults [11],
    \gpio_defaults_block_4/gpio_defaults [10],
    \gpio_defaults_block_4/gpio_defaults [9],
    \gpio_defaults_block_4/gpio_defaults [8],
    \gpio_defaults_block_4/gpio_defaults [7],
    \gpio_defaults_block_4/gpio_defaults [6],
    \gpio_defaults_block_4/gpio_defaults [5],
    \gpio_defaults_block_4/gpio_defaults [4],
    \gpio_defaults_block_4/gpio_defaults [3],
    \gpio_defaults_block_4/gpio_defaults [2],
    \gpio_defaults_block_4/gpio_defaults [1],
    \gpio_defaults_block_4/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [14],
    \padframe/mprj_io_dm [13],
    \padframe/mprj_io_dm [12]}));
 gpio_control_block \gpio_control_in_2[15]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [34]),
    .mgmt_gpio_oeb(\gpio_control_in_2[15]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [34]),
    .one(\gpio_control_in_2[15]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [34]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [34]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [34]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [34]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [34]),
    .pad_gpio_in(\padframe/mprj_io_in [34]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [34]),
    .pad_gpio_out(\padframe/mprj_io_out [34]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [34]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [34]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [34]),
    .resetn(\gpio_control_in_2[15]/resetn ),
    .resetn_out(\gpio_control_in_2[14]/resetn ),
    .serial_clock(\gpio_control_in_2[15]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[14]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[15]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[14]/serial_data_in ),
    .serial_load(\gpio_control_in_2[15]/serial_load ),
    .serial_load_out(\gpio_control_in_2[14]/serial_load ),
    .user_gpio_in(\mprj/io_in [34]),
    .user_gpio_oeb(\mprj/io_oeb [34]),
    .user_gpio_out(\mprj/io_out [34]),
    .zero(\gpio_control_in_2[15]/zero ),
    .gpio_defaults({\gpio_control_in_2[15]/gpio_defaults [12],
    \gpio_control_in_2[15]/gpio_defaults [11],
    \gpio_control_in_2[15]/gpio_defaults [10],
    \gpio_control_in_2[15]/gpio_defaults [9],
    \gpio_control_in_2[15]/gpio_defaults [8],
    \gpio_control_in_2[15]/gpio_defaults [7],
    \gpio_control_in_2[15]/gpio_defaults [6],
    \gpio_control_in_2[15]/gpio_defaults [5],
    \gpio_control_in_2[15]/gpio_defaults [4],
    \gpio_control_in_2[15]/gpio_defaults [3],
    \gpio_control_in_2[15]/gpio_defaults [2],
    \gpio_control_in_2[15]/gpio_defaults [1],
    \gpio_control_in_2[15]/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [104],
    \padframe/mprj_io_dm [103],
    \padframe/mprj_io_dm [102]}));
 gpio_control_block \gpio_control_in_2[14]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [33]),
    .mgmt_gpio_oeb(\gpio_control_in_2[14]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [33]),
    .one(\gpio_control_in_2[14]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [33]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [33]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [33]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [33]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [33]),
    .pad_gpio_in(\padframe/mprj_io_in [33]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [33]),
    .pad_gpio_out(\padframe/mprj_io_out [33]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [33]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [33]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [33]),
    .resetn(\gpio_control_in_2[14]/resetn ),
    .resetn_out(\gpio_control_in_2[13]/resetn ),
    .serial_clock(\gpio_control_in_2[14]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[13]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[14]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[13]/serial_data_in ),
    .serial_load(\gpio_control_in_2[14]/serial_load ),
    .serial_load_out(\gpio_control_in_2[13]/serial_load ),
    .user_gpio_in(\mprj/io_in [33]),
    .user_gpio_oeb(\mprj/io_oeb [33]),
    .user_gpio_out(\mprj/io_out [33]),
    .zero(\gpio_control_in_2[14]/zero ),
    .gpio_defaults({\gpio_defaults_block_33/gpio_defaults [12],
    \gpio_defaults_block_33/gpio_defaults [11],
    \gpio_defaults_block_33/gpio_defaults [10],
    \gpio_defaults_block_33/gpio_defaults [9],
    \gpio_defaults_block_33/gpio_defaults [8],
    \gpio_defaults_block_33/gpio_defaults [7],
    \gpio_defaults_block_33/gpio_defaults [6],
    \gpio_defaults_block_33/gpio_defaults [5],
    \gpio_defaults_block_33/gpio_defaults [4],
    \gpio_defaults_block_33/gpio_defaults [3],
    \gpio_defaults_block_33/gpio_defaults [2],
    \gpio_defaults_block_33/gpio_defaults [1],
    \gpio_defaults_block_33/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [101],
    \padframe/mprj_io_dm [100],
    \padframe/mprj_io_dm [99]}));
 gpio_control_block \gpio_control_in_2[13]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [32]),
    .mgmt_gpio_oeb(\gpio_control_in_2[13]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [32]),
    .one(\gpio_control_in_2[13]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [32]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [32]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [32]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [32]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [32]),
    .pad_gpio_in(\padframe/mprj_io_in [32]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [32]),
    .pad_gpio_out(\padframe/mprj_io_out [32]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [32]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [32]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [32]),
    .resetn(\gpio_control_in_2[13]/resetn ),
    .resetn_out(\gpio_control_in_2[12]/resetn ),
    .serial_clock(\gpio_control_in_2[13]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[12]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[13]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[12]/serial_data_in ),
    .serial_load(\gpio_control_in_2[13]/serial_load ),
    .serial_load_out(\gpio_control_in_2[12]/serial_load ),
    .user_gpio_in(\mprj/io_in [32]),
    .user_gpio_oeb(\mprj/io_oeb [32]),
    .user_gpio_out(\mprj/io_out [32]),
    .zero(\gpio_control_in_2[13]/zero ),
    .gpio_defaults({\gpio_defaults_block_32/gpio_defaults [12],
    \gpio_defaults_block_32/gpio_defaults [11],
    \gpio_defaults_block_32/gpio_defaults [10],
    \gpio_defaults_block_32/gpio_defaults [9],
    \gpio_defaults_block_32/gpio_defaults [8],
    \gpio_defaults_block_32/gpio_defaults [7],
    \gpio_defaults_block_32/gpio_defaults [6],
    \gpio_defaults_block_32/gpio_defaults [5],
    \gpio_defaults_block_32/gpio_defaults [4],
    \gpio_defaults_block_32/gpio_defaults [3],
    \gpio_defaults_block_32/gpio_defaults [2],
    \gpio_defaults_block_32/gpio_defaults [1],
    \gpio_defaults_block_32/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [98],
    \padframe/mprj_io_dm [97],
    \padframe/mprj_io_dm [96]}));
 gpio_defaults_block gpio_defaults_defaults_block_34 (.gpio_defaults({\gpio_control_in_2[15]/gpio_defaults [12],
    \gpio_control_in_2[15]/gpio_defaults [11],
    \gpio_control_in_2[15]/gpio_defaults [10],
    \gpio_control_in_2[15]/gpio_defaults [9],
    \gpio_control_in_2[15]/gpio_defaults [8],
    \gpio_control_in_2[15]/gpio_defaults [7],
    \gpio_control_in_2[15]/gpio_defaults [6],
    \gpio_control_in_2[15]/gpio_defaults [5],
    \gpio_control_in_2[15]/gpio_defaults [4],
    \gpio_control_in_2[15]/gpio_defaults [3],
    \gpio_control_in_2[15]/gpio_defaults [2],
    \gpio_control_in_2[15]/gpio_defaults [1],
    \gpio_control_in_2[15]/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_33 (.gpio_defaults({\gpio_defaults_block_33/gpio_defaults [12],
    \gpio_defaults_block_33/gpio_defaults [11],
    \gpio_defaults_block_33/gpio_defaults [10],
    \gpio_defaults_block_33/gpio_defaults [9],
    \gpio_defaults_block_33/gpio_defaults [8],
    \gpio_defaults_block_33/gpio_defaults [7],
    \gpio_defaults_block_33/gpio_defaults [6],
    \gpio_defaults_block_33/gpio_defaults [5],
    \gpio_defaults_block_33/gpio_defaults [4],
    \gpio_defaults_block_33/gpio_defaults [3],
    \gpio_defaults_block_33/gpio_defaults [2],
    \gpio_defaults_block_33/gpio_defaults [1],
    \gpio_defaults_block_33/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_32 (.gpio_defaults({\gpio_defaults_block_32/gpio_defaults [12],
    \gpio_defaults_block_32/gpio_defaults [11],
    \gpio_defaults_block_32/gpio_defaults [10],
    \gpio_defaults_block_32/gpio_defaults [9],
    \gpio_defaults_block_32/gpio_defaults [8],
    \gpio_defaults_block_32/gpio_defaults [7],
    \gpio_defaults_block_32/gpio_defaults [6],
    \gpio_defaults_block_32/gpio_defaults [5],
    \gpio_defaults_block_32/gpio_defaults [4],
    \gpio_defaults_block_32/gpio_defaults [3],
    \gpio_defaults_block_32/gpio_defaults [2],
    \gpio_defaults_block_32/gpio_defaults [1],
    \gpio_defaults_block_32/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1a[5]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [7]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[5]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [7]),
    .one(\gpio_control_in_1a[5]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [7]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [7]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [7]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [7]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [7]),
    .pad_gpio_in(\padframe/mprj_io_in [7]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [7]),
    .pad_gpio_out(\padframe/mprj_io_out [7]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [7]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [7]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [7]),
    .resetn(\gpio_control_in_1a[5]/resetn ),
    .resetn_out(\gpio_control_in_1[0]/resetn ),
    .serial_clock(\gpio_control_in_1a[5]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[0]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[5]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[0]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[5]/serial_load ),
    .serial_load_out(\gpio_control_in_1[0]/serial_load ),
    .user_gpio_in(\mprj/io_in [7]),
    .user_gpio_oeb(\mprj/io_oeb [7]),
    .user_gpio_out(\mprj/io_out [7]),
    .zero(\gpio_control_in_1a[5]/zero ),
    .gpio_defaults({\gpio_defaults_block_7/gpio_defaults [12],
    \gpio_defaults_block_7/gpio_defaults [11],
    \gpio_defaults_block_7/gpio_defaults [10],
    \gpio_defaults_block_7/gpio_defaults [9],
    \gpio_defaults_block_7/gpio_defaults [8],
    \gpio_defaults_block_7/gpio_defaults [7],
    \gpio_defaults_block_7/gpio_defaults [6],
    \gpio_defaults_block_7/gpio_defaults [5],
    \gpio_defaults_block_7/gpio_defaults [4],
    \gpio_defaults_block_7/gpio_defaults [3],
    \gpio_defaults_block_7/gpio_defaults [2],
    \gpio_defaults_block_7/gpio_defaults [1],
    \gpio_defaults_block_7/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [23],
    \padframe/mprj_io_dm [22],
    \padframe/mprj_io_dm [21]}));
 gpio_control_block \gpio_control_in_1a[4]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [6]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[4]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [6]),
    .one(\gpio_control_in_1a[4]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [6]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [6]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [6]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [6]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [6]),
    .pad_gpio_in(\padframe/mprj_io_in [6]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [6]),
    .pad_gpio_out(\padframe/mprj_io_out [6]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [6]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [6]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [6]),
    .resetn(\gpio_control_in_1a[4]/resetn ),
    .resetn_out(\gpio_control_in_1a[5]/resetn ),
    .serial_clock(\gpio_control_in_1a[4]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[5]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[4]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[5]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[4]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[5]/serial_load ),
    .user_gpio_in(\mprj/io_in [6]),
    .user_gpio_oeb(\mprj/io_oeb [6]),
    .user_gpio_out(\mprj/io_out [6]),
    .zero(\gpio_control_in_1a[4]/zero ),
    .gpio_defaults({\gpio_defaults_block_6/gpio_defaults [12],
    \gpio_defaults_block_6/gpio_defaults [11],
    \gpio_defaults_block_6/gpio_defaults [10],
    \gpio_defaults_block_6/gpio_defaults [9],
    \gpio_defaults_block_6/gpio_defaults [8],
    \gpio_defaults_block_6/gpio_defaults [7],
    \gpio_defaults_block_6/gpio_defaults [6],
    \gpio_defaults_block_6/gpio_defaults [5],
    \gpio_defaults_block_6/gpio_defaults [4],
    \gpio_defaults_block_6/gpio_defaults [3],
    \gpio_defaults_block_6/gpio_defaults [2],
    \gpio_defaults_block_6/gpio_defaults [1],
    \gpio_defaults_block_6/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [20],
    \padframe/mprj_io_dm [19],
    \padframe/mprj_io_dm [18]}));
 gpio_control_block \gpio_control_in_1a[3]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [5]),
    .mgmt_gpio_oeb(\gpio_control_in_1a[3]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [5]),
    .one(\gpio_control_in_1a[3]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [5]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [5]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [5]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [5]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [5]),
    .pad_gpio_in(\padframe/mprj_io_in [5]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [5]),
    .pad_gpio_out(\padframe/mprj_io_out [5]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [5]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [5]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [5]),
    .resetn(\gpio_control_in_1a[3]/resetn ),
    .resetn_out(\gpio_control_in_1a[4]/resetn ),
    .serial_clock(\gpio_control_in_1a[3]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1a[4]/serial_clock ),
    .serial_data_in(\gpio_control_in_1a[3]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1a[4]/serial_data_in ),
    .serial_load(\gpio_control_in_1a[3]/serial_load ),
    .serial_load_out(\gpio_control_in_1a[4]/serial_load ),
    .user_gpio_in(\mprj/io_in [5]),
    .user_gpio_oeb(\mprj/io_oeb [5]),
    .user_gpio_out(\mprj/io_out [5]),
    .zero(\gpio_control_in_1a[3]/zero ),
    .gpio_defaults({\gpio_defaults_block_5/gpio_defaults [12],
    \gpio_defaults_block_5/gpio_defaults [11],
    \gpio_defaults_block_5/gpio_defaults [10],
    \gpio_defaults_block_5/gpio_defaults [9],
    \gpio_defaults_block_5/gpio_defaults [8],
    \gpio_defaults_block_5/gpio_defaults [7],
    \gpio_defaults_block_5/gpio_defaults [6],
    \gpio_defaults_block_5/gpio_defaults [5],
    \gpio_defaults_block_5/gpio_defaults [4],
    \gpio_defaults_block_5/gpio_defaults [3],
    \gpio_defaults_block_5/gpio_defaults [2],
    \gpio_defaults_block_5/gpio_defaults [1],
    \gpio_defaults_block_5/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [17],
    \padframe/mprj_io_dm [16],
    \padframe/mprj_io_dm [15]}));
 gpio_defaults_block gpio_defaults_block_7 (.gpio_defaults({\gpio_defaults_block_7/gpio_defaults [12],
    \gpio_defaults_block_7/gpio_defaults [11],
    \gpio_defaults_block_7/gpio_defaults [10],
    \gpio_defaults_block_7/gpio_defaults [9],
    \gpio_defaults_block_7/gpio_defaults [8],
    \gpio_defaults_block_7/gpio_defaults [7],
    \gpio_defaults_block_7/gpio_defaults [6],
    \gpio_defaults_block_7/gpio_defaults [5],
    \gpio_defaults_block_7/gpio_defaults [4],
    \gpio_defaults_block_7/gpio_defaults [3],
    \gpio_defaults_block_7/gpio_defaults [2],
    \gpio_defaults_block_7/gpio_defaults [1],
    \gpio_defaults_block_7/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_5 (.gpio_defaults({\gpio_defaults_block_5/gpio_defaults [12],
    \gpio_defaults_block_5/gpio_defaults [11],
    \gpio_defaults_block_5/gpio_defaults [10],
    \gpio_defaults_block_5/gpio_defaults [9],
    \gpio_defaults_block_5/gpio_defaults [8],
    \gpio_defaults_block_5/gpio_defaults [7],
    \gpio_defaults_block_5/gpio_defaults [6],
    \gpio_defaults_block_5/gpio_defaults [5],
    \gpio_defaults_block_5/gpio_defaults [4],
    \gpio_defaults_block_5/gpio_defaults [3],
    \gpio_defaults_block_5/gpio_defaults [2],
    \gpio_defaults_block_5/gpio_defaults [1],
    \gpio_defaults_block_5/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_6 (.gpio_defaults({\gpio_defaults_block_6/gpio_defaults [12],
    \gpio_defaults_block_6/gpio_defaults [11],
    \gpio_defaults_block_6/gpio_defaults [10],
    \gpio_defaults_block_6/gpio_defaults [9],
    \gpio_defaults_block_6/gpio_defaults [8],
    \gpio_defaults_block_6/gpio_defaults [7],
    \gpio_defaults_block_6/gpio_defaults [6],
    \gpio_defaults_block_6/gpio_defaults [5],
    \gpio_defaults_block_6/gpio_defaults [4],
    \gpio_defaults_block_6/gpio_defaults [3],
    \gpio_defaults_block_6/gpio_defaults [2],
    \gpio_defaults_block_6/gpio_defaults [1],
    \gpio_defaults_block_6/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_30 (.gpio_defaults({\gpio_defaults_block_30/gpio_defaults [12],
    \gpio_defaults_block_30/gpio_defaults [11],
    \gpio_defaults_block_30/gpio_defaults [10],
    \gpio_defaults_block_30/gpio_defaults [9],
    \gpio_defaults_block_30/gpio_defaults [8],
    \gpio_defaults_block_30/gpio_defaults [7],
    \gpio_defaults_block_30/gpio_defaults [6],
    \gpio_defaults_block_30/gpio_defaults [5],
    \gpio_defaults_block_30/gpio_defaults [4],
    \gpio_defaults_block_30/gpio_defaults [3],
    \gpio_defaults_block_30/gpio_defaults [2],
    \gpio_defaults_block_30/gpio_defaults [1],
    \gpio_defaults_block_30/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_31 (.gpio_defaults({\gpio_defaults_block_31/gpio_defaults [12],
    \gpio_defaults_block_31/gpio_defaults [11],
    \gpio_defaults_block_31/gpio_defaults [10],
    \gpio_defaults_block_31/gpio_defaults [9],
    \gpio_defaults_block_31/gpio_defaults [8],
    \gpio_defaults_block_31/gpio_defaults [7],
    \gpio_defaults_block_31/gpio_defaults [6],
    \gpio_defaults_block_31/gpio_defaults [5],
    \gpio_defaults_block_31/gpio_defaults [4],
    \gpio_defaults_block_31/gpio_defaults [3],
    \gpio_defaults_block_31/gpio_defaults [2],
    \gpio_defaults_block_31/gpio_defaults [1],
    \gpio_defaults_block_31/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[12]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [31]),
    .mgmt_gpio_oeb(\gpio_control_in_2[12]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [31]),
    .one(\gpio_control_in_2[12]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [31]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [31]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [31]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [31]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [31]),
    .pad_gpio_in(\padframe/mprj_io_in [31]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [31]),
    .pad_gpio_out(\padframe/mprj_io_out [31]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [31]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [31]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [31]),
    .resetn(\gpio_control_in_2[12]/resetn ),
    .resetn_out(\gpio_control_in_2[11]/resetn ),
    .serial_clock(\gpio_control_in_2[12]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[11]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[12]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[11]/serial_data_in ),
    .serial_load(\gpio_control_in_2[12]/serial_load ),
    .serial_load_out(\gpio_control_in_2[11]/serial_load ),
    .user_gpio_in(\mprj/io_in [31]),
    .user_gpio_oeb(\mprj/io_oeb [31]),
    .user_gpio_out(\mprj/io_out [31]),
    .zero(\gpio_control_in_2[12]/zero ),
    .gpio_defaults({\gpio_defaults_block_31/gpio_defaults [12],
    \gpio_defaults_block_31/gpio_defaults [11],
    \gpio_defaults_block_31/gpio_defaults [10],
    \gpio_defaults_block_31/gpio_defaults [9],
    \gpio_defaults_block_31/gpio_defaults [8],
    \gpio_defaults_block_31/gpio_defaults [7],
    \gpio_defaults_block_31/gpio_defaults [6],
    \gpio_defaults_block_31/gpio_defaults [5],
    \gpio_defaults_block_31/gpio_defaults [4],
    \gpio_defaults_block_31/gpio_defaults [3],
    \gpio_defaults_block_31/gpio_defaults [2],
    \gpio_defaults_block_31/gpio_defaults [1],
    \gpio_defaults_block_31/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [95],
    \padframe/mprj_io_dm [94],
    \padframe/mprj_io_dm [93]}));
 gpio_control_block \gpio_control_in_2[11]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [30]),
    .mgmt_gpio_oeb(\gpio_control_in_2[11]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [30]),
    .one(\gpio_control_in_2[11]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [30]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [30]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [30]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [30]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [30]),
    .pad_gpio_in(\padframe/mprj_io_in [30]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [30]),
    .pad_gpio_out(\padframe/mprj_io_out [30]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [30]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [30]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [30]),
    .resetn(\gpio_control_in_2[11]/resetn ),
    .resetn_out(\gpio_control_in_2[10]/resetn ),
    .serial_clock(\gpio_control_in_2[11]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[10]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[11]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[10]/serial_data_in ),
    .serial_load(\gpio_control_in_2[11]/serial_load ),
    .serial_load_out(\gpio_control_in_2[10]/serial_load ),
    .user_gpio_in(\mprj/io_in [30]),
    .user_gpio_oeb(\mprj/io_oeb [30]),
    .user_gpio_out(\mprj/io_out [30]),
    .zero(\gpio_control_in_2[11]/zero ),
    .gpio_defaults({\gpio_defaults_block_30/gpio_defaults [12],
    \gpio_defaults_block_30/gpio_defaults [11],
    \gpio_defaults_block_30/gpio_defaults [10],
    \gpio_defaults_block_30/gpio_defaults [9],
    \gpio_defaults_block_30/gpio_defaults [8],
    \gpio_defaults_block_30/gpio_defaults [7],
    \gpio_defaults_block_30/gpio_defaults [6],
    \gpio_defaults_block_30/gpio_defaults [5],
    \gpio_defaults_block_30/gpio_defaults [4],
    \gpio_defaults_block_30/gpio_defaults [3],
    \gpio_defaults_block_30/gpio_defaults [2],
    \gpio_defaults_block_30/gpio_defaults [1],
    \gpio_defaults_block_30/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [92],
    \padframe/mprj_io_dm [91],
    \padframe/mprj_io_dm [90]}));
 gpio_defaults_block gpio_defaults_block_9 (.gpio_defaults({\gpio_defaults_block_9/gpio_defaults [12],
    \gpio_defaults_block_9/gpio_defaults [11],
    \gpio_defaults_block_9/gpio_defaults [10],
    \gpio_defaults_block_9/gpio_defaults [9],
    \gpio_defaults_block_9/gpio_defaults [8],
    \gpio_defaults_block_9/gpio_defaults [7],
    \gpio_defaults_block_9/gpio_defaults [6],
    \gpio_defaults_block_9/gpio_defaults [5],
    \gpio_defaults_block_9/gpio_defaults [4],
    \gpio_defaults_block_9/gpio_defaults [3],
    \gpio_defaults_block_9/gpio_defaults [2],
    \gpio_defaults_block_9/gpio_defaults [1],
    \gpio_defaults_block_9/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_8 (.gpio_defaults({\gpio_defaults_block_8/gpio_defaults [12],
    \gpio_defaults_block_8/gpio_defaults [11],
    \gpio_defaults_block_8/gpio_defaults [10],
    \gpio_defaults_block_8/gpio_defaults [9],
    \gpio_defaults_block_8/gpio_defaults [8],
    \gpio_defaults_block_8/gpio_defaults [7],
    \gpio_defaults_block_8/gpio_defaults [6],
    \gpio_defaults_block_8/gpio_defaults [5],
    \gpio_defaults_block_8/gpio_defaults [4],
    \gpio_defaults_block_8/gpio_defaults [3],
    \gpio_defaults_block_8/gpio_defaults [2],
    \gpio_defaults_block_8/gpio_defaults [1],
    \gpio_defaults_block_8/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[1]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [9]),
    .mgmt_gpio_oeb(\gpio_control_in_1[1]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [9]),
    .one(\gpio_control_in_1[1]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [9]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [9]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [9]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [9]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [9]),
    .pad_gpio_in(\padframe/mprj_io_in [9]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [9]),
    .pad_gpio_out(\padframe/mprj_io_out [9]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [9]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [9]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [9]),
    .resetn(\gpio_control_in_1[1]/resetn ),
    .resetn_out(\gpio_control_in_1[2]/resetn ),
    .serial_clock(\gpio_control_in_1[1]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[2]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[1]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[2]/serial_data_in ),
    .serial_load(\gpio_control_in_1[1]/serial_load ),
    .serial_load_out(\gpio_control_in_1[2]/serial_load ),
    .user_gpio_in(\mprj/io_in [9]),
    .user_gpio_oeb(\mprj/io_oeb [9]),
    .user_gpio_out(\mprj/io_out [9]),
    .zero(\gpio_control_in_1[1]/zero ),
    .gpio_defaults({\gpio_defaults_block_9/gpio_defaults [12],
    \gpio_defaults_block_9/gpio_defaults [11],
    \gpio_defaults_block_9/gpio_defaults [10],
    \gpio_defaults_block_9/gpio_defaults [9],
    \gpio_defaults_block_9/gpio_defaults [8],
    \gpio_defaults_block_9/gpio_defaults [7],
    \gpio_defaults_block_9/gpio_defaults [6],
    \gpio_defaults_block_9/gpio_defaults [5],
    \gpio_defaults_block_9/gpio_defaults [4],
    \gpio_defaults_block_9/gpio_defaults [3],
    \gpio_defaults_block_9/gpio_defaults [2],
    \gpio_defaults_block_9/gpio_defaults [1],
    \gpio_defaults_block_9/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [29],
    \padframe/mprj_io_dm [28],
    \padframe/mprj_io_dm [27]}));
 gpio_control_block \gpio_control_in_1[0]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [8]),
    .mgmt_gpio_oeb(\gpio_control_in_1[0]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [8]),
    .one(\gpio_control_in_1[0]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [8]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [8]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [8]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [8]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [8]),
    .pad_gpio_in(\padframe/mprj_io_in [8]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [8]),
    .pad_gpio_out(\padframe/mprj_io_out [8]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [8]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [8]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [8]),
    .resetn(\gpio_control_in_1[0]/resetn ),
    .resetn_out(\gpio_control_in_1[1]/resetn ),
    .serial_clock(\gpio_control_in_1[0]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[1]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[0]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[1]/serial_data_in ),
    .serial_load(\gpio_control_in_1[0]/serial_load ),
    .serial_load_out(\gpio_control_in_1[1]/serial_load ),
    .user_gpio_in(\mprj/io_in [8]),
    .user_gpio_oeb(\mprj/io_oeb [8]),
    .user_gpio_out(\mprj/io_out [8]),
    .zero(\gpio_control_in_1[0]/zero ),
    .gpio_defaults({\gpio_defaults_block_8/gpio_defaults [12],
    \gpio_defaults_block_8/gpio_defaults [11],
    \gpio_defaults_block_8/gpio_defaults [10],
    \gpio_defaults_block_8/gpio_defaults [9],
    \gpio_defaults_block_8/gpio_defaults [8],
    \gpio_defaults_block_8/gpio_defaults [7],
    \gpio_defaults_block_8/gpio_defaults [6],
    \gpio_defaults_block_8/gpio_defaults [5],
    \gpio_defaults_block_8/gpio_defaults [4],
    \gpio_defaults_block_8/gpio_defaults [3],
    \gpio_defaults_block_8/gpio_defaults [2],
    \gpio_defaults_block_8/gpio_defaults [1],
    \gpio_defaults_block_8/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [26],
    \padframe/mprj_io_dm [25],
    \padframe/mprj_io_dm [24]}));
 gpio_defaults_block gpio_defaults_block_28 (.gpio_defaults({\gpio_defaults_block_28/gpio_defaults [12],
    \gpio_defaults_block_28/gpio_defaults [11],
    \gpio_defaults_block_28/gpio_defaults [10],
    \gpio_defaults_block_28/gpio_defaults [9],
    \gpio_defaults_block_28/gpio_defaults [8],
    \gpio_defaults_block_28/gpio_defaults [7],
    \gpio_defaults_block_28/gpio_defaults [6],
    \gpio_defaults_block_28/gpio_defaults [5],
    \gpio_defaults_block_28/gpio_defaults [4],
    \gpio_defaults_block_28/gpio_defaults [3],
    \gpio_defaults_block_28/gpio_defaults [2],
    \gpio_defaults_block_28/gpio_defaults [1],
    \gpio_defaults_block_28/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_29 (.gpio_defaults({\gpio_defaults_block_29/gpio_defaults [12],
    \gpio_defaults_block_29/gpio_defaults [11],
    \gpio_defaults_block_29/gpio_defaults [10],
    \gpio_defaults_block_29/gpio_defaults [9],
    \gpio_defaults_block_29/gpio_defaults [8],
    \gpio_defaults_block_29/gpio_defaults [7],
    \gpio_defaults_block_29/gpio_defaults [6],
    \gpio_defaults_block_29/gpio_defaults [5],
    \gpio_defaults_block_29/gpio_defaults [4],
    \gpio_defaults_block_29/gpio_defaults [3],
    \gpio_defaults_block_29/gpio_defaults [2],
    \gpio_defaults_block_29/gpio_defaults [1],
    \gpio_defaults_block_29/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[9]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [28]),
    .mgmt_gpio_oeb(\gpio_control_in_2[9]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [28]),
    .one(\gpio_control_in_2[9]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [28]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [28]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [28]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [28]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [28]),
    .pad_gpio_in(\padframe/mprj_io_in [28]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [28]),
    .pad_gpio_out(\padframe/mprj_io_out [28]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [28]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [28]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [28]),
    .resetn(\gpio_control_in_2[9]/resetn ),
    .resetn_out(\gpio_control_in_2[8]/resetn ),
    .serial_clock(\gpio_control_in_2[9]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[8]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[9]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[8]/serial_data_in ),
    .serial_load(\gpio_control_in_2[9]/serial_load ),
    .serial_load_out(\gpio_control_in_2[8]/serial_load ),
    .user_gpio_in(\mprj/io_in [28]),
    .user_gpio_oeb(\mprj/io_oeb [28]),
    .user_gpio_out(\mprj/io_out [28]),
    .zero(\gpio_control_in_2[9]/zero ),
    .gpio_defaults({\gpio_defaults_block_28/gpio_defaults [12],
    \gpio_defaults_block_28/gpio_defaults [11],
    \gpio_defaults_block_28/gpio_defaults [10],
    \gpio_defaults_block_28/gpio_defaults [9],
    \gpio_defaults_block_28/gpio_defaults [8],
    \gpio_defaults_block_28/gpio_defaults [7],
    \gpio_defaults_block_28/gpio_defaults [6],
    \gpio_defaults_block_28/gpio_defaults [5],
    \gpio_defaults_block_28/gpio_defaults [4],
    \gpio_defaults_block_28/gpio_defaults [3],
    \gpio_defaults_block_28/gpio_defaults [2],
    \gpio_defaults_block_28/gpio_defaults [1],
    \gpio_defaults_block_28/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [86],
    \padframe/mprj_io_dm [85],
    \padframe/mprj_io_dm [84]}));
 gpio_control_block \gpio_control_in_2[10]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [29]),
    .mgmt_gpio_oeb(\gpio_control_in_2[10]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [29]),
    .one(\gpio_control_in_2[10]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [29]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [29]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [29]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [29]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [29]),
    .pad_gpio_in(\padframe/mprj_io_in [29]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [29]),
    .pad_gpio_out(\padframe/mprj_io_out [29]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [29]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [29]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [29]),
    .resetn(\gpio_control_in_2[10]/resetn ),
    .resetn_out(\gpio_control_in_2[9]/resetn ),
    .serial_clock(\gpio_control_in_2[10]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[9]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[10]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[9]/serial_data_in ),
    .serial_load(\gpio_control_in_2[10]/serial_load ),
    .serial_load_out(\gpio_control_in_2[9]/serial_load ),
    .user_gpio_in(\mprj/io_in [29]),
    .user_gpio_oeb(\mprj/io_oeb [29]),
    .user_gpio_out(\mprj/io_out [29]),
    .zero(\gpio_control_in_2[10]/zero ),
    .gpio_defaults({\gpio_defaults_block_29/gpio_defaults [12],
    \gpio_defaults_block_29/gpio_defaults [11],
    \gpio_defaults_block_29/gpio_defaults [10],
    \gpio_defaults_block_29/gpio_defaults [9],
    \gpio_defaults_block_29/gpio_defaults [8],
    \gpio_defaults_block_29/gpio_defaults [7],
    \gpio_defaults_block_29/gpio_defaults [6],
    \gpio_defaults_block_29/gpio_defaults [5],
    \gpio_defaults_block_29/gpio_defaults [4],
    \gpio_defaults_block_29/gpio_defaults [3],
    \gpio_defaults_block_29/gpio_defaults [2],
    \gpio_defaults_block_29/gpio_defaults [1],
    \gpio_defaults_block_29/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [89],
    \padframe/mprj_io_dm [88],
    \padframe/mprj_io_dm [87]}));
 gpio_defaults_block gpio_defaults_block_11 (.gpio_defaults({\gpio_defaults_block_11/gpio_defaults [12],
    \gpio_defaults_block_11/gpio_defaults [11],
    \gpio_defaults_block_11/gpio_defaults [10],
    \gpio_defaults_block_11/gpio_defaults [9],
    \gpio_defaults_block_11/gpio_defaults [8],
    \gpio_defaults_block_11/gpio_defaults [7],
    \gpio_defaults_block_11/gpio_defaults [6],
    \gpio_defaults_block_11/gpio_defaults [5],
    \gpio_defaults_block_11/gpio_defaults [4],
    \gpio_defaults_block_11/gpio_defaults [3],
    \gpio_defaults_block_11/gpio_defaults [2],
    \gpio_defaults_block_11/gpio_defaults [1],
    \gpio_defaults_block_11/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_10 (.gpio_defaults({\gpio_defaults_block_10/gpio_defaults [12],
    \gpio_defaults_block_10/gpio_defaults [11],
    \gpio_defaults_block_10/gpio_defaults [10],
    \gpio_defaults_block_10/gpio_defaults [9],
    \gpio_defaults_block_10/gpio_defaults [8],
    \gpio_defaults_block_10/gpio_defaults [7],
    \gpio_defaults_block_10/gpio_defaults [6],
    \gpio_defaults_block_10/gpio_defaults [5],
    \gpio_defaults_block_10/gpio_defaults [4],
    \gpio_defaults_block_10/gpio_defaults [3],
    \gpio_defaults_block_10/gpio_defaults [2],
    \gpio_defaults_block_10/gpio_defaults [1],
    \gpio_defaults_block_10/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[3]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [11]),
    .mgmt_gpio_oeb(\gpio_control_in_1[3]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [11]),
    .one(\gpio_control_in_1[3]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [11]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [11]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [11]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [11]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [11]),
    .pad_gpio_in(\padframe/mprj_io_in [11]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [11]),
    .pad_gpio_out(\padframe/mprj_io_out [11]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [11]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [11]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [11]),
    .resetn(\gpio_control_in_1[3]/resetn ),
    .resetn_out(\gpio_control_in_1[4]/resetn ),
    .serial_clock(\gpio_control_in_1[3]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[4]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[3]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[4]/serial_data_in ),
    .serial_load(\gpio_control_in_1[3]/serial_load ),
    .serial_load_out(\gpio_control_in_1[4]/serial_load ),
    .user_gpio_in(\mprj/io_in [11]),
    .user_gpio_oeb(\mprj/io_oeb [11]),
    .user_gpio_out(\mprj/io_out [11]),
    .zero(\gpio_control_in_1[3]/zero ),
    .gpio_defaults({\gpio_defaults_block_11/gpio_defaults [12],
    \gpio_defaults_block_11/gpio_defaults [11],
    \gpio_defaults_block_11/gpio_defaults [10],
    \gpio_defaults_block_11/gpio_defaults [9],
    \gpio_defaults_block_11/gpio_defaults [8],
    \gpio_defaults_block_11/gpio_defaults [7],
    \gpio_defaults_block_11/gpio_defaults [6],
    \gpio_defaults_block_11/gpio_defaults [5],
    \gpio_defaults_block_11/gpio_defaults [4],
    \gpio_defaults_block_11/gpio_defaults [3],
    \gpio_defaults_block_11/gpio_defaults [2],
    \gpio_defaults_block_11/gpio_defaults [1],
    \gpio_defaults_block_11/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [35],
    \padframe/mprj_io_dm [34],
    \padframe/mprj_io_dm [33]}));
 gpio_control_block \gpio_control_in_1[2]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [10]),
    .mgmt_gpio_oeb(\gpio_control_in_1[2]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [10]),
    .one(\gpio_control_in_1[2]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [10]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [10]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [10]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [10]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [10]),
    .pad_gpio_in(\padframe/mprj_io_in [10]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [10]),
    .pad_gpio_out(\padframe/mprj_io_out [10]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [10]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [10]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [10]),
    .resetn(\gpio_control_in_1[2]/resetn ),
    .resetn_out(\gpio_control_in_1[3]/resetn ),
    .serial_clock(\gpio_control_in_1[2]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[3]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[2]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[3]/serial_data_in ),
    .serial_load(\gpio_control_in_1[2]/serial_load ),
    .serial_load_out(\gpio_control_in_1[3]/serial_load ),
    .user_gpio_in(\mprj/io_in [10]),
    .user_gpio_oeb(\mprj/io_oeb [10]),
    .user_gpio_out(\mprj/io_out [10]),
    .zero(\gpio_control_in_1[2]/zero ),
    .gpio_defaults({\gpio_defaults_block_10/gpio_defaults [12],
    \gpio_defaults_block_10/gpio_defaults [11],
    \gpio_defaults_block_10/gpio_defaults [10],
    \gpio_defaults_block_10/gpio_defaults [9],
    \gpio_defaults_block_10/gpio_defaults [8],
    \gpio_defaults_block_10/gpio_defaults [7],
    \gpio_defaults_block_10/gpio_defaults [6],
    \gpio_defaults_block_10/gpio_defaults [5],
    \gpio_defaults_block_10/gpio_defaults [4],
    \gpio_defaults_block_10/gpio_defaults [3],
    \gpio_defaults_block_10/gpio_defaults [2],
    \gpio_defaults_block_10/gpio_defaults [1],
    \gpio_defaults_block_10/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [32],
    \padframe/mprj_io_dm [31],
    \padframe/mprj_io_dm [30]}));
 gpio_defaults_block gpio_defaults_block_26 (.gpio_defaults({\gpio_defaults_block_26/gpio_defaults [12],
    \gpio_defaults_block_26/gpio_defaults [11],
    \gpio_defaults_block_26/gpio_defaults [10],
    \gpio_defaults_block_26/gpio_defaults [9],
    \gpio_defaults_block_26/gpio_defaults [8],
    \gpio_defaults_block_26/gpio_defaults [7],
    \gpio_defaults_block_26/gpio_defaults [6],
    \gpio_defaults_block_26/gpio_defaults [5],
    \gpio_defaults_block_26/gpio_defaults [4],
    \gpio_defaults_block_26/gpio_defaults [3],
    \gpio_defaults_block_26/gpio_defaults [2],
    \gpio_defaults_block_26/gpio_defaults [1],
    \gpio_defaults_block_26/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_27 (.gpio_defaults({\gpio_defaults_block_27/gpio_defaults [12],
    \gpio_defaults_block_27/gpio_defaults [11],
    \gpio_defaults_block_27/gpio_defaults [10],
    \gpio_defaults_block_27/gpio_defaults [9],
    \gpio_defaults_block_27/gpio_defaults [8],
    \gpio_defaults_block_27/gpio_defaults [7],
    \gpio_defaults_block_27/gpio_defaults [6],
    \gpio_defaults_block_27/gpio_defaults [5],
    \gpio_defaults_block_27/gpio_defaults [4],
    \gpio_defaults_block_27/gpio_defaults [3],
    \gpio_defaults_block_27/gpio_defaults [2],
    \gpio_defaults_block_27/gpio_defaults [1],
    \gpio_defaults_block_27/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[8]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [27]),
    .mgmt_gpio_oeb(\gpio_control_in_2[8]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [27]),
    .one(\gpio_control_in_2[8]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [27]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [27]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [27]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [27]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [27]),
    .pad_gpio_in(\padframe/mprj_io_in [27]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [27]),
    .pad_gpio_out(\padframe/mprj_io_out [27]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [27]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [27]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [27]),
    .resetn(\gpio_control_in_2[8]/resetn ),
    .resetn_out(\gpio_control_in_2[7]/resetn ),
    .serial_clock(\gpio_control_in_2[8]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[7]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[8]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[7]/serial_data_in ),
    .serial_load(\gpio_control_in_2[8]/serial_load ),
    .serial_load_out(\gpio_control_in_2[7]/serial_load ),
    .user_gpio_in(\mprj/io_in [27]),
    .user_gpio_oeb(\mprj/io_oeb [27]),
    .user_gpio_out(\mprj/io_out [27]),
    .zero(\gpio_control_in_2[8]/zero ),
    .gpio_defaults({\gpio_defaults_block_27/gpio_defaults [12],
    \gpio_defaults_block_27/gpio_defaults [11],
    \gpio_defaults_block_27/gpio_defaults [10],
    \gpio_defaults_block_27/gpio_defaults [9],
    \gpio_defaults_block_27/gpio_defaults [8],
    \gpio_defaults_block_27/gpio_defaults [7],
    \gpio_defaults_block_27/gpio_defaults [6],
    \gpio_defaults_block_27/gpio_defaults [5],
    \gpio_defaults_block_27/gpio_defaults [4],
    \gpio_defaults_block_27/gpio_defaults [3],
    \gpio_defaults_block_27/gpio_defaults [2],
    \gpio_defaults_block_27/gpio_defaults [1],
    \gpio_defaults_block_27/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [83],
    \padframe/mprj_io_dm [82],
    \padframe/mprj_io_dm [81]}));
 gpio_control_block \gpio_control_in_2[7]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [26]),
    .mgmt_gpio_oeb(\gpio_control_in_2[7]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [26]),
    .one(\gpio_control_in_2[7]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [26]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [26]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [26]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [26]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [26]),
    .pad_gpio_in(\padframe/mprj_io_in [26]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [26]),
    .pad_gpio_out(\padframe/mprj_io_out [26]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [26]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [26]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [26]),
    .resetn(\gpio_control_in_2[7]/resetn ),
    .resetn_out(\gpio_control_in_2[6]/resetn ),
    .serial_clock(\gpio_control_in_2[7]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[6]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[7]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[6]/serial_data_in ),
    .serial_load(\gpio_control_in_2[7]/serial_load ),
    .serial_load_out(\gpio_control_in_2[6]/serial_load ),
    .user_gpio_in(\mprj/io_in [26]),
    .user_gpio_oeb(\mprj/io_oeb [26]),
    .user_gpio_out(\mprj/io_out [26]),
    .zero(\gpio_control_in_2[7]/zero ),
    .gpio_defaults({\gpio_defaults_block_26/gpio_defaults [12],
    \gpio_defaults_block_26/gpio_defaults [11],
    \gpio_defaults_block_26/gpio_defaults [10],
    \gpio_defaults_block_26/gpio_defaults [9],
    \gpio_defaults_block_26/gpio_defaults [8],
    \gpio_defaults_block_26/gpio_defaults [7],
    \gpio_defaults_block_26/gpio_defaults [6],
    \gpio_defaults_block_26/gpio_defaults [5],
    \gpio_defaults_block_26/gpio_defaults [4],
    \gpio_defaults_block_26/gpio_defaults [3],
    \gpio_defaults_block_26/gpio_defaults [2],
    \gpio_defaults_block_26/gpio_defaults [1],
    \gpio_defaults_block_26/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [80],
    \padframe/mprj_io_dm [79],
    \padframe/mprj_io_dm [78]}));
 gpio_defaults_block gpio_defaults_block_13 (.gpio_defaults({\gpio_defaults_block_13/gpio_defaults [12],
    \gpio_defaults_block_13/gpio_defaults [11],
    \gpio_defaults_block_13/gpio_defaults [10],
    \gpio_defaults_block_13/gpio_defaults [9],
    \gpio_defaults_block_13/gpio_defaults [8],
    \gpio_defaults_block_13/gpio_defaults [7],
    \gpio_defaults_block_13/gpio_defaults [6],
    \gpio_defaults_block_13/gpio_defaults [5],
    \gpio_defaults_block_13/gpio_defaults [4],
    \gpio_defaults_block_13/gpio_defaults [3],
    \gpio_defaults_block_13/gpio_defaults [2],
    \gpio_defaults_block_13/gpio_defaults [1],
    \gpio_defaults_block_13/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_12 (.gpio_defaults({\gpio_defaults_block_12/gpio_defaults [12],
    \gpio_defaults_block_12/gpio_defaults [11],
    \gpio_defaults_block_12/gpio_defaults [10],
    \gpio_defaults_block_12/gpio_defaults [9],
    \gpio_defaults_block_12/gpio_defaults [8],
    \gpio_defaults_block_12/gpio_defaults [7],
    \gpio_defaults_block_12/gpio_defaults [6],
    \gpio_defaults_block_12/gpio_defaults [5],
    \gpio_defaults_block_12/gpio_defaults [4],
    \gpio_defaults_block_12/gpio_defaults [3],
    \gpio_defaults_block_12/gpio_defaults [2],
    \gpio_defaults_block_12/gpio_defaults [1],
    \gpio_defaults_block_12/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[5]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [13]),
    .mgmt_gpio_oeb(\gpio_control_in_1[5]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [13]),
    .one(\gpio_control_in_1[5]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [13]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [13]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [13]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [13]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [13]),
    .pad_gpio_in(\padframe/mprj_io_in [13]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [13]),
    .pad_gpio_out(\padframe/mprj_io_out [13]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [13]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [13]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [13]),
    .resetn(\gpio_control_in_1[5]/resetn ),
    .resetn_out(\gpio_control_in_1[6]/resetn ),
    .serial_clock(\gpio_control_in_1[5]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[6]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[5]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[6]/serial_data_in ),
    .serial_load(\gpio_control_in_1[5]/serial_load ),
    .serial_load_out(\gpio_control_in_1[6]/serial_load ),
    .user_gpio_in(\mprj/io_in [13]),
    .user_gpio_oeb(\mprj/io_oeb [13]),
    .user_gpio_out(\mprj/io_out [13]),
    .zero(\gpio_control_in_1[5]/zero ),
    .gpio_defaults({\gpio_defaults_block_13/gpio_defaults [12],
    \gpio_defaults_block_13/gpio_defaults [11],
    \gpio_defaults_block_13/gpio_defaults [10],
    \gpio_defaults_block_13/gpio_defaults [9],
    \gpio_defaults_block_13/gpio_defaults [8],
    \gpio_defaults_block_13/gpio_defaults [7],
    \gpio_defaults_block_13/gpio_defaults [6],
    \gpio_defaults_block_13/gpio_defaults [5],
    \gpio_defaults_block_13/gpio_defaults [4],
    \gpio_defaults_block_13/gpio_defaults [3],
    \gpio_defaults_block_13/gpio_defaults [2],
    \gpio_defaults_block_13/gpio_defaults [1],
    \gpio_defaults_block_13/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [41],
    \padframe/mprj_io_dm [40],
    \padframe/mprj_io_dm [39]}));
 gpio_control_block \gpio_control_in_1[4]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [12]),
    .mgmt_gpio_oeb(\gpio_control_in_1[4]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [12]),
    .one(\gpio_control_in_1[4]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [12]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [12]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [12]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [12]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [12]),
    .pad_gpio_in(\padframe/mprj_io_in [12]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [12]),
    .pad_gpio_out(\padframe/mprj_io_out [12]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [12]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [12]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [12]),
    .resetn(\gpio_control_in_1[4]/resetn ),
    .resetn_out(\gpio_control_in_1[5]/resetn ),
    .serial_clock(\gpio_control_in_1[4]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[5]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[4]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[5]/serial_data_in ),
    .serial_load(\gpio_control_in_1[4]/serial_load ),
    .serial_load_out(\gpio_control_in_1[5]/serial_load ),
    .user_gpio_in(\mprj/io_in [12]),
    .user_gpio_oeb(\mprj/io_oeb [12]),
    .user_gpio_out(\mprj/io_out [12]),
    .zero(\gpio_control_in_1[4]/zero ),
    .gpio_defaults({\gpio_defaults_block_12/gpio_defaults [12],
    \gpio_defaults_block_12/gpio_defaults [11],
    \gpio_defaults_block_12/gpio_defaults [10],
    \gpio_defaults_block_12/gpio_defaults [9],
    \gpio_defaults_block_12/gpio_defaults [8],
    \gpio_defaults_block_12/gpio_defaults [7],
    \gpio_defaults_block_12/gpio_defaults [6],
    \gpio_defaults_block_12/gpio_defaults [5],
    \gpio_defaults_block_12/gpio_defaults [4],
    \gpio_defaults_block_12/gpio_defaults [3],
    \gpio_defaults_block_12/gpio_defaults [2],
    \gpio_defaults_block_12/gpio_defaults [1],
    \gpio_defaults_block_12/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [38],
    \padframe/mprj_io_dm [37],
    \padframe/mprj_io_dm [36]}));
 gpio_defaults_block gpio_defaults_block_25 (.gpio_defaults({\gpio_defaults_block_25/gpio_defaults [12],
    \gpio_defaults_block_25/gpio_defaults [11],
    \gpio_defaults_block_25/gpio_defaults [10],
    \gpio_defaults_block_25/gpio_defaults [9],
    \gpio_defaults_block_25/gpio_defaults [8],
    \gpio_defaults_block_25/gpio_defaults [7],
    \gpio_defaults_block_25/gpio_defaults [6],
    \gpio_defaults_block_25/gpio_defaults [5],
    \gpio_defaults_block_25/gpio_defaults [4],
    \gpio_defaults_block_25/gpio_defaults [3],
    \gpio_defaults_block_25/gpio_defaults [2],
    \gpio_defaults_block_25/gpio_defaults [1],
    \gpio_defaults_block_25/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[6]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [25]),
    .mgmt_gpio_oeb(\gpio_control_in_2[6]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [25]),
    .one(\gpio_control_in_2[6]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [25]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [25]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [25]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [25]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [25]),
    .pad_gpio_in(\padframe/mprj_io_in [25]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [25]),
    .pad_gpio_out(\padframe/mprj_io_out [25]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [25]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [25]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [25]),
    .resetn(\gpio_control_in_2[6]/resetn ),
    .resetn_out(\gpio_control_in_2[5]/resetn ),
    .serial_clock(\gpio_control_in_2[6]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[5]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[6]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[5]/serial_data_in ),
    .serial_load(\gpio_control_in_2[6]/serial_load ),
    .serial_load_out(\gpio_control_in_2[5]/serial_load ),
    .user_gpio_in(\mprj/io_in [25]),
    .user_gpio_oeb(\mprj/io_oeb [25]),
    .user_gpio_out(\mprj/io_out [25]),
    .zero(\gpio_control_in_2[6]/zero ),
    .gpio_defaults({\gpio_defaults_block_25/gpio_defaults [12],
    \gpio_defaults_block_25/gpio_defaults [11],
    \gpio_defaults_block_25/gpio_defaults [10],
    \gpio_defaults_block_25/gpio_defaults [9],
    \gpio_defaults_block_25/gpio_defaults [8],
    \gpio_defaults_block_25/gpio_defaults [7],
    \gpio_defaults_block_25/gpio_defaults [6],
    \gpio_defaults_block_25/gpio_defaults [5],
    \gpio_defaults_block_25/gpio_defaults [4],
    \gpio_defaults_block_25/gpio_defaults [3],
    \gpio_defaults_block_25/gpio_defaults [2],
    \gpio_defaults_block_25/gpio_defaults [1],
    \gpio_defaults_block_25/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [77],
    \padframe/mprj_io_dm [76],
    \padframe/mprj_io_dm [75]}));
 gpio_defaults_block gpio_defaults_block_24 (.gpio_defaults({\gpio_defaults_block_24/gpio_defaults [12],
    \gpio_defaults_block_24/gpio_defaults [11],
    \gpio_defaults_block_24/gpio_defaults [10],
    \gpio_defaults_block_24/gpio_defaults [9],
    \gpio_defaults_block_24/gpio_defaults [8],
    \gpio_defaults_block_24/gpio_defaults [7],
    \gpio_defaults_block_24/gpio_defaults [6],
    \gpio_defaults_block_24/gpio_defaults [5],
    \gpio_defaults_block_24/gpio_defaults [4],
    \gpio_defaults_block_24/gpio_defaults [3],
    \gpio_defaults_block_24/gpio_defaults [2],
    \gpio_defaults_block_24/gpio_defaults [1],
    \gpio_defaults_block_24/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[5]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [24]),
    .mgmt_gpio_oeb(\gpio_control_in_2[5]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [24]),
    .one(\gpio_control_in_2[5]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [24]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [24]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [24]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [24]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [24]),
    .pad_gpio_in(\padframe/mprj_io_in [24]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [24]),
    .pad_gpio_out(\padframe/mprj_io_out [24]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [24]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [24]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [24]),
    .resetn(\gpio_control_in_2[5]/resetn ),
    .resetn_out(\gpio_control_in_2[4]/resetn ),
    .serial_clock(\gpio_control_in_2[5]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[4]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[5]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[4]/serial_data_in ),
    .serial_load(\gpio_control_in_2[5]/serial_load ),
    .serial_load_out(\gpio_control_in_2[4]/serial_load ),
    .user_gpio_in(\mprj/io_in [24]),
    .user_gpio_oeb(\mprj/io_oeb [24]),
    .user_gpio_out(\mprj/io_out [24]),
    .zero(\gpio_control_in_2[5]/zero ),
    .gpio_defaults({\gpio_defaults_block_24/gpio_defaults [12],
    \gpio_defaults_block_24/gpio_defaults [11],
    \gpio_defaults_block_24/gpio_defaults [10],
    \gpio_defaults_block_24/gpio_defaults [9],
    \gpio_defaults_block_24/gpio_defaults [8],
    \gpio_defaults_block_24/gpio_defaults [7],
    \gpio_defaults_block_24/gpio_defaults [6],
    \gpio_defaults_block_24/gpio_defaults [5],
    \gpio_defaults_block_24/gpio_defaults [4],
    \gpio_defaults_block_24/gpio_defaults [3],
    \gpio_defaults_block_24/gpio_defaults [2],
    \gpio_defaults_block_24/gpio_defaults [1],
    \gpio_defaults_block_24/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [74],
    \padframe/mprj_io_dm [73],
    \padframe/mprj_io_dm [72]}));
 gpio_defaults_block gpio_defaults_block_14 (.gpio_defaults({\gpio_defaults_block_14/gpio_defaults [12],
    \gpio_defaults_block_14/gpio_defaults [11],
    \gpio_defaults_block_14/gpio_defaults [10],
    \gpio_defaults_block_14/gpio_defaults [9],
    \gpio_defaults_block_14/gpio_defaults [8],
    \gpio_defaults_block_14/gpio_defaults [7],
    \gpio_defaults_block_14/gpio_defaults [6],
    \gpio_defaults_block_14/gpio_defaults [5],
    \gpio_defaults_block_14/gpio_defaults [4],
    \gpio_defaults_block_14/gpio_defaults [3],
    \gpio_defaults_block_14/gpio_defaults [2],
    \gpio_defaults_block_14/gpio_defaults [1],
    \gpio_defaults_block_14/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[6]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [14]),
    .mgmt_gpio_oeb(\gpio_control_in_1[6]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [14]),
    .one(\gpio_control_in_1[6]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [14]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [14]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [14]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [14]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [14]),
    .pad_gpio_in(\padframe/mprj_io_in [14]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [14]),
    .pad_gpio_out(\padframe/mprj_io_out [14]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [14]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [14]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [14]),
    .resetn(\gpio_control_in_1[6]/resetn ),
    .resetn_out(\gpio_control_in_1[7]/resetn ),
    .serial_clock(\gpio_control_in_1[6]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[7]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[6]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[7]/serial_data_in ),
    .serial_load(\gpio_control_in_1[6]/serial_load ),
    .serial_load_out(\gpio_control_in_1[7]/serial_load ),
    .user_gpio_in(\mprj/io_in [14]),
    .user_gpio_oeb(\mprj/io_oeb [14]),
    .user_gpio_out(\mprj/io_out [14]),
    .zero(\gpio_control_in_1[6]/zero ),
    .gpio_defaults({\gpio_defaults_block_14/gpio_defaults [12],
    \gpio_defaults_block_14/gpio_defaults [11],
    \gpio_defaults_block_14/gpio_defaults [10],
    \gpio_defaults_block_14/gpio_defaults [9],
    \gpio_defaults_block_14/gpio_defaults [8],
    \gpio_defaults_block_14/gpio_defaults [7],
    \gpio_defaults_block_14/gpio_defaults [6],
    \gpio_defaults_block_14/gpio_defaults [5],
    \gpio_defaults_block_14/gpio_defaults [4],
    \gpio_defaults_block_14/gpio_defaults [3],
    \gpio_defaults_block_14/gpio_defaults [2],
    \gpio_defaults_block_14/gpio_defaults [1],
    \gpio_defaults_block_14/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [44],
    \padframe/mprj_io_dm [43],
    \padframe/mprj_io_dm [42]}));
 gpio_defaults_block gpio_defaults_block_22 (.gpio_defaults({\gpio_defaults_block_22/gpio_defaults [12],
    \gpio_defaults_block_22/gpio_defaults [11],
    \gpio_defaults_block_22/gpio_defaults [10],
    \gpio_defaults_block_22/gpio_defaults [9],
    \gpio_defaults_block_22/gpio_defaults [8],
    \gpio_defaults_block_22/gpio_defaults [7],
    \gpio_defaults_block_22/gpio_defaults [6],
    \gpio_defaults_block_22/gpio_defaults [5],
    \gpio_defaults_block_22/gpio_defaults [4],
    \gpio_defaults_block_22/gpio_defaults [3],
    \gpio_defaults_block_22/gpio_defaults [2],
    \gpio_defaults_block_22/gpio_defaults [1],
    \gpio_defaults_block_22/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_23 (.gpio_defaults({\gpio_defaults_block_23/gpio_defaults [12],
    \gpio_defaults_block_23/gpio_defaults [11],
    \gpio_defaults_block_23/gpio_defaults [10],
    \gpio_defaults_block_23/gpio_defaults [9],
    \gpio_defaults_block_23/gpio_defaults [8],
    \gpio_defaults_block_23/gpio_defaults [7],
    \gpio_defaults_block_23/gpio_defaults [6],
    \gpio_defaults_block_23/gpio_defaults [5],
    \gpio_defaults_block_23/gpio_defaults [4],
    \gpio_defaults_block_23/gpio_defaults [3],
    \gpio_defaults_block_23/gpio_defaults [2],
    \gpio_defaults_block_23/gpio_defaults [1],
    \gpio_defaults_block_23/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[4]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [23]),
    .mgmt_gpio_oeb(\gpio_control_in_2[4]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [23]),
    .one(\gpio_control_in_2[4]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [23]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [23]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [23]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [23]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [23]),
    .pad_gpio_in(\padframe/mprj_io_in [23]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [23]),
    .pad_gpio_out(\padframe/mprj_io_out [23]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [23]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [23]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [23]),
    .resetn(\gpio_control_in_2[4]/resetn ),
    .resetn_out(\gpio_control_in_2[3]/resetn ),
    .serial_clock(\gpio_control_in_2[4]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[3]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[4]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[3]/serial_data_in ),
    .serial_load(\gpio_control_in_2[4]/serial_load ),
    .serial_load_out(\gpio_control_in_2[3]/serial_load ),
    .user_gpio_in(\mprj/io_in [23]),
    .user_gpio_oeb(\mprj/io_oeb [23]),
    .user_gpio_out(\mprj/io_out [23]),
    .zero(\gpio_control_in_2[4]/zero ),
    .gpio_defaults({\gpio_defaults_block_23/gpio_defaults [12],
    \gpio_defaults_block_23/gpio_defaults [11],
    \gpio_defaults_block_23/gpio_defaults [10],
    \gpio_defaults_block_23/gpio_defaults [9],
    \gpio_defaults_block_23/gpio_defaults [8],
    \gpio_defaults_block_23/gpio_defaults [7],
    \gpio_defaults_block_23/gpio_defaults [6],
    \gpio_defaults_block_23/gpio_defaults [5],
    \gpio_defaults_block_23/gpio_defaults [4],
    \gpio_defaults_block_23/gpio_defaults [3],
    \gpio_defaults_block_23/gpio_defaults [2],
    \gpio_defaults_block_23/gpio_defaults [1],
    \gpio_defaults_block_23/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [71],
    \padframe/mprj_io_dm [70],
    \padframe/mprj_io_dm [69]}));
 gpio_control_block \gpio_control_in_2[3]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [22]),
    .mgmt_gpio_oeb(\gpio_control_in_2[3]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [22]),
    .one(\gpio_control_in_2[3]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [22]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [22]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [22]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [22]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [22]),
    .pad_gpio_in(\padframe/mprj_io_in [22]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [22]),
    .pad_gpio_out(\padframe/mprj_io_out [22]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [22]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [22]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [22]),
    .resetn(\gpio_control_in_2[3]/resetn ),
    .resetn_out(\gpio_control_in_2[2]/resetn ),
    .serial_clock(\gpio_control_in_2[3]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[2]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[3]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[2]/serial_data_in ),
    .serial_load(\gpio_control_in_2[3]/serial_load ),
    .serial_load_out(\gpio_control_in_2[2]/serial_load ),
    .user_gpio_in(\mprj/io_in [22]),
    .user_gpio_oeb(\mprj/io_oeb [22]),
    .user_gpio_out(\mprj/io_out [22]),
    .zero(\gpio_control_in_2[3]/zero ),
    .gpio_defaults({\gpio_defaults_block_22/gpio_defaults [12],
    \gpio_defaults_block_22/gpio_defaults [11],
    \gpio_defaults_block_22/gpio_defaults [10],
    \gpio_defaults_block_22/gpio_defaults [9],
    \gpio_defaults_block_22/gpio_defaults [8],
    \gpio_defaults_block_22/gpio_defaults [7],
    \gpio_defaults_block_22/gpio_defaults [6],
    \gpio_defaults_block_22/gpio_defaults [5],
    \gpio_defaults_block_22/gpio_defaults [4],
    \gpio_defaults_block_22/gpio_defaults [3],
    \gpio_defaults_block_22/gpio_defaults [2],
    \gpio_defaults_block_22/gpio_defaults [1],
    \gpio_defaults_block_22/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [68],
    \padframe/mprj_io_dm [67],
    \padframe/mprj_io_dm [66]}));
 gpio_defaults_block gpio_defaults_block_21 (.gpio_defaults({\gpio_defaults_block_21/gpio_defaults [12],
    \gpio_defaults_block_21/gpio_defaults [11],
    \gpio_defaults_block_21/gpio_defaults [10],
    \gpio_defaults_block_21/gpio_defaults [9],
    \gpio_defaults_block_21/gpio_defaults [8],
    \gpio_defaults_block_21/gpio_defaults [7],
    \gpio_defaults_block_21/gpio_defaults [6],
    \gpio_defaults_block_21/gpio_defaults [5],
    \gpio_defaults_block_21/gpio_defaults [4],
    \gpio_defaults_block_21/gpio_defaults [3],
    \gpio_defaults_block_21/gpio_defaults [2],
    \gpio_defaults_block_21/gpio_defaults [1],
    \gpio_defaults_block_21/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[2]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [21]),
    .mgmt_gpio_oeb(\gpio_control_in_2[2]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [21]),
    .one(\gpio_control_in_2[2]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [21]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [21]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [21]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [21]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [21]),
    .pad_gpio_in(\padframe/mprj_io_in [21]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [21]),
    .pad_gpio_out(\padframe/mprj_io_out [21]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [21]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [21]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [21]),
    .resetn(\gpio_control_in_2[2]/resetn ),
    .resetn_out(\gpio_control_in_2[1]/resetn ),
    .serial_clock(\gpio_control_in_2[2]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[1]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[2]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[1]/serial_data_in ),
    .serial_load(\gpio_control_in_2[2]/serial_load ),
    .serial_load_out(\gpio_control_in_2[1]/serial_load ),
    .user_gpio_in(\mprj/io_in [21]),
    .user_gpio_oeb(\mprj/io_oeb [21]),
    .user_gpio_out(\mprj/io_out [21]),
    .zero(\gpio_control_in_2[2]/zero ),
    .gpio_defaults({\gpio_defaults_block_21/gpio_defaults [12],
    \gpio_defaults_block_21/gpio_defaults [11],
    \gpio_defaults_block_21/gpio_defaults [10],
    \gpio_defaults_block_21/gpio_defaults [9],
    \gpio_defaults_block_21/gpio_defaults [8],
    \gpio_defaults_block_21/gpio_defaults [7],
    \gpio_defaults_block_21/gpio_defaults [6],
    \gpio_defaults_block_21/gpio_defaults [5],
    \gpio_defaults_block_21/gpio_defaults [4],
    \gpio_defaults_block_21/gpio_defaults [3],
    \gpio_defaults_block_21/gpio_defaults [2],
    \gpio_defaults_block_21/gpio_defaults [1],
    \gpio_defaults_block_21/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [65],
    \padframe/mprj_io_dm [64],
    \padframe/mprj_io_dm [63]}));
 gpio_control_block \gpio_control_in_2[1]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [20]),
    .mgmt_gpio_oeb(\gpio_control_in_2[1]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [20]),
    .one(\gpio_control_in_2[1]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [20]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [20]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [20]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [20]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [20]),
    .pad_gpio_in(\padframe/mprj_io_in [20]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [20]),
    .pad_gpio_out(\padframe/mprj_io_out [20]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [20]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [20]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [20]),
    .resetn(\gpio_control_in_2[1]/resetn ),
    .resetn_out(\gpio_control_in_2[0]/resetn ),
    .serial_clock(\gpio_control_in_2[1]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[0]/serial_clock ),
    .serial_data_in(\gpio_control_in_2[1]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[0]/serial_data_in ),
    .serial_load(\gpio_control_in_2[1]/serial_load ),
    .serial_load_out(\gpio_control_in_2[0]/serial_load ),
    .user_gpio_in(\mprj/io_in [20]),
    .user_gpio_oeb(\mprj/io_oeb [20]),
    .user_gpio_out(\mprj/io_out [20]),
    .zero(\gpio_control_in_2[1]/zero ),
    .gpio_defaults({\gpio_defaults_block_20/gpio_defaults [12],
    \gpio_defaults_block_20/gpio_defaults [11],
    \gpio_defaults_block_20/gpio_defaults [10],
    \gpio_defaults_block_20/gpio_defaults [9],
    \gpio_defaults_block_20/gpio_defaults [8],
    \gpio_defaults_block_20/gpio_defaults [7],
    \gpio_defaults_block_20/gpio_defaults [6],
    \gpio_defaults_block_20/gpio_defaults [5],
    \gpio_defaults_block_20/gpio_defaults [4],
    \gpio_defaults_block_20/gpio_defaults [3],
    \gpio_defaults_block_20/gpio_defaults [2],
    \gpio_defaults_block_20/gpio_defaults [1],
    \gpio_defaults_block_20/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [62],
    \padframe/mprj_io_dm [61],
    \padframe/mprj_io_dm [60]}));
 gpio_defaults_block gpio_defaults_block_19 (.gpio_defaults({\gpio_defaults_block_19/gpio_defaults [12],
    \gpio_defaults_block_19/gpio_defaults [11],
    \gpio_defaults_block_19/gpio_defaults [10],
    \gpio_defaults_block_19/gpio_defaults [9],
    \gpio_defaults_block_19/gpio_defaults [8],
    \gpio_defaults_block_19/gpio_defaults [7],
    \gpio_defaults_block_19/gpio_defaults [6],
    \gpio_defaults_block_19/gpio_defaults [5],
    \gpio_defaults_block_19/gpio_defaults [4],
    \gpio_defaults_block_19/gpio_defaults [3],
    \gpio_defaults_block_19/gpio_defaults [2],
    \gpio_defaults_block_19/gpio_defaults [1],
    \gpio_defaults_block_19/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_20 (.gpio_defaults({\gpio_defaults_block_20/gpio_defaults [12],
    \gpio_defaults_block_20/gpio_defaults [11],
    \gpio_defaults_block_20/gpio_defaults [10],
    \gpio_defaults_block_20/gpio_defaults [9],
    \gpio_defaults_block_20/gpio_defaults [8],
    \gpio_defaults_block_20/gpio_defaults [7],
    \gpio_defaults_block_20/gpio_defaults [6],
    \gpio_defaults_block_20/gpio_defaults [5],
    \gpio_defaults_block_20/gpio_defaults [4],
    \gpio_defaults_block_20/gpio_defaults [3],
    \gpio_defaults_block_20/gpio_defaults [2],
    \gpio_defaults_block_20/gpio_defaults [1],
    \gpio_defaults_block_20/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_2[0]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [19]),
    .mgmt_gpio_oeb(\gpio_control_in_2[0]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [19]),
    .one(\gpio_control_in_2[0]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [19]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [19]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [19]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [19]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [19]),
    .pad_gpio_in(\padframe/mprj_io_in [19]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [19]),
    .pad_gpio_out(\padframe/mprj_io_out [19]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [19]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [19]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [19]),
    .resetn(\gpio_control_in_2[0]/resetn ),
    .resetn_out(\gpio_control_in_2[0]/resetn_out ),
    .serial_clock(\gpio_control_in_2[0]/serial_clock ),
    .serial_clock_out(\gpio_control_in_2[0]/serial_clock_out ),
    .serial_data_in(\gpio_control_in_2[0]/serial_data_in ),
    .serial_data_out(\gpio_control_in_2[0]/serial_data_out ),
    .serial_load(\gpio_control_in_2[0]/serial_load ),
    .serial_load_out(\gpio_control_in_2[0]/serial_load_out ),
    .user_gpio_in(\mprj/io_in [19]),
    .user_gpio_oeb(\mprj/io_oeb [19]),
    .user_gpio_out(\mprj/io_out [19]),
    .zero(\gpio_control_in_2[0]/zero ),
    .gpio_defaults({\gpio_defaults_block_19/gpio_defaults [12],
    \gpio_defaults_block_19/gpio_defaults [11],
    \gpio_defaults_block_19/gpio_defaults [10],
    \gpio_defaults_block_19/gpio_defaults [9],
    \gpio_defaults_block_19/gpio_defaults [8],
    \gpio_defaults_block_19/gpio_defaults [7],
    \gpio_defaults_block_19/gpio_defaults [6],
    \gpio_defaults_block_19/gpio_defaults [5],
    \gpio_defaults_block_19/gpio_defaults [4],
    \gpio_defaults_block_19/gpio_defaults [3],
    \gpio_defaults_block_19/gpio_defaults [2],
    \gpio_defaults_block_19/gpio_defaults [1],
    \gpio_defaults_block_19/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [59],
    \padframe/mprj_io_dm [58],
    \padframe/mprj_io_dm [57]}));
 gpio_defaults_block gpio_defaults_block_17 (.gpio_defaults({\gpio_defaults_block_17/gpio_defaults [12],
    \gpio_defaults_block_17/gpio_defaults [11],
    \gpio_defaults_block_17/gpio_defaults [10],
    \gpio_defaults_block_17/gpio_defaults [9],
    \gpio_defaults_block_17/gpio_defaults [8],
    \gpio_defaults_block_17/gpio_defaults [7],
    \gpio_defaults_block_17/gpio_defaults [6],
    \gpio_defaults_block_17/gpio_defaults [5],
    \gpio_defaults_block_17/gpio_defaults [4],
    \gpio_defaults_block_17/gpio_defaults [3],
    \gpio_defaults_block_17/gpio_defaults [2],
    \gpio_defaults_block_17/gpio_defaults [1],
    \gpio_defaults_block_17/gpio_defaults [0]}));
 gpio_defaults_block gpio_defaults_block_18 (.gpio_defaults({\gpio_defaults_block_18/gpio_defaults [12],
    \gpio_defaults_block_18/gpio_defaults [11],
    \gpio_defaults_block_18/gpio_defaults [10],
    \gpio_defaults_block_18/gpio_defaults [9],
    \gpio_defaults_block_18/gpio_defaults [8],
    \gpio_defaults_block_18/gpio_defaults [7],
    \gpio_defaults_block_18/gpio_defaults [6],
    \gpio_defaults_block_18/gpio_defaults [5],
    \gpio_defaults_block_18/gpio_defaults [4],
    \gpio_defaults_block_18/gpio_defaults [3],
    \gpio_defaults_block_18/gpio_defaults [2],
    \gpio_defaults_block_18/gpio_defaults [1],
    \gpio_defaults_block_18/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[9]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [17]),
    .mgmt_gpio_oeb(\gpio_control_in_1[9]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [17]),
    .one(\gpio_control_in_1[9]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [17]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [17]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [17]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [17]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [17]),
    .pad_gpio_in(\padframe/mprj_io_in [17]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [17]),
    .pad_gpio_out(\padframe/mprj_io_out [17]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [17]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [17]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [17]),
    .resetn(\gpio_control_in_1[9]/resetn ),
    .resetn_out(\gpio_control_in_1[10]/resetn ),
    .serial_clock(\gpio_control_in_1[9]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[10]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[9]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[9]/serial_data_out ),
    .serial_load(\gpio_control_in_1[9]/serial_load ),
    .serial_load_out(\gpio_control_in_1[10]/serial_load ),
    .user_gpio_in(\mprj/io_in [17]),
    .user_gpio_oeb(\mprj/io_oeb [17]),
    .user_gpio_out(\mprj/io_out [17]),
    .zero(\gpio_control_in_1[9]/zero ),
    .gpio_defaults({\gpio_defaults_block_17/gpio_defaults [12],
    \gpio_defaults_block_17/gpio_defaults [11],
    \gpio_defaults_block_17/gpio_defaults [10],
    \gpio_defaults_block_17/gpio_defaults [9],
    \gpio_defaults_block_17/gpio_defaults [8],
    \gpio_defaults_block_17/gpio_defaults [7],
    \gpio_defaults_block_17/gpio_defaults [6],
    \gpio_defaults_block_17/gpio_defaults [5],
    \gpio_defaults_block_17/gpio_defaults [4],
    \gpio_defaults_block_17/gpio_defaults [3],
    \gpio_defaults_block_17/gpio_defaults [2],
    \gpio_defaults_block_17/gpio_defaults [1],
    \gpio_defaults_block_17/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [53],
    \padframe/mprj_io_dm [52],
    \padframe/mprj_io_dm [51]}));
 gpio_control_block \gpio_control_in_1[10]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [18]),
    .mgmt_gpio_oeb(\gpio_control_in_1[10]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [18]),
    .one(\gpio_control_in_1[10]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [18]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [18]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [18]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [18]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [18]),
    .pad_gpio_in(\padframe/mprj_io_in [18]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [18]),
    .pad_gpio_out(\padframe/mprj_io_out [18]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [18]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [18]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [18]),
    .resetn(\gpio_control_in_1[10]/resetn ),
    .resetn_out(\gpio_control_in_1[10]/resetn_out ),
    .serial_clock(\gpio_control_in_1[10]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[10]/serial_clock_out ),
    .serial_data_in(\gpio_control_in_1[9]/serial_data_out ),
    .serial_data_out(\gpio_control_in_1[10]/serial_data_out ),
    .serial_load(\gpio_control_in_1[10]/serial_load ),
    .serial_load_out(\gpio_control_in_1[10]/serial_load_out ),
    .user_gpio_in(\mprj/io_in [18]),
    .user_gpio_oeb(\mprj/io_oeb [18]),
    .user_gpio_out(\mprj/io_out [18]),
    .zero(\gpio_control_in_1[10]/zero ),
    .gpio_defaults({\gpio_defaults_block_18/gpio_defaults [12],
    \gpio_defaults_block_18/gpio_defaults [11],
    \gpio_defaults_block_18/gpio_defaults [10],
    \gpio_defaults_block_18/gpio_defaults [9],
    \gpio_defaults_block_18/gpio_defaults [8],
    \gpio_defaults_block_18/gpio_defaults [7],
    \gpio_defaults_block_18/gpio_defaults [6],
    \gpio_defaults_block_18/gpio_defaults [5],
    \gpio_defaults_block_18/gpio_defaults [4],
    \gpio_defaults_block_18/gpio_defaults [3],
    \gpio_defaults_block_18/gpio_defaults [2],
    \gpio_defaults_block_18/gpio_defaults [1],
    \gpio_defaults_block_18/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [56],
    \padframe/mprj_io_dm [55],
    \padframe/mprj_io_dm [54]}));
 gpio_defaults_block gpio_defaults_block_16 (.gpio_defaults({\gpio_defaults_block_16/gpio_defaults [12],
    \gpio_defaults_block_16/gpio_defaults [11],
    \gpio_defaults_block_16/gpio_defaults [10],
    \gpio_defaults_block_16/gpio_defaults [9],
    \gpio_defaults_block_16/gpio_defaults [8],
    \gpio_defaults_block_16/gpio_defaults [7],
    \gpio_defaults_block_16/gpio_defaults [6],
    \gpio_defaults_block_16/gpio_defaults [5],
    \gpio_defaults_block_16/gpio_defaults [4],
    \gpio_defaults_block_16/gpio_defaults [3],
    \gpio_defaults_block_16/gpio_defaults [2],
    \gpio_defaults_block_16/gpio_defaults [1],
    \gpio_defaults_block_16/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[8]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [16]),
    .mgmt_gpio_oeb(\gpio_control_in_1[8]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [16]),
    .one(\gpio_control_in_1[8]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [16]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [16]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [16]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [16]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [16]),
    .pad_gpio_in(\padframe/mprj_io_in [16]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [16]),
    .pad_gpio_out(\padframe/mprj_io_out [16]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [16]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [16]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [16]),
    .resetn(\gpio_control_in_1[8]/resetn ),
    .resetn_out(\gpio_control_in_1[9]/resetn ),
    .serial_clock(\gpio_control_in_1[8]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[9]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[8]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[9]/serial_data_in ),
    .serial_load(\gpio_control_in_1[8]/serial_load ),
    .serial_load_out(\gpio_control_in_1[9]/serial_load ),
    .user_gpio_in(\mprj/io_in [16]),
    .user_gpio_oeb(\mprj/io_oeb [16]),
    .user_gpio_out(\mprj/io_out [16]),
    .zero(\gpio_control_in_1[8]/zero ),
    .gpio_defaults({\gpio_defaults_block_16/gpio_defaults [12],
    \gpio_defaults_block_16/gpio_defaults [11],
    \gpio_defaults_block_16/gpio_defaults [10],
    \gpio_defaults_block_16/gpio_defaults [9],
    \gpio_defaults_block_16/gpio_defaults [8],
    \gpio_defaults_block_16/gpio_defaults [7],
    \gpio_defaults_block_16/gpio_defaults [6],
    \gpio_defaults_block_16/gpio_defaults [5],
    \gpio_defaults_block_16/gpio_defaults [4],
    \gpio_defaults_block_16/gpio_defaults [3],
    \gpio_defaults_block_16/gpio_defaults [2],
    \gpio_defaults_block_16/gpio_defaults [1],
    \gpio_defaults_block_16/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [50],
    \padframe/mprj_io_dm [49],
    \padframe/mprj_io_dm [48]}));
 gpio_defaults_block gpio_defaults_block_15 (.gpio_defaults({\gpio_defaults_block_15/gpio_defaults [12],
    \gpio_defaults_block_15/gpio_defaults [11],
    \gpio_defaults_block_15/gpio_defaults [10],
    \gpio_defaults_block_15/gpio_defaults [9],
    \gpio_defaults_block_15/gpio_defaults [8],
    \gpio_defaults_block_15/gpio_defaults [7],
    \gpio_defaults_block_15/gpio_defaults [6],
    \gpio_defaults_block_15/gpio_defaults [5],
    \gpio_defaults_block_15/gpio_defaults [4],
    \gpio_defaults_block_15/gpio_defaults [3],
    \gpio_defaults_block_15/gpio_defaults [2],
    \gpio_defaults_block_15/gpio_defaults [1],
    \gpio_defaults_block_15/gpio_defaults [0]}));
 gpio_control_block \gpio_control_in_1[7]  (.mgmt_gpio_in(\housekeeping/mgmt_gpio_in [15]),
    .mgmt_gpio_oeb(\gpio_control_in_1[7]/one ),
    .mgmt_gpio_out(\housekeeping/mgmt_gpio_in [15]),
    .one(\gpio_control_in_1[7]/one ),
    .pad_gpio_ana_en(\padframe/mprj_io_analog_en [15]),
    .pad_gpio_ana_pol(\padframe/mprj_io_analog_pol [15]),
    .pad_gpio_ana_sel(\padframe/mprj_io_analog_sel [15]),
    .pad_gpio_holdover(\padframe/mprj_io_holdover [15]),
    .pad_gpio_ib_mode_sel(\padframe/mprj_io_ib_mode_sel [15]),
    .pad_gpio_in(\padframe/mprj_io_in [15]),
    .pad_gpio_inenb(\padframe/mprj_io_inp_dis [15]),
    .pad_gpio_out(\padframe/mprj_io_out [15]),
    .pad_gpio_outenb(\padframe/mprj_io_oeb [15]),
    .pad_gpio_slow_sel(\padframe/mprj_io_slow_sel [15]),
    .pad_gpio_vtrip_sel(\padframe/mprj_io_vtrip_sel [15]),
    .resetn(\gpio_control_in_1[7]/resetn ),
    .resetn_out(\gpio_control_in_1[8]/resetn ),
    .serial_clock(\gpio_control_in_1[7]/serial_clock ),
    .serial_clock_out(\gpio_control_in_1[8]/serial_clock ),
    .serial_data_in(\gpio_control_in_1[7]/serial_data_in ),
    .serial_data_out(\gpio_control_in_1[8]/serial_data_in ),
    .serial_load(\gpio_control_in_1[7]/serial_load ),
    .serial_load_out(\gpio_control_in_1[8]/serial_load ),
    .user_gpio_in(\mprj/io_in [15]),
    .user_gpio_oeb(\mprj/io_oeb [15]),
    .user_gpio_out(\mprj/io_out [15]),
    .zero(\gpio_control_in_1[7]/zero ),
    .gpio_defaults({\gpio_defaults_block_15/gpio_defaults [12],
    \gpio_defaults_block_15/gpio_defaults [11],
    \gpio_defaults_block_15/gpio_defaults [10],
    \gpio_defaults_block_15/gpio_defaults [9],
    \gpio_defaults_block_15/gpio_defaults [8],
    \gpio_defaults_block_15/gpio_defaults [7],
    \gpio_defaults_block_15/gpio_defaults [6],
    \gpio_defaults_block_15/gpio_defaults [5],
    \gpio_defaults_block_15/gpio_defaults [4],
    \gpio_defaults_block_15/gpio_defaults [3],
    \gpio_defaults_block_15/gpio_defaults [2],
    \gpio_defaults_block_15/gpio_defaults [1],
    \gpio_defaults_block_15/gpio_defaults [0]}),
    .pad_gpio_dm({\padframe/mprj_io_dm [47],
    \padframe/mprj_io_dm [46],
    \padframe/mprj_io_dm [45]}));
 user_project_wrapper mprj (.user_clock2(\mprj/user_clock2 ),
    .wb_clk_i(\mprj/wb_clk_i ),
    .wb_rst_i(\mprj/wb_rst_i ),
    .wbs_ack_o(\mprj/wbs_ack_o ),
    .wbs_cyc_i(\mprj/wbs_cyc_i ),
    .wbs_stb_i(\mprj/wbs_stb_i ),
    .wbs_we_i(\mprj/wbs_we_i ),
    .analog_io({\mprj/analog_io [28],
    \mprj/analog_io [27],
    \mprj/analog_io [26],
    \mprj/analog_io [25],
    \mprj/analog_io [24],
    \mprj/analog_io [23],
    \mprj/analog_io [22],
    \mprj/analog_io [21],
    \mprj/analog_io [20],
    \mprj/analog_io [19],
    \mprj/analog_io [18],
    \mprj/analog_io [17],
    \mprj/analog_io [16],
    \mprj/analog_io [15],
    \mprj/analog_io [14],
    \mprj/analog_io [13],
    \mprj/analog_io [12],
    \mprj/analog_io [11],
    \mprj/analog_io [10],
    \mprj/analog_io [9],
    \mprj/analog_io [8],
    \mprj/analog_io [7],
    \mprj/analog_io [6],
    \mprj/analog_io [5],
    \mprj/analog_io [4],
    \mprj/analog_io [3],
    \mprj/analog_io [2],
    \mprj/analog_io [1],
    \mprj/analog_io [0]}),
    .io_in({\mprj/io_in [37],
    \mprj/io_in [36],
    \mprj/io_in [35],
    \mprj/io_in [34],
    \mprj/io_in [33],
    \mprj/io_in [32],
    \mprj/io_in [31],
    \mprj/io_in [30],
    \mprj/io_in [29],
    \mprj/io_in [28],
    \mprj/io_in [27],
    \mprj/io_in [26],
    \mprj/io_in [25],
    \mprj/io_in [24],
    \mprj/io_in [23],
    \mprj/io_in [22],
    \mprj/io_in [21],
    \mprj/io_in [20],
    \mprj/io_in [19],
    \mprj/io_in [18],
    \mprj/io_in [17],
    \mprj/io_in [16],
    \mprj/io_in [15],
    \mprj/io_in [14],
    \mprj/io_in [13],
    \mprj/io_in [12],
    \mprj/io_in [11],
    \mprj/io_in [10],
    \mprj/io_in [9],
    \mprj/io_in [8],
    \mprj/io_in [7],
    \mprj/io_in [6],
    \mprj/io_in [5],
    \mprj/io_in [4],
    \mprj/io_in [3],
    \mprj/io_in [2],
    \mprj/io_in [1],
    \mprj/io_in [0]}),
    .io_oeb({\mprj/io_oeb [37],
    \mprj/io_oeb [36],
    \mprj/io_oeb [35],
    \mprj/io_oeb [34],
    \mprj/io_oeb [33],
    \mprj/io_oeb [32],
    \mprj/io_oeb [31],
    \mprj/io_oeb [30],
    \mprj/io_oeb [29],
    \mprj/io_oeb [28],
    \mprj/io_oeb [27],
    \mprj/io_oeb [26],
    \mprj/io_oeb [25],
    \mprj/io_oeb [24],
    \mprj/io_oeb [23],
    \mprj/io_oeb [22],
    \mprj/io_oeb [21],
    \mprj/io_oeb [20],
    \mprj/io_oeb [19],
    \mprj/io_oeb [18],
    \mprj/io_oeb [17],
    \mprj/io_oeb [16],
    \mprj/io_oeb [15],
    \mprj/io_oeb [14],
    \mprj/io_oeb [13],
    \mprj/io_oeb [12],
    \mprj/io_oeb [11],
    \mprj/io_oeb [10],
    \mprj/io_oeb [9],
    \mprj/io_oeb [8],
    \mprj/io_oeb [7],
    \mprj/io_oeb [6],
    \mprj/io_oeb [5],
    \mprj/io_oeb [4],
    \mprj/io_oeb [3],
    \mprj/io_oeb [2],
    \mprj/io_oeb [1],
    \mprj/io_oeb [0]}),
    .io_out({\mprj/io_out [37],
    \mprj/io_out [36],
    \mprj/io_out [35],
    \mprj/io_out [34],
    \mprj/io_out [33],
    \mprj/io_out [32],
    \mprj/io_out [31],
    \mprj/io_out [30],
    \mprj/io_out [29],
    \mprj/io_out [28],
    \mprj/io_out [27],
    \mprj/io_out [26],
    \mprj/io_out [25],
    \mprj/io_out [24],
    \mprj/io_out [23],
    \mprj/io_out [22],
    \mprj/io_out [21],
    \mprj/io_out [20],
    \mprj/io_out [19],
    \mprj/io_out [18],
    \mprj/io_out [17],
    \mprj/io_out [16],
    \mprj/io_out [15],
    \mprj/io_out [14],
    \mprj/io_out [13],
    \mprj/io_out [12],
    \mprj/io_out [11],
    \mprj/io_out [10],
    \mprj/io_out [9],
    \mprj/io_out [8],
    \mprj/io_out [7],
    \mprj/io_out [6],
    \mprj/io_out [5],
    \mprj/io_out [4],
    \mprj/io_out [3],
    \mprj/io_out [2],
    \mprj/io_out [1],
    \mprj/io_out [0]}),
    .la_data_in({\mprj/la_data_in [127],
    \mprj/la_data_in [126],
    \mprj/la_data_in [125],
    \mprj/la_data_in [124],
    \mprj/la_data_in [123],
    \mprj/la_data_in [122],
    \mprj/la_data_in [121],
    \mprj/la_data_in [120],
    \mprj/la_data_in [119],
    \mprj/la_data_in [118],
    \mprj/la_data_in [117],
    \mprj/la_data_in [116],
    \mprj/la_data_in [115],
    \mprj/la_data_in [114],
    \mprj/la_data_in [113],
    \mprj/la_data_in [112],
    \mprj/la_data_in [111],
    \mprj/la_data_in [110],
    \mprj/la_data_in [109],
    \mprj/la_data_in [108],
    \mprj/la_data_in [107],
    \mprj/la_data_in [106],
    \mprj/la_data_in [105],
    \mprj/la_data_in [104],
    \mprj/la_data_in [103],
    \mprj/la_data_in [102],
    \mprj/la_data_in [101],
    \mprj/la_data_in [100],
    \mprj/la_data_in [99],
    \mprj/la_data_in [98],
    \mprj/la_data_in [97],
    \mprj/la_data_in [96],
    \mprj/la_data_in [95],
    \mprj/la_data_in [94],
    \mprj/la_data_in [93],
    \mprj/la_data_in [92],
    \mprj/la_data_in [91],
    \mprj/la_data_in [90],
    \mprj/la_data_in [89],
    \mprj/la_data_in [88],
    \mprj/la_data_in [87],
    \mprj/la_data_in [86],
    \mprj/la_data_in [85],
    \mprj/la_data_in [84],
    \mprj/la_data_in [83],
    \mprj/la_data_in [82],
    \mprj/la_data_in [81],
    \mprj/la_data_in [80],
    \mprj/la_data_in [79],
    \mprj/la_data_in [78],
    \mprj/la_data_in [77],
    \mprj/la_data_in [76],
    \mprj/la_data_in [75],
    \mprj/la_data_in [74],
    \mprj/la_data_in [73],
    \mprj/la_data_in [72],
    \mprj/la_data_in [71],
    \mprj/la_data_in [70],
    \mprj/la_data_in [69],
    \mprj/la_data_in [68],
    \mprj/la_data_in [67],
    \mprj/la_data_in [66],
    \mprj/la_data_in [65],
    \mprj/la_data_in [64],
    \mprj/la_data_in [63],
    \mprj/la_data_in [62],
    \mprj/la_data_in [61],
    \mprj/la_data_in [60],
    \mprj/la_data_in [59],
    \mprj/la_data_in [58],
    \mprj/la_data_in [57],
    \mprj/la_data_in [56],
    \mprj/la_data_in [55],
    \mprj/la_data_in [54],
    \mprj/la_data_in [53],
    \mprj/la_data_in [52],
    \mprj/la_data_in [51],
    \mprj/la_data_in [50],
    \mprj/la_data_in [49],
    \mprj/la_data_in [48],
    \mprj/la_data_in [47],
    \mprj/la_data_in [46],
    \mprj/la_data_in [45],
    \mprj/la_data_in [44],
    \mprj/la_data_in [43],
    \mprj/la_data_in [42],
    \mprj/la_data_in [41],
    \mprj/la_data_in [40],
    \mprj/la_data_in [39],
    \mprj/la_data_in [38],
    \mprj/la_data_in [37],
    \mprj/la_data_in [36],
    \mprj/la_data_in [35],
    \mprj/la_data_in [34],
    \mprj/la_data_in [33],
    \mprj/la_data_in [32],
    \mprj/la_data_in [31],
    \mprj/la_data_in [30],
    \mprj/la_data_in [29],
    \mprj/la_data_in [28],
    \mprj/la_data_in [27],
    \mprj/la_data_in [26],
    \mprj/la_data_in [25],
    \mprj/la_data_in [24],
    \mprj/la_data_in [23],
    \mprj/la_data_in [22],
    \mprj/la_data_in [21],
    \mprj/la_data_in [20],
    \mprj/la_data_in [19],
    \mprj/la_data_in [18],
    \mprj/la_data_in [17],
    \mprj/la_data_in [16],
    \mprj/la_data_in [15],
    \mprj/la_data_in [14],
    \mprj/la_data_in [13],
    \mprj/la_data_in [12],
    \mprj/la_data_in [11],
    \mprj/la_data_in [10],
    \mprj/la_data_in [9],
    \mprj/la_data_in [8],
    \mprj/la_data_in [7],
    \mprj/la_data_in [6],
    \mprj/la_data_in [5],
    \mprj/la_data_in [4],
    \mprj/la_data_in [3],
    \mprj/la_data_in [2],
    \mprj/la_data_in [1],
    \mprj/la_data_in [0]}),
    .la_data_out({\mprj/la_data_out [127],
    \mprj/la_data_out [126],
    \mprj/la_data_out [125],
    \mprj/la_data_out [124],
    \mprj/la_data_out [123],
    \mprj/la_data_out [122],
    \mprj/la_data_out [121],
    \mprj/la_data_out [120],
    \mprj/la_data_out [119],
    \mprj/la_data_out [118],
    \mprj/la_data_out [117],
    \mprj/la_data_out [116],
    \mprj/la_data_out [115],
    \mprj/la_data_out [114],
    \mprj/la_data_out [113],
    \mprj/la_data_out [112],
    \mprj/la_data_out [111],
    \mprj/la_data_out [110],
    \mprj/la_data_out [109],
    \mprj/la_data_out [108],
    \mprj/la_data_out [107],
    \mprj/la_data_out [106],
    \mprj/la_data_out [105],
    \mprj/la_data_out [104],
    \mprj/la_data_out [103],
    \mprj/la_data_out [102],
    \mprj/la_data_out [101],
    \mprj/la_data_out [100],
    \mprj/la_data_out [99],
    \mprj/la_data_out [98],
    \mprj/la_data_out [97],
    \mprj/la_data_out [96],
    \mprj/la_data_out [95],
    \mprj/la_data_out [94],
    \mprj/la_data_out [93],
    \mprj/la_data_out [92],
    \mprj/la_data_out [91],
    \mprj/la_data_out [90],
    \mprj/la_data_out [89],
    \mprj/la_data_out [88],
    \mprj/la_data_out [87],
    \mprj/la_data_out [86],
    \mprj/la_data_out [85],
    \mprj/la_data_out [84],
    \mprj/la_data_out [83],
    \mprj/la_data_out [82],
    \mprj/la_data_out [81],
    \mprj/la_data_out [80],
    \mprj/la_data_out [79],
    \mprj/la_data_out [78],
    \mprj/la_data_out [77],
    \mprj/la_data_out [76],
    \mprj/la_data_out [75],
    \mprj/la_data_out [74],
    \mprj/la_data_out [73],
    \mprj/la_data_out [72],
    \mprj/la_data_out [71],
    \mprj/la_data_out [70],
    \mprj/la_data_out [69],
    \mprj/la_data_out [68],
    \mprj/la_data_out [67],
    \mprj/la_data_out [66],
    \mprj/la_data_out [65],
    \mprj/la_data_out [64],
    \mprj/la_data_out [63],
    \mprj/la_data_out [62],
    \mprj/la_data_out [61],
    \mprj/la_data_out [60],
    \mprj/la_data_out [59],
    \mprj/la_data_out [58],
    \mprj/la_data_out [57],
    \mprj/la_data_out [56],
    \mprj/la_data_out [55],
    \mprj/la_data_out [54],
    \mprj/la_data_out [53],
    \mprj/la_data_out [52],
    \mprj/la_data_out [51],
    \mprj/la_data_out [50],
    \mprj/la_data_out [49],
    \mprj/la_data_out [48],
    \mprj/la_data_out [47],
    \mprj/la_data_out [46],
    \mprj/la_data_out [45],
    \mprj/la_data_out [44],
    \mprj/la_data_out [43],
    \mprj/la_data_out [42],
    \mprj/la_data_out [41],
    \mprj/la_data_out [40],
    \mprj/la_data_out [39],
    \mprj/la_data_out [38],
    \mprj/la_data_out [37],
    \mprj/la_data_out [36],
    \mprj/la_data_out [35],
    \mprj/la_data_out [34],
    \mprj/la_data_out [33],
    \mprj/la_data_out [32],
    \mprj/la_data_out [31],
    \mprj/la_data_out [30],
    \mprj/la_data_out [29],
    \mprj/la_data_out [28],
    \mprj/la_data_out [27],
    \mprj/la_data_out [26],
    \mprj/la_data_out [25],
    \mprj/la_data_out [24],
    \mprj/la_data_out [23],
    \mprj/la_data_out [22],
    \mprj/la_data_out [21],
    \mprj/la_data_out [20],
    \mprj/la_data_out [19],
    \mprj/la_data_out [18],
    \mprj/la_data_out [17],
    \mprj/la_data_out [16],
    \mprj/la_data_out [15],
    \mprj/la_data_out [14],
    \mprj/la_data_out [13],
    \mprj/la_data_out [12],
    \mprj/la_data_out [11],
    \mprj/la_data_out [10],
    \mprj/la_data_out [9],
    \mprj/la_data_out [8],
    \mprj/la_data_out [7],
    \mprj/la_data_out [6],
    \mprj/la_data_out [5],
    \mprj/la_data_out [4],
    \mprj/la_data_out [3],
    \mprj/la_data_out [2],
    \mprj/la_data_out [1],
    \mprj/la_data_out [0]}),
    .la_oenb({\mprj/la_oenb [127],
    \mprj/la_oenb [126],
    \mprj/la_oenb [125],
    \mprj/la_oenb [124],
    \mprj/la_oenb [123],
    \mprj/la_oenb [122],
    \mprj/la_oenb [121],
    \mprj/la_oenb [120],
    \mprj/la_oenb [119],
    \mprj/la_oenb [118],
    \mprj/la_oenb [117],
    \mprj/la_oenb [116],
    \mprj/la_oenb [115],
    \mprj/la_oenb [114],
    \mprj/la_oenb [113],
    \mprj/la_oenb [112],
    \mprj/la_oenb [111],
    \mprj/la_oenb [110],
    \mprj/la_oenb [109],
    \mprj/la_oenb [108],
    \mprj/la_oenb [107],
    \mprj/la_oenb [106],
    \mprj/la_oenb [105],
    \mprj/la_oenb [104],
    \mprj/la_oenb [103],
    \mprj/la_oenb [102],
    \mprj/la_oenb [101],
    \mprj/la_oenb [100],
    \mprj/la_oenb [99],
    \mprj/la_oenb [98],
    \mprj/la_oenb [97],
    \mprj/la_oenb [96],
    \mprj/la_oenb [95],
    \mprj/la_oenb [94],
    \mprj/la_oenb [93],
    \mprj/la_oenb [92],
    \mprj/la_oenb [91],
    \mprj/la_oenb [90],
    \mprj/la_oenb [89],
    \mprj/la_oenb [88],
    \mprj/la_oenb [87],
    \mprj/la_oenb [86],
    \mprj/la_oenb [85],
    \mprj/la_oenb [84],
    \mprj/la_oenb [83],
    \mprj/la_oenb [82],
    \mprj/la_oenb [81],
    \mprj/la_oenb [80],
    \mprj/la_oenb [79],
    \mprj/la_oenb [78],
    \mprj/la_oenb [77],
    \mprj/la_oenb [76],
    \mprj/la_oenb [75],
    \mprj/la_oenb [74],
    \mprj/la_oenb [73],
    \mprj/la_oenb [72],
    \mprj/la_oenb [71],
    \mprj/la_oenb [70],
    \mprj/la_oenb [69],
    \mprj/la_oenb [68],
    \mprj/la_oenb [67],
    \mprj/la_oenb [66],
    \mprj/la_oenb [65],
    \mprj/la_oenb [64],
    \mprj/la_oenb [63],
    \mprj/la_oenb [62],
    \mprj/la_oenb [61],
    \mprj/la_oenb [60],
    \mprj/la_oenb [59],
    \mprj/la_oenb [58],
    \mprj/la_oenb [57],
    \mprj/la_oenb [56],
    \mprj/la_oenb [55],
    \mprj/la_oenb [54],
    \mprj/la_oenb [53],
    \mprj/la_oenb [52],
    \mprj/la_oenb [51],
    \mprj/la_oenb [50],
    \mprj/la_oenb [49],
    \mprj/la_oenb [48],
    \mprj/la_oenb [47],
    \mprj/la_oenb [46],
    \mprj/la_oenb [45],
    \mprj/la_oenb [44],
    \mprj/la_oenb [43],
    \mprj/la_oenb [42],
    \mprj/la_oenb [41],
    \mprj/la_oenb [40],
    \mprj/la_oenb [39],
    \mprj/la_oenb [38],
    \mprj/la_oenb [37],
    \mprj/la_oenb [36],
    \mprj/la_oenb [35],
    \mprj/la_oenb [34],
    \mprj/la_oenb [33],
    \mprj/la_oenb [32],
    \mprj/la_oenb [31],
    \mprj/la_oenb [30],
    \mprj/la_oenb [29],
    \mprj/la_oenb [28],
    \mprj/la_oenb [27],
    \mprj/la_oenb [26],
    \mprj/la_oenb [25],
    \mprj/la_oenb [24],
    \mprj/la_oenb [23],
    \mprj/la_oenb [22],
    \mprj/la_oenb [21],
    \mprj/la_oenb [20],
    \mprj/la_oenb [19],
    \mprj/la_oenb [18],
    \mprj/la_oenb [17],
    \mprj/la_oenb [16],
    \mprj/la_oenb [15],
    \mprj/la_oenb [14],
    \mprj/la_oenb [13],
    \mprj/la_oenb [12],
    \mprj/la_oenb [11],
    \mprj/la_oenb [10],
    \mprj/la_oenb [9],
    \mprj/la_oenb [8],
    \mprj/la_oenb [7],
    \mprj/la_oenb [6],
    \mprj/la_oenb [5],
    \mprj/la_oenb [4],
    \mprj/la_oenb [3],
    \mprj/la_oenb [2],
    \mprj/la_oenb [1],
    \mprj/la_oenb [0]}),
    .user_irq({\mprj/user_irq [2],
    \mprj/user_irq [1],
    \mprj/user_irq [0]}),
    .wbs_adr_i({\mprj/wbs_adr_i [31],
    \mprj/wbs_adr_i [30],
    \mprj/wbs_adr_i [29],
    \mprj/wbs_adr_i [28],
    \mprj/wbs_adr_i [27],
    \mprj/wbs_adr_i [26],
    \mprj/wbs_adr_i [25],
    \mprj/wbs_adr_i [24],
    \mprj/wbs_adr_i [23],
    \mprj/wbs_adr_i [22],
    \mprj/wbs_adr_i [21],
    \mprj/wbs_adr_i [20],
    \mprj/wbs_adr_i [19],
    \mprj/wbs_adr_i [18],
    \mprj/wbs_adr_i [17],
    \mprj/wbs_adr_i [16],
    \mprj/wbs_adr_i [15],
    \mprj/wbs_adr_i [14],
    \mprj/wbs_adr_i [13],
    \mprj/wbs_adr_i [12],
    \mprj/wbs_adr_i [11],
    \mprj/wbs_adr_i [10],
    \mprj/wbs_adr_i [9],
    \mprj/wbs_adr_i [8],
    \mprj/wbs_adr_i [7],
    \mprj/wbs_adr_i [6],
    \mprj/wbs_adr_i [5],
    \mprj/wbs_adr_i [4],
    \mprj/wbs_adr_i [3],
    \mprj/wbs_adr_i [2],
    \mprj/wbs_adr_i [1],
    \mprj/wbs_adr_i [0]}),
    .wbs_dat_i({\mprj/wbs_dat_i [31],
    \mprj/wbs_dat_i [30],
    \mprj/wbs_dat_i [29],
    \mprj/wbs_dat_i [28],
    \mprj/wbs_dat_i [27],
    \mprj/wbs_dat_i [26],
    \mprj/wbs_dat_i [25],
    \mprj/wbs_dat_i [24],
    \mprj/wbs_dat_i [23],
    \mprj/wbs_dat_i [22],
    \mprj/wbs_dat_i [21],
    \mprj/wbs_dat_i [20],
    \mprj/wbs_dat_i [19],
    \mprj/wbs_dat_i [18],
    \mprj/wbs_dat_i [17],
    \mprj/wbs_dat_i [16],
    \mprj/wbs_dat_i [15],
    \mprj/wbs_dat_i [14],
    \mprj/wbs_dat_i [13],
    \mprj/wbs_dat_i [12],
    \mprj/wbs_dat_i [11],
    \mprj/wbs_dat_i [10],
    \mprj/wbs_dat_i [9],
    \mprj/wbs_dat_i [8],
    \mprj/wbs_dat_i [7],
    \mprj/wbs_dat_i [6],
    \mprj/wbs_dat_i [5],
    \mprj/wbs_dat_i [4],
    \mprj/wbs_dat_i [3],
    \mprj/wbs_dat_i [2],
    \mprj/wbs_dat_i [1],
    \mprj/wbs_dat_i [0]}),
    .wbs_dat_o({\mprj/wbs_dat_o [31],
    \mprj/wbs_dat_o [30],
    \mprj/wbs_dat_o [29],
    \mprj/wbs_dat_o [28],
    \mprj/wbs_dat_o [27],
    \mprj/wbs_dat_o [26],
    \mprj/wbs_dat_o [25],
    \mprj/wbs_dat_o [24],
    \mprj/wbs_dat_o [23],
    \mprj/wbs_dat_o [22],
    \mprj/wbs_dat_o [21],
    \mprj/wbs_dat_o [20],
    \mprj/wbs_dat_o [19],
    \mprj/wbs_dat_o [18],
    \mprj/wbs_dat_o [17],
    \mprj/wbs_dat_o [16],
    \mprj/wbs_dat_o [15],
    \mprj/wbs_dat_o [14],
    \mprj/wbs_dat_o [13],
    \mprj/wbs_dat_o [12],
    \mprj/wbs_dat_o [11],
    \mprj/wbs_dat_o [10],
    \mprj/wbs_dat_o [9],
    \mprj/wbs_dat_o [8],
    \mprj/wbs_dat_o [7],
    \mprj/wbs_dat_o [6],
    \mprj/wbs_dat_o [5],
    \mprj/wbs_dat_o [4],
    \mprj/wbs_dat_o [3],
    \mprj/wbs_dat_o [2],
    \mprj/wbs_dat_o [1],
    \mprj/wbs_dat_o [0]}),
    .wbs_sel_i({\mprj/wbs_sel_i [3],
    \mprj/wbs_sel_i [2],
    \mprj/wbs_sel_i [1],
    \mprj/wbs_sel_i [0]}));
 chip_io padframe (.clock(clock),
    .clock_core(\pll/osc ),
    .por(\por/por_l ),
    .flash_clk(flash_clk),
    .flash_clk_core(\padframe/flash_clk_core ),
    .flash_clk_ieb_core(\padframe/flash_clk_ieb_core ),
    .flash_clk_oeb_core(\padframe/flash_clk_oeb_core ),
    .flash_csb(flash_csb),
    .flash_csb_core(\padframe/flash_csb_core ),
    .flash_csb_ieb_core(\padframe/flash_csb_ieb_core ),
    .flash_csb_oeb_core(\padframe/flash_csb_oeb_core ),
    .flash_io0(flash_io0),
    .flash_io0_di_core(\padframe/flash_io0_di_core ),
    .flash_io0_do_core(\padframe/flash_io0_do_core ),
    .flash_io0_ieb_core(\padframe/flash_io0_ieb_core ),
    .flash_io0_oeb_core(\padframe/flash_io0_oeb_core ),
    .flash_io1(flash_io1),
    .flash_io1_di_core(\padframe/flash_io1_di_core ),
    .flash_io1_do_core(\padframe/flash_io1_do_core ),
    .flash_io1_ieb_core(\padframe/flash_io1_ieb_core ),
    .flash_io1_oeb_core(\padframe/flash_io1_oeb_core ),
    .gpio(gpio),
    .gpio_in_core(\soc/gpio_in_pad ),
    .gpio_inenb_core(\soc/gpio_inenb_pad ),
    .gpio_mode0_core(\soc/gpio_mode0_pad ),
    .gpio_mode1_core(\soc/gpio_mode1_pad ),
    .gpio_out_core(\soc/gpio_out_pad ),
    .gpio_outenb_core(\soc/gpio_outenb_pad ),
    .porb_h(\por/porb_h ),
    .resetb(resetb),
    .resetb_core_h(\rstb_level/A ),
    .mprj_analog_io({\mprj/analog_io [28],
    \mprj/analog_io [27],
    \mprj/analog_io [26],
    \mprj/analog_io [25],
    \mprj/analog_io [24],
    \mprj/analog_io [23],
    \mprj/analog_io [22],
    \mprj/analog_io [21],
    \mprj/analog_io [20],
    \mprj/analog_io [19],
    \mprj/analog_io [18],
    \mprj/analog_io [17],
    \mprj/analog_io [16],
    \mprj/analog_io [15],
    \mprj/analog_io [14],
    \mprj/analog_io [13],
    \mprj/analog_io [12],
    \mprj/analog_io [11],
    \mprj/analog_io [10],
    \mprj/analog_io [9],
    \mprj/analog_io [8],
    \mprj/analog_io [7],
    \mprj/analog_io [6],
    \mprj/analog_io [5],
    \mprj/analog_io [4],
    \mprj/analog_io [3],
    \mprj/analog_io [2],
    \mprj/analog_io [1],
    \mprj/analog_io [0]}),
    .mprj_io({mprj_io[37],
    mprj_io[36],
    mprj_io[35],
    mprj_io[34],
    mprj_io[33],
    mprj_io[32],
    mprj_io[31],
    mprj_io[30],
    mprj_io[29],
    mprj_io[28],
    mprj_io[27],
    mprj_io[26],
    mprj_io[25],
    mprj_io[24],
    mprj_io[23],
    mprj_io[22],
    mprj_io[21],
    mprj_io[20],
    mprj_io[19],
    mprj_io[18],
    mprj_io[17],
    mprj_io[16],
    mprj_io[15],
    mprj_io[14],
    mprj_io[13],
    mprj_io[12],
    mprj_io[11],
    mprj_io[10],
    mprj_io[9],
    mprj_io[8],
    mprj_io[7],
    mprj_io[6],
    mprj_io[5],
    mprj_io[4],
    mprj_io[3],
    mprj_io[2],
    mprj_io[1],
    mprj_io[0]}),
    .mprj_io_analog_en({\padframe/mprj_io_analog_en [37],
    \padframe/mprj_io_analog_en [36],
    \padframe/mprj_io_analog_en [35],
    \padframe/mprj_io_analog_en [34],
    \padframe/mprj_io_analog_en [33],
    \padframe/mprj_io_analog_en [32],
    \padframe/mprj_io_analog_en [31],
    \padframe/mprj_io_analog_en [30],
    \padframe/mprj_io_analog_en [29],
    \padframe/mprj_io_analog_en [28],
    \padframe/mprj_io_analog_en [27],
    \padframe/mprj_io_analog_en [26],
    \padframe/mprj_io_analog_en [25],
    \padframe/mprj_io_analog_en [24],
    \padframe/mprj_io_analog_en [23],
    \padframe/mprj_io_analog_en [22],
    \padframe/mprj_io_analog_en [21],
    \padframe/mprj_io_analog_en [20],
    \padframe/mprj_io_analog_en [19],
    \padframe/mprj_io_analog_en [18],
    \padframe/mprj_io_analog_en [17],
    \padframe/mprj_io_analog_en [16],
    \padframe/mprj_io_analog_en [15],
    \padframe/mprj_io_analog_en [14],
    \padframe/mprj_io_analog_en [13],
    \padframe/mprj_io_analog_en [12],
    \padframe/mprj_io_analog_en [11],
    \padframe/mprj_io_analog_en [10],
    \padframe/mprj_io_analog_en [9],
    \padframe/mprj_io_analog_en [8],
    \padframe/mprj_io_analog_en [7],
    \padframe/mprj_io_analog_en [6],
    \padframe/mprj_io_analog_en [5],
    \padframe/mprj_io_analog_en [4],
    \padframe/mprj_io_analog_en [3],
    \padframe/mprj_io_analog_en [2],
    \padframe/mprj_io_analog_en [1],
    \padframe/mprj_io_analog_en [0]}),
    .mprj_io_analog_pol({\padframe/mprj_io_analog_pol [37],
    \padframe/mprj_io_analog_pol [36],
    \padframe/mprj_io_analog_pol [35],
    \padframe/mprj_io_analog_pol [34],
    \padframe/mprj_io_analog_pol [33],
    \padframe/mprj_io_analog_pol [32],
    \padframe/mprj_io_analog_pol [31],
    \padframe/mprj_io_analog_pol [30],
    \padframe/mprj_io_analog_pol [29],
    \padframe/mprj_io_analog_pol [28],
    \padframe/mprj_io_analog_pol [27],
    \padframe/mprj_io_analog_pol [26],
    \padframe/mprj_io_analog_pol [25],
    \padframe/mprj_io_analog_pol [24],
    \padframe/mprj_io_analog_pol [23],
    \padframe/mprj_io_analog_pol [22],
    \padframe/mprj_io_analog_pol [21],
    \padframe/mprj_io_analog_pol [20],
    \padframe/mprj_io_analog_pol [19],
    \padframe/mprj_io_analog_pol [18],
    \padframe/mprj_io_analog_pol [17],
    \padframe/mprj_io_analog_pol [16],
    \padframe/mprj_io_analog_pol [15],
    \padframe/mprj_io_analog_pol [14],
    \padframe/mprj_io_analog_pol [13],
    \padframe/mprj_io_analog_pol [12],
    \padframe/mprj_io_analog_pol [11],
    \padframe/mprj_io_analog_pol [10],
    \padframe/mprj_io_analog_pol [9],
    \padframe/mprj_io_analog_pol [8],
    \padframe/mprj_io_analog_pol [7],
    \padframe/mprj_io_analog_pol [6],
    \padframe/mprj_io_analog_pol [5],
    \padframe/mprj_io_analog_pol [4],
    \padframe/mprj_io_analog_pol [3],
    \padframe/mprj_io_analog_pol [2],
    \padframe/mprj_io_analog_pol [1],
    \padframe/mprj_io_analog_pol [0]}),
    .mprj_io_analog_sel({\padframe/mprj_io_analog_sel [37],
    \padframe/mprj_io_analog_sel [36],
    \padframe/mprj_io_analog_sel [35],
    \padframe/mprj_io_analog_sel [34],
    \padframe/mprj_io_analog_sel [33],
    \padframe/mprj_io_analog_sel [32],
    \padframe/mprj_io_analog_sel [31],
    \padframe/mprj_io_analog_sel [30],
    \padframe/mprj_io_analog_sel [29],
    \padframe/mprj_io_analog_sel [28],
    \padframe/mprj_io_analog_sel [27],
    \padframe/mprj_io_analog_sel [26],
    \padframe/mprj_io_analog_sel [25],
    \padframe/mprj_io_analog_sel [24],
    \padframe/mprj_io_analog_sel [23],
    \padframe/mprj_io_analog_sel [22],
    \padframe/mprj_io_analog_sel [21],
    \padframe/mprj_io_analog_sel [20],
    \padframe/mprj_io_analog_sel [19],
    \padframe/mprj_io_analog_sel [18],
    \padframe/mprj_io_analog_sel [17],
    \padframe/mprj_io_analog_sel [16],
    \padframe/mprj_io_analog_sel [15],
    \padframe/mprj_io_analog_sel [14],
    \padframe/mprj_io_analog_sel [13],
    \padframe/mprj_io_analog_sel [12],
    \padframe/mprj_io_analog_sel [11],
    \padframe/mprj_io_analog_sel [10],
    \padframe/mprj_io_analog_sel [9],
    \padframe/mprj_io_analog_sel [8],
    \padframe/mprj_io_analog_sel [7],
    \padframe/mprj_io_analog_sel [6],
    \padframe/mprj_io_analog_sel [5],
    \padframe/mprj_io_analog_sel [4],
    \padframe/mprj_io_analog_sel [3],
    \padframe/mprj_io_analog_sel [2],
    \padframe/mprj_io_analog_sel [1],
    \padframe/mprj_io_analog_sel [0]}),
    .mprj_io_dm({\padframe/mprj_io_dm [113],
    \padframe/mprj_io_dm [112],
    \padframe/mprj_io_dm [111],
    \padframe/mprj_io_dm [110],
    \padframe/mprj_io_dm [109],
    \padframe/mprj_io_dm [108],
    \padframe/mprj_io_dm [107],
    \padframe/mprj_io_dm [106],
    \padframe/mprj_io_dm [105],
    \padframe/mprj_io_dm [104],
    \padframe/mprj_io_dm [103],
    \padframe/mprj_io_dm [102],
    \padframe/mprj_io_dm [101],
    \padframe/mprj_io_dm [100],
    \padframe/mprj_io_dm [99],
    \padframe/mprj_io_dm [98],
    \padframe/mprj_io_dm [97],
    \padframe/mprj_io_dm [96],
    \padframe/mprj_io_dm [95],
    \padframe/mprj_io_dm [94],
    \padframe/mprj_io_dm [93],
    \padframe/mprj_io_dm [92],
    \padframe/mprj_io_dm [91],
    \padframe/mprj_io_dm [90],
    \padframe/mprj_io_dm [89],
    \padframe/mprj_io_dm [88],
    \padframe/mprj_io_dm [87],
    \padframe/mprj_io_dm [86],
    \padframe/mprj_io_dm [85],
    \padframe/mprj_io_dm [84],
    \padframe/mprj_io_dm [83],
    \padframe/mprj_io_dm [82],
    \padframe/mprj_io_dm [81],
    \padframe/mprj_io_dm [80],
    \padframe/mprj_io_dm [79],
    \padframe/mprj_io_dm [78],
    \padframe/mprj_io_dm [77],
    \padframe/mprj_io_dm [76],
    \padframe/mprj_io_dm [75],
    \padframe/mprj_io_dm [74],
    \padframe/mprj_io_dm [73],
    \padframe/mprj_io_dm [72],
    \padframe/mprj_io_dm [71],
    \padframe/mprj_io_dm [70],
    \padframe/mprj_io_dm [69],
    \padframe/mprj_io_dm [68],
    \padframe/mprj_io_dm [67],
    \padframe/mprj_io_dm [66],
    \padframe/mprj_io_dm [65],
    \padframe/mprj_io_dm [64],
    \padframe/mprj_io_dm [63],
    \padframe/mprj_io_dm [62],
    \padframe/mprj_io_dm [61],
    \padframe/mprj_io_dm [60],
    \padframe/mprj_io_dm [59],
    \padframe/mprj_io_dm [58],
    \padframe/mprj_io_dm [57],
    \padframe/mprj_io_dm [56],
    \padframe/mprj_io_dm [55],
    \padframe/mprj_io_dm [54],
    \padframe/mprj_io_dm [53],
    \padframe/mprj_io_dm [52],
    \padframe/mprj_io_dm [51],
    \padframe/mprj_io_dm [50],
    \padframe/mprj_io_dm [49],
    \padframe/mprj_io_dm [48],
    \padframe/mprj_io_dm [47],
    \padframe/mprj_io_dm [46],
    \padframe/mprj_io_dm [45],
    \padframe/mprj_io_dm [44],
    \padframe/mprj_io_dm [43],
    \padframe/mprj_io_dm [42],
    \padframe/mprj_io_dm [41],
    \padframe/mprj_io_dm [40],
    \padframe/mprj_io_dm [39],
    \padframe/mprj_io_dm [38],
    \padframe/mprj_io_dm [37],
    \padframe/mprj_io_dm [36],
    \padframe/mprj_io_dm [35],
    \padframe/mprj_io_dm [34],
    \padframe/mprj_io_dm [33],
    \padframe/mprj_io_dm [32],
    \padframe/mprj_io_dm [31],
    \padframe/mprj_io_dm [30],
    \padframe/mprj_io_dm [29],
    \padframe/mprj_io_dm [28],
    \padframe/mprj_io_dm [27],
    \padframe/mprj_io_dm [26],
    \padframe/mprj_io_dm [25],
    \padframe/mprj_io_dm [24],
    \padframe/mprj_io_dm [23],
    \padframe/mprj_io_dm [22],
    \padframe/mprj_io_dm [21],
    \padframe/mprj_io_dm [20],
    \padframe/mprj_io_dm [19],
    \padframe/mprj_io_dm [18],
    \padframe/mprj_io_dm [17],
    \padframe/mprj_io_dm [16],
    \padframe/mprj_io_dm [15],
    \padframe/mprj_io_dm [14],
    \padframe/mprj_io_dm [13],
    \padframe/mprj_io_dm [12],
    \padframe/mprj_io_dm [11],
    \padframe/mprj_io_dm [10],
    \padframe/mprj_io_dm [9],
    \padframe/mprj_io_dm [8],
    \padframe/mprj_io_dm [7],
    \padframe/mprj_io_dm [6],
    \padframe/mprj_io_dm [5],
    \padframe/mprj_io_dm [4],
    \padframe/mprj_io_dm [3],
    \padframe/mprj_io_dm [2],
    \padframe/mprj_io_dm [1],
    \padframe/mprj_io_dm [0]}),
    .mprj_io_holdover({\padframe/mprj_io_holdover [37],
    \padframe/mprj_io_holdover [36],
    \padframe/mprj_io_holdover [35],
    \padframe/mprj_io_holdover [34],
    \padframe/mprj_io_holdover [33],
    \padframe/mprj_io_holdover [32],
    \padframe/mprj_io_holdover [31],
    \padframe/mprj_io_holdover [30],
    \padframe/mprj_io_holdover [29],
    \padframe/mprj_io_holdover [28],
    \padframe/mprj_io_holdover [27],
    \padframe/mprj_io_holdover [26],
    \padframe/mprj_io_holdover [25],
    \padframe/mprj_io_holdover [24],
    \padframe/mprj_io_holdover [23],
    \padframe/mprj_io_holdover [22],
    \padframe/mprj_io_holdover [21],
    \padframe/mprj_io_holdover [20],
    \padframe/mprj_io_holdover [19],
    \padframe/mprj_io_holdover [18],
    \padframe/mprj_io_holdover [17],
    \padframe/mprj_io_holdover [16],
    \padframe/mprj_io_holdover [15],
    \padframe/mprj_io_holdover [14],
    \padframe/mprj_io_holdover [13],
    \padframe/mprj_io_holdover [12],
    \padframe/mprj_io_holdover [11],
    \padframe/mprj_io_holdover [10],
    \padframe/mprj_io_holdover [9],
    \padframe/mprj_io_holdover [8],
    \padframe/mprj_io_holdover [7],
    \padframe/mprj_io_holdover [6],
    \padframe/mprj_io_holdover [5],
    \padframe/mprj_io_holdover [4],
    \padframe/mprj_io_holdover [3],
    \padframe/mprj_io_holdover [2],
    \padframe/mprj_io_holdover [1],
    \padframe/mprj_io_holdover [0]}),
    .mprj_io_ib_mode_sel({\padframe/mprj_io_ib_mode_sel [37],
    \padframe/mprj_io_ib_mode_sel [36],
    \padframe/mprj_io_ib_mode_sel [35],
    \padframe/mprj_io_ib_mode_sel [34],
    \padframe/mprj_io_ib_mode_sel [33],
    \padframe/mprj_io_ib_mode_sel [32],
    \padframe/mprj_io_ib_mode_sel [31],
    \padframe/mprj_io_ib_mode_sel [30],
    \padframe/mprj_io_ib_mode_sel [29],
    \padframe/mprj_io_ib_mode_sel [28],
    \padframe/mprj_io_ib_mode_sel [27],
    \padframe/mprj_io_ib_mode_sel [26],
    \padframe/mprj_io_ib_mode_sel [25],
    \padframe/mprj_io_ib_mode_sel [24],
    \padframe/mprj_io_ib_mode_sel [23],
    \padframe/mprj_io_ib_mode_sel [22],
    \padframe/mprj_io_ib_mode_sel [21],
    \padframe/mprj_io_ib_mode_sel [20],
    \padframe/mprj_io_ib_mode_sel [19],
    \padframe/mprj_io_ib_mode_sel [18],
    \padframe/mprj_io_ib_mode_sel [17],
    \padframe/mprj_io_ib_mode_sel [16],
    \padframe/mprj_io_ib_mode_sel [15],
    \padframe/mprj_io_ib_mode_sel [14],
    \padframe/mprj_io_ib_mode_sel [13],
    \padframe/mprj_io_ib_mode_sel [12],
    \padframe/mprj_io_ib_mode_sel [11],
    \padframe/mprj_io_ib_mode_sel [10],
    \padframe/mprj_io_ib_mode_sel [9],
    \padframe/mprj_io_ib_mode_sel [8],
    \padframe/mprj_io_ib_mode_sel [7],
    \padframe/mprj_io_ib_mode_sel [6],
    \padframe/mprj_io_ib_mode_sel [5],
    \padframe/mprj_io_ib_mode_sel [4],
    \padframe/mprj_io_ib_mode_sel [3],
    \padframe/mprj_io_ib_mode_sel [2],
    \padframe/mprj_io_ib_mode_sel [1],
    \padframe/mprj_io_ib_mode_sel [0]}),
    .mprj_io_in({\padframe/mprj_io_in [37],
    \padframe/mprj_io_in [36],
    \padframe/mprj_io_in [35],
    \padframe/mprj_io_in [34],
    \padframe/mprj_io_in [33],
    \padframe/mprj_io_in [32],
    \padframe/mprj_io_in [31],
    \padframe/mprj_io_in [30],
    \padframe/mprj_io_in [29],
    \padframe/mprj_io_in [28],
    \padframe/mprj_io_in [27],
    \padframe/mprj_io_in [26],
    \padframe/mprj_io_in [25],
    \padframe/mprj_io_in [24],
    \padframe/mprj_io_in [23],
    \padframe/mprj_io_in [22],
    \padframe/mprj_io_in [21],
    \padframe/mprj_io_in [20],
    \padframe/mprj_io_in [19],
    \padframe/mprj_io_in [18],
    \padframe/mprj_io_in [17],
    \padframe/mprj_io_in [16],
    \padframe/mprj_io_in [15],
    \padframe/mprj_io_in [14],
    \padframe/mprj_io_in [13],
    \padframe/mprj_io_in [12],
    \padframe/mprj_io_in [11],
    \padframe/mprj_io_in [10],
    \padframe/mprj_io_in [9],
    \padframe/mprj_io_in [8],
    \padframe/mprj_io_in [7],
    \padframe/mprj_io_in [6],
    \padframe/mprj_io_in [5],
    \padframe/mprj_io_in [4],
    \padframe/mprj_io_in [3],
    \padframe/mprj_io_in [2],
    \padframe/mprj_io_in [1],
    \padframe/mprj_io_in [0]}),
    .mprj_io_inp_dis({\padframe/mprj_io_inp_dis [37],
    \padframe/mprj_io_inp_dis [36],
    \padframe/mprj_io_inp_dis [35],
    \padframe/mprj_io_inp_dis [34],
    \padframe/mprj_io_inp_dis [33],
    \padframe/mprj_io_inp_dis [32],
    \padframe/mprj_io_inp_dis [31],
    \padframe/mprj_io_inp_dis [30],
    \padframe/mprj_io_inp_dis [29],
    \padframe/mprj_io_inp_dis [28],
    \padframe/mprj_io_inp_dis [27],
    \padframe/mprj_io_inp_dis [26],
    \padframe/mprj_io_inp_dis [25],
    \padframe/mprj_io_inp_dis [24],
    \padframe/mprj_io_inp_dis [23],
    \padframe/mprj_io_inp_dis [22],
    \padframe/mprj_io_inp_dis [21],
    \padframe/mprj_io_inp_dis [20],
    \padframe/mprj_io_inp_dis [19],
    \padframe/mprj_io_inp_dis [18],
    \padframe/mprj_io_inp_dis [17],
    \padframe/mprj_io_inp_dis [16],
    \padframe/mprj_io_inp_dis [15],
    \padframe/mprj_io_inp_dis [14],
    \padframe/mprj_io_inp_dis [13],
    \padframe/mprj_io_inp_dis [12],
    \padframe/mprj_io_inp_dis [11],
    \padframe/mprj_io_inp_dis [10],
    \padframe/mprj_io_inp_dis [9],
    \padframe/mprj_io_inp_dis [8],
    \padframe/mprj_io_inp_dis [7],
    \padframe/mprj_io_inp_dis [6],
    \padframe/mprj_io_inp_dis [5],
    \padframe/mprj_io_inp_dis [4],
    \padframe/mprj_io_inp_dis [3],
    \padframe/mprj_io_inp_dis [2],
    \padframe/mprj_io_inp_dis [1],
    \padframe/mprj_io_inp_dis [0]}),
    .mprj_io_oeb({\padframe/mprj_io_oeb [37],
    \padframe/mprj_io_oeb [36],
    \padframe/mprj_io_oeb [35],
    \padframe/mprj_io_oeb [34],
    \padframe/mprj_io_oeb [33],
    \padframe/mprj_io_oeb [32],
    \padframe/mprj_io_oeb [31],
    \padframe/mprj_io_oeb [30],
    \padframe/mprj_io_oeb [29],
    \padframe/mprj_io_oeb [28],
    \padframe/mprj_io_oeb [27],
    \padframe/mprj_io_oeb [26],
    \padframe/mprj_io_oeb [25],
    \padframe/mprj_io_oeb [24],
    \padframe/mprj_io_oeb [23],
    \padframe/mprj_io_oeb [22],
    \padframe/mprj_io_oeb [21],
    \padframe/mprj_io_oeb [20],
    \padframe/mprj_io_oeb [19],
    \padframe/mprj_io_oeb [18],
    \padframe/mprj_io_oeb [17],
    \padframe/mprj_io_oeb [16],
    \padframe/mprj_io_oeb [15],
    \padframe/mprj_io_oeb [14],
    \padframe/mprj_io_oeb [13],
    \padframe/mprj_io_oeb [12],
    \padframe/mprj_io_oeb [11],
    \padframe/mprj_io_oeb [10],
    \padframe/mprj_io_oeb [9],
    \padframe/mprj_io_oeb [8],
    \padframe/mprj_io_oeb [7],
    \padframe/mprj_io_oeb [6],
    \padframe/mprj_io_oeb [5],
    \padframe/mprj_io_oeb [4],
    \padframe/mprj_io_oeb [3],
    \padframe/mprj_io_oeb [2],
    \padframe/mprj_io_oeb [1],
    \padframe/mprj_io_oeb [0]}),
    .mprj_io_out({\padframe/mprj_io_out [37],
    \padframe/mprj_io_out [36],
    \padframe/mprj_io_out [35],
    \padframe/mprj_io_out [34],
    \padframe/mprj_io_out [33],
    \padframe/mprj_io_out [32],
    \padframe/mprj_io_out [31],
    \padframe/mprj_io_out [30],
    \padframe/mprj_io_out [29],
    \padframe/mprj_io_out [28],
    \padframe/mprj_io_out [27],
    \padframe/mprj_io_out [26],
    \padframe/mprj_io_out [25],
    \padframe/mprj_io_out [24],
    \padframe/mprj_io_out [23],
    \padframe/mprj_io_out [22],
    \padframe/mprj_io_out [21],
    \padframe/mprj_io_out [20],
    \padframe/mprj_io_out [19],
    \padframe/mprj_io_out [18],
    \padframe/mprj_io_out [17],
    \padframe/mprj_io_out [16],
    \padframe/mprj_io_out [15],
    \padframe/mprj_io_out [14],
    \padframe/mprj_io_out [13],
    \padframe/mprj_io_out [12],
    \padframe/mprj_io_out [11],
    \padframe/mprj_io_out [10],
    \padframe/mprj_io_out [9],
    \padframe/mprj_io_out [8],
    \padframe/mprj_io_out [7],
    \padframe/mprj_io_out [6],
    \padframe/mprj_io_out [5],
    \padframe/mprj_io_out [4],
    \padframe/mprj_io_out [3],
    \padframe/mprj_io_out [2],
    \padframe/mprj_io_out [1],
    \padframe/mprj_io_out [0]}),
    .mprj_io_slow_sel({\padframe/mprj_io_slow_sel [37],
    \padframe/mprj_io_slow_sel [36],
    \padframe/mprj_io_slow_sel [35],
    \padframe/mprj_io_slow_sel [34],
    \padframe/mprj_io_slow_sel [33],
    \padframe/mprj_io_slow_sel [32],
    \padframe/mprj_io_slow_sel [31],
    \padframe/mprj_io_slow_sel [30],
    \padframe/mprj_io_slow_sel [29],
    \padframe/mprj_io_slow_sel [28],
    \padframe/mprj_io_slow_sel [27],
    \padframe/mprj_io_slow_sel [26],
    \padframe/mprj_io_slow_sel [25],
    \padframe/mprj_io_slow_sel [24],
    \padframe/mprj_io_slow_sel [23],
    \padframe/mprj_io_slow_sel [22],
    \padframe/mprj_io_slow_sel [21],
    \padframe/mprj_io_slow_sel [20],
    \padframe/mprj_io_slow_sel [19],
    \padframe/mprj_io_slow_sel [18],
    \padframe/mprj_io_slow_sel [17],
    \padframe/mprj_io_slow_sel [16],
    \padframe/mprj_io_slow_sel [15],
    \padframe/mprj_io_slow_sel [14],
    \padframe/mprj_io_slow_sel [13],
    \padframe/mprj_io_slow_sel [12],
    \padframe/mprj_io_slow_sel [11],
    \padframe/mprj_io_slow_sel [10],
    \padframe/mprj_io_slow_sel [9],
    \padframe/mprj_io_slow_sel [8],
    \padframe/mprj_io_slow_sel [7],
    \padframe/mprj_io_slow_sel [6],
    \padframe/mprj_io_slow_sel [5],
    \padframe/mprj_io_slow_sel [4],
    \padframe/mprj_io_slow_sel [3],
    \padframe/mprj_io_slow_sel [2],
    \padframe/mprj_io_slow_sel [1],
    \padframe/mprj_io_slow_sel [0]}),
    .mprj_io_vtrip_sel({\padframe/mprj_io_vtrip_sel [37],
    \padframe/mprj_io_vtrip_sel [36],
    \padframe/mprj_io_vtrip_sel [35],
    \padframe/mprj_io_vtrip_sel [34],
    \padframe/mprj_io_vtrip_sel [33],
    \padframe/mprj_io_vtrip_sel [32],
    \padframe/mprj_io_vtrip_sel [31],
    \padframe/mprj_io_vtrip_sel [30],
    \padframe/mprj_io_vtrip_sel [29],
    \padframe/mprj_io_vtrip_sel [28],
    \padframe/mprj_io_vtrip_sel [27],
    \padframe/mprj_io_vtrip_sel [26],
    \padframe/mprj_io_vtrip_sel [25],
    \padframe/mprj_io_vtrip_sel [24],
    \padframe/mprj_io_vtrip_sel [23],
    \padframe/mprj_io_vtrip_sel [22],
    \padframe/mprj_io_vtrip_sel [21],
    \padframe/mprj_io_vtrip_sel [20],
    \padframe/mprj_io_vtrip_sel [19],
    \padframe/mprj_io_vtrip_sel [18],
    \padframe/mprj_io_vtrip_sel [17],
    \padframe/mprj_io_vtrip_sel [16],
    \padframe/mprj_io_vtrip_sel [15],
    \padframe/mprj_io_vtrip_sel [14],
    \padframe/mprj_io_vtrip_sel [13],
    \padframe/mprj_io_vtrip_sel [12],
    \padframe/mprj_io_vtrip_sel [11],
    \padframe/mprj_io_vtrip_sel [10],
    \padframe/mprj_io_vtrip_sel [9],
    \padframe/mprj_io_vtrip_sel [8],
    \padframe/mprj_io_vtrip_sel [7],
    \padframe/mprj_io_vtrip_sel [6],
    \padframe/mprj_io_vtrip_sel [5],
    \padframe/mprj_io_vtrip_sel [4],
    \padframe/mprj_io_vtrip_sel [3],
    \padframe/mprj_io_vtrip_sel [2],
    \padframe/mprj_io_vtrip_sel [1],
    \padframe/mprj_io_vtrip_sel [0]}));
endmodule
