magic
tech sky130A
magscale 1 2
timestamp 1638030917
<< locali >>
rect 7941 7395 7975 8177
rect 7941 5491 7975 7157
rect 7941 119 7975 2805
<< viali >>
rect 7941 8177 7975 8211
rect 6929 7361 6963 7395
rect 7941 7361 7975 7395
rect 7021 7157 7055 7191
rect 7941 7157 7975 7191
rect 6469 6953 6503 6987
rect 1593 6817 1627 6851
rect 4169 6817 4203 6851
rect 6929 6817 6963 6851
rect 2237 6749 2271 6783
rect 2789 6749 2823 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 5825 6749 5859 6783
rect 5733 6613 5767 6647
rect 1593 6273 1627 6307
rect 1869 6273 1903 6307
rect 3249 6273 3283 6307
rect 6653 6273 6687 6307
rect 1501 6205 1535 6239
rect 2329 6205 2363 6239
rect 7021 5865 7055 5899
rect 1593 5661 1627 5695
rect 6745 5661 6779 5695
rect 6469 5593 6503 5627
rect 6561 5525 6595 5559
rect 7941 5457 7975 5491
rect 6469 4981 6503 5015
rect 1777 4777 1811 4811
rect 6469 4777 6503 4811
rect 6929 4777 6963 4811
rect 2421 4573 2455 4607
rect 1501 4165 1535 4199
rect 1593 4165 1627 4199
rect 1777 4097 1811 4131
rect 2605 4097 2639 4131
rect 6837 4097 6871 4131
rect 7113 4097 7147 4131
rect 5825 4029 5859 4063
rect 6837 3961 6871 3995
rect 2053 3893 2087 3927
rect 6469 3689 6503 3723
rect 1593 3485 1627 3519
rect 3985 3145 4019 3179
rect 2329 3009 2363 3043
rect 3801 3009 3835 3043
rect 7113 3009 7147 3043
rect 1961 2941 1995 2975
rect 4261 2805 4295 2839
rect 7021 2805 7055 2839
rect 7941 2805 7975 2839
rect 5181 2601 5215 2635
rect 2237 2465 2271 2499
rect 1593 2397 1627 2431
rect 2881 2397 2915 2431
rect 5825 2397 5859 2431
rect 6929 2397 6963 2431
rect 7021 2261 7055 2295
rect 2605 1921 2639 1955
rect 4077 1921 4111 1955
rect 6377 1921 6411 1955
rect 6561 1921 6595 1955
rect 2237 1853 2271 1887
rect 5273 1853 5307 1887
rect 6745 1853 6779 1887
rect 4261 1785 4295 1819
rect 4537 1785 4571 1819
rect 1593 1717 1627 1751
rect 3249 1513 3283 1547
rect 5181 1513 5215 1547
rect 3985 1377 4019 1411
rect 7113 1377 7147 1411
rect 7941 85 7975 119
<< metal1 >>
rect 7926 8208 7932 8220
rect 7887 8180 7932 8208
rect 7926 8168 7932 8180
rect 7984 8168 7990 8220
rect 1104 7642 7820 7664
rect 1104 7590 3150 7642
rect 3202 7590 3214 7642
rect 3266 7590 3278 7642
rect 3330 7590 3342 7642
rect 3394 7590 3406 7642
rect 3458 7590 7150 7642
rect 7202 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7820 7642
rect 1104 7568 7820 7590
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6512 7364 6929 7392
rect 6512 7352 6518 7364
rect 6917 7361 6929 7364
rect 6963 7392 6975 7395
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 6963 7364 7941 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 7055 7160 7941 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7929 7157 7941 7160
rect 7975 7157 7987 7191
rect 7929 7151 7987 7157
rect 1104 7098 7820 7120
rect 1104 7046 1150 7098
rect 1202 7046 1214 7098
rect 1266 7046 1278 7098
rect 1330 7046 1342 7098
rect 1394 7046 1406 7098
rect 1458 7046 5150 7098
rect 5202 7046 5214 7098
rect 5266 7046 5278 7098
rect 5330 7046 5342 7098
rect 5394 7046 5406 7098
rect 5458 7046 7820 7098
rect 1104 7024 7820 7046
rect 6454 6984 6460 6996
rect 6415 6956 6460 6984
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 4154 6848 4160 6860
rect 3108 6820 4016 6848
rect 4115 6820 4160 6848
rect 3108 6808 3114 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2590 6780 2596 6792
rect 2271 6752 2596 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2590 6740 2596 6752
rect 2648 6780 2654 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2648 6752 2789 6780
rect 2648 6740 2654 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 3786 6780 3792 6792
rect 3747 6752 3792 6780
rect 2777 6743 2835 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3988 6789 4016 6820
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6880 6820 6929 6848
rect 6880 6808 6886 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 8386 6780 8392 6792
rect 5859 6752 8392 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 6932 6724 6960 6752
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 6914 6672 6920 6724
rect 6972 6672 6978 6724
rect 5718 6644 5724 6656
rect 5679 6616 5724 6644
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 1104 6554 7820 6576
rect 1104 6502 3150 6554
rect 3202 6502 3214 6554
rect 3266 6502 3278 6554
rect 3330 6502 3342 6554
rect 3394 6502 3406 6554
rect 3458 6502 7150 6554
rect 7202 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7820 6554
rect 1104 6480 7820 6502
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 1486 6236 1492 6248
rect 1447 6208 1492 6236
rect 1486 6196 1492 6208
rect 1544 6196 1550 6248
rect 1872 6236 1900 6267
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3108 6276 3249 6304
rect 3108 6264 3114 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 6914 6304 6920 6316
rect 6687 6276 6920 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 1872 6208 2329 6236
rect 2317 6205 2329 6208
rect 2363 6236 2375 6239
rect 4798 6236 4804 6248
rect 2363 6208 4804 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 1104 6010 7820 6032
rect 1104 5958 1150 6010
rect 1202 5958 1214 6010
rect 1266 5958 1278 6010
rect 1330 5958 1342 6010
rect 1394 5958 1406 6010
rect 1458 5958 5150 6010
rect 5202 5958 5214 6010
rect 5266 5958 5278 6010
rect 5330 5958 5342 6010
rect 5394 5958 5406 6010
rect 5458 5958 7820 6010
rect 1104 5936 7820 5958
rect 7006 5896 7012 5908
rect 6967 5868 7012 5896
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 6822 5692 6828 5704
rect 6779 5664 6828 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6454 5624 6460 5636
rect 6415 5596 6460 5624
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6420 5528 6561 5556
rect 6420 5516 6426 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 7926 5488 7932 5500
rect 1104 5466 7820 5488
rect 1104 5414 3150 5466
rect 3202 5414 3214 5466
rect 3266 5414 3278 5466
rect 3330 5414 3342 5466
rect 3394 5414 3406 5466
rect 3458 5414 7150 5466
rect 7202 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7820 5466
rect 7887 5460 7932 5488
rect 7926 5448 7932 5460
rect 7984 5448 7990 5500
rect 1104 5392 7820 5414
rect 14 5312 20 5364
rect 72 5352 78 5364
rect 5718 5352 5724 5364
rect 72 5324 5724 5352
rect 72 5312 78 5324
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6420 4984 6469 5012
rect 6420 4972 6426 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 1104 4922 7820 4944
rect 1104 4870 1150 4922
rect 1202 4870 1214 4922
rect 1266 4870 1278 4922
rect 1330 4870 1342 4922
rect 1394 4870 1406 4922
rect 1458 4870 5150 4922
rect 5202 4870 5214 4922
rect 5266 4870 5278 4922
rect 5330 4870 5342 4922
rect 5394 4870 5406 4922
rect 5458 4870 7820 4922
rect 1104 4848 7820 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1946 4808 1952 4820
rect 1811 4780 1952 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7742 4808 7748 4820
rect 6972 4780 7748 4808
rect 6972 4768 6978 4780
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 1544 4576 2421 4604
rect 1544 4564 1550 4576
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 1104 4378 7820 4400
rect 1104 4326 3150 4378
rect 3202 4326 3214 4378
rect 3266 4326 3278 4378
rect 3330 4326 3342 4378
rect 3394 4326 3406 4378
rect 3458 4326 7150 4378
rect 7202 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7820 4378
rect 1104 4304 7820 4326
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 5810 4264 5816 4276
rect 4948 4236 5816 4264
rect 4948 4224 4954 4236
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 658 4156 664 4208
rect 716 4196 722 4208
rect 1486 4196 1492 4208
rect 716 4168 1492 4196
rect 716 4156 722 4168
rect 1486 4156 1492 4168
rect 1544 4156 1550 4208
rect 1581 4199 1639 4205
rect 1581 4165 1593 4199
rect 1627 4196 1639 4199
rect 2866 4196 2872 4208
rect 1627 4168 2872 4196
rect 1627 4165 1639 4168
rect 1581 4159 1639 4165
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 6454 4196 6460 4208
rect 4120 4168 6460 4196
rect 4120 4156 4126 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6914 4196 6920 4208
rect 6840 4168 6920 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 1946 4128 1952 4140
rect 1811 4100 1952 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2774 4128 2780 4140
rect 2639 4100 2780 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2774 4088 2780 4100
rect 2832 4128 2838 4140
rect 3786 4128 3792 4140
rect 2832 4100 3792 4128
rect 2832 4088 2838 4100
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 6840 4137 6868 4168
rect 6914 4156 6920 4168
rect 6972 4156 6978 4208
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 6825 4091 6883 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 7116 4060 7144 4088
rect 5859 4032 7144 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 1026 3952 1032 4004
rect 1084 3992 1090 4004
rect 6825 3995 6883 4001
rect 6825 3992 6837 3995
rect 1084 3964 6837 3992
rect 1084 3952 1090 3964
rect 6825 3961 6837 3964
rect 6871 3961 6883 3995
rect 6825 3955 6883 3961
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 4982 3924 4988 3936
rect 2087 3896 4988 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 1104 3834 7820 3856
rect 1104 3782 1150 3834
rect 1202 3782 1214 3834
rect 1266 3782 1278 3834
rect 1330 3782 1342 3834
rect 1394 3782 1406 3834
rect 1458 3782 5150 3834
rect 5202 3782 5214 3834
rect 5266 3782 5278 3834
rect 5330 3782 5342 3834
rect 5394 3782 5406 3834
rect 5458 3782 7820 3834
rect 1104 3760 7820 3782
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 14 3544 20 3596
rect 72 3584 78 3596
rect 6362 3584 6368 3596
rect 72 3556 6368 3584
rect 72 3544 78 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2866 3516 2872 3528
rect 1627 3488 2872 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 1104 3290 7820 3312
rect 1104 3238 3150 3290
rect 3202 3238 3214 3290
rect 3266 3238 3278 3290
rect 3330 3238 3342 3290
rect 3394 3238 3406 3290
rect 3458 3238 7150 3290
rect 7202 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7820 3290
rect 1104 3216 7820 3238
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4522 3176 4528 3188
rect 4019 3148 4528 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 2774 3068 2780 3120
rect 2832 3068 2838 3120
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 1636 3012 2329 3040
rect 1636 3000 1642 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 5074 3040 5080 3052
rect 3835 3012 5080 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 7742 3040 7748 3052
rect 7147 3012 7748 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 4212 2808 4261 2836
rect 4212 2796 4218 2808
rect 4249 2805 4261 2808
rect 4295 2805 4307 2839
rect 4249 2799 4307 2805
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7929 2839 7987 2845
rect 7929 2836 7941 2839
rect 7055 2808 7941 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7929 2805 7941 2808
rect 7975 2805 7987 2839
rect 7929 2799 7987 2805
rect 1104 2746 7820 2768
rect 1104 2694 1150 2746
rect 1202 2694 1214 2746
rect 1266 2694 1278 2746
rect 1330 2694 1342 2746
rect 1394 2694 1406 2746
rect 1458 2694 5150 2746
rect 5202 2694 5214 2746
rect 5266 2694 5278 2746
rect 5330 2694 5342 2746
rect 5394 2694 5406 2746
rect 5458 2694 7820 2746
rect 1104 2672 7820 2694
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 5132 2604 5181 2632
rect 5132 2592 5138 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 2004 2468 2237 2496
rect 2004 2456 2010 2468
rect 2225 2465 2237 2468
rect 2271 2496 2283 2499
rect 4246 2496 4252 2508
rect 2271 2468 4252 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2832 2400 2881 2428
rect 2832 2388 2838 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 2869 2391 2927 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6512 2400 6929 2428
rect 6512 2388 6518 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7009 2295 7067 2301
rect 7009 2261 7021 2295
rect 7055 2292 7067 2295
rect 8386 2292 8392 2304
rect 7055 2264 8392 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 1104 2202 7820 2224
rect 1104 2150 3150 2202
rect 3202 2150 3214 2202
rect 3266 2150 3278 2202
rect 3330 2150 3342 2202
rect 3394 2150 3406 2202
rect 3458 2150 7150 2202
rect 7202 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7820 2202
rect 1104 2128 7820 2150
rect 4890 2088 4896 2100
rect 2332 2060 4896 2088
rect 2332 1952 2360 2060
rect 4890 2048 4896 2060
rect 4948 2048 4954 2100
rect 3234 1980 3240 2032
rect 3292 1980 3298 2032
rect 5810 1980 5816 2032
rect 5868 2020 5874 2032
rect 5868 1992 6592 2020
rect 5868 1980 5874 1992
rect 2593 1955 2651 1961
rect 2593 1952 2605 1955
rect 2332 1924 2605 1952
rect 2593 1921 2605 1924
rect 2639 1921 2651 1955
rect 2593 1915 2651 1921
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 4065 1955 4123 1961
rect 4065 1952 4077 1955
rect 3936 1924 4077 1952
rect 3936 1912 3942 1924
rect 4065 1921 4077 1924
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 4430 1912 4436 1964
rect 4488 1952 4494 1964
rect 6564 1961 6592 1992
rect 6365 1955 6423 1961
rect 6365 1952 6377 1955
rect 4488 1924 6377 1952
rect 4488 1912 4494 1924
rect 6365 1921 6377 1924
rect 6411 1921 6423 1955
rect 6365 1915 6423 1921
rect 6549 1955 6607 1961
rect 6549 1921 6561 1955
rect 6595 1921 6607 1955
rect 6549 1915 6607 1921
rect 2225 1887 2283 1893
rect 2225 1884 2237 1887
rect 1596 1856 2237 1884
rect 658 1708 664 1760
rect 716 1748 722 1760
rect 1596 1757 1624 1856
rect 2225 1853 2237 1856
rect 2271 1853 2283 1887
rect 2225 1847 2283 1853
rect 4890 1844 4896 1896
rect 4948 1884 4954 1896
rect 5261 1887 5319 1893
rect 5261 1884 5273 1887
rect 4948 1856 5273 1884
rect 4948 1844 4954 1856
rect 5261 1853 5273 1856
rect 5307 1853 5319 1887
rect 6730 1884 6736 1896
rect 6691 1856 6736 1884
rect 5261 1847 5319 1853
rect 6730 1844 6736 1856
rect 6788 1844 6794 1896
rect 4249 1819 4307 1825
rect 4249 1785 4261 1819
rect 4295 1816 4307 1819
rect 4338 1816 4344 1828
rect 4295 1788 4344 1816
rect 4295 1785 4307 1788
rect 4249 1779 4307 1785
rect 4338 1776 4344 1788
rect 4396 1776 4402 1828
rect 4525 1819 4583 1825
rect 4525 1785 4537 1819
rect 4571 1816 4583 1819
rect 6454 1816 6460 1828
rect 4571 1788 6460 1816
rect 4571 1785 4583 1788
rect 4525 1779 4583 1785
rect 6454 1776 6460 1788
rect 6512 1776 6518 1828
rect 1581 1751 1639 1757
rect 1581 1748 1593 1751
rect 716 1720 1593 1748
rect 716 1708 722 1720
rect 1581 1717 1593 1720
rect 1627 1717 1639 1751
rect 1581 1711 1639 1717
rect 1104 1658 7820 1680
rect 1104 1606 1150 1658
rect 1202 1606 1214 1658
rect 1266 1606 1278 1658
rect 1330 1606 1342 1658
rect 1394 1606 1406 1658
rect 1458 1606 5150 1658
rect 5202 1606 5214 1658
rect 5266 1606 5278 1658
rect 5330 1606 5342 1658
rect 5394 1606 5406 1658
rect 5458 1606 7820 1658
rect 1104 1584 7820 1606
rect 3234 1544 3240 1556
rect 3195 1516 3240 1544
rect 3234 1504 3240 1516
rect 3292 1504 3298 1556
rect 4430 1504 4436 1556
rect 4488 1544 4494 1556
rect 5169 1547 5227 1553
rect 5169 1544 5181 1547
rect 4488 1516 5181 1544
rect 4488 1504 4494 1516
rect 5169 1513 5181 1516
rect 5215 1513 5227 1547
rect 5169 1507 5227 1513
rect 3878 1368 3884 1420
rect 3936 1408 3942 1420
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 3936 1380 3985 1408
rect 3936 1368 3942 1380
rect 3973 1377 3985 1380
rect 4019 1377 4031 1411
rect 3973 1371 4031 1377
rect 7101 1411 7159 1417
rect 7101 1377 7113 1411
rect 7147 1408 7159 1411
rect 7742 1408 7748 1420
rect 7147 1380 7748 1408
rect 7147 1377 7159 1380
rect 7101 1371 7159 1377
rect 7742 1368 7748 1380
rect 7800 1368 7806 1420
rect 1104 1114 7820 1136
rect 1104 1062 3150 1114
rect 3202 1062 3214 1114
rect 3266 1062 3278 1114
rect 3330 1062 3342 1114
rect 3394 1062 3406 1114
rect 3458 1062 7150 1114
rect 7202 1062 7214 1114
rect 7266 1062 7278 1114
rect 7330 1062 7342 1114
rect 7394 1062 7406 1114
rect 7458 1062 7820 1114
rect 1104 1040 7820 1062
rect 7926 116 7932 128
rect 7887 88 7932 116
rect 7926 76 7932 88
rect 7984 76 7990 128
<< via1 >>
rect 7932 8211 7984 8220
rect 7932 8177 7941 8211
rect 7941 8177 7975 8211
rect 7975 8177 7984 8211
rect 7932 8168 7984 8177
rect 3150 7590 3202 7642
rect 3214 7590 3266 7642
rect 3278 7590 3330 7642
rect 3342 7590 3394 7642
rect 3406 7590 3458 7642
rect 7150 7590 7202 7642
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 6460 7352 6512 7404
rect 1150 7046 1202 7098
rect 1214 7046 1266 7098
rect 1278 7046 1330 7098
rect 1342 7046 1394 7098
rect 1406 7046 1458 7098
rect 5150 7046 5202 7098
rect 5214 7046 5266 7098
rect 5278 7046 5330 7098
rect 5342 7046 5394 7098
rect 5406 7046 5458 7098
rect 6460 6987 6512 6996
rect 6460 6953 6469 6987
rect 6469 6953 6503 6987
rect 6503 6953 6512 6987
rect 6460 6944 6512 6953
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 3056 6808 3108 6860
rect 4160 6851 4212 6860
rect 2596 6740 2648 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 6828 6808 6880 6860
rect 8392 6740 8444 6792
rect 6920 6672 6972 6724
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 3150 6502 3202 6554
rect 3214 6502 3266 6554
rect 3278 6502 3330 6554
rect 3342 6502 3394 6554
rect 3406 6502 3458 6554
rect 7150 6502 7202 6554
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 3056 6264 3108 6316
rect 6920 6264 6972 6316
rect 4804 6196 4856 6248
rect 1150 5958 1202 6010
rect 1214 5958 1266 6010
rect 1278 5958 1330 6010
rect 1342 5958 1394 6010
rect 1406 5958 1458 6010
rect 5150 5958 5202 6010
rect 5214 5958 5266 6010
rect 5278 5958 5330 6010
rect 5342 5958 5394 6010
rect 5406 5958 5458 6010
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 6828 5652 6880 5704
rect 6460 5627 6512 5636
rect 6460 5593 6469 5627
rect 6469 5593 6503 5627
rect 6503 5593 6512 5627
rect 6460 5584 6512 5593
rect 6368 5516 6420 5568
rect 7932 5491 7984 5500
rect 3150 5414 3202 5466
rect 3214 5414 3266 5466
rect 3278 5414 3330 5466
rect 3342 5414 3394 5466
rect 3406 5414 3458 5466
rect 7150 5414 7202 5466
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 7932 5457 7941 5491
rect 7941 5457 7975 5491
rect 7975 5457 7984 5491
rect 7932 5448 7984 5457
rect 20 5312 72 5364
rect 5724 5312 5776 5364
rect 6368 4972 6420 5024
rect 1150 4870 1202 4922
rect 1214 4870 1266 4922
rect 1278 4870 1330 4922
rect 1342 4870 1394 4922
rect 1406 4870 1458 4922
rect 5150 4870 5202 4922
rect 5214 4870 5266 4922
rect 5278 4870 5330 4922
rect 5342 4870 5394 4922
rect 5406 4870 5458 4922
rect 1952 4768 2004 4820
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 7748 4768 7800 4820
rect 1492 4564 1544 4616
rect 3150 4326 3202 4378
rect 3214 4326 3266 4378
rect 3278 4326 3330 4378
rect 3342 4326 3394 4378
rect 3406 4326 3458 4378
rect 7150 4326 7202 4378
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 4896 4224 4948 4276
rect 5816 4224 5868 4276
rect 664 4156 716 4208
rect 1492 4199 1544 4208
rect 1492 4165 1501 4199
rect 1501 4165 1535 4199
rect 1535 4165 1544 4199
rect 1492 4156 1544 4165
rect 2872 4156 2924 4208
rect 4068 4156 4120 4208
rect 6460 4156 6512 4208
rect 1952 4088 2004 4140
rect 2780 4088 2832 4140
rect 3792 4088 3844 4140
rect 6920 4156 6972 4208
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 1032 3952 1084 4004
rect 4988 3884 5040 3936
rect 1150 3782 1202 3834
rect 1214 3782 1266 3834
rect 1278 3782 1330 3834
rect 1342 3782 1394 3834
rect 1406 3782 1458 3834
rect 5150 3782 5202 3834
rect 5214 3782 5266 3834
rect 5278 3782 5330 3834
rect 5342 3782 5394 3834
rect 5406 3782 5458 3834
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 20 3544 72 3596
rect 6368 3544 6420 3596
rect 2872 3476 2924 3528
rect 3150 3238 3202 3290
rect 3214 3238 3266 3290
rect 3278 3238 3330 3290
rect 3342 3238 3394 3290
rect 3406 3238 3458 3290
rect 7150 3238 7202 3290
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 4528 3136 4580 3188
rect 2780 3068 2832 3120
rect 1584 3000 1636 3052
rect 5080 3000 5132 3052
rect 7748 3000 7800 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 4160 2796 4212 2848
rect 1150 2694 1202 2746
rect 1214 2694 1266 2746
rect 1278 2694 1330 2746
rect 1342 2694 1394 2746
rect 1406 2694 1458 2746
rect 5150 2694 5202 2746
rect 5214 2694 5266 2746
rect 5278 2694 5330 2746
rect 5342 2694 5394 2746
rect 5406 2694 5458 2746
rect 5080 2592 5132 2644
rect 1952 2456 2004 2508
rect 4252 2456 4304 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2780 2388 2832 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6460 2388 6512 2440
rect 8392 2252 8444 2304
rect 3150 2150 3202 2202
rect 3214 2150 3266 2202
rect 3278 2150 3330 2202
rect 3342 2150 3394 2202
rect 3406 2150 3458 2202
rect 7150 2150 7202 2202
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 4896 2048 4948 2100
rect 3240 1980 3292 2032
rect 5816 1980 5868 2032
rect 3884 1912 3936 1964
rect 4436 1912 4488 1964
rect 664 1708 716 1760
rect 4896 1844 4948 1896
rect 6736 1887 6788 1896
rect 6736 1853 6745 1887
rect 6745 1853 6779 1887
rect 6779 1853 6788 1887
rect 6736 1844 6788 1853
rect 4344 1776 4396 1828
rect 6460 1776 6512 1828
rect 1150 1606 1202 1658
rect 1214 1606 1266 1658
rect 1278 1606 1330 1658
rect 1342 1606 1394 1658
rect 1406 1606 1458 1658
rect 5150 1606 5202 1658
rect 5214 1606 5266 1658
rect 5278 1606 5330 1658
rect 5342 1606 5394 1658
rect 5406 1606 5458 1658
rect 3240 1547 3292 1556
rect 3240 1513 3249 1547
rect 3249 1513 3283 1547
rect 3283 1513 3292 1547
rect 3240 1504 3292 1513
rect 4436 1504 4488 1556
rect 3884 1368 3936 1420
rect 7748 1368 7800 1420
rect 3150 1062 3202 1114
rect 3214 1062 3266 1114
rect 3278 1062 3330 1114
rect 3342 1062 3394 1114
rect 3406 1062 3458 1114
rect 7150 1062 7202 1114
rect 7214 1062 7266 1114
rect 7278 1062 7330 1114
rect 7342 1062 7394 1114
rect 7406 1062 7458 1114
rect 7932 119 7984 128
rect 7932 85 7941 119
rect 7941 85 7975 119
rect 7975 85 7984 119
rect 7932 76 7984 85
<< metal2 >>
rect 18 8200 74 9000
rect 662 8200 718 9000
rect 1950 8200 2006 9000
rect 2594 8200 2650 9000
rect 3238 8200 3294 9000
rect 4066 8936 4122 8945
rect 4122 8894 4292 8922
rect 4066 8871 4122 8880
rect 32 5370 60 8200
rect 20 5364 72 5370
rect 20 5306 72 5312
rect 676 4214 704 8200
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1150 7100 1458 7120
rect 1150 7098 1156 7100
rect 1212 7098 1236 7100
rect 1292 7098 1316 7100
rect 1372 7098 1396 7100
rect 1452 7098 1458 7100
rect 1212 7046 1214 7098
rect 1394 7046 1396 7098
rect 1150 7044 1156 7046
rect 1212 7044 1236 7046
rect 1292 7044 1316 7046
rect 1372 7044 1396 7046
rect 1452 7044 1458 7046
rect 1150 7024 1458 7044
rect 1596 6866 1624 7511
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1492 6248 1544 6254
rect 1490 6216 1492 6225
rect 1544 6216 1546 6225
rect 1490 6151 1546 6160
rect 1150 6012 1458 6032
rect 1150 6010 1156 6012
rect 1212 6010 1236 6012
rect 1292 6010 1316 6012
rect 1372 6010 1396 6012
rect 1452 6010 1458 6012
rect 1212 5958 1214 6010
rect 1394 5958 1396 6010
rect 1150 5956 1156 5958
rect 1212 5956 1236 5958
rect 1292 5956 1316 5958
rect 1372 5956 1396 5958
rect 1452 5956 1458 5958
rect 1150 5936 1458 5956
rect 1596 5710 1624 6258
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5137 1624 5646
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1150 4924 1458 4944
rect 1150 4922 1156 4924
rect 1212 4922 1236 4924
rect 1292 4922 1316 4924
rect 1372 4922 1396 4924
rect 1452 4922 1458 4924
rect 1212 4870 1214 4922
rect 1394 4870 1396 4922
rect 1150 4868 1156 4870
rect 1212 4868 1236 4870
rect 1292 4868 1316 4870
rect 1372 4868 1396 4870
rect 1452 4868 1458 4870
rect 1150 4848 1458 4868
rect 1964 4826 1992 8200
rect 2608 6798 2636 8200
rect 3252 7834 3280 8200
rect 3068 7806 3280 7834
rect 3068 6866 3096 7806
rect 3150 7644 3458 7664
rect 3150 7642 3156 7644
rect 3212 7642 3236 7644
rect 3292 7642 3316 7644
rect 3372 7642 3396 7644
rect 3452 7642 3458 7644
rect 3212 7590 3214 7642
rect 3394 7590 3396 7642
rect 3150 7588 3156 7590
rect 3212 7588 3236 7590
rect 3292 7588 3316 7590
rect 3372 7588 3396 7590
rect 3452 7588 3458 7590
rect 3150 7568 3458 7588
rect 4264 6914 4292 8894
rect 4526 8200 4582 9000
rect 4816 8214 5120 8242
rect 4158 6896 4214 6905
rect 3056 6860 3108 6866
rect 4264 6886 4476 6914
rect 4158 6831 4160 6840
rect 3056 6802 3108 6808
rect 4212 6831 4214 6840
rect 4160 6802 4212 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 3068 6322 3096 6802
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 4342 6760 4398 6769
rect 3150 6556 3458 6576
rect 3150 6554 3156 6556
rect 3212 6554 3236 6556
rect 3292 6554 3316 6556
rect 3372 6554 3396 6556
rect 3452 6554 3458 6556
rect 3212 6502 3214 6554
rect 3394 6502 3396 6554
rect 3150 6500 3156 6502
rect 3212 6500 3236 6502
rect 3292 6500 3316 6502
rect 3372 6500 3396 6502
rect 3452 6500 3458 6502
rect 3150 6480 3458 6500
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3150 5468 3458 5488
rect 3150 5466 3156 5468
rect 3212 5466 3236 5468
rect 3292 5466 3316 5468
rect 3372 5466 3396 5468
rect 3452 5466 3458 5468
rect 3212 5414 3214 5466
rect 3394 5414 3396 5466
rect 3150 5412 3156 5414
rect 3212 5412 3236 5414
rect 3292 5412 3316 5414
rect 3372 5412 3396 5414
rect 3452 5412 3458 5414
rect 3150 5392 3458 5412
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1504 4214 1532 4558
rect 664 4208 716 4214
rect 664 4150 716 4156
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1964 4146 1992 4762
rect 3150 4380 3458 4400
rect 3150 4378 3156 4380
rect 3212 4378 3236 4380
rect 3292 4378 3316 4380
rect 3372 4378 3396 4380
rect 3452 4378 3458 4380
rect 3212 4326 3214 4378
rect 3394 4326 3396 4378
rect 3150 4324 3156 4326
rect 3212 4324 3236 4326
rect 3292 4324 3316 4326
rect 3372 4324 3396 4326
rect 3452 4324 3458 4326
rect 3150 4304 3458 4324
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 1032 4004 1084 4010
rect 1032 3946 1084 3952
rect 20 3596 72 3602
rect 20 3538 72 3544
rect 32 800 60 3538
rect 664 1760 716 1766
rect 664 1702 716 1708
rect 676 800 704 1702
rect 18 0 74 800
rect 662 0 718 800
rect 1044 762 1072 3946
rect 1150 3836 1458 3856
rect 1150 3834 1156 3836
rect 1212 3834 1236 3836
rect 1292 3834 1316 3836
rect 1372 3834 1396 3836
rect 1452 3834 1458 3836
rect 1212 3782 1214 3834
rect 1394 3782 1396 3834
rect 1150 3780 1156 3782
rect 1212 3780 1236 3782
rect 1292 3780 1316 3782
rect 1372 3780 1396 3782
rect 1452 3780 1458 3782
rect 1150 3760 1458 3780
rect 2792 3505 2820 4082
rect 2884 3534 2912 4150
rect 3804 4146 3832 6734
rect 4342 6695 4398 6704
rect 4068 4208 4120 4214
rect 4066 4176 4068 4185
rect 4120 4176 4122 4185
rect 3792 4140 3844 4146
rect 4066 4111 4122 4120
rect 3792 4082 3844 4088
rect 2872 3528 2924 3534
rect 2778 3496 2834 3505
rect 2872 3470 2924 3476
rect 2778 3431 2834 3440
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1150 2748 1458 2768
rect 1150 2746 1156 2748
rect 1212 2746 1236 2748
rect 1292 2746 1316 2748
rect 1372 2746 1396 2748
rect 1452 2746 1458 2748
rect 1212 2694 1214 2746
rect 1394 2694 1396 2746
rect 1150 2692 1156 2694
rect 1212 2692 1236 2694
rect 1292 2692 1316 2694
rect 1372 2692 1396 2694
rect 1452 2692 1458 2694
rect 1150 2672 1458 2692
rect 1596 2446 1624 2994
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1964 2514 1992 2926
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2792 2446 2820 3062
rect 1584 2440 1636 2446
rect 2780 2440 2832 2446
rect 1584 2382 1636 2388
rect 2608 2388 2780 2394
rect 2608 2382 2832 2388
rect 1150 1660 1458 1680
rect 1150 1658 1156 1660
rect 1212 1658 1236 1660
rect 1292 1658 1316 1660
rect 1372 1658 1396 1660
rect 1452 1658 1458 1660
rect 1212 1606 1214 1658
rect 1394 1606 1396 1658
rect 1150 1604 1156 1606
rect 1212 1604 1236 1606
rect 1292 1604 1316 1606
rect 1372 1604 1396 1606
rect 1452 1604 1458 1606
rect 1150 1584 1458 1604
rect 1228 870 1348 898
rect 1228 762 1256 870
rect 1320 800 1348 870
rect 1044 734 1256 762
rect 1306 0 1362 800
rect 1596 785 1624 2382
rect 2608 2366 2820 2382
rect 2608 800 2636 2366
rect 2884 1465 2912 3470
rect 3150 3292 3458 3312
rect 3150 3290 3156 3292
rect 3212 3290 3236 3292
rect 3292 3290 3316 3292
rect 3372 3290 3396 3292
rect 3452 3290 3458 3292
rect 3212 3238 3214 3290
rect 3394 3238 3396 3290
rect 3150 3236 3156 3238
rect 3212 3236 3236 3238
rect 3292 3236 3316 3238
rect 3372 3236 3396 3238
rect 3452 3236 3458 3238
rect 3150 3216 3458 3236
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3150 2204 3458 2224
rect 3150 2202 3156 2204
rect 3212 2202 3236 2204
rect 3292 2202 3316 2204
rect 3372 2202 3396 2204
rect 3452 2202 3458 2204
rect 3212 2150 3214 2202
rect 3394 2150 3396 2202
rect 3150 2148 3156 2150
rect 3212 2148 3236 2150
rect 3292 2148 3316 2150
rect 3372 2148 3396 2150
rect 3452 2148 3458 2150
rect 3150 2128 3458 2148
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 4066 2000 4122 2009
rect 3252 1562 3280 1974
rect 3884 1964 3936 1970
rect 4172 1986 4200 2790
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4264 2417 4292 2450
rect 4250 2408 4306 2417
rect 4250 2343 4306 2352
rect 4122 1958 4200 1986
rect 4066 1935 4122 1944
rect 3884 1906 3936 1912
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 1306 3280 1498
rect 3896 1426 3924 1906
rect 4356 1834 4384 6695
rect 4448 1970 4476 6886
rect 4540 3194 4568 8200
rect 4816 6254 4844 8214
rect 5092 8106 5120 8214
rect 5170 8200 5226 9000
rect 5814 8200 5870 9000
rect 7102 8200 7158 9000
rect 7746 8200 7802 9000
rect 7930 8256 7986 8265
rect 8390 8200 8446 9000
rect 5184 8106 5212 8200
rect 5092 8078 5212 8106
rect 5150 7100 5458 7120
rect 5150 7098 5156 7100
rect 5212 7098 5236 7100
rect 5292 7098 5316 7100
rect 5372 7098 5396 7100
rect 5452 7098 5458 7100
rect 5212 7046 5214 7098
rect 5394 7046 5396 7098
rect 5150 7044 5156 7046
rect 5212 7044 5236 7046
rect 5292 7044 5316 7046
rect 5372 7044 5396 7046
rect 5452 7044 5458 7046
rect 5150 7024 5458 7044
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5150 6012 5458 6032
rect 5150 6010 5156 6012
rect 5212 6010 5236 6012
rect 5292 6010 5316 6012
rect 5372 6010 5396 6012
rect 5452 6010 5458 6012
rect 5212 5958 5214 6010
rect 5394 5958 5396 6010
rect 5150 5956 5156 5958
rect 5212 5956 5236 5958
rect 5292 5956 5316 5958
rect 5372 5956 5396 5958
rect 5452 5956 5458 5958
rect 5150 5936 5458 5956
rect 5736 5370 5764 6598
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5150 4924 5458 4944
rect 5150 4922 5156 4924
rect 5212 4922 5236 4924
rect 5292 4922 5316 4924
rect 5372 4922 5396 4924
rect 5452 4922 5458 4924
rect 5212 4870 5214 4922
rect 5394 4870 5396 4922
rect 5150 4868 5156 4870
rect 5212 4868 5236 4870
rect 5292 4868 5316 4870
rect 5372 4868 5396 4870
rect 5452 4868 5458 4870
rect 5150 4848 5458 4868
rect 5828 4282 5856 8200
rect 7116 7834 7144 8200
rect 7024 7806 7144 7834
rect 6826 7440 6882 7449
rect 6460 7404 6512 7410
rect 6826 7375 6882 7384
rect 6460 7346 6512 7352
rect 6472 7002 6500 7346
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6840 6866 6868 7375
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 5710 6868 6802
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6322 6960 6666
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7024 5914 7052 7806
rect 7150 7644 7458 7664
rect 7150 7642 7156 7644
rect 7212 7642 7236 7644
rect 7292 7642 7316 7644
rect 7372 7642 7396 7644
rect 7452 7642 7458 7644
rect 7212 7590 7214 7642
rect 7394 7590 7396 7642
rect 7150 7588 7156 7590
rect 7212 7588 7236 7590
rect 7292 7588 7316 7590
rect 7372 7588 7396 7590
rect 7452 7588 7458 7590
rect 7150 7568 7458 7588
rect 7150 6556 7458 6576
rect 7150 6554 7156 6556
rect 7212 6554 7236 6556
rect 7292 6554 7316 6556
rect 7372 6554 7396 6556
rect 7452 6554 7458 6556
rect 7212 6502 7214 6554
rect 7394 6502 7396 6554
rect 7150 6500 7156 6502
rect 7212 6500 7236 6502
rect 7292 6500 7316 6502
rect 7372 6500 7396 6502
rect 7452 6500 7458 6502
rect 7150 6480 7458 6500
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 5030 6408 5510
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4908 2106 4936 4218
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4344 1828 4396 1834
rect 4344 1770 4396 1776
rect 4448 1562 4476 1906
rect 4908 1902 4936 2042
rect 4896 1896 4948 1902
rect 4896 1838 4948 1844
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 5000 1442 5028 3878
rect 5150 3836 5458 3856
rect 5150 3834 5156 3836
rect 5212 3834 5236 3836
rect 5292 3834 5316 3836
rect 5372 3834 5396 3836
rect 5452 3834 5458 3836
rect 5212 3782 5214 3834
rect 5394 3782 5396 3834
rect 5150 3780 5156 3782
rect 5212 3780 5236 3782
rect 5292 3780 5316 3782
rect 5372 3780 5396 3782
rect 5452 3780 5458 3782
rect 5150 3760 5458 3780
rect 6380 3602 6408 4966
rect 6472 4865 6500 5578
rect 7150 5468 7458 5488
rect 7150 5466 7156 5468
rect 7212 5466 7236 5468
rect 7292 5466 7316 5468
rect 7372 5466 7396 5468
rect 7452 5466 7458 5468
rect 7212 5414 7214 5466
rect 7394 5414 7396 5466
rect 7150 5412 7156 5414
rect 7212 5412 7236 5414
rect 7292 5412 7316 5414
rect 7372 5412 7396 5414
rect 7452 5412 7458 5414
rect 7150 5392 7458 5412
rect 6458 4856 6514 4865
rect 7760 4826 7788 8200
rect 7930 8191 7932 8200
rect 7984 8191 7986 8200
rect 7932 8162 7984 8168
rect 8404 6798 8432 8200
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 7930 5536 7986 5545
rect 7930 5471 7932 5480
rect 7984 5471 7986 5480
rect 7932 5442 7984 5448
rect 6458 4791 6460 4800
rect 6512 4791 6514 4800
rect 6920 4820 6972 4826
rect 6460 4762 6512 4768
rect 6920 4762 6972 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 6472 4731 6500 4762
rect 6932 4214 6960 4762
rect 7150 4380 7458 4400
rect 7150 4378 7156 4380
rect 7212 4378 7236 4380
rect 7292 4378 7316 4380
rect 7372 4378 7396 4380
rect 7452 4378 7458 4380
rect 7212 4326 7214 4378
rect 7394 4326 7396 4378
rect 7150 4324 7156 4326
rect 7212 4324 7236 4326
rect 7292 4324 7316 4326
rect 7372 4324 7396 4326
rect 7452 4324 7458 4326
rect 7150 4304 7458 4324
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 7102 4176 7158 4185
rect 6472 3738 6500 4150
rect 7102 4111 7104 4120
rect 7156 4111 7158 4120
rect 7104 4082 7156 4088
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5092 2961 5120 2994
rect 5078 2952 5134 2961
rect 5078 2887 5134 2896
rect 5092 2650 5120 2887
rect 5150 2748 5458 2768
rect 5150 2746 5156 2748
rect 5212 2746 5236 2748
rect 5292 2746 5316 2748
rect 5372 2746 5396 2748
rect 5452 2746 5458 2748
rect 5212 2694 5214 2746
rect 5394 2694 5396 2746
rect 5150 2692 5156 2694
rect 5212 2692 5236 2694
rect 5292 2692 5316 2694
rect 5372 2692 5396 2694
rect 5452 2692 5458 2694
rect 5150 2672 5458 2692
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 6472 2446 6500 3674
rect 7150 3292 7458 3312
rect 7150 3290 7156 3292
rect 7212 3290 7236 3292
rect 7292 3290 7316 3292
rect 7372 3290 7396 3292
rect 7452 3290 7458 3292
rect 7212 3238 7214 3290
rect 7394 3238 7396 3290
rect 7150 3236 7156 3238
rect 7212 3236 7236 3238
rect 7292 3236 7316 3238
rect 7372 3236 7396 3238
rect 7452 3236 7458 3238
rect 7150 3216 7458 3236
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 5828 2038 5856 2382
rect 7150 2204 7458 2224
rect 7150 2202 7156 2204
rect 7212 2202 7236 2204
rect 7292 2202 7316 2204
rect 7372 2202 7396 2204
rect 7452 2202 7458 2204
rect 7212 2150 7214 2202
rect 7394 2150 7396 2202
rect 7150 2148 7156 2150
rect 7212 2148 7236 2150
rect 7292 2148 7316 2150
rect 7372 2148 7396 2150
rect 7452 2148 7458 2150
rect 7150 2128 7458 2148
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 5150 1660 5458 1680
rect 5150 1658 5156 1660
rect 5212 1658 5236 1660
rect 5292 1658 5316 1660
rect 5372 1658 5396 1660
rect 5452 1658 5458 1660
rect 5212 1606 5214 1658
rect 5394 1606 5396 1658
rect 5150 1604 5156 1606
rect 5212 1604 5236 1606
rect 5292 1604 5316 1606
rect 5372 1604 5396 1606
rect 5452 1604 5458 1606
rect 5150 1584 5458 1604
rect 3884 1420 3936 1426
rect 5000 1414 5212 1442
rect 3884 1362 3936 1368
rect 3068 1278 3280 1306
rect 3068 898 3096 1278
rect 3150 1116 3458 1136
rect 3150 1114 3156 1116
rect 3212 1114 3236 1116
rect 3292 1114 3316 1116
rect 3372 1114 3396 1116
rect 3452 1114 3458 1116
rect 3212 1062 3214 1114
rect 3394 1062 3396 1114
rect 3150 1060 3156 1062
rect 3212 1060 3236 1062
rect 3292 1060 3316 1062
rect 3372 1060 3396 1062
rect 3452 1060 3458 1062
rect 3150 1040 3458 1060
rect 3068 870 3280 898
rect 3252 800 3280 870
rect 3896 800 3924 1362
rect 5184 800 5212 1414
rect 5828 800 5856 1974
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6460 1828 6512 1834
rect 6460 1770 6512 1776
rect 6472 800 6500 1770
rect 6748 1465 6776 1838
rect 6734 1456 6790 1465
rect 7760 1426 7788 2994
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 6734 1391 6790 1400
rect 7748 1420 7800 1426
rect 7748 1362 7800 1368
rect 7150 1116 7458 1136
rect 7150 1114 7156 1116
rect 7212 1114 7236 1116
rect 7292 1114 7316 1116
rect 7372 1114 7396 1116
rect 7452 1114 7458 1116
rect 7212 1062 7214 1114
rect 7394 1062 7396 1114
rect 7150 1060 7156 1062
rect 7212 1060 7236 1062
rect 7292 1060 7316 1062
rect 7372 1060 7396 1062
rect 7452 1060 7458 1062
rect 7150 1040 7458 1060
rect 7760 800 7788 1362
rect 8404 800 8432 2246
rect 1582 776 1638 785
rect 1582 711 1638 720
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 7932 128 7984 134
rect 7930 96 7932 105
rect 7984 96 7986 105
rect 7930 31 7986 40
rect 8390 0 8446 800
<< via2 >>
rect 4066 8880 4122 8936
rect 1582 7520 1638 7576
rect 1156 7098 1212 7100
rect 1236 7098 1292 7100
rect 1316 7098 1372 7100
rect 1396 7098 1452 7100
rect 1156 7046 1202 7098
rect 1202 7046 1212 7098
rect 1236 7046 1266 7098
rect 1266 7046 1278 7098
rect 1278 7046 1292 7098
rect 1316 7046 1330 7098
rect 1330 7046 1342 7098
rect 1342 7046 1372 7098
rect 1396 7046 1406 7098
rect 1406 7046 1452 7098
rect 1156 7044 1212 7046
rect 1236 7044 1292 7046
rect 1316 7044 1372 7046
rect 1396 7044 1452 7046
rect 1490 6196 1492 6216
rect 1492 6196 1544 6216
rect 1544 6196 1546 6216
rect 1490 6160 1546 6196
rect 1156 6010 1212 6012
rect 1236 6010 1292 6012
rect 1316 6010 1372 6012
rect 1396 6010 1452 6012
rect 1156 5958 1202 6010
rect 1202 5958 1212 6010
rect 1236 5958 1266 6010
rect 1266 5958 1278 6010
rect 1278 5958 1292 6010
rect 1316 5958 1330 6010
rect 1330 5958 1342 6010
rect 1342 5958 1372 6010
rect 1396 5958 1406 6010
rect 1406 5958 1452 6010
rect 1156 5956 1212 5958
rect 1236 5956 1292 5958
rect 1316 5956 1372 5958
rect 1396 5956 1452 5958
rect 1582 5072 1638 5128
rect 1156 4922 1212 4924
rect 1236 4922 1292 4924
rect 1316 4922 1372 4924
rect 1396 4922 1452 4924
rect 1156 4870 1202 4922
rect 1202 4870 1212 4922
rect 1236 4870 1266 4922
rect 1266 4870 1278 4922
rect 1278 4870 1292 4922
rect 1316 4870 1330 4922
rect 1330 4870 1342 4922
rect 1342 4870 1372 4922
rect 1396 4870 1406 4922
rect 1406 4870 1452 4922
rect 1156 4868 1212 4870
rect 1236 4868 1292 4870
rect 1316 4868 1372 4870
rect 1396 4868 1452 4870
rect 3156 7642 3212 7644
rect 3236 7642 3292 7644
rect 3316 7642 3372 7644
rect 3396 7642 3452 7644
rect 3156 7590 3202 7642
rect 3202 7590 3212 7642
rect 3236 7590 3266 7642
rect 3266 7590 3278 7642
rect 3278 7590 3292 7642
rect 3316 7590 3330 7642
rect 3330 7590 3342 7642
rect 3342 7590 3372 7642
rect 3396 7590 3406 7642
rect 3406 7590 3452 7642
rect 3156 7588 3212 7590
rect 3236 7588 3292 7590
rect 3316 7588 3372 7590
rect 3396 7588 3452 7590
rect 4158 6860 4214 6896
rect 4158 6840 4160 6860
rect 4160 6840 4212 6860
rect 4212 6840 4214 6860
rect 3156 6554 3212 6556
rect 3236 6554 3292 6556
rect 3316 6554 3372 6556
rect 3396 6554 3452 6556
rect 3156 6502 3202 6554
rect 3202 6502 3212 6554
rect 3236 6502 3266 6554
rect 3266 6502 3278 6554
rect 3278 6502 3292 6554
rect 3316 6502 3330 6554
rect 3330 6502 3342 6554
rect 3342 6502 3372 6554
rect 3396 6502 3406 6554
rect 3406 6502 3452 6554
rect 3156 6500 3212 6502
rect 3236 6500 3292 6502
rect 3316 6500 3372 6502
rect 3396 6500 3452 6502
rect 3156 5466 3212 5468
rect 3236 5466 3292 5468
rect 3316 5466 3372 5468
rect 3396 5466 3452 5468
rect 3156 5414 3202 5466
rect 3202 5414 3212 5466
rect 3236 5414 3266 5466
rect 3266 5414 3278 5466
rect 3278 5414 3292 5466
rect 3316 5414 3330 5466
rect 3330 5414 3342 5466
rect 3342 5414 3372 5466
rect 3396 5414 3406 5466
rect 3406 5414 3452 5466
rect 3156 5412 3212 5414
rect 3236 5412 3292 5414
rect 3316 5412 3372 5414
rect 3396 5412 3452 5414
rect 3156 4378 3212 4380
rect 3236 4378 3292 4380
rect 3316 4378 3372 4380
rect 3396 4378 3452 4380
rect 3156 4326 3202 4378
rect 3202 4326 3212 4378
rect 3236 4326 3266 4378
rect 3266 4326 3278 4378
rect 3278 4326 3292 4378
rect 3316 4326 3330 4378
rect 3330 4326 3342 4378
rect 3342 4326 3372 4378
rect 3396 4326 3406 4378
rect 3406 4326 3452 4378
rect 3156 4324 3212 4326
rect 3236 4324 3292 4326
rect 3316 4324 3372 4326
rect 3396 4324 3452 4326
rect 1156 3834 1212 3836
rect 1236 3834 1292 3836
rect 1316 3834 1372 3836
rect 1396 3834 1452 3836
rect 1156 3782 1202 3834
rect 1202 3782 1212 3834
rect 1236 3782 1266 3834
rect 1266 3782 1278 3834
rect 1278 3782 1292 3834
rect 1316 3782 1330 3834
rect 1330 3782 1342 3834
rect 1342 3782 1372 3834
rect 1396 3782 1406 3834
rect 1406 3782 1452 3834
rect 1156 3780 1212 3782
rect 1236 3780 1292 3782
rect 1316 3780 1372 3782
rect 1396 3780 1452 3782
rect 4342 6704 4398 6760
rect 4066 4156 4068 4176
rect 4068 4156 4120 4176
rect 4120 4156 4122 4176
rect 4066 4120 4122 4156
rect 2778 3440 2834 3496
rect 1156 2746 1212 2748
rect 1236 2746 1292 2748
rect 1316 2746 1372 2748
rect 1396 2746 1452 2748
rect 1156 2694 1202 2746
rect 1202 2694 1212 2746
rect 1236 2694 1266 2746
rect 1266 2694 1278 2746
rect 1278 2694 1292 2746
rect 1316 2694 1330 2746
rect 1330 2694 1342 2746
rect 1342 2694 1372 2746
rect 1396 2694 1406 2746
rect 1406 2694 1452 2746
rect 1156 2692 1212 2694
rect 1236 2692 1292 2694
rect 1316 2692 1372 2694
rect 1396 2692 1452 2694
rect 1156 1658 1212 1660
rect 1236 1658 1292 1660
rect 1316 1658 1372 1660
rect 1396 1658 1452 1660
rect 1156 1606 1202 1658
rect 1202 1606 1212 1658
rect 1236 1606 1266 1658
rect 1266 1606 1278 1658
rect 1278 1606 1292 1658
rect 1316 1606 1330 1658
rect 1330 1606 1342 1658
rect 1342 1606 1372 1658
rect 1396 1606 1406 1658
rect 1406 1606 1452 1658
rect 1156 1604 1212 1606
rect 1236 1604 1292 1606
rect 1316 1604 1372 1606
rect 1396 1604 1452 1606
rect 3156 3290 3212 3292
rect 3236 3290 3292 3292
rect 3316 3290 3372 3292
rect 3396 3290 3452 3292
rect 3156 3238 3202 3290
rect 3202 3238 3212 3290
rect 3236 3238 3266 3290
rect 3266 3238 3278 3290
rect 3278 3238 3292 3290
rect 3316 3238 3330 3290
rect 3330 3238 3342 3290
rect 3342 3238 3372 3290
rect 3396 3238 3406 3290
rect 3406 3238 3452 3290
rect 3156 3236 3212 3238
rect 3236 3236 3292 3238
rect 3316 3236 3372 3238
rect 3396 3236 3452 3238
rect 3156 2202 3212 2204
rect 3236 2202 3292 2204
rect 3316 2202 3372 2204
rect 3396 2202 3452 2204
rect 3156 2150 3202 2202
rect 3202 2150 3212 2202
rect 3236 2150 3266 2202
rect 3266 2150 3278 2202
rect 3278 2150 3292 2202
rect 3316 2150 3330 2202
rect 3330 2150 3342 2202
rect 3342 2150 3372 2202
rect 3396 2150 3406 2202
rect 3406 2150 3452 2202
rect 3156 2148 3212 2150
rect 3236 2148 3292 2150
rect 3316 2148 3372 2150
rect 3396 2148 3452 2150
rect 4066 1944 4122 2000
rect 4250 2352 4306 2408
rect 2870 1400 2926 1456
rect 7930 8220 7986 8256
rect 7930 8200 7932 8220
rect 7932 8200 7984 8220
rect 7984 8200 7986 8220
rect 5156 7098 5212 7100
rect 5236 7098 5292 7100
rect 5316 7098 5372 7100
rect 5396 7098 5452 7100
rect 5156 7046 5202 7098
rect 5202 7046 5212 7098
rect 5236 7046 5266 7098
rect 5266 7046 5278 7098
rect 5278 7046 5292 7098
rect 5316 7046 5330 7098
rect 5330 7046 5342 7098
rect 5342 7046 5372 7098
rect 5396 7046 5406 7098
rect 5406 7046 5452 7098
rect 5156 7044 5212 7046
rect 5236 7044 5292 7046
rect 5316 7044 5372 7046
rect 5396 7044 5452 7046
rect 5156 6010 5212 6012
rect 5236 6010 5292 6012
rect 5316 6010 5372 6012
rect 5396 6010 5452 6012
rect 5156 5958 5202 6010
rect 5202 5958 5212 6010
rect 5236 5958 5266 6010
rect 5266 5958 5278 6010
rect 5278 5958 5292 6010
rect 5316 5958 5330 6010
rect 5330 5958 5342 6010
rect 5342 5958 5372 6010
rect 5396 5958 5406 6010
rect 5406 5958 5452 6010
rect 5156 5956 5212 5958
rect 5236 5956 5292 5958
rect 5316 5956 5372 5958
rect 5396 5956 5452 5958
rect 5156 4922 5212 4924
rect 5236 4922 5292 4924
rect 5316 4922 5372 4924
rect 5396 4922 5452 4924
rect 5156 4870 5202 4922
rect 5202 4870 5212 4922
rect 5236 4870 5266 4922
rect 5266 4870 5278 4922
rect 5278 4870 5292 4922
rect 5316 4870 5330 4922
rect 5330 4870 5342 4922
rect 5342 4870 5372 4922
rect 5396 4870 5406 4922
rect 5406 4870 5452 4922
rect 5156 4868 5212 4870
rect 5236 4868 5292 4870
rect 5316 4868 5372 4870
rect 5396 4868 5452 4870
rect 6826 7384 6882 7440
rect 7156 7642 7212 7644
rect 7236 7642 7292 7644
rect 7316 7642 7372 7644
rect 7396 7642 7452 7644
rect 7156 7590 7202 7642
rect 7202 7590 7212 7642
rect 7236 7590 7266 7642
rect 7266 7590 7278 7642
rect 7278 7590 7292 7642
rect 7316 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7372 7642
rect 7396 7590 7406 7642
rect 7406 7590 7452 7642
rect 7156 7588 7212 7590
rect 7236 7588 7292 7590
rect 7316 7588 7372 7590
rect 7396 7588 7452 7590
rect 7156 6554 7212 6556
rect 7236 6554 7292 6556
rect 7316 6554 7372 6556
rect 7396 6554 7452 6556
rect 7156 6502 7202 6554
rect 7202 6502 7212 6554
rect 7236 6502 7266 6554
rect 7266 6502 7278 6554
rect 7278 6502 7292 6554
rect 7316 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7372 6554
rect 7396 6502 7406 6554
rect 7406 6502 7452 6554
rect 7156 6500 7212 6502
rect 7236 6500 7292 6502
rect 7316 6500 7372 6502
rect 7396 6500 7452 6502
rect 5156 3834 5212 3836
rect 5236 3834 5292 3836
rect 5316 3834 5372 3836
rect 5396 3834 5452 3836
rect 5156 3782 5202 3834
rect 5202 3782 5212 3834
rect 5236 3782 5266 3834
rect 5266 3782 5278 3834
rect 5278 3782 5292 3834
rect 5316 3782 5330 3834
rect 5330 3782 5342 3834
rect 5342 3782 5372 3834
rect 5396 3782 5406 3834
rect 5406 3782 5452 3834
rect 5156 3780 5212 3782
rect 5236 3780 5292 3782
rect 5316 3780 5372 3782
rect 5396 3780 5452 3782
rect 7156 5466 7212 5468
rect 7236 5466 7292 5468
rect 7316 5466 7372 5468
rect 7396 5466 7452 5468
rect 7156 5414 7202 5466
rect 7202 5414 7212 5466
rect 7236 5414 7266 5466
rect 7266 5414 7278 5466
rect 7278 5414 7292 5466
rect 7316 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7372 5466
rect 7396 5414 7406 5466
rect 7406 5414 7452 5466
rect 7156 5412 7212 5414
rect 7236 5412 7292 5414
rect 7316 5412 7372 5414
rect 7396 5412 7452 5414
rect 6458 4820 6514 4856
rect 7930 5500 7986 5536
rect 7930 5480 7932 5500
rect 7932 5480 7984 5500
rect 7984 5480 7986 5500
rect 6458 4800 6460 4820
rect 6460 4800 6512 4820
rect 6512 4800 6514 4820
rect 7156 4378 7212 4380
rect 7236 4378 7292 4380
rect 7316 4378 7372 4380
rect 7396 4378 7452 4380
rect 7156 4326 7202 4378
rect 7202 4326 7212 4378
rect 7236 4326 7266 4378
rect 7266 4326 7278 4378
rect 7278 4326 7292 4378
rect 7316 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7372 4378
rect 7396 4326 7406 4378
rect 7406 4326 7452 4378
rect 7156 4324 7212 4326
rect 7236 4324 7292 4326
rect 7316 4324 7372 4326
rect 7396 4324 7452 4326
rect 7102 4140 7158 4176
rect 7102 4120 7104 4140
rect 7104 4120 7156 4140
rect 7156 4120 7158 4140
rect 5078 2896 5134 2952
rect 5156 2746 5212 2748
rect 5236 2746 5292 2748
rect 5316 2746 5372 2748
rect 5396 2746 5452 2748
rect 5156 2694 5202 2746
rect 5202 2694 5212 2746
rect 5236 2694 5266 2746
rect 5266 2694 5278 2746
rect 5278 2694 5292 2746
rect 5316 2694 5330 2746
rect 5330 2694 5342 2746
rect 5342 2694 5372 2746
rect 5396 2694 5406 2746
rect 5406 2694 5452 2746
rect 5156 2692 5212 2694
rect 5236 2692 5292 2694
rect 5316 2692 5372 2694
rect 5396 2692 5452 2694
rect 7156 3290 7212 3292
rect 7236 3290 7292 3292
rect 7316 3290 7372 3292
rect 7396 3290 7452 3292
rect 7156 3238 7202 3290
rect 7202 3238 7212 3290
rect 7236 3238 7266 3290
rect 7266 3238 7278 3290
rect 7278 3238 7292 3290
rect 7316 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7372 3290
rect 7396 3238 7406 3290
rect 7406 3238 7452 3290
rect 7156 3236 7212 3238
rect 7236 3236 7292 3238
rect 7316 3236 7372 3238
rect 7396 3236 7452 3238
rect 7156 2202 7212 2204
rect 7236 2202 7292 2204
rect 7316 2202 7372 2204
rect 7396 2202 7452 2204
rect 7156 2150 7202 2202
rect 7202 2150 7212 2202
rect 7236 2150 7266 2202
rect 7266 2150 7278 2202
rect 7278 2150 7292 2202
rect 7316 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7372 2202
rect 7396 2150 7406 2202
rect 7406 2150 7452 2202
rect 7156 2148 7212 2150
rect 7236 2148 7292 2150
rect 7316 2148 7372 2150
rect 7396 2148 7452 2150
rect 5156 1658 5212 1660
rect 5236 1658 5292 1660
rect 5316 1658 5372 1660
rect 5396 1658 5452 1660
rect 5156 1606 5202 1658
rect 5202 1606 5212 1658
rect 5236 1606 5266 1658
rect 5266 1606 5278 1658
rect 5278 1606 5292 1658
rect 5316 1606 5330 1658
rect 5330 1606 5342 1658
rect 5342 1606 5372 1658
rect 5396 1606 5406 1658
rect 5406 1606 5452 1658
rect 5156 1604 5212 1606
rect 5236 1604 5292 1606
rect 5316 1604 5372 1606
rect 5396 1604 5452 1606
rect 3156 1114 3212 1116
rect 3236 1114 3292 1116
rect 3316 1114 3372 1116
rect 3396 1114 3452 1116
rect 3156 1062 3202 1114
rect 3202 1062 3212 1114
rect 3236 1062 3266 1114
rect 3266 1062 3278 1114
rect 3278 1062 3292 1114
rect 3316 1062 3330 1114
rect 3330 1062 3342 1114
rect 3342 1062 3372 1114
rect 3396 1062 3406 1114
rect 3406 1062 3452 1114
rect 3156 1060 3212 1062
rect 3236 1060 3292 1062
rect 3316 1060 3372 1062
rect 3396 1060 3452 1062
rect 6734 1400 6790 1456
rect 7156 1114 7212 1116
rect 7236 1114 7292 1116
rect 7316 1114 7372 1116
rect 7396 1114 7452 1116
rect 7156 1062 7202 1114
rect 7202 1062 7212 1114
rect 7236 1062 7266 1114
rect 7266 1062 7278 1114
rect 7278 1062 7292 1114
rect 7316 1062 7330 1114
rect 7330 1062 7342 1114
rect 7342 1062 7372 1114
rect 7396 1062 7406 1114
rect 7406 1062 7452 1114
rect 7156 1060 7212 1062
rect 7236 1060 7292 1062
rect 7316 1060 7372 1062
rect 7396 1060 7452 1062
rect 1582 720 1638 776
rect 7930 76 7932 96
rect 7932 76 7984 96
rect 7984 76 7986 96
rect 7930 40 7986 76
<< metal3 >>
rect 0 8938 800 8968
rect 4061 8938 4127 8941
rect 0 8936 4127 8938
rect 0 8880 4066 8936
rect 4122 8880 4127 8936
rect 0 8878 4127 8880
rect 0 8848 800 8878
rect 4061 8875 4127 8878
rect 7925 8258 7991 8261
rect 8200 8258 9000 8288
rect 7925 8256 9000 8258
rect 7925 8200 7930 8256
rect 7986 8200 9000 8256
rect 7925 8198 9000 8200
rect 7925 8195 7991 8198
rect 8200 8168 9000 8198
rect 3144 7648 3464 7649
rect 0 7578 800 7608
rect 3144 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3464 7648
rect 3144 7583 3464 7584
rect 7144 7648 7464 7649
rect 7144 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7464 7648
rect 7144 7583 7464 7584
rect 1577 7578 1643 7581
rect 8200 7578 9000 7608
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 7606 7518 9000 7578
rect 6821 7442 6887 7445
rect 7606 7442 7666 7518
rect 8200 7488 9000 7518
rect 6821 7440 7666 7442
rect 6821 7384 6826 7440
rect 6882 7384 7666 7440
rect 6821 7382 7666 7384
rect 6821 7379 6887 7382
rect 1144 7104 1464 7105
rect 1144 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1464 7104
rect 1144 7039 1464 7040
rect 5144 7104 5464 7105
rect 5144 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5464 7104
rect 5144 7039 5464 7040
rect 0 6898 800 6928
rect 4153 6898 4219 6901
rect 8200 6898 9000 6928
rect 0 6838 3986 6898
rect 0 6808 800 6838
rect 3926 6762 3986 6838
rect 4153 6896 9000 6898
rect 4153 6840 4158 6896
rect 4214 6840 9000 6896
rect 4153 6838 9000 6840
rect 4153 6835 4219 6838
rect 8200 6808 9000 6838
rect 4337 6762 4403 6765
rect 3926 6760 4403 6762
rect 3926 6704 4342 6760
rect 4398 6704 4403 6760
rect 3926 6702 4403 6704
rect 4337 6699 4403 6702
rect 3144 6560 3464 6561
rect 3144 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3464 6560
rect 3144 6495 3464 6496
rect 7144 6560 7464 6561
rect 7144 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7464 6560
rect 7144 6495 7464 6496
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 1144 6016 1464 6017
rect 1144 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1464 6016
rect 1144 5951 1464 5952
rect 5144 6016 5464 6017
rect 5144 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5464 6016
rect 5144 5951 5464 5952
rect 7925 5538 7991 5541
rect 8200 5538 9000 5568
rect 7925 5536 9000 5538
rect 7925 5480 7930 5536
rect 7986 5480 9000 5536
rect 7925 5478 9000 5480
rect 7925 5475 7991 5478
rect 3144 5472 3464 5473
rect 3144 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3464 5472
rect 3144 5407 3464 5408
rect 7144 5472 7464 5473
rect 7144 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7464 5472
rect 8200 5448 9000 5478
rect 7144 5407 7464 5408
rect 1577 5130 1643 5133
rect 982 5128 1643 5130
rect 982 5072 1582 5128
rect 1638 5072 1643 5128
rect 982 5070 1643 5072
rect 0 4858 800 4888
rect 982 4858 1042 5070
rect 1577 5067 1643 5070
rect 1144 4928 1464 4929
rect 1144 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1464 4928
rect 1144 4863 1464 4864
rect 5144 4928 5464 4929
rect 5144 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5464 4928
rect 5144 4863 5464 4864
rect 0 4798 1042 4858
rect 6453 4858 6519 4861
rect 8200 4858 9000 4888
rect 6453 4856 9000 4858
rect 6453 4800 6458 4856
rect 6514 4800 9000 4856
rect 6453 4798 9000 4800
rect 0 4768 800 4798
rect 6453 4795 6519 4798
rect 8200 4768 9000 4798
rect 3144 4384 3464 4385
rect 3144 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3464 4384
rect 3144 4319 3464 4320
rect 7144 4384 7464 4385
rect 7144 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7464 4384
rect 7144 4319 7464 4320
rect 0 4178 800 4208
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4088 800 4118
rect 4061 4115 4127 4118
rect 7097 4178 7163 4181
rect 8200 4178 9000 4208
rect 7097 4176 9000 4178
rect 7097 4120 7102 4176
rect 7158 4120 9000 4176
rect 7097 4118 9000 4120
rect 7097 4115 7163 4118
rect 8200 4088 9000 4118
rect 1144 3840 1464 3841
rect 1144 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1464 3840
rect 1144 3775 1464 3776
rect 5144 3840 5464 3841
rect 5144 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5464 3840
rect 5144 3775 5464 3776
rect 0 3498 800 3528
rect 2773 3498 2839 3501
rect 0 3496 2839 3498
rect 0 3440 2778 3496
rect 2834 3440 2839 3496
rect 0 3438 2839 3440
rect 0 3408 800 3438
rect 2773 3435 2839 3438
rect 3144 3296 3464 3297
rect 3144 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3464 3296
rect 3144 3231 3464 3232
rect 7144 3296 7464 3297
rect 7144 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7464 3296
rect 7144 3231 7464 3232
rect 5073 2954 5139 2957
rect 5073 2952 6930 2954
rect 5073 2896 5078 2952
rect 5134 2896 6930 2952
rect 5073 2894 6930 2896
rect 5073 2891 5139 2894
rect 6870 2818 6930 2894
rect 8200 2818 9000 2848
rect 6870 2758 9000 2818
rect 1144 2752 1464 2753
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1144 2687 1464 2688
rect 5144 2752 5464 2753
rect 5144 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5464 2752
rect 8200 2728 9000 2758
rect 5144 2687 5464 2688
rect 4245 2410 4311 2413
rect 4245 2408 7666 2410
rect 4245 2352 4250 2408
rect 4306 2352 7666 2408
rect 4245 2350 7666 2352
rect 4245 2347 4311 2350
rect 3144 2208 3464 2209
rect 0 2138 800 2168
rect 3144 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3464 2208
rect 3144 2143 3464 2144
rect 7144 2208 7464 2209
rect 7144 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7464 2208
rect 7144 2143 7464 2144
rect 7606 2138 7666 2350
rect 8200 2138 9000 2168
rect 0 2078 2146 2138
rect 7606 2078 9000 2138
rect 0 2048 800 2078
rect 2086 2002 2146 2078
rect 8200 2048 9000 2078
rect 4061 2002 4127 2005
rect 2086 2000 4127 2002
rect 2086 1944 4066 2000
rect 4122 1944 4127 2000
rect 2086 1942 4127 1944
rect 4061 1939 4127 1942
rect 1144 1664 1464 1665
rect 1144 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1464 1664
rect 1144 1599 1464 1600
rect 5144 1664 5464 1665
rect 5144 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5464 1664
rect 5144 1599 5464 1600
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 6729 1458 6795 1461
rect 8200 1458 9000 1488
rect 6729 1456 9000 1458
rect 6729 1400 6734 1456
rect 6790 1400 9000 1456
rect 6729 1398 9000 1400
rect 6729 1395 6795 1398
rect 8200 1368 9000 1398
rect 3144 1120 3464 1121
rect 3144 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3464 1120
rect 3144 1055 3464 1056
rect 7144 1120 7464 1121
rect 7144 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7464 1120
rect 7144 1055 7464 1056
rect 0 778 800 808
rect 1577 778 1643 781
rect 0 776 1643 778
rect 0 720 1582 776
rect 1638 720 1643 776
rect 0 718 1643 720
rect 0 688 800 718
rect 1577 715 1643 718
rect 7925 98 7991 101
rect 8200 98 9000 128
rect 7925 96 9000 98
rect 7925 40 7930 96
rect 7986 40 9000 96
rect 7925 38 9000 40
rect 7925 35 7991 38
rect 8200 8 9000 38
<< via3 >>
rect 3152 7644 3216 7648
rect 3152 7588 3156 7644
rect 3156 7588 3212 7644
rect 3212 7588 3216 7644
rect 3152 7584 3216 7588
rect 3232 7644 3296 7648
rect 3232 7588 3236 7644
rect 3236 7588 3292 7644
rect 3292 7588 3296 7644
rect 3232 7584 3296 7588
rect 3312 7644 3376 7648
rect 3312 7588 3316 7644
rect 3316 7588 3372 7644
rect 3372 7588 3376 7644
rect 3312 7584 3376 7588
rect 3392 7644 3456 7648
rect 3392 7588 3396 7644
rect 3396 7588 3452 7644
rect 3452 7588 3456 7644
rect 3392 7584 3456 7588
rect 7152 7644 7216 7648
rect 7152 7588 7156 7644
rect 7156 7588 7212 7644
rect 7212 7588 7216 7644
rect 7152 7584 7216 7588
rect 7232 7644 7296 7648
rect 7232 7588 7236 7644
rect 7236 7588 7292 7644
rect 7292 7588 7296 7644
rect 7232 7584 7296 7588
rect 7312 7644 7376 7648
rect 7312 7588 7316 7644
rect 7316 7588 7372 7644
rect 7372 7588 7376 7644
rect 7312 7584 7376 7588
rect 7392 7644 7456 7648
rect 7392 7588 7396 7644
rect 7396 7588 7452 7644
rect 7452 7588 7456 7644
rect 7392 7584 7456 7588
rect 1152 7100 1216 7104
rect 1152 7044 1156 7100
rect 1156 7044 1212 7100
rect 1212 7044 1216 7100
rect 1152 7040 1216 7044
rect 1232 7100 1296 7104
rect 1232 7044 1236 7100
rect 1236 7044 1292 7100
rect 1292 7044 1296 7100
rect 1232 7040 1296 7044
rect 1312 7100 1376 7104
rect 1312 7044 1316 7100
rect 1316 7044 1372 7100
rect 1372 7044 1376 7100
rect 1312 7040 1376 7044
rect 1392 7100 1456 7104
rect 1392 7044 1396 7100
rect 1396 7044 1452 7100
rect 1452 7044 1456 7100
rect 1392 7040 1456 7044
rect 5152 7100 5216 7104
rect 5152 7044 5156 7100
rect 5156 7044 5212 7100
rect 5212 7044 5216 7100
rect 5152 7040 5216 7044
rect 5232 7100 5296 7104
rect 5232 7044 5236 7100
rect 5236 7044 5292 7100
rect 5292 7044 5296 7100
rect 5232 7040 5296 7044
rect 5312 7100 5376 7104
rect 5312 7044 5316 7100
rect 5316 7044 5372 7100
rect 5372 7044 5376 7100
rect 5312 7040 5376 7044
rect 5392 7100 5456 7104
rect 5392 7044 5396 7100
rect 5396 7044 5452 7100
rect 5452 7044 5456 7100
rect 5392 7040 5456 7044
rect 3152 6556 3216 6560
rect 3152 6500 3156 6556
rect 3156 6500 3212 6556
rect 3212 6500 3216 6556
rect 3152 6496 3216 6500
rect 3232 6556 3296 6560
rect 3232 6500 3236 6556
rect 3236 6500 3292 6556
rect 3292 6500 3296 6556
rect 3232 6496 3296 6500
rect 3312 6556 3376 6560
rect 3312 6500 3316 6556
rect 3316 6500 3372 6556
rect 3372 6500 3376 6556
rect 3312 6496 3376 6500
rect 3392 6556 3456 6560
rect 3392 6500 3396 6556
rect 3396 6500 3452 6556
rect 3452 6500 3456 6556
rect 3392 6496 3456 6500
rect 7152 6556 7216 6560
rect 7152 6500 7156 6556
rect 7156 6500 7212 6556
rect 7212 6500 7216 6556
rect 7152 6496 7216 6500
rect 7232 6556 7296 6560
rect 7232 6500 7236 6556
rect 7236 6500 7292 6556
rect 7292 6500 7296 6556
rect 7232 6496 7296 6500
rect 7312 6556 7376 6560
rect 7312 6500 7316 6556
rect 7316 6500 7372 6556
rect 7372 6500 7376 6556
rect 7312 6496 7376 6500
rect 7392 6556 7456 6560
rect 7392 6500 7396 6556
rect 7396 6500 7452 6556
rect 7452 6500 7456 6556
rect 7392 6496 7456 6500
rect 1152 6012 1216 6016
rect 1152 5956 1156 6012
rect 1156 5956 1212 6012
rect 1212 5956 1216 6012
rect 1152 5952 1216 5956
rect 1232 6012 1296 6016
rect 1232 5956 1236 6012
rect 1236 5956 1292 6012
rect 1292 5956 1296 6012
rect 1232 5952 1296 5956
rect 1312 6012 1376 6016
rect 1312 5956 1316 6012
rect 1316 5956 1372 6012
rect 1372 5956 1376 6012
rect 1312 5952 1376 5956
rect 1392 6012 1456 6016
rect 1392 5956 1396 6012
rect 1396 5956 1452 6012
rect 1452 5956 1456 6012
rect 1392 5952 1456 5956
rect 5152 6012 5216 6016
rect 5152 5956 5156 6012
rect 5156 5956 5212 6012
rect 5212 5956 5216 6012
rect 5152 5952 5216 5956
rect 5232 6012 5296 6016
rect 5232 5956 5236 6012
rect 5236 5956 5292 6012
rect 5292 5956 5296 6012
rect 5232 5952 5296 5956
rect 5312 6012 5376 6016
rect 5312 5956 5316 6012
rect 5316 5956 5372 6012
rect 5372 5956 5376 6012
rect 5312 5952 5376 5956
rect 5392 6012 5456 6016
rect 5392 5956 5396 6012
rect 5396 5956 5452 6012
rect 5452 5956 5456 6012
rect 5392 5952 5456 5956
rect 3152 5468 3216 5472
rect 3152 5412 3156 5468
rect 3156 5412 3212 5468
rect 3212 5412 3216 5468
rect 3152 5408 3216 5412
rect 3232 5468 3296 5472
rect 3232 5412 3236 5468
rect 3236 5412 3292 5468
rect 3292 5412 3296 5468
rect 3232 5408 3296 5412
rect 3312 5468 3376 5472
rect 3312 5412 3316 5468
rect 3316 5412 3372 5468
rect 3372 5412 3376 5468
rect 3312 5408 3376 5412
rect 3392 5468 3456 5472
rect 3392 5412 3396 5468
rect 3396 5412 3452 5468
rect 3452 5412 3456 5468
rect 3392 5408 3456 5412
rect 7152 5468 7216 5472
rect 7152 5412 7156 5468
rect 7156 5412 7212 5468
rect 7212 5412 7216 5468
rect 7152 5408 7216 5412
rect 7232 5468 7296 5472
rect 7232 5412 7236 5468
rect 7236 5412 7292 5468
rect 7292 5412 7296 5468
rect 7232 5408 7296 5412
rect 7312 5468 7376 5472
rect 7312 5412 7316 5468
rect 7316 5412 7372 5468
rect 7372 5412 7376 5468
rect 7312 5408 7376 5412
rect 7392 5468 7456 5472
rect 7392 5412 7396 5468
rect 7396 5412 7452 5468
rect 7452 5412 7456 5468
rect 7392 5408 7456 5412
rect 1152 4924 1216 4928
rect 1152 4868 1156 4924
rect 1156 4868 1212 4924
rect 1212 4868 1216 4924
rect 1152 4864 1216 4868
rect 1232 4924 1296 4928
rect 1232 4868 1236 4924
rect 1236 4868 1292 4924
rect 1292 4868 1296 4924
rect 1232 4864 1296 4868
rect 1312 4924 1376 4928
rect 1312 4868 1316 4924
rect 1316 4868 1372 4924
rect 1372 4868 1376 4924
rect 1312 4864 1376 4868
rect 1392 4924 1456 4928
rect 1392 4868 1396 4924
rect 1396 4868 1452 4924
rect 1452 4868 1456 4924
rect 1392 4864 1456 4868
rect 5152 4924 5216 4928
rect 5152 4868 5156 4924
rect 5156 4868 5212 4924
rect 5212 4868 5216 4924
rect 5152 4864 5216 4868
rect 5232 4924 5296 4928
rect 5232 4868 5236 4924
rect 5236 4868 5292 4924
rect 5292 4868 5296 4924
rect 5232 4864 5296 4868
rect 5312 4924 5376 4928
rect 5312 4868 5316 4924
rect 5316 4868 5372 4924
rect 5372 4868 5376 4924
rect 5312 4864 5376 4868
rect 5392 4924 5456 4928
rect 5392 4868 5396 4924
rect 5396 4868 5452 4924
rect 5452 4868 5456 4924
rect 5392 4864 5456 4868
rect 3152 4380 3216 4384
rect 3152 4324 3156 4380
rect 3156 4324 3212 4380
rect 3212 4324 3216 4380
rect 3152 4320 3216 4324
rect 3232 4380 3296 4384
rect 3232 4324 3236 4380
rect 3236 4324 3292 4380
rect 3292 4324 3296 4380
rect 3232 4320 3296 4324
rect 3312 4380 3376 4384
rect 3312 4324 3316 4380
rect 3316 4324 3372 4380
rect 3372 4324 3376 4380
rect 3312 4320 3376 4324
rect 3392 4380 3456 4384
rect 3392 4324 3396 4380
rect 3396 4324 3452 4380
rect 3452 4324 3456 4380
rect 3392 4320 3456 4324
rect 7152 4380 7216 4384
rect 7152 4324 7156 4380
rect 7156 4324 7212 4380
rect 7212 4324 7216 4380
rect 7152 4320 7216 4324
rect 7232 4380 7296 4384
rect 7232 4324 7236 4380
rect 7236 4324 7292 4380
rect 7292 4324 7296 4380
rect 7232 4320 7296 4324
rect 7312 4380 7376 4384
rect 7312 4324 7316 4380
rect 7316 4324 7372 4380
rect 7372 4324 7376 4380
rect 7312 4320 7376 4324
rect 7392 4380 7456 4384
rect 7392 4324 7396 4380
rect 7396 4324 7452 4380
rect 7452 4324 7456 4380
rect 7392 4320 7456 4324
rect 1152 3836 1216 3840
rect 1152 3780 1156 3836
rect 1156 3780 1212 3836
rect 1212 3780 1216 3836
rect 1152 3776 1216 3780
rect 1232 3836 1296 3840
rect 1232 3780 1236 3836
rect 1236 3780 1292 3836
rect 1292 3780 1296 3836
rect 1232 3776 1296 3780
rect 1312 3836 1376 3840
rect 1312 3780 1316 3836
rect 1316 3780 1372 3836
rect 1372 3780 1376 3836
rect 1312 3776 1376 3780
rect 1392 3836 1456 3840
rect 1392 3780 1396 3836
rect 1396 3780 1452 3836
rect 1452 3780 1456 3836
rect 1392 3776 1456 3780
rect 5152 3836 5216 3840
rect 5152 3780 5156 3836
rect 5156 3780 5212 3836
rect 5212 3780 5216 3836
rect 5152 3776 5216 3780
rect 5232 3836 5296 3840
rect 5232 3780 5236 3836
rect 5236 3780 5292 3836
rect 5292 3780 5296 3836
rect 5232 3776 5296 3780
rect 5312 3836 5376 3840
rect 5312 3780 5316 3836
rect 5316 3780 5372 3836
rect 5372 3780 5376 3836
rect 5312 3776 5376 3780
rect 5392 3836 5456 3840
rect 5392 3780 5396 3836
rect 5396 3780 5452 3836
rect 5452 3780 5456 3836
rect 5392 3776 5456 3780
rect 3152 3292 3216 3296
rect 3152 3236 3156 3292
rect 3156 3236 3212 3292
rect 3212 3236 3216 3292
rect 3152 3232 3216 3236
rect 3232 3292 3296 3296
rect 3232 3236 3236 3292
rect 3236 3236 3292 3292
rect 3292 3236 3296 3292
rect 3232 3232 3296 3236
rect 3312 3292 3376 3296
rect 3312 3236 3316 3292
rect 3316 3236 3372 3292
rect 3372 3236 3376 3292
rect 3312 3232 3376 3236
rect 3392 3292 3456 3296
rect 3392 3236 3396 3292
rect 3396 3236 3452 3292
rect 3452 3236 3456 3292
rect 3392 3232 3456 3236
rect 7152 3292 7216 3296
rect 7152 3236 7156 3292
rect 7156 3236 7212 3292
rect 7212 3236 7216 3292
rect 7152 3232 7216 3236
rect 7232 3292 7296 3296
rect 7232 3236 7236 3292
rect 7236 3236 7292 3292
rect 7292 3236 7296 3292
rect 7232 3232 7296 3236
rect 7312 3292 7376 3296
rect 7312 3236 7316 3292
rect 7316 3236 7372 3292
rect 7372 3236 7376 3292
rect 7312 3232 7376 3236
rect 7392 3292 7456 3296
rect 7392 3236 7396 3292
rect 7396 3236 7452 3292
rect 7452 3236 7456 3292
rect 7392 3232 7456 3236
rect 1152 2748 1216 2752
rect 1152 2692 1156 2748
rect 1156 2692 1212 2748
rect 1212 2692 1216 2748
rect 1152 2688 1216 2692
rect 1232 2748 1296 2752
rect 1232 2692 1236 2748
rect 1236 2692 1292 2748
rect 1292 2692 1296 2748
rect 1232 2688 1296 2692
rect 1312 2748 1376 2752
rect 1312 2692 1316 2748
rect 1316 2692 1372 2748
rect 1372 2692 1376 2748
rect 1312 2688 1376 2692
rect 1392 2748 1456 2752
rect 1392 2692 1396 2748
rect 1396 2692 1452 2748
rect 1452 2692 1456 2748
rect 1392 2688 1456 2692
rect 5152 2748 5216 2752
rect 5152 2692 5156 2748
rect 5156 2692 5212 2748
rect 5212 2692 5216 2748
rect 5152 2688 5216 2692
rect 5232 2748 5296 2752
rect 5232 2692 5236 2748
rect 5236 2692 5292 2748
rect 5292 2692 5296 2748
rect 5232 2688 5296 2692
rect 5312 2748 5376 2752
rect 5312 2692 5316 2748
rect 5316 2692 5372 2748
rect 5372 2692 5376 2748
rect 5312 2688 5376 2692
rect 5392 2748 5456 2752
rect 5392 2692 5396 2748
rect 5396 2692 5452 2748
rect 5452 2692 5456 2748
rect 5392 2688 5456 2692
rect 3152 2204 3216 2208
rect 3152 2148 3156 2204
rect 3156 2148 3212 2204
rect 3212 2148 3216 2204
rect 3152 2144 3216 2148
rect 3232 2204 3296 2208
rect 3232 2148 3236 2204
rect 3236 2148 3292 2204
rect 3292 2148 3296 2204
rect 3232 2144 3296 2148
rect 3312 2204 3376 2208
rect 3312 2148 3316 2204
rect 3316 2148 3372 2204
rect 3372 2148 3376 2204
rect 3312 2144 3376 2148
rect 3392 2204 3456 2208
rect 3392 2148 3396 2204
rect 3396 2148 3452 2204
rect 3452 2148 3456 2204
rect 3392 2144 3456 2148
rect 7152 2204 7216 2208
rect 7152 2148 7156 2204
rect 7156 2148 7212 2204
rect 7212 2148 7216 2204
rect 7152 2144 7216 2148
rect 7232 2204 7296 2208
rect 7232 2148 7236 2204
rect 7236 2148 7292 2204
rect 7292 2148 7296 2204
rect 7232 2144 7296 2148
rect 7312 2204 7376 2208
rect 7312 2148 7316 2204
rect 7316 2148 7372 2204
rect 7372 2148 7376 2204
rect 7312 2144 7376 2148
rect 7392 2204 7456 2208
rect 7392 2148 7396 2204
rect 7396 2148 7452 2204
rect 7452 2148 7456 2204
rect 7392 2144 7456 2148
rect 1152 1660 1216 1664
rect 1152 1604 1156 1660
rect 1156 1604 1212 1660
rect 1212 1604 1216 1660
rect 1152 1600 1216 1604
rect 1232 1660 1296 1664
rect 1232 1604 1236 1660
rect 1236 1604 1292 1660
rect 1292 1604 1296 1660
rect 1232 1600 1296 1604
rect 1312 1660 1376 1664
rect 1312 1604 1316 1660
rect 1316 1604 1372 1660
rect 1372 1604 1376 1660
rect 1312 1600 1376 1604
rect 1392 1660 1456 1664
rect 1392 1604 1396 1660
rect 1396 1604 1452 1660
rect 1452 1604 1456 1660
rect 1392 1600 1456 1604
rect 5152 1660 5216 1664
rect 5152 1604 5156 1660
rect 5156 1604 5212 1660
rect 5212 1604 5216 1660
rect 5152 1600 5216 1604
rect 5232 1660 5296 1664
rect 5232 1604 5236 1660
rect 5236 1604 5292 1660
rect 5292 1604 5296 1660
rect 5232 1600 5296 1604
rect 5312 1660 5376 1664
rect 5312 1604 5316 1660
rect 5316 1604 5372 1660
rect 5372 1604 5376 1660
rect 5312 1600 5376 1604
rect 5392 1660 5456 1664
rect 5392 1604 5396 1660
rect 5396 1604 5452 1660
rect 5452 1604 5456 1660
rect 5392 1600 5456 1604
rect 3152 1116 3216 1120
rect 3152 1060 3156 1116
rect 3156 1060 3212 1116
rect 3212 1060 3216 1116
rect 3152 1056 3216 1060
rect 3232 1116 3296 1120
rect 3232 1060 3236 1116
rect 3236 1060 3292 1116
rect 3292 1060 3296 1116
rect 3232 1056 3296 1060
rect 3312 1116 3376 1120
rect 3312 1060 3316 1116
rect 3316 1060 3372 1116
rect 3372 1060 3376 1116
rect 3312 1056 3376 1060
rect 3392 1116 3456 1120
rect 3392 1060 3396 1116
rect 3396 1060 3452 1116
rect 3452 1060 3456 1116
rect 3392 1056 3456 1060
rect 7152 1116 7216 1120
rect 7152 1060 7156 1116
rect 7156 1060 7212 1116
rect 7212 1060 7216 1116
rect 7152 1056 7216 1060
rect 7232 1116 7296 1120
rect 7232 1060 7236 1116
rect 7236 1060 7292 1116
rect 7292 1060 7296 1116
rect 7232 1056 7296 1060
rect 7312 1116 7376 1120
rect 7312 1060 7316 1116
rect 7316 1060 7372 1116
rect 7372 1060 7376 1116
rect 7312 1056 7376 1060
rect 7392 1116 7456 1120
rect 7392 1060 7396 1116
rect 7396 1060 7452 1116
rect 7452 1060 7456 1116
rect 7392 1056 7456 1060
<< metal4 >>
rect 1144 7104 1464 7664
rect 1144 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1464 7104
rect 1144 6016 1464 7040
rect 1144 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1464 6016
rect 1144 5558 1464 5952
rect 1144 5322 1186 5558
rect 1422 5322 1464 5558
rect 1144 4928 1464 5322
rect 1144 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1464 4928
rect 1144 3840 1464 4864
rect 1144 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1464 3840
rect 1144 2752 1464 3776
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1144 1664 1464 2688
rect 1144 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1464 1664
rect 1144 1558 1464 1600
rect 1144 1322 1186 1558
rect 1422 1322 1464 1558
rect 1144 1040 1464 1322
rect 3144 7648 3464 7664
rect 3144 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3464 7648
rect 3144 6560 3464 7584
rect 3144 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3464 6560
rect 3144 5472 3464 6496
rect 3144 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3464 5472
rect 3144 4384 3464 5408
rect 3144 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3464 4384
rect 3144 3558 3464 4320
rect 3144 3322 3186 3558
rect 3422 3322 3464 3558
rect 3144 3296 3464 3322
rect 3144 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3464 3296
rect 3144 2208 3464 3232
rect 3144 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3464 2208
rect 3144 1120 3464 2144
rect 3144 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3464 1120
rect 3144 1040 3464 1056
rect 5144 7104 5464 7664
rect 5144 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5464 7104
rect 5144 6016 5464 7040
rect 5144 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5464 6016
rect 5144 5558 5464 5952
rect 5144 5322 5186 5558
rect 5422 5322 5464 5558
rect 5144 4928 5464 5322
rect 5144 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5464 4928
rect 5144 3840 5464 4864
rect 5144 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5464 3840
rect 5144 2752 5464 3776
rect 5144 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5464 2752
rect 5144 1664 5464 2688
rect 5144 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5464 1664
rect 5144 1558 5464 1600
rect 5144 1322 5186 1558
rect 5422 1322 5464 1558
rect 5144 1040 5464 1322
rect 7144 7648 7464 7664
rect 7144 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7464 7648
rect 7144 6560 7464 7584
rect 7144 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7464 6560
rect 7144 5472 7464 6496
rect 7144 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7464 5472
rect 7144 4384 7464 5408
rect 7144 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7464 4384
rect 7144 3558 7464 4320
rect 7144 3322 7186 3558
rect 7422 3322 7464 3558
rect 7144 3296 7464 3322
rect 7144 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7464 3296
rect 7144 2208 7464 3232
rect 7144 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7464 2208
rect 7144 1120 7464 2144
rect 7144 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7464 1120
rect 7144 1040 7464 1056
<< via4 >>
rect 1186 5322 1422 5558
rect 1186 1322 1422 1558
rect 3186 3322 3422 3558
rect 5186 5322 5422 5558
rect 5186 1322 5422 1558
rect 7186 3322 7422 3558
<< metal5 >>
rect 1104 5558 7820 5600
rect 1104 5322 1186 5558
rect 1422 5322 5186 5558
rect 5422 5322 7820 5558
rect 1104 5280 7820 5322
rect 1104 3558 7820 3600
rect 1104 3322 3186 3558
rect 3422 3322 7186 3558
rect 7422 3322 7820 3558
rect 1104 3280 7820 3322
rect 1104 1558 7820 1600
rect 1104 1322 1186 1558
rect 1422 1322 5186 1558
rect 5422 1322 7820 1558
rect 1104 1280 7820 1322
use sky130_fd_sc_hd__fill_2  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[22\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 1840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1638025753
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2484 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[24\]
timestamp 1638025753
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1638025753
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[1\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2208 0 -1 2176
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 4232 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1638025753
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[26\]
timestamp 1638025753
transform -1 0 4232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1638025753
transform 1 0 4968 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_38
timestamp 1638025753
transform 1 0 4600 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[8\]
timestamp 1638025753
transform -1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 5152 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1638025753
transform 1 0 5520 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1638025753
transform 1 0 5428 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[20\]
timestamp 1638025753
transform -1 0 5520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[1\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 6348 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1638025753
transform 1 0 6808 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1638025753
transform 1 0 6348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1638025753
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1638025753
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1638025753
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[1\]
timestamp 1638025753
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1638025753
transform -1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1638025753
transform -1 0 7820 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1638025753
transform 1 0 7176 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1638025753
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1638025753
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1638025753
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[19\]
timestamp 1638025753
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[21\]
timestamp 1638025753
transform -1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[23\]
timestamp 1638025753
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1638025753
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1638025753
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1638025753
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp 1638025753
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1638025753
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1638025753
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[25\]
timestamp 1638025753
transform -1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[6\]
timestamp 1638025753
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_62
timestamp 1638025753
transform 1 0 6808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1638025753
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1638025753
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_54
timestamp 1638025753
transform 1 0 6072 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1638025753
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1638025753
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[0\]
timestamp 1638025753
transform 1 0 1932 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_12  FILLER_3_35
timestamp 1638025753
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1638025753
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1638025753
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1638025753
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1638025753
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1638025753
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1638025753
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[1\]
timestamp 1638025753
transform -1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1638025753
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_8
timestamp 1638025753
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[16\]
timestamp 1638025753
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1638025753
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1638025753
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1638025753
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1638025753
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1638025753
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1638025753
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1638025753
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1638025753
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1638025753
transform -1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[0\]
timestamp 1638025753
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_61
timestamp 1638025753
transform 1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1638025753
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1638025753
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1638025753
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[7\]
timestamp 1638025753
transform -1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[1\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 2208 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1638025753
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1638025753
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[9\]
timestamp 1638025753
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp 1638025753
transform 1 0 5060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1638025753
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1638025753
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1638025753
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1638025753
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform -1 0 7176 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[14\]
timestamp 1638025753
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1638025753
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1638025753
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1638025753
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1638025753
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1638025753
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1638025753
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[18\]
timestamp 1638025753
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1638025753
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1638025753
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1638025753
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp 1638025753
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1638025753
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1638025753
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1638025753
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1638025753
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1638025753
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_61
timestamp 1638025753
transform 1 0 6716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[17\]
timestamp 1638025753
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[15\]
timestamp 1638025753
transform -1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1638025753
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_59
timestamp 1638025753
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1638025753
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1638025753
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[11\]
timestamp 1638025753
transform -1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1638025753
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1638025753
transform -1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1638025753
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp 1638025753
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1638025753
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_8
timestamp 1638025753
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[12\]
timestamp 1638025753
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1638025753
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1638025753
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1638025753
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1638025753
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1638025753
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1638025753
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1638025753
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1638025753
transform -1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[0\]
timestamp 1638025753
transform -1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_20
timestamp 1638025753
transform 1 0 2944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1638025753
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1638025753
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1638025753
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1638025753
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_24
timestamp 1638025753
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[10\]
timestamp 1638025753
transform -1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[5\]
timestamp 1638025753
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[1\]
timestamp 1638025753
transform -1 0 1932 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_9_36
timestamp 1638025753
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1638025753
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_69
timestamp 1638025753
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1638025753
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1638025753
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1638025753
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[3\]
timestamp 1638025753
transform -1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_63
timestamp 1638025753
transform 1 0 6900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1638025753
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1638025753
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[4\]
timestamp 1638025753
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1638025753
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1638025753
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  spare_logic_biginv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1638025753
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1638025753
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_46
timestamp 1638025753
transform 1 0 5336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_34
timestamp 1638025753
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1638025753
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[0\]
timestamp 1638025753
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[3\]
timestamp 1638025753
transform -1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_59
timestamp 1638025753
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1638025753
transform 1 0 7176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1638025753
transform -1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[13\]
timestamp 1638025753
transform -1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[2\]
timestamp 1638025753
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1638025753
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1638025753
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1638025753
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1638025753
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1638025753
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1638025753
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1638025753
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1638025753
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1638025753
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1638025753
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1638025753
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1638025753
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[2\]
timestamp 1638025753
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 2048 800 2168 6 spare_xfq[0]
port 0 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 spare_xfq[1]
port 1 nsew signal tristate
rlabel metal2 s 4526 8200 4582 9000 6 spare_xfqn[0]
port 2 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 spare_xfqn[1]
port 3 nsew signal tristate
rlabel metal2 s 8390 0 8446 800 6 spare_xi[0]
port 4 nsew signal tristate
rlabel metal3 s 8200 8 9000 128 6 spare_xi[1]
port 5 nsew signal tristate
rlabel metal3 s 8200 5448 9000 5568 6 spare_xi[2]
port 6 nsew signal tristate
rlabel metal2 s 18 8200 74 9000 6 spare_xi[3]
port 7 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 spare_xib
port 8 nsew signal tristate
rlabel metal2 s 7102 8200 7158 9000 6 spare_xmx[0]
port 9 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 spare_xmx[1]
port 10 nsew signal tristate
rlabel metal3 s 8200 6808 9000 6928 6 spare_xna[0]
port 11 nsew signal tristate
rlabel metal3 s 8200 1368 9000 1488 6 spare_xna[1]
port 12 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 spare_xno[0]
port 13 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 spare_xno[1]
port 14 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 spare_xz[0]
port 15 nsew signal tristate
rlabel metal2 s 5170 8200 5226 9000 6 spare_xz[10]
port 16 nsew signal tristate
rlabel metal2 s 7746 8200 7802 9000 6 spare_xz[11]
port 17 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 spare_xz[12]
port 18 nsew signal tristate
rlabel metal3 s 8200 7488 9000 7608 6 spare_xz[13]
port 19 nsew signal tristate
rlabel metal2 s 1950 8200 2006 9000 6 spare_xz[14]
port 20 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 spare_xz[15]
port 21 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 spare_xz[16]
port 22 nsew signal tristate
rlabel metal3 s 8200 4768 9000 4888 6 spare_xz[17]
port 23 nsew signal tristate
rlabel metal2 s 662 8200 718 9000 6 spare_xz[18]
port 24 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 spare_xz[19]
port 25 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 spare_xz[1]
port 26 nsew signal tristate
rlabel metal2 s 5814 8200 5870 9000 6 spare_xz[20]
port 27 nsew signal tristate
rlabel metal3 s 8200 2048 9000 2168 6 spare_xz[21]
port 28 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 spare_xz[22]
port 29 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 spare_xz[23]
port 30 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 spare_xz[24]
port 31 nsew signal tristate
rlabel metal3 s 8200 2728 9000 2848 6 spare_xz[25]
port 32 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 spare_xz[26]
port 33 nsew signal tristate
rlabel metal3 s 8200 8168 9000 8288 6 spare_xz[2]
port 34 nsew signal tristate
rlabel metal2 s 8390 8200 8446 9000 6 spare_xz[3]
port 35 nsew signal tristate
rlabel metal2 s 2594 8200 2650 9000 6 spare_xz[4]
port 36 nsew signal tristate
rlabel metal2 s 3238 8200 3294 9000 6 spare_xz[5]
port 37 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 spare_xz[6]
port 38 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 spare_xz[7]
port 39 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 spare_xz[8]
port 40 nsew signal tristate
rlabel metal3 s 8200 4088 9000 4208 6 spare_xz[9]
port 41 nsew signal tristate
rlabel metal5 s 1104 1280 7820 1600 6 vccd
port 42 nsew power input
rlabel metal5 s 1104 5280 7820 5600 6 vccd
port 42 nsew power input
rlabel metal4 s 1144 1040 1464 7664 6 vccd
port 42 nsew power input
rlabel metal4 s 5144 1040 5464 7664 6 vccd
port 42 nsew power input
rlabel metal5 s 1104 3280 7820 3600 6 vssd
port 43 nsew ground input
rlabel metal4 s 3144 1040 3464 7664 6 vssd
port 43 nsew ground input
rlabel metal4 s 7144 1040 7464 7664 6 vssd
port 43 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 9000 9000
<< end >>
