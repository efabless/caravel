module caravan_motto ();
endmodule
