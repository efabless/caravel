magic
tech sky130A
magscale 1 2
timestamp 1665254080
<< viali >>
rect 581 1853 615 1887
rect 1409 1717 1443 1751
rect 765 1513 799 1547
rect 581 1173 615 1207
rect 949 833 983 867
rect 581 765 615 799
<< metal1 >>
rect 92 2202 2668 2224
rect 92 2150 234 2202
rect 286 2150 298 2202
rect 350 2150 1234 2202
rect 1286 2150 1298 2202
rect 1350 2150 2234 2202
rect 2286 2150 2298 2202
rect 2350 2150 2668 2202
rect 92 2128 2668 2150
rect 566 1884 572 1896
rect 527 1856 572 1884
rect 566 1844 572 1856
rect 624 1844 630 1896
rect 1394 1748 1400 1760
rect 1355 1720 1400 1748
rect 1394 1708 1400 1720
rect 1452 1708 1458 1760
rect 92 1658 2668 1680
rect 92 1606 734 1658
rect 786 1606 798 1658
rect 850 1606 1734 1658
rect 1786 1606 1798 1658
rect 1850 1606 2668 1658
rect 92 1584 2668 1606
rect 566 1504 572 1556
rect 624 1544 630 1556
rect 753 1547 811 1553
rect 753 1544 765 1547
rect 624 1516 765 1544
rect 624 1504 630 1516
rect 753 1513 765 1516
rect 799 1513 811 1547
rect 753 1507 811 1513
rect 566 1204 572 1216
rect 527 1176 572 1204
rect 566 1164 572 1176
rect 624 1164 630 1216
rect 92 1114 2668 1136
rect 92 1062 234 1114
rect 286 1062 298 1114
rect 350 1062 1234 1114
rect 1286 1062 1298 1114
rect 1350 1062 2234 1114
rect 2286 1062 2298 1114
rect 2350 1062 2668 1114
rect 92 1040 2668 1062
rect 934 864 940 876
rect 895 836 940 864
rect 934 824 940 836
rect 992 824 998 876
rect 566 796 572 808
rect 527 768 572 796
rect 566 756 572 768
rect 624 756 630 808
rect 92 570 2668 592
rect 92 518 734 570
rect 786 518 798 570
rect 850 518 1734 570
rect 1786 518 1798 570
rect 1850 518 2668 570
rect 92 496 2668 518
<< via1 >>
rect 234 2150 286 2202
rect 298 2150 350 2202
rect 1234 2150 1286 2202
rect 1298 2150 1350 2202
rect 2234 2150 2286 2202
rect 2298 2150 2350 2202
rect 572 1887 624 1896
rect 572 1853 581 1887
rect 581 1853 615 1887
rect 615 1853 624 1887
rect 572 1844 624 1853
rect 1400 1751 1452 1760
rect 1400 1717 1409 1751
rect 1409 1717 1443 1751
rect 1443 1717 1452 1751
rect 1400 1708 1452 1717
rect 734 1606 786 1658
rect 798 1606 850 1658
rect 1734 1606 1786 1658
rect 1798 1606 1850 1658
rect 572 1504 624 1556
rect 572 1207 624 1216
rect 572 1173 581 1207
rect 581 1173 615 1207
rect 615 1173 624 1207
rect 572 1164 624 1173
rect 234 1062 286 1114
rect 298 1062 350 1114
rect 1234 1062 1286 1114
rect 1298 1062 1350 1114
rect 2234 1062 2286 1114
rect 2298 1062 2350 1114
rect 940 867 992 876
rect 940 833 949 867
rect 949 833 983 867
rect 983 833 992 867
rect 940 824 992 833
rect 572 799 624 808
rect 572 765 581 799
rect 581 765 615 799
rect 615 765 624 799
rect 572 756 624 765
rect 734 518 786 570
rect 798 518 850 570
rect 1734 518 1786 570
rect 1798 518 1850 570
<< metal2 >>
rect 224 2204 360 2213
rect 280 2202 304 2204
rect 286 2150 298 2202
rect 280 2148 304 2150
rect 224 2139 360 2148
rect 1224 2204 1360 2213
rect 1280 2202 1304 2204
rect 1286 2150 1298 2202
rect 1280 2148 1304 2150
rect 1224 2139 1360 2148
rect 2224 2204 2360 2213
rect 2280 2202 2304 2204
rect 2286 2150 2298 2202
rect 2280 2148 2304 2150
rect 2224 2139 2360 2148
rect 572 1896 624 1902
rect 572 1838 624 1844
rect 584 1562 612 1838
rect 1400 1760 1452 1766
rect 1400 1702 1452 1708
rect 724 1660 860 1669
rect 780 1658 804 1660
rect 786 1606 798 1658
rect 780 1604 804 1606
rect 724 1595 860 1604
rect 572 1556 624 1562
rect 572 1498 624 1504
rect 1412 1329 1440 1702
rect 1724 1660 1860 1669
rect 1780 1658 1804 1660
rect 1786 1606 1798 1658
rect 1780 1604 1804 1606
rect 1724 1595 1860 1604
rect 938 1320 994 1329
rect 938 1255 994 1264
rect 1398 1320 1454 1329
rect 1398 1255 1454 1264
rect 572 1216 624 1222
rect 572 1158 624 1164
rect 224 1116 360 1125
rect 280 1114 304 1116
rect 286 1062 298 1114
rect 280 1060 304 1062
rect 224 1051 360 1060
rect 584 814 612 1158
rect 952 882 980 1255
rect 1224 1116 1360 1125
rect 1280 1114 1304 1116
rect 1286 1062 1298 1114
rect 1280 1060 1304 1062
rect 1224 1051 1360 1060
rect 2224 1116 2360 1125
rect 2280 1114 2304 1116
rect 2286 1062 2298 1114
rect 2280 1060 2304 1062
rect 2224 1051 2360 1060
rect 940 876 992 882
rect 940 818 992 824
rect 572 808 624 814
rect 572 750 624 756
rect 724 572 860 581
rect 780 570 804 572
rect 786 518 798 570
rect 780 516 804 518
rect 724 507 860 516
rect 1724 572 1860 581
rect 1780 570 1804 572
rect 1786 518 1798 570
rect 1780 516 1804 518
rect 1724 507 1860 516
<< via2 >>
rect 224 2202 280 2204
rect 304 2202 360 2204
rect 224 2150 234 2202
rect 234 2150 280 2202
rect 304 2150 350 2202
rect 350 2150 360 2202
rect 224 2148 280 2150
rect 304 2148 360 2150
rect 1224 2202 1280 2204
rect 1304 2202 1360 2204
rect 1224 2150 1234 2202
rect 1234 2150 1280 2202
rect 1304 2150 1350 2202
rect 1350 2150 1360 2202
rect 1224 2148 1280 2150
rect 1304 2148 1360 2150
rect 2224 2202 2280 2204
rect 2304 2202 2360 2204
rect 2224 2150 2234 2202
rect 2234 2150 2280 2202
rect 2304 2150 2350 2202
rect 2350 2150 2360 2202
rect 2224 2148 2280 2150
rect 2304 2148 2360 2150
rect 724 1658 780 1660
rect 804 1658 860 1660
rect 724 1606 734 1658
rect 734 1606 780 1658
rect 804 1606 850 1658
rect 850 1606 860 1658
rect 724 1604 780 1606
rect 804 1604 860 1606
rect 1724 1658 1780 1660
rect 1804 1658 1860 1660
rect 1724 1606 1734 1658
rect 1734 1606 1780 1658
rect 1804 1606 1850 1658
rect 1850 1606 1860 1658
rect 1724 1604 1780 1606
rect 1804 1604 1860 1606
rect 938 1264 994 1320
rect 1398 1264 1454 1320
rect 224 1114 280 1116
rect 304 1114 360 1116
rect 224 1062 234 1114
rect 234 1062 280 1114
rect 304 1062 350 1114
rect 350 1062 360 1114
rect 224 1060 280 1062
rect 304 1060 360 1062
rect 1224 1114 1280 1116
rect 1304 1114 1360 1116
rect 1224 1062 1234 1114
rect 1234 1062 1280 1114
rect 1304 1062 1350 1114
rect 1350 1062 1360 1114
rect 1224 1060 1280 1062
rect 1304 1060 1360 1062
rect 2224 1114 2280 1116
rect 2304 1114 2360 1116
rect 2224 1062 2234 1114
rect 2234 1062 2280 1114
rect 2304 1062 2350 1114
rect 2350 1062 2360 1114
rect 2224 1060 2280 1062
rect 2304 1060 2360 1062
rect 724 570 780 572
rect 804 570 860 572
rect 724 518 734 570
rect 734 518 780 570
rect 804 518 850 570
rect 850 518 860 570
rect 724 516 780 518
rect 804 516 860 518
rect 1724 570 1780 572
rect 1804 570 1860 572
rect 1724 518 1734 570
rect 1734 518 1780 570
rect 1804 518 1850 570
rect 1850 518 1860 570
rect 1724 516 1780 518
rect 1804 516 1860 518
<< metal3 >>
rect 214 2208 370 2209
rect 214 2144 220 2208
rect 284 2144 300 2208
rect 364 2144 370 2208
rect 214 2143 370 2144
rect 1214 2208 1370 2209
rect 1214 2144 1220 2208
rect 1284 2144 1300 2208
rect 1364 2144 1370 2208
rect 1214 2143 1370 2144
rect 2214 2208 2370 2209
rect 2214 2144 2220 2208
rect 2284 2144 2300 2208
rect 2364 2144 2370 2208
rect 2214 2143 2370 2144
rect 714 1664 870 1665
rect 714 1600 720 1664
rect 784 1600 800 1664
rect 864 1600 870 1664
rect 714 1599 870 1600
rect 1714 1664 1870 1665
rect 1714 1600 1720 1664
rect 1784 1600 1800 1664
rect 1864 1600 1870 1664
rect 1714 1599 1870 1600
rect 0 1322 800 1352
rect 933 1322 999 1325
rect 0 1320 999 1322
rect 0 1264 938 1320
rect 994 1264 999 1320
rect 0 1262 999 1264
rect 0 1232 800 1262
rect 933 1259 999 1262
rect 1393 1322 1459 1325
rect 2000 1322 2800 1352
rect 1393 1320 2800 1322
rect 1393 1264 1398 1320
rect 1454 1264 2800 1320
rect 1393 1262 2800 1264
rect 1393 1259 1459 1262
rect 2000 1232 2800 1262
rect 214 1120 370 1121
rect 214 1056 220 1120
rect 284 1056 300 1120
rect 364 1056 370 1120
rect 214 1055 370 1056
rect 1214 1120 1370 1121
rect 1214 1056 1220 1120
rect 1284 1056 1300 1120
rect 1364 1056 1370 1120
rect 1214 1055 1370 1056
rect 2214 1120 2370 1121
rect 2214 1056 2220 1120
rect 2284 1056 2300 1120
rect 2364 1056 2370 1120
rect 2214 1055 2370 1056
rect 714 576 870 577
rect 714 512 720 576
rect 784 512 800 576
rect 864 512 870 576
rect 714 511 870 512
rect 1714 576 1870 577
rect 1714 512 1720 576
rect 1784 512 1800 576
rect 1864 512 1870 576
rect 1714 511 1870 512
<< via3 >>
rect 220 2204 284 2208
rect 220 2148 224 2204
rect 224 2148 280 2204
rect 280 2148 284 2204
rect 220 2144 284 2148
rect 300 2204 364 2208
rect 300 2148 304 2204
rect 304 2148 360 2204
rect 360 2148 364 2204
rect 300 2144 364 2148
rect 1220 2204 1284 2208
rect 1220 2148 1224 2204
rect 1224 2148 1280 2204
rect 1280 2148 1284 2204
rect 1220 2144 1284 2148
rect 1300 2204 1364 2208
rect 1300 2148 1304 2204
rect 1304 2148 1360 2204
rect 1360 2148 1364 2204
rect 1300 2144 1364 2148
rect 2220 2204 2284 2208
rect 2220 2148 2224 2204
rect 2224 2148 2280 2204
rect 2280 2148 2284 2204
rect 2220 2144 2284 2148
rect 2300 2204 2364 2208
rect 2300 2148 2304 2204
rect 2304 2148 2360 2204
rect 2360 2148 2364 2204
rect 2300 2144 2364 2148
rect 720 1660 784 1664
rect 720 1604 724 1660
rect 724 1604 780 1660
rect 780 1604 784 1660
rect 720 1600 784 1604
rect 800 1660 864 1664
rect 800 1604 804 1660
rect 804 1604 860 1660
rect 860 1604 864 1660
rect 800 1600 864 1604
rect 1720 1660 1784 1664
rect 1720 1604 1724 1660
rect 1724 1604 1780 1660
rect 1780 1604 1784 1660
rect 1720 1600 1784 1604
rect 1800 1660 1864 1664
rect 1800 1604 1804 1660
rect 1804 1604 1860 1660
rect 1860 1604 1864 1660
rect 1800 1600 1864 1604
rect 220 1116 284 1120
rect 220 1060 224 1116
rect 224 1060 280 1116
rect 280 1060 284 1116
rect 220 1056 284 1060
rect 300 1116 364 1120
rect 300 1060 304 1116
rect 304 1060 360 1116
rect 360 1060 364 1116
rect 300 1056 364 1060
rect 1220 1116 1284 1120
rect 1220 1060 1224 1116
rect 1224 1060 1280 1116
rect 1280 1060 1284 1116
rect 1220 1056 1284 1060
rect 1300 1116 1364 1120
rect 1300 1060 1304 1116
rect 1304 1060 1360 1116
rect 1360 1060 1364 1116
rect 1300 1056 1364 1060
rect 2220 1116 2284 1120
rect 2220 1060 2224 1116
rect 2224 1060 2280 1116
rect 2280 1060 2284 1116
rect 2220 1056 2284 1060
rect 2300 1116 2364 1120
rect 2300 1060 2304 1116
rect 2304 1060 2360 1116
rect 2360 1060 2364 1116
rect 2300 1056 2364 1060
rect 720 572 784 576
rect 720 516 724 572
rect 724 516 780 572
rect 780 516 784 572
rect 720 512 784 516
rect 800 572 864 576
rect 800 516 804 572
rect 804 516 860 572
rect 860 516 864 572
rect 800 512 864 516
rect 1720 572 1784 576
rect 1720 516 1724 572
rect 1724 516 1780 572
rect 1780 516 1784 572
rect 1720 512 1784 516
rect 1800 572 1864 576
rect 1800 516 1804 572
rect 1804 516 1860 572
rect 1860 516 1864 572
rect 1800 512 1864 516
<< metal4 >>
rect 202 2208 382 2224
rect 202 2144 220 2208
rect 284 2144 300 2208
rect 364 2144 382 2208
rect 202 1120 382 2144
rect 202 1056 220 1120
rect 284 1056 300 1120
rect 364 1056 382 1120
rect 202 496 382 1056
rect 702 1664 882 2224
rect 702 1600 720 1664
rect 784 1600 800 1664
rect 864 1600 882 1664
rect 702 576 882 1600
rect 702 512 720 576
rect 784 512 800 576
rect 864 512 882 576
rect 702 496 882 512
rect 1202 2208 1382 2224
rect 1202 2144 1220 2208
rect 1284 2144 1300 2208
rect 1364 2144 1382 2208
rect 1202 1120 1382 2144
rect 1202 1056 1220 1120
rect 1284 1056 1300 1120
rect 1364 1056 1382 1120
rect 1202 496 1382 1056
rect 1702 1664 1882 2224
rect 1702 1600 1720 1664
rect 1784 1600 1800 1664
rect 1864 1600 1882 1664
rect 1702 576 1882 1600
rect 1702 512 1720 576
rect 1784 512 1800 576
rect 1864 512 1882 576
rect 1702 496 1882 512
rect 2202 2208 2382 2224
rect 2202 2144 2220 2208
rect 2284 2144 2300 2208
rect 2364 2144 2382 2208
rect 2202 1120 2382 2144
rect 2202 1056 2220 1120
rect 2284 1056 2300 1120
rect 2364 1056 2382 1120
rect 2202 496 2382 1056
use sky130_fd_sc_hd__fill_2  FILLER_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 92 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1663720911
transform 1 0 2300 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 92 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4
timestamp 1663720911
transform 1 0 460 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 828 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_16
timestamp 1663720911
transform 1 0 1564 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_24
timestamp 1663720911
transform 1 0 2300 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_0
timestamp 1663720911
transform 1 0 92 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1663720911
transform 1 0 2300 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1663720911
transform 1 0 2576 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 2484 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1
timestamp 1663720911
transform 1 0 2484 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__buf_16  const_one_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform 1 0 276 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663720911
transform -1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_16  const_zero_buf
timestamp 1663720911
transform 1 0 276 0 1 544
box -38 -48 2062 592
<< labels >>
flabel metal3 s 2000 1232 2800 1352 0 FreeSans 480 0 0 0 one
port 0 nsew signal tristate
flabel metal4 s 202 496 382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal4 s 1202 496 1382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal4 s 2202 496 2382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal4 s 702 496 882 2224 0 FreeSans 960 90 0 0 vssd
port 2 nsew ground bidirectional
flabel metal4 s 1702 496 1882 2224 0 FreeSans 960 90 0 0 vssd
port 2 nsew ground bidirectional
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 zero
port 3 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 2800 2600
<< end >>
