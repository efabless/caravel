magic
tech sky130A
magscale 1 2
timestamp 1665957051
<< locali >>
rect 416588 996667 416806 996673
rect 661989 996585 662207 996591
rect 663185 996585 663403 996591
rect 664381 996585 664599 996591
rect 665577 996585 665795 996591
rect 167978 996342 168196 996348
rect 169174 996342 169392 996348
rect 170370 996342 170588 996348
rect 41236 891200 41242 891418
rect 41236 890004 41242 890222
rect 41236 888808 41242 889026
rect 41236 887612 41242 887830
rect 41236 886416 41242 886634
rect 676332 727440 676338 727658
rect 676332 726244 676338 726462
rect 676332 725048 676338 725266
rect 676332 723852 676338 724070
rect 676332 722656 676338 722874
rect 676332 721460 676338 721678
rect 41261 609954 41267 610172
rect 41261 608758 41267 608976
rect 41261 607562 41267 607780
rect 41261 606366 41267 606584
rect 41261 605170 41267 605388
rect 41261 603974 41267 604192
rect 41261 602778 41267 602996
rect 41261 601582 41267 601800
rect 41261 600386 41267 600604
rect 41261 599190 41267 599408
rect 41261 597994 41267 598212
rect 676332 453416 676338 453634
rect 676332 452220 676338 452438
rect 676332 451024 676338 451242
rect 676332 449828 676338 450046
rect 676332 448632 676338 448850
rect 676332 447436 676338 447654
rect 676332 446240 676338 446458
rect 676332 445044 676338 445262
rect 676332 443848 676338 444066
rect 676332 442652 676338 442870
rect 676332 441456 676338 441674
rect 676332 440260 676338 440478
rect 41283 352373 41289 352591
rect 41283 351177 41289 351395
rect 41283 349981 41289 350199
rect 41283 348785 41289 349003
rect 41283 347589 41289 347807
rect 41283 346393 41289 346611
rect 41283 345197 41289 345415
rect 41283 344001 41289 344219
rect 41283 342805 41289 343023
rect 41283 341609 41289 341827
rect 41283 340413 41289 340631
rect 41283 339217 41289 339435
rect 41283 338021 41289 338239
rect 41283 336825 41289 337043
rect 41283 335629 41289 335847
rect 134848 43204 135066 43210
rect 136044 43204 136262 43210
rect 137240 43204 137458 43210
rect 138436 43204 138654 43210
rect 139632 43204 139850 43210
rect 140828 43204 141046 43210
rect 142024 43204 142242 43210
rect 143220 43204 143438 43210
rect 144416 43204 144634 43210
rect 145612 43204 145830 43210
rect 146808 43204 147026 43210
rect 148004 43204 148222 43210
rect 149200 43204 149418 43210
rect 150396 43204 150614 43210
rect 151592 43204 151810 43210
rect 152788 43204 153006 43210
rect 153984 43204 154202 43210
rect 155180 43204 155398 43210
rect 156376 43204 156594 43210
rect 157572 43204 157790 43210
rect 158768 43204 158986 43210
rect 430248 43204 430466 43210
rect 431444 43204 431662 43210
rect 432640 43204 432858 43210
rect 433836 43204 434054 43210
rect 435032 43204 435250 43210
rect 436228 43204 436446 43210
rect 437424 43204 437642 43210
rect 438620 43204 438838 43210
rect 439816 43204 440034 43210
rect 441012 43204 441230 43210
rect 442208 43204 442426 43210
rect 443404 43204 443622 43210
rect 444600 43204 444818 43210
rect 445796 43204 446014 43210
rect 446992 43204 447210 43210
rect 448188 43204 448406 43210
rect 449384 43204 449602 43210
rect 450580 43204 450798 43210
rect 451776 43204 451994 43210
rect 452972 43204 453190 43210
rect 454168 43204 454386 43210
<< viali >>
rect 416870 997217 416904 997387
rect 417514 997285 417732 997319
rect 662271 997135 662305 997305
rect 662915 997203 663133 997237
rect 663467 997135 663501 997305
rect 664111 997203 664329 997237
rect 664663 997135 664697 997305
rect 665307 997203 665525 997237
rect 665859 997135 665893 997305
rect 666503 997203 666721 997237
rect 167052 996960 167270 996994
rect 167880 996892 167914 997062
rect 168248 996960 168466 996994
rect 169076 996892 169110 997062
rect 169444 996960 169662 996994
rect 170272 996892 170306 997062
rect 416588 996673 416806 996707
rect 417516 996605 417550 996775
rect 661989 996591 662207 996625
rect 662917 996523 662951 996693
rect 663185 996591 663403 996625
rect 664113 996523 664147 996693
rect 664381 996591 664599 996625
rect 665309 996523 665343 996693
rect 665577 996591 665795 996625
rect 666505 996523 666539 996693
rect 167234 996280 167268 996450
rect 167978 996348 168196 996382
rect 168430 996280 168464 996450
rect 169174 996348 169392 996382
rect 169626 996280 169660 996450
rect 170370 996348 170588 996382
rect 41202 891200 41236 891418
rect 40522 891102 40692 891136
rect 40590 890274 40624 890492
rect 41134 890456 41304 890490
rect 41202 890004 41236 890222
rect 40522 889906 40692 889940
rect 40590 889078 40624 889296
rect 41134 889260 41304 889294
rect 41202 888808 41236 889026
rect 40522 888710 40692 888744
rect 40590 887882 40624 888100
rect 41134 888064 41304 888098
rect 41202 887612 41236 887830
rect 40522 887514 40692 887548
rect 40590 886686 40624 886904
rect 41134 886868 41304 886902
rect 41202 886416 41236 886634
rect 40522 886318 40692 886352
rect 40590 885490 40624 885708
rect 41134 885672 41304 885706
rect 676338 727440 676372 727658
rect 676882 727342 677052 727376
rect 676270 726696 676440 726730
rect 676950 726514 676984 726732
rect 676338 726244 676372 726462
rect 676882 726146 677052 726180
rect 676270 725500 676440 725534
rect 676950 725318 676984 725536
rect 676338 725048 676372 725266
rect 676882 724950 677052 724984
rect 676270 724304 676440 724338
rect 676950 724122 676984 724340
rect 676338 723852 676372 724070
rect 676882 723754 677052 723788
rect 676270 723108 676440 723142
rect 676950 722926 676984 723144
rect 676338 722656 676372 722874
rect 676882 722558 677052 722592
rect 676270 721912 676440 721946
rect 676950 721730 676984 721948
rect 676338 721460 676372 721678
rect 676882 721362 677052 721396
rect 676270 720716 676440 720750
rect 676950 720534 676984 720752
rect 41227 609954 41261 610172
rect 40547 609856 40717 609890
rect 40615 609028 40649 609246
rect 41159 609210 41329 609244
rect 41227 608758 41261 608976
rect 40547 608660 40717 608694
rect 40615 607832 40649 608050
rect 41159 608014 41329 608048
rect 41227 607562 41261 607780
rect 40547 607464 40717 607498
rect 40615 606636 40649 606854
rect 41159 606818 41329 606852
rect 41227 606366 41261 606584
rect 40547 606268 40717 606302
rect 40615 605440 40649 605658
rect 41159 605622 41329 605656
rect 41227 605170 41261 605388
rect 40547 605072 40717 605106
rect 40615 604244 40649 604462
rect 41159 604426 41329 604460
rect 41227 603974 41261 604192
rect 40547 603876 40717 603910
rect 40615 603048 40649 603266
rect 41159 603230 41329 603264
rect 41227 602778 41261 602996
rect 40547 602680 40717 602714
rect 40615 601852 40649 602070
rect 41159 602034 41329 602068
rect 41227 601582 41261 601800
rect 40547 601484 40717 601518
rect 40615 600656 40649 600874
rect 41159 600838 41329 600872
rect 41227 600386 41261 600604
rect 40547 600288 40717 600322
rect 40615 599460 40649 599678
rect 41159 599642 41329 599676
rect 41227 599190 41261 599408
rect 40547 599092 40717 599126
rect 40615 598264 40649 598482
rect 41159 598446 41329 598480
rect 41227 597994 41261 598212
rect 40547 597896 40717 597930
rect 40615 597068 40649 597286
rect 41159 597250 41329 597284
rect 676338 453416 676372 453634
rect 676882 453318 677052 453352
rect 676270 452672 676440 452706
rect 676950 452490 676984 452708
rect 676338 452220 676372 452438
rect 676882 452122 677052 452156
rect 676270 451476 676440 451510
rect 676950 451294 676984 451512
rect 676338 451024 676372 451242
rect 676882 450926 677052 450960
rect 676270 450280 676440 450314
rect 676950 450098 676984 450316
rect 676338 449828 676372 450046
rect 676882 449730 677052 449764
rect 676270 449084 676440 449118
rect 676950 448902 676984 449120
rect 676338 448632 676372 448850
rect 676882 448534 677052 448568
rect 676270 447888 676440 447922
rect 676950 447706 676984 447924
rect 676338 447436 676372 447654
rect 676882 447338 677052 447372
rect 676270 446692 676440 446726
rect 676950 446510 676984 446728
rect 676338 446240 676372 446458
rect 676882 446142 677052 446176
rect 676270 445496 676440 445530
rect 676950 445314 676984 445532
rect 676338 445044 676372 445262
rect 676882 444946 677052 444980
rect 676270 444300 676440 444334
rect 676950 444118 676984 444336
rect 676338 443848 676372 444066
rect 676882 443750 677052 443784
rect 676270 443104 676440 443138
rect 676950 442922 676984 443140
rect 676338 442652 676372 442870
rect 676882 442554 677052 442588
rect 676270 441908 676440 441942
rect 676950 441726 676984 441944
rect 676338 441456 676372 441674
rect 676882 441358 677052 441392
rect 676270 440712 676440 440746
rect 676950 440530 676984 440748
rect 676338 440260 676372 440478
rect 676882 440162 677052 440196
rect 676270 439516 676440 439550
rect 676950 439334 676984 439552
rect 41249 352373 41283 352591
rect 40569 352275 40739 352309
rect 40637 351447 40671 351665
rect 41181 351629 41351 351663
rect 41249 351177 41283 351395
rect 40569 351079 40739 351113
rect 40637 350251 40671 350469
rect 41171 350433 41341 350467
rect 41249 349981 41283 350199
rect 40569 349883 40739 349917
rect 40637 349055 40671 349273
rect 41181 349237 41351 349271
rect 41249 348785 41283 349003
rect 40569 348687 40739 348721
rect 40637 347859 40671 348077
rect 41181 348041 41351 348075
rect 41249 347589 41283 347807
rect 40569 347491 40739 347525
rect 40637 346663 40671 346881
rect 41181 346845 41351 346879
rect 41249 346393 41283 346611
rect 40569 346295 40739 346329
rect 40637 345467 40671 345685
rect 41181 345649 41351 345683
rect 41249 345197 41283 345415
rect 40569 345099 40739 345133
rect 40637 344271 40671 344489
rect 41181 344453 41351 344487
rect 41249 344001 41283 344219
rect 40569 343903 40739 343937
rect 40637 343075 40671 343293
rect 41181 343257 41351 343291
rect 41249 342805 41283 343023
rect 40569 342707 40739 342741
rect 40637 341879 40671 342097
rect 41181 342061 41351 342095
rect 41249 341609 41283 341827
rect 40569 341511 40739 341545
rect 40637 340683 40671 340901
rect 41181 340865 41351 340899
rect 41249 340413 41283 340631
rect 40569 340315 40739 340349
rect 40637 339487 40671 339705
rect 41181 339669 41351 339703
rect 41249 339217 41283 339435
rect 40569 339119 40739 339153
rect 40637 338291 40671 338509
rect 41181 338473 41351 338507
rect 41249 338021 41283 338239
rect 40569 337923 40739 337957
rect 40637 337095 40671 337313
rect 41181 337277 41351 337311
rect 41249 336825 41283 337043
rect 40569 336727 40739 336761
rect 40637 335899 40671 336117
rect 41181 336081 41351 336115
rect 41249 335629 41283 335847
rect 40569 335531 40739 335565
rect 40637 334703 40671 334921
rect 41181 334885 41351 334919
rect 134104 43102 134138 43272
rect 134848 43170 135066 43204
rect 135300 43102 135334 43272
rect 136044 43170 136262 43204
rect 136496 43102 136530 43272
rect 137240 43170 137458 43204
rect 137692 43102 137726 43272
rect 138436 43170 138654 43204
rect 138888 43102 138922 43272
rect 139632 43170 139850 43204
rect 140084 43102 140118 43272
rect 140828 43170 141046 43204
rect 141280 43102 141314 43272
rect 142024 43170 142242 43204
rect 142476 43102 142510 43272
rect 143220 43170 143438 43204
rect 143672 43102 143706 43272
rect 144416 43170 144634 43204
rect 144868 43102 144902 43272
rect 145612 43170 145830 43204
rect 146064 43102 146098 43272
rect 146808 43170 147026 43204
rect 147260 43102 147294 43272
rect 148004 43170 148222 43204
rect 148456 43102 148490 43272
rect 149200 43170 149418 43204
rect 149652 43102 149686 43272
rect 150396 43170 150614 43204
rect 150848 43102 150882 43272
rect 151592 43170 151810 43204
rect 152044 43102 152078 43272
rect 152788 43170 153006 43204
rect 153240 43102 153274 43272
rect 153984 43170 154202 43204
rect 154436 43102 154470 43272
rect 155180 43170 155398 43204
rect 155632 43102 155666 43272
rect 156376 43170 156594 43204
rect 156828 43102 156862 43272
rect 157572 43170 157790 43204
rect 158024 43102 158058 43272
rect 158768 43170 158986 43204
rect 429504 43102 429538 43272
rect 430248 43170 430466 43204
rect 430700 43102 430734 43272
rect 431444 43170 431662 43204
rect 431896 43102 431930 43272
rect 432640 43170 432858 43204
rect 433092 43102 433126 43272
rect 433836 43170 434054 43204
rect 434288 43102 434322 43272
rect 435032 43170 435250 43204
rect 435484 43102 435518 43272
rect 436228 43170 436446 43204
rect 436680 43102 436714 43272
rect 437424 43170 437642 43204
rect 437876 43102 437910 43272
rect 438620 43170 438838 43204
rect 439072 43102 439106 43272
rect 439816 43170 440034 43204
rect 440268 43102 440302 43272
rect 441012 43170 441230 43204
rect 441464 43102 441498 43272
rect 442208 43170 442426 43204
rect 442660 43102 442694 43272
rect 443404 43170 443622 43204
rect 443856 43102 443890 43272
rect 444600 43170 444818 43204
rect 445052 43102 445086 43272
rect 445796 43170 446014 43204
rect 446248 43102 446282 43272
rect 446992 43170 447210 43204
rect 447444 43102 447478 43272
rect 448188 43170 448406 43204
rect 448640 43102 448674 43272
rect 449384 43170 449602 43204
rect 449836 43102 449870 43272
rect 450580 43170 450798 43204
rect 451032 43102 451066 43272
rect 451776 43170 451994 43204
rect 452228 43102 452262 43272
rect 452972 43170 453190 43204
rect 453424 43102 453458 43272
rect 454168 43170 454386 43204
rect 135118 42558 135336 42592
rect 135946 42490 135980 42660
rect 136314 42558 136532 42592
rect 137142 42490 137176 42660
rect 137510 42558 137728 42592
rect 138338 42490 138372 42660
rect 138706 42558 138924 42592
rect 139534 42490 139568 42660
rect 139902 42558 140120 42592
rect 140730 42490 140764 42660
rect 141098 42558 141316 42592
rect 141926 42490 141960 42660
rect 142294 42558 142512 42592
rect 143122 42490 143156 42660
rect 143490 42558 143708 42592
rect 144318 42490 144352 42660
rect 144686 42558 144904 42592
rect 145514 42490 145548 42660
rect 145882 42558 146100 42592
rect 146710 42490 146744 42660
rect 147078 42558 147296 42592
rect 147906 42490 147940 42660
rect 148274 42558 148492 42592
rect 149102 42490 149136 42660
rect 149470 42558 149688 42592
rect 150298 42490 150332 42660
rect 150666 42558 150884 42592
rect 151494 42490 151528 42660
rect 151862 42558 152080 42592
rect 152690 42490 152724 42660
rect 153058 42558 153276 42592
rect 153886 42490 153920 42660
rect 154254 42558 154472 42592
rect 155082 42490 155116 42660
rect 155450 42558 155668 42592
rect 156278 42490 156312 42660
rect 156646 42558 156864 42592
rect 157474 42490 157508 42660
rect 158024 42490 158058 42660
rect 158668 42558 158886 42592
rect 430518 42558 430736 42592
rect 431346 42490 431380 42660
rect 431714 42558 431932 42592
rect 432542 42490 432576 42660
rect 432910 42558 433128 42592
rect 433738 42490 433772 42660
rect 434106 42558 434324 42592
rect 434934 42490 434968 42660
rect 435302 42558 435520 42592
rect 436130 42490 436164 42660
rect 436498 42558 436716 42592
rect 437326 42490 437360 42660
rect 437694 42558 437912 42592
rect 438522 42490 438556 42660
rect 438890 42558 439108 42592
rect 439718 42490 439752 42660
rect 440086 42558 440304 42592
rect 440914 42490 440948 42660
rect 441282 42558 441500 42592
rect 442110 42490 442144 42660
rect 442478 42558 442696 42592
rect 443306 42490 443340 42660
rect 443674 42558 443892 42592
rect 444502 42490 444536 42660
rect 444870 42558 445088 42592
rect 445698 42490 445732 42660
rect 446066 42558 446284 42592
rect 446894 42490 446928 42660
rect 447262 42558 447480 42592
rect 448090 42490 448124 42660
rect 448458 42558 448676 42592
rect 449286 42490 449320 42660
rect 449654 42558 449872 42592
rect 450482 42490 450516 42660
rect 450850 42558 451068 42592
rect 451678 42490 451712 42660
rect 452046 42558 452264 42592
rect 452874 42490 452908 42660
rect 453424 42490 453458 42660
rect 454068 42558 454286 42592
<< metal1 >>
rect 416862 997387 416914 997399
rect 417502 997275 417514 997327
rect 417732 997275 417744 997327
rect 662263 997305 662315 997317
rect 416862 997205 416914 997217
rect 663459 997305 663511 997317
rect 662903 997193 662915 997245
rect 663133 997193 663145 997245
rect 662263 997123 662315 997135
rect 664655 997305 664707 997317
rect 664099 997193 664111 997245
rect 664329 997193 664341 997245
rect 663459 997123 663511 997135
rect 665851 997305 665903 997317
rect 665295 997193 665307 997245
rect 665525 997193 665537 997245
rect 664655 997123 664707 997135
rect 666491 997193 666503 997245
rect 666721 997193 666733 997245
rect 665851 997123 665903 997135
rect 167870 997062 167922 997074
rect 167040 996950 167052 997002
rect 167270 996950 167282 997002
rect 169066 997062 169118 997074
rect 168236 996950 168248 997002
rect 168466 996950 168478 997002
rect 167870 996880 167922 996892
rect 170262 997062 170314 997074
rect 169432 996950 169444 997002
rect 169662 996950 169674 997002
rect 169066 996880 169118 996892
rect 417844 997026 418598 997044
rect 417844 996966 418223 997026
rect 418580 996966 418598 997026
rect 417844 996948 418598 996966
rect 170262 996880 170314 996892
rect 417508 996775 417560 996787
rect 416576 996663 416588 996715
rect 416806 996663 416818 996715
rect 662909 996693 662961 996705
rect 417508 996593 417560 996605
rect 661977 996581 661989 996633
rect 662207 996581 662219 996633
rect 664105 996693 664157 996705
rect 663173 996581 663185 996633
rect 663403 996581 663415 996633
rect 662909 996511 662961 996523
rect 665301 996693 665353 996705
rect 664369 996581 664381 996633
rect 664599 996581 664611 996633
rect 664105 996511 664157 996523
rect 666497 996693 666549 996705
rect 665565 996581 665577 996633
rect 665795 996581 665807 996633
rect 665301 996511 665353 996523
rect 666497 996511 666549 996523
rect 167224 996450 167276 996462
rect 168420 996450 168472 996462
rect 167966 996338 167978 996390
rect 168196 996338 168208 996390
rect 167224 996268 167276 996280
rect 169616 996450 169668 996462
rect 169162 996338 169174 996390
rect 169392 996338 169404 996390
rect 168420 996268 168472 996280
rect 170358 996338 170370 996390
rect 170588 996338 170600 996390
rect 169616 996268 169668 996280
rect 417852 995938 418598 995956
rect 417852 995878 418223 995938
rect 418580 995878 418598 995938
rect 417852 995860 418598 995878
rect 42235 995429 169626 995457
rect 41194 891418 41246 891430
rect 42235 891357 42263 995429
rect 169620 995405 169626 995429
rect 169678 995405 169684 995457
rect 170463 995401 170469 995453
rect 170521 995429 170527 995453
rect 170521 995401 172109 995429
rect 42211 891351 42263 891357
rect 42211 891293 42263 891299
rect 42291 995373 169502 995401
rect 41194 891188 41246 891200
rect 42291 891163 42319 995373
rect 169496 995349 169502 995373
rect 169554 995349 169560 995401
rect 416649 995387 416655 995411
rect 415907 995359 416655 995387
rect 416707 995359 416713 995411
rect 662050 995359 662056 995383
rect 170269 995289 170275 995341
rect 170327 995317 170333 995341
rect 170327 995289 171909 995317
rect 417492 995307 417498 995359
rect 417550 995331 662056 995359
rect 662108 995331 662114 995383
rect 662893 995335 662899 995387
rect 662951 995359 675332 995387
rect 662951 995335 662957 995359
rect 417550 995307 417556 995331
rect 662244 995303 662250 995327
rect 416843 995275 416849 995299
rect 416107 995247 416849 995275
rect 416901 995247 416907 995299
rect 417611 995275 417622 995303
rect 417616 995251 417622 995275
rect 417674 995275 662250 995303
rect 662302 995275 662308 995327
rect 663017 995279 663023 995331
rect 663075 995303 675276 995331
rect 663075 995279 663081 995303
rect 417674 995251 417680 995275
rect 42267 891157 42319 891163
rect 40510 891092 40522 891144
rect 40692 891092 40704 891144
rect 42267 891099 42319 891105
rect 42459 995205 168430 995233
rect 42207 890508 42259 890514
rect 40582 890492 40634 890504
rect 41122 890446 41134 890498
rect 41304 890446 41316 890498
rect 42207 890450 42259 890456
rect 40582 890262 40634 890274
rect 41194 890222 41246 890234
rect 41194 889992 41246 890004
rect 40510 889896 40522 889948
rect 40692 889896 40704 889948
rect 40582 889296 40634 889308
rect 41122 889250 41134 889302
rect 41304 889250 41316 889302
rect 40582 889066 40634 889078
rect 41194 889026 41246 889038
rect 41194 888796 41246 888808
rect 40510 888700 40522 888752
rect 40692 888700 40704 888752
rect 40582 888100 40634 888112
rect 41122 888054 41134 888106
rect 41304 888054 41316 888106
rect 40582 887870 40634 887882
rect 41194 887830 41246 887842
rect 41194 887600 41246 887612
rect 40510 887504 40522 887556
rect 40692 887504 40704 887556
rect 40582 886904 40634 886916
rect 41122 886858 41134 886910
rect 41304 886858 41316 886910
rect 40582 886674 40634 886686
rect 41194 886634 41246 886646
rect 41194 886404 41246 886416
rect 40510 886308 40522 886360
rect 40692 886308 40704 886360
rect 40582 885708 40634 885720
rect 41122 885662 41134 885714
rect 41304 885662 41316 885714
rect 40582 885478 40634 885490
rect 41219 610172 41271 610184
rect 42207 610111 42235 890450
rect 42183 610105 42235 610111
rect 42183 610047 42235 610053
rect 42263 890384 42315 890390
rect 42263 890326 42315 890332
rect 41219 609942 41271 609954
rect 42263 609917 42291 890326
rect 42459 890137 42487 995205
rect 168424 995181 168430 995205
rect 168482 995181 168488 995233
rect 169243 995177 169249 995229
rect 169301 995205 169307 995229
rect 169301 995177 171711 995205
rect 42435 890131 42487 890137
rect 42435 890073 42487 890079
rect 42515 995149 168306 995177
rect 42515 889967 42543 995149
rect 168300 995125 168306 995149
rect 168358 995125 168364 995177
rect 169073 995121 169079 995173
rect 169131 995149 169137 995173
rect 169131 995121 170871 995149
rect 663246 995135 663252 995159
rect 170843 995093 170871 995121
rect 660323 995107 663252 995135
rect 663304 995107 663310 995159
rect 664089 995111 664095 995163
rect 664147 995135 675080 995163
rect 664147 995111 664153 995135
rect 170843 995065 171511 995093
rect 663440 995079 663446 995103
rect 661224 995051 663446 995079
rect 663498 995051 663504 995103
rect 664213 995055 664219 995107
rect 664271 995079 675024 995107
rect 664271 995055 664277 995079
rect 661224 995023 661252 995051
rect 42491 889961 42543 889967
rect 42491 889903 42543 889909
rect 42683 994981 167234 995009
rect 42239 609911 42291 609917
rect 40535 609846 40547 609898
rect 40717 609846 40729 609898
rect 42239 609853 42291 609859
rect 42431 889312 42483 889318
rect 42431 889254 42483 889260
rect 42179 609262 42231 609268
rect 40607 609246 40659 609258
rect 41147 609200 41159 609252
rect 41329 609200 41341 609252
rect 42179 609204 42231 609210
rect 40607 609016 40659 609028
rect 41219 608976 41271 608988
rect 41219 608746 41271 608758
rect 40535 608650 40547 608702
rect 40717 608650 40729 608702
rect 40607 608050 40659 608062
rect 41147 608004 41159 608056
rect 41329 608004 41341 608056
rect 40607 607820 40659 607832
rect 41219 607780 41271 607792
rect 41219 607550 41271 607562
rect 40535 607454 40547 607506
rect 40717 607454 40729 607506
rect 40607 606854 40659 606866
rect 41147 606808 41159 606860
rect 41329 606808 41341 606860
rect 40607 606624 40659 606636
rect 41219 606584 41271 606596
rect 41219 606354 41271 606366
rect 40535 606258 40547 606310
rect 40717 606258 40729 606310
rect 40607 605658 40659 605670
rect 41147 605612 41159 605664
rect 41329 605612 41341 605664
rect 40607 605428 40659 605440
rect 41219 605388 41271 605400
rect 41219 605158 41271 605170
rect 40535 605062 40547 605114
rect 40717 605062 40729 605114
rect 40607 604462 40659 604474
rect 41147 604416 41159 604468
rect 41329 604416 41341 604468
rect 40607 604232 40659 604244
rect 41219 604192 41271 604204
rect 41219 603962 41271 603974
rect 40535 603866 40547 603918
rect 40717 603866 40729 603918
rect 40607 603266 40659 603278
rect 41147 603220 41159 603272
rect 41329 603220 41341 603272
rect 40607 603036 40659 603048
rect 41219 602996 41271 603008
rect 41219 602766 41271 602778
rect 40535 602670 40547 602722
rect 40717 602670 40729 602722
rect 40607 602070 40659 602082
rect 41147 602024 41159 602076
rect 41329 602024 41341 602076
rect 40607 601840 40659 601852
rect 41219 601800 41271 601812
rect 41219 601570 41271 601582
rect 40535 601474 40547 601526
rect 40717 601474 40729 601526
rect 40607 600874 40659 600886
rect 41147 600828 41159 600880
rect 41329 600828 41341 600880
rect 40607 600644 40659 600656
rect 41219 600604 41271 600616
rect 41219 600374 41271 600386
rect 40535 600278 40547 600330
rect 40717 600278 40729 600330
rect 40607 599678 40659 599690
rect 41147 599632 41159 599684
rect 41329 599632 41341 599684
rect 40607 599448 40659 599460
rect 41219 599408 41271 599420
rect 41219 599178 41271 599190
rect 40535 599082 40547 599134
rect 40717 599082 40729 599134
rect 40607 598482 40659 598494
rect 41147 598436 41159 598488
rect 41329 598436 41341 598488
rect 40607 598252 40659 598264
rect 41219 598212 41271 598224
rect 41219 597982 41271 597994
rect 40535 597886 40547 597938
rect 40717 597886 40729 597938
rect 40607 597286 40659 597298
rect 41147 597240 41159 597292
rect 41329 597240 41341 597292
rect 40607 597056 40659 597068
rect 41241 352591 41293 352603
rect 42179 352530 42207 609204
rect 42155 352524 42207 352530
rect 42155 352466 42207 352472
rect 42235 609138 42287 609144
rect 42235 609080 42287 609086
rect 41241 352361 41293 352373
rect 42235 352336 42263 609080
rect 42431 608891 42459 889254
rect 42407 608885 42459 608891
rect 42407 608827 42459 608833
rect 42487 889188 42539 889194
rect 42487 889130 42539 889136
rect 42487 608721 42515 889130
rect 42683 888965 42711 994981
rect 167228 994957 167234 994981
rect 167286 994957 167292 995009
rect 168071 994953 168077 995005
rect 168129 994981 168135 995005
rect 660523 994995 661252 995023
rect 168129 994953 171310 994981
rect 42659 888959 42711 888965
rect 42659 888901 42711 888907
rect 42739 994925 167110 994953
rect 42739 888771 42767 994925
rect 167104 994901 167110 994925
rect 167162 994901 167168 994953
rect 167877 994897 167883 994949
rect 167935 994925 167941 994949
rect 167935 994897 170441 994925
rect 664442 994911 664448 994935
rect 170413 994869 170441 994897
rect 660723 994883 664448 994911
rect 664500 994883 664506 994935
rect 665285 994887 665291 994939
rect 665343 994911 674856 994939
rect 665343 994887 665349 994911
rect 170413 994841 171110 994869
rect 664636 994855 664642 994879
rect 661670 994827 664642 994855
rect 664694 994827 664700 994879
rect 665409 994831 665415 994883
rect 665467 994855 674800 994883
rect 665467 994831 665473 994855
rect 661670 994799 661698 994827
rect 660923 994771 661698 994799
rect 665638 994687 665644 994711
rect 661123 994659 665644 994687
rect 665696 994659 665702 994711
rect 666481 994663 666487 994715
rect 666539 994687 674632 994715
rect 666539 994663 666545 994687
rect 665832 994631 665838 994655
rect 662034 994603 665838 994631
rect 665890 994603 665896 994655
rect 666600 994631 666611 994659
rect 666605 994607 666611 994631
rect 666663 994631 674576 994659
rect 666663 994607 666669 994631
rect 662034 994575 662062 994603
rect 661323 994547 662062 994575
rect 42851 892083 42879 892517
rect 42851 892055 42935 892083
rect 42715 888765 42767 888771
rect 42715 888707 42767 888713
rect 42463 608715 42515 608721
rect 42463 608657 42515 608663
rect 42655 888116 42707 888122
rect 42655 888058 42707 888064
rect 42211 352330 42263 352336
rect 40557 352265 40569 352317
rect 40739 352265 40751 352317
rect 42211 352272 42263 352278
rect 42403 608066 42455 608072
rect 42403 608008 42455 608014
rect 42151 351681 42203 351687
rect 40629 351665 40681 351677
rect 41169 351619 41181 351671
rect 41351 351619 41363 351671
rect 42151 351623 42203 351629
rect 40629 351435 40681 351447
rect 41241 351395 41293 351407
rect 41241 351165 41293 351177
rect 40557 351069 40569 351121
rect 40739 351069 40751 351121
rect 40629 350469 40681 350481
rect 41159 350423 41171 350475
rect 41341 350423 41353 350475
rect 40629 350239 40681 350251
rect 41241 350199 41293 350211
rect 41241 349969 41293 349981
rect 40557 349873 40569 349925
rect 40739 349873 40751 349925
rect 40629 349273 40681 349285
rect 41169 349227 41181 349279
rect 41351 349227 41363 349279
rect 40629 349043 40681 349055
rect 41241 349003 41293 349015
rect 41241 348773 41293 348785
rect 40557 348677 40569 348729
rect 40739 348677 40751 348729
rect 40629 348077 40681 348089
rect 41169 348031 41181 348083
rect 41351 348031 41363 348083
rect 40629 347847 40681 347859
rect 41241 347807 41293 347819
rect 41241 347577 41293 347589
rect 40557 347481 40569 347533
rect 40739 347481 40751 347533
rect 40629 346881 40681 346893
rect 41169 346835 41181 346887
rect 41351 346835 41363 346887
rect 40629 346651 40681 346663
rect 41241 346611 41293 346623
rect 41241 346381 41293 346393
rect 40557 346285 40569 346337
rect 40739 346285 40751 346337
rect 40629 345685 40681 345697
rect 41169 345639 41181 345691
rect 41351 345639 41363 345691
rect 40629 345455 40681 345467
rect 41241 345415 41293 345427
rect 41241 345185 41293 345197
rect 40557 345089 40569 345141
rect 40739 345089 40751 345141
rect 40629 344489 40681 344501
rect 41169 344443 41181 344495
rect 41351 344443 41363 344495
rect 40629 344259 40681 344271
rect 41241 344219 41293 344231
rect 41241 343989 41293 344001
rect 40557 343893 40569 343945
rect 40739 343893 40751 343945
rect 40629 343293 40681 343305
rect 41169 343247 41181 343299
rect 41351 343247 41363 343299
rect 40629 343133 40637 343161
rect 40671 343133 40681 343161
rect 40629 343063 40681 343075
rect 41241 343023 41293 343035
rect 41241 342793 41293 342805
rect 40557 342697 40569 342749
rect 40739 342697 40751 342749
rect 40629 342097 40681 342109
rect 41169 342051 41181 342103
rect 41351 342051 41363 342103
rect 40629 341867 40681 341879
rect 41241 341827 41293 341839
rect 41241 341597 41293 341609
rect 40557 341501 40569 341553
rect 40739 341501 40751 341553
rect 40629 340901 40681 340913
rect 41169 340855 41181 340907
rect 41351 340855 41363 340907
rect 40629 340671 40681 340683
rect 41241 340631 41293 340643
rect 41241 340401 41293 340413
rect 40557 340305 40569 340357
rect 40739 340305 40751 340357
rect 40629 339705 40681 339717
rect 41169 339659 41181 339711
rect 41351 339659 41363 339711
rect 40629 339475 40681 339487
rect 41241 339435 41293 339447
rect 41241 339205 41293 339217
rect 40557 339109 40569 339161
rect 40739 339109 40751 339161
rect 40629 338509 40681 338521
rect 41169 338463 41181 338515
rect 41351 338463 41363 338515
rect 40629 338279 40681 338291
rect 41241 338239 41293 338251
rect 41241 338009 41293 338021
rect 40557 337913 40569 337965
rect 40739 337913 40751 337965
rect 40629 337313 40681 337325
rect 41169 337267 41181 337319
rect 41351 337267 41363 337319
rect 40629 337083 40681 337095
rect 41241 337043 41293 337055
rect 41241 336813 41293 336825
rect 40557 336717 40569 336769
rect 40739 336717 40751 336769
rect 40629 336117 40681 336129
rect 41169 336071 41181 336123
rect 41351 336071 41363 336123
rect 40629 335887 40681 335899
rect 41241 335847 41293 335859
rect 41241 335617 41293 335629
rect 40557 335521 40569 335573
rect 40739 335521 40751 335573
rect 40629 334921 40681 334933
rect 41169 334875 41181 334927
rect 41351 334875 41363 334927
rect 40629 334691 40681 334703
rect 42151 45188 42179 351623
rect 42207 351557 42259 351563
rect 42207 351499 42259 351505
rect 42207 45244 42235 351499
rect 42403 351310 42431 608008
rect 42379 351304 42431 351310
rect 42379 351246 42431 351252
rect 42459 607942 42511 607948
rect 42459 607884 42511 607890
rect 42459 351140 42487 607884
rect 42655 607719 42683 888058
rect 42631 607713 42683 607719
rect 42631 607655 42683 607661
rect 42711 887992 42763 887998
rect 42711 887934 42763 887940
rect 42711 607525 42739 887934
rect 42907 887745 42935 892055
rect 42883 887739 42935 887745
rect 42883 887681 42935 887687
rect 42963 887575 42991 892317
rect 43075 891676 43103 892117
rect 43075 891648 43159 891676
rect 42939 887569 42991 887575
rect 42939 887511 42991 887517
rect 42687 607519 42739 607525
rect 42687 607461 42739 607467
rect 42879 886920 42931 886926
rect 42879 886862 42931 886868
rect 42435 351134 42487 351140
rect 42435 351076 42487 351082
rect 42627 606870 42679 606876
rect 42627 606812 42679 606818
rect 42375 350485 42427 350491
rect 42375 350427 42427 350433
rect 42375 45356 42403 350427
rect 42431 350361 42483 350367
rect 42431 350303 42483 350309
rect 42431 45412 42459 350303
rect 42627 350138 42655 606812
rect 42603 350132 42655 350138
rect 42603 350074 42655 350080
rect 42683 606746 42735 606752
rect 42683 606688 42735 606694
rect 42683 349944 42711 606688
rect 42879 606499 42907 886862
rect 42855 606493 42907 606499
rect 42855 606435 42907 606441
rect 42935 886796 42987 886802
rect 42935 886738 42987 886744
rect 42935 606329 42963 886738
rect 43131 886573 43159 891648
rect 43107 886567 43159 886573
rect 43107 886509 43159 886515
rect 43187 886379 43215 891917
rect 43163 886373 43215 886379
rect 43163 886315 43215 886321
rect 42911 606323 42963 606329
rect 42911 606265 42963 606271
rect 43103 885724 43155 885730
rect 43103 885666 43155 885672
rect 42659 349938 42711 349944
rect 42659 349880 42711 349886
rect 42851 605674 42903 605680
rect 42851 605616 42903 605622
rect 42599 349289 42651 349295
rect 42599 349231 42651 349237
rect 42599 45524 42627 349231
rect 42655 349165 42707 349171
rect 42655 349107 42707 349113
rect 42655 45580 42683 349107
rect 42851 348918 42879 605616
rect 42827 348912 42879 348918
rect 42827 348854 42879 348860
rect 42907 605550 42959 605556
rect 42907 605492 42959 605498
rect 42907 348748 42935 605492
rect 43103 605327 43131 885666
rect 43079 605321 43131 605327
rect 43079 605263 43131 605269
rect 43159 885600 43211 885606
rect 43159 885542 43211 885548
rect 43159 605133 43187 885542
rect 674044 727608 674072 728121
rect 674044 727580 674128 727608
rect 674100 721423 674128 727580
rect 674156 721617 674184 728321
rect 674268 727990 674296 728521
rect 674268 727962 674352 727990
rect 674324 722619 674352 727962
rect 674380 722813 674408 728721
rect 674548 723815 674576 994631
rect 674604 724009 674632 994687
rect 674772 725011 674800 994855
rect 674828 725205 674856 994911
rect 674996 726207 675024 995079
rect 675052 726401 675080 995135
rect 675248 727403 675276 995303
rect 675304 727573 675332 995359
rect 676328 727658 676380 727670
rect 675304 727567 675356 727573
rect 675304 727509 675356 727515
rect 676328 727428 676380 727440
rect 675248 727397 675300 727403
rect 675248 727339 675300 727345
rect 676870 727332 676882 727384
rect 677052 727332 677064 727384
rect 675308 726748 675360 726754
rect 675308 726690 675360 726696
rect 675252 726624 675304 726630
rect 675252 726566 675304 726572
rect 675052 726395 675104 726401
rect 675052 726337 675104 726343
rect 674996 726201 675048 726207
rect 674996 726143 675048 726149
rect 675056 725552 675108 725558
rect 675056 725494 675108 725500
rect 675000 725428 675052 725434
rect 675000 725370 675052 725376
rect 674828 725199 674880 725205
rect 674828 725141 674880 725147
rect 674772 725005 674824 725011
rect 674772 724947 674824 724953
rect 674832 724356 674884 724362
rect 674832 724298 674884 724304
rect 674776 724232 674828 724238
rect 674776 724174 674828 724180
rect 674604 724003 674656 724009
rect 674604 723945 674656 723951
rect 674548 723809 674600 723815
rect 674548 723751 674600 723757
rect 674608 723160 674660 723166
rect 674608 723102 674660 723108
rect 674552 723036 674604 723042
rect 674552 722978 674604 722984
rect 674380 722807 674432 722813
rect 674380 722749 674432 722755
rect 674324 722613 674376 722619
rect 674324 722555 674376 722561
rect 674384 721964 674436 721970
rect 674384 721906 674436 721912
rect 674328 721840 674380 721846
rect 674328 721782 674380 721788
rect 674156 721611 674208 721617
rect 674156 721553 674208 721559
rect 674100 721417 674152 721423
rect 674100 721359 674152 721365
rect 674160 720768 674212 720774
rect 674160 720710 674212 720716
rect 674128 720650 674156 720655
rect 674104 720644 674156 720650
rect 674104 720586 674156 720592
rect 43271 612349 43299 612956
rect 43271 612321 43355 612349
rect 43135 605127 43187 605133
rect 43135 605069 43187 605075
rect 42883 348742 42935 348748
rect 42883 348684 42935 348690
rect 43075 604478 43127 604484
rect 43075 604420 43127 604426
rect 42823 348093 42875 348099
rect 42823 348035 42875 348041
rect 42823 45692 42851 348035
rect 42879 347969 42931 347975
rect 42879 347911 42931 347917
rect 42879 45748 42907 347911
rect 43075 347746 43103 604420
rect 43051 347740 43103 347746
rect 43051 347682 43103 347688
rect 43131 604354 43183 604360
rect 43131 604296 43183 604302
rect 43131 347552 43159 604296
rect 43327 604131 43355 612321
rect 43303 604125 43355 604131
rect 43303 604067 43355 604073
rect 43383 603937 43411 612756
rect 43495 611937 43523 612556
rect 43495 611909 43579 611937
rect 43359 603931 43411 603937
rect 43359 603873 43411 603879
rect 43107 347546 43159 347552
rect 43107 347488 43159 347494
rect 43299 603282 43351 603288
rect 43299 603224 43351 603230
rect 43047 346897 43099 346903
rect 43047 346839 43099 346845
rect 43047 45860 43075 346839
rect 43103 346773 43155 346779
rect 43103 346715 43155 346721
rect 43103 45916 43131 346715
rect 43299 346550 43327 603224
rect 43275 346544 43327 346550
rect 43275 346486 43327 346492
rect 43355 603158 43407 603164
rect 43355 603100 43407 603106
rect 43355 346356 43383 603100
rect 43551 602935 43579 611909
rect 43527 602929 43579 602935
rect 43527 602871 43579 602877
rect 43607 602741 43635 612356
rect 43719 611534 43747 612156
rect 43719 611506 43803 611534
rect 43583 602735 43635 602741
rect 43583 602677 43635 602683
rect 43331 346350 43383 346356
rect 43331 346292 43383 346298
rect 43523 602086 43575 602092
rect 43523 602028 43575 602034
rect 43271 345701 43323 345707
rect 43271 345643 43323 345649
rect 43271 46028 43299 345643
rect 43327 345577 43379 345583
rect 43327 345519 43379 345525
rect 43327 46084 43355 345519
rect 43523 345354 43551 602028
rect 43499 345348 43551 345354
rect 43499 345290 43551 345296
rect 43579 601962 43631 601968
rect 43579 601904 43631 601910
rect 43579 345160 43607 601904
rect 43775 601739 43803 611506
rect 43751 601733 43803 601739
rect 43751 601675 43803 601681
rect 43831 601545 43859 611956
rect 43943 611157 43971 611756
rect 43943 611129 44027 611157
rect 43807 601539 43859 601545
rect 43807 601481 43859 601487
rect 43555 345154 43607 345160
rect 43555 345096 43607 345102
rect 43747 600890 43799 600896
rect 43747 600832 43799 600838
rect 43495 344505 43547 344511
rect 43495 344447 43547 344453
rect 43495 46196 43523 344447
rect 43551 344381 43603 344387
rect 43551 344323 43603 344329
rect 43551 46252 43579 344323
rect 43747 344158 43775 600832
rect 43723 344152 43775 344158
rect 43723 344094 43775 344100
rect 43803 600766 43855 600772
rect 43803 600708 43855 600714
rect 43803 343964 43831 600708
rect 43999 600543 44027 611129
rect 43975 600537 44027 600543
rect 43975 600479 44027 600485
rect 44055 600349 44083 611556
rect 44167 610759 44195 611356
rect 44167 610731 44251 610759
rect 44031 600343 44083 600349
rect 44031 600285 44083 600291
rect 43779 343958 43831 343964
rect 43779 343900 43831 343906
rect 43971 599694 44023 599700
rect 43971 599636 44023 599642
rect 43719 343309 43771 343315
rect 43719 343251 43771 343257
rect 43719 46364 43747 343251
rect 43775 343185 43827 343191
rect 43775 343127 43827 343133
rect 43775 46420 43803 343127
rect 43971 342962 43999 599636
rect 43947 342956 43999 342962
rect 43947 342898 43999 342904
rect 44027 599570 44079 599576
rect 44027 599512 44079 599518
rect 44027 342768 44055 599512
rect 44223 599347 44251 610731
rect 44199 599341 44251 599347
rect 44199 599283 44251 599289
rect 44279 599153 44307 611156
rect 44391 610321 44419 610956
rect 44391 610293 44475 610321
rect 44255 599147 44307 599153
rect 44255 599089 44307 599095
rect 44003 342762 44055 342768
rect 44003 342704 44055 342710
rect 44195 598498 44247 598504
rect 44195 598440 44247 598446
rect 43943 342113 43995 342119
rect 43943 342055 43995 342061
rect 43943 46532 43971 342055
rect 43999 341989 44051 341995
rect 43999 341931 44051 341937
rect 43999 46588 44027 341931
rect 44195 341766 44223 598440
rect 44171 341760 44223 341766
rect 44171 341702 44223 341708
rect 44251 598374 44303 598380
rect 44251 598316 44303 598322
rect 44251 341572 44279 598316
rect 44447 598151 44475 610293
rect 44423 598145 44475 598151
rect 44423 598087 44475 598093
rect 44503 597957 44531 610756
rect 44479 597951 44531 597957
rect 44479 597893 44531 597899
rect 44227 341566 44279 341572
rect 44227 341508 44279 341514
rect 44419 597302 44471 597308
rect 44419 597244 44471 597250
rect 44167 340917 44219 340923
rect 44167 340859 44219 340865
rect 44167 46700 44195 340859
rect 44223 340793 44275 340799
rect 44223 340735 44275 340741
rect 44223 46756 44251 340735
rect 44419 340570 44447 597244
rect 44395 340564 44447 340570
rect 44395 340506 44447 340512
rect 44475 597178 44527 597184
rect 44475 597120 44527 597126
rect 44475 340376 44503 597120
rect 672728 453370 672756 454055
rect 672728 453342 672812 453370
rect 672784 440223 672812 453342
rect 672840 440417 672868 454255
rect 672952 453758 672980 454455
rect 672952 453730 673036 453758
rect 673008 441419 673036 453730
rect 673064 441613 673092 454655
rect 673176 454180 673204 454855
rect 673176 454152 673260 454180
rect 673232 442615 673260 454152
rect 673288 442809 673316 455055
rect 673400 454622 673428 455255
rect 673400 454594 673484 454622
rect 673456 443811 673484 454594
rect 673512 444005 673540 455455
rect 673624 455002 673652 455655
rect 673624 454974 673708 455002
rect 673680 445007 673708 454974
rect 673736 445201 673764 455855
rect 673848 455378 673876 456055
rect 673848 455350 673932 455378
rect 673904 446203 673932 455350
rect 673960 446397 673988 456255
rect 674128 447399 674156 720586
rect 674184 447593 674212 720710
rect 674352 448595 674380 721782
rect 674408 448789 674436 721906
rect 674576 449791 674604 722978
rect 674632 449961 674660 723102
rect 674800 450987 674828 724174
rect 674856 451181 674884 724298
rect 675024 452183 675052 725370
rect 675080 452353 675108 725494
rect 675276 453379 675304 726566
rect 675332 453573 675360 726690
rect 676258 726686 676270 726738
rect 676440 726686 676452 726738
rect 676940 726732 676992 726744
rect 676940 726502 676992 726514
rect 676328 726462 676380 726474
rect 676328 726232 676380 726244
rect 676870 726136 676882 726188
rect 677052 726136 677064 726188
rect 676258 725490 676270 725542
rect 676440 725490 676452 725542
rect 676940 725536 676992 725548
rect 676940 725306 676992 725318
rect 676328 725266 676380 725278
rect 676328 725036 676380 725048
rect 676870 724940 676882 724992
rect 677052 724940 677064 724992
rect 676258 724294 676270 724346
rect 676440 724294 676452 724346
rect 676940 724340 676992 724352
rect 676940 724110 676992 724122
rect 676328 724070 676380 724082
rect 676328 723840 676380 723852
rect 676870 723744 676882 723796
rect 677052 723744 677064 723796
rect 676258 723098 676270 723150
rect 676440 723098 676452 723150
rect 676940 723144 676992 723156
rect 676940 722914 676992 722926
rect 676328 722874 676380 722886
rect 676328 722644 676380 722656
rect 676870 722548 676882 722600
rect 677052 722548 677064 722600
rect 676258 721902 676270 721954
rect 676440 721902 676452 721954
rect 676940 721948 676992 721960
rect 676940 721718 676992 721730
rect 676328 721678 676380 721690
rect 676328 721448 676380 721460
rect 676870 721352 676882 721404
rect 677052 721352 677064 721404
rect 676258 720706 676270 720758
rect 676440 720706 676452 720758
rect 676940 720752 676992 720764
rect 676940 720522 676992 720534
rect 676328 453634 676380 453646
rect 675332 453567 675384 453573
rect 675332 453509 675384 453515
rect 676328 453404 676380 453416
rect 675276 453373 675328 453379
rect 675276 453315 675328 453321
rect 676870 453308 676882 453360
rect 677052 453308 677064 453360
rect 675336 452724 675388 452730
rect 675336 452666 675388 452672
rect 675280 452600 675332 452606
rect 675280 452542 675332 452548
rect 675080 452347 675132 452353
rect 675080 452289 675132 452295
rect 675024 452177 675076 452183
rect 675024 452119 675076 452125
rect 675084 451528 675136 451534
rect 675084 451470 675136 451476
rect 675028 451404 675080 451410
rect 675028 451346 675080 451352
rect 674856 451175 674908 451181
rect 674856 451117 674908 451123
rect 674800 450981 674852 450987
rect 674800 450923 674852 450929
rect 674860 450332 674912 450338
rect 674860 450274 674912 450280
rect 674804 450208 674856 450214
rect 674804 450150 674856 450156
rect 674632 449955 674684 449961
rect 674632 449897 674684 449903
rect 674576 449785 674628 449791
rect 674576 449727 674628 449733
rect 674636 449136 674688 449142
rect 674636 449078 674688 449084
rect 674580 449012 674632 449018
rect 674580 448954 674632 448960
rect 674408 448783 674460 448789
rect 674408 448725 674460 448731
rect 674352 448589 674404 448595
rect 674352 448531 674404 448537
rect 674412 447940 674464 447946
rect 674412 447882 674464 447888
rect 674356 447816 674408 447822
rect 674356 447758 674408 447764
rect 674184 447587 674236 447593
rect 674184 447529 674236 447535
rect 674128 447393 674180 447399
rect 674128 447335 674180 447341
rect 674188 446744 674240 446750
rect 674188 446686 674240 446692
rect 674132 446620 674184 446626
rect 674132 446562 674184 446568
rect 673960 446391 674012 446397
rect 673960 446333 674012 446339
rect 673904 446197 673956 446203
rect 673904 446139 673956 446145
rect 673964 445548 674016 445554
rect 673964 445490 674016 445496
rect 673908 445424 673960 445430
rect 673908 445366 673960 445372
rect 673736 445195 673788 445201
rect 673736 445137 673788 445143
rect 673680 445001 673732 445007
rect 673680 444943 673732 444949
rect 673740 444352 673792 444358
rect 673740 444294 673792 444300
rect 673684 444228 673736 444234
rect 673684 444170 673736 444176
rect 673512 443999 673564 444005
rect 673512 443941 673564 443947
rect 673456 443805 673508 443811
rect 673456 443747 673508 443753
rect 673516 443156 673568 443162
rect 673516 443098 673568 443104
rect 673460 443032 673512 443038
rect 673460 442974 673512 442980
rect 673288 442803 673340 442809
rect 673288 442745 673340 442751
rect 673232 442609 673284 442615
rect 673232 442551 673284 442557
rect 673292 441960 673344 441966
rect 673292 441902 673344 441908
rect 673236 441836 673288 441842
rect 673236 441778 673288 441784
rect 673064 441607 673116 441613
rect 673064 441549 673116 441555
rect 673008 441413 673060 441419
rect 673008 441355 673060 441361
rect 673068 440764 673120 440770
rect 673068 440706 673120 440712
rect 673012 440640 673064 440646
rect 673012 440582 673064 440588
rect 672840 440411 672892 440417
rect 672840 440353 672892 440359
rect 672784 440217 672836 440223
rect 672784 440159 672836 440165
rect 672844 439568 672896 439574
rect 672844 439510 672896 439516
rect 672788 439444 672840 439450
rect 672788 439386 672840 439392
rect 44587 354170 44615 354730
rect 44587 354142 44671 354170
rect 44451 340370 44503 340376
rect 44451 340312 44503 340318
rect 44391 339721 44443 339727
rect 44391 339663 44443 339669
rect 44391 46868 44419 339663
rect 44447 339597 44499 339603
rect 44447 339539 44499 339545
rect 44447 46924 44475 339539
rect 44643 339374 44671 354142
rect 44619 339368 44671 339374
rect 44619 339310 44671 339316
rect 44699 339180 44727 354530
rect 44811 353795 44839 354330
rect 44811 353767 44895 353795
rect 44675 339174 44727 339180
rect 44675 339116 44727 339122
rect 44615 338525 44667 338531
rect 44615 338467 44667 338473
rect 44615 47036 44643 338467
rect 44671 338401 44723 338407
rect 44671 338343 44723 338349
rect 44671 47092 44699 338343
rect 44867 338178 44895 353767
rect 44843 338172 44895 338178
rect 44843 338114 44895 338120
rect 44923 337984 44951 354130
rect 45035 353383 45063 353930
rect 45035 353355 45119 353383
rect 44899 337978 44951 337984
rect 44899 337920 44951 337926
rect 44839 337329 44891 337335
rect 44839 337271 44891 337277
rect 44839 47204 44867 337271
rect 44895 337205 44947 337211
rect 44895 337147 44947 337153
rect 44895 47260 44923 337147
rect 45091 336958 45119 353355
rect 45067 336952 45119 336958
rect 45067 336894 45119 336900
rect 45147 336788 45175 353730
rect 45259 352982 45287 353530
rect 45259 352954 45343 352982
rect 45123 336782 45175 336788
rect 45123 336724 45175 336730
rect 45063 336133 45115 336139
rect 45063 336075 45115 336081
rect 45063 47372 45091 336075
rect 45119 336009 45171 336015
rect 45119 335951 45171 335957
rect 45119 47428 45147 335951
rect 45315 335786 45343 352954
rect 45291 335780 45343 335786
rect 45291 335722 45343 335728
rect 45371 335592 45399 353330
rect 45347 335586 45399 335592
rect 45347 335528 45399 335534
rect 45287 334937 45339 334943
rect 45287 334879 45339 334885
rect 45287 47540 45315 334879
rect 45343 334813 45395 334819
rect 45343 334755 45395 334761
rect 45343 47596 45371 334755
rect 672812 238848 672840 439386
rect 672756 238820 672840 238848
rect 672756 238050 672784 238820
rect 672868 237850 672896 439510
rect 673036 238360 673064 440582
rect 672980 238332 673064 238360
rect 672980 237650 673008 238332
rect 673092 237450 673120 440706
rect 673260 238014 673288 441778
rect 673204 237986 673288 238014
rect 673204 237250 673232 237986
rect 673316 237050 673344 441902
rect 673484 237648 673512 442974
rect 673428 237620 673512 237648
rect 673428 236850 673456 237620
rect 673540 236650 673568 443098
rect 673708 237204 673736 444170
rect 673652 237176 673736 237204
rect 673652 236450 673680 237176
rect 673764 236250 673792 444294
rect 673932 236798 673960 445366
rect 673876 236770 673960 236798
rect 673876 236050 673904 236770
rect 673988 235850 674016 445490
rect 674156 236400 674184 446562
rect 674100 236372 674184 236400
rect 674100 235650 674128 236372
rect 674212 235450 674240 446686
rect 674380 236022 674408 447758
rect 674324 235994 674408 236022
rect 674324 235250 674352 235994
rect 674436 235050 674464 447882
rect 674604 235640 674632 448954
rect 674548 235612 674632 235640
rect 674548 234850 674576 235612
rect 674660 234650 674688 449078
rect 674828 235254 674856 450150
rect 674772 235226 674856 235254
rect 674772 234450 674800 235226
rect 674884 234250 674912 450274
rect 675052 234836 675080 451346
rect 674996 234808 675080 234836
rect 674996 234050 675024 234808
rect 675108 233850 675136 451470
rect 675304 234436 675332 452542
rect 675248 234408 675332 234436
rect 675248 233650 675276 234408
rect 675360 233450 675388 452666
rect 676258 452662 676270 452714
rect 676440 452662 676452 452714
rect 676940 452708 676992 452720
rect 676940 452478 676992 452490
rect 676328 452438 676380 452450
rect 676328 452208 676380 452220
rect 676870 452112 676882 452164
rect 677052 452112 677064 452164
rect 676258 451466 676270 451518
rect 676440 451466 676452 451518
rect 676940 451512 676992 451524
rect 676940 451282 676992 451294
rect 676328 451242 676380 451254
rect 676328 451012 676380 451024
rect 676870 450916 676882 450968
rect 677052 450916 677064 450968
rect 676258 450270 676270 450322
rect 676440 450270 676452 450322
rect 676940 450316 676992 450328
rect 676940 450086 676992 450098
rect 676328 450046 676380 450058
rect 676328 449816 676380 449828
rect 676870 449720 676882 449772
rect 677052 449720 677064 449772
rect 676258 449074 676270 449126
rect 676440 449074 676452 449126
rect 676940 449120 676992 449132
rect 676940 448890 676992 448902
rect 676328 448850 676380 448862
rect 676328 448620 676380 448632
rect 676870 448524 676882 448576
rect 677052 448524 677064 448576
rect 676258 447878 676270 447930
rect 676440 447878 676452 447930
rect 676940 447924 676992 447936
rect 676940 447694 676992 447706
rect 676328 447654 676380 447666
rect 676328 447424 676380 447436
rect 676870 447328 676882 447380
rect 677052 447328 677064 447380
rect 676258 446682 676270 446734
rect 676440 446682 676452 446734
rect 676940 446728 676992 446740
rect 676940 446498 676992 446510
rect 676328 446458 676380 446470
rect 676328 446228 676380 446240
rect 676870 446132 676882 446184
rect 677052 446132 677064 446184
rect 676258 445486 676270 445538
rect 676440 445486 676452 445538
rect 676940 445532 676992 445544
rect 676940 445302 676992 445314
rect 676328 445262 676380 445274
rect 676328 445032 676380 445044
rect 676870 444936 676882 444988
rect 677052 444936 677064 444988
rect 676258 444290 676270 444342
rect 676440 444290 676452 444342
rect 676940 444336 676992 444348
rect 676940 444106 676992 444118
rect 676328 444066 676380 444078
rect 676328 443836 676380 443848
rect 676870 443740 676882 443792
rect 677052 443740 677064 443792
rect 676258 443094 676270 443146
rect 676440 443094 676452 443146
rect 676940 443140 676992 443152
rect 676940 442910 676992 442922
rect 676328 442870 676380 442882
rect 676328 442640 676380 442652
rect 676870 442544 676882 442596
rect 677052 442544 677064 442596
rect 676258 441898 676270 441950
rect 676440 441898 676452 441950
rect 676940 441944 676992 441956
rect 676940 441714 676992 441726
rect 676328 441674 676380 441686
rect 676328 441444 676380 441456
rect 676870 441348 676882 441400
rect 677052 441348 677064 441400
rect 676258 440702 676270 440754
rect 676440 440702 676452 440754
rect 676940 440748 676992 440760
rect 676940 440518 676992 440530
rect 676328 440478 676380 440490
rect 676328 440248 676380 440260
rect 676870 440152 676882 440204
rect 677052 440152 677064 440204
rect 676258 439506 676270 439558
rect 676440 439506 676452 439558
rect 676940 439552 676992 439564
rect 676940 439322 676992 439334
rect 429498 47624 429504 47648
rect 134098 47596 134104 47620
rect 45343 47568 134104 47596
rect 134156 47568 134162 47620
rect 134941 47572 134947 47624
rect 134999 47596 141269 47624
rect 134999 47572 135005 47596
rect 135170 47540 135176 47564
rect 45287 47512 135176 47540
rect 135228 47512 135234 47564
rect 135943 47516 135949 47568
rect 136001 47540 141213 47568
rect 136001 47516 136007 47540
rect 135294 47428 135300 47452
rect 45119 47400 135300 47428
rect 135352 47400 135358 47452
rect 136137 47404 136143 47456
rect 136195 47428 141101 47456
rect 136195 47404 136201 47428
rect 136366 47372 136372 47396
rect 45063 47344 136372 47372
rect 136424 47344 136430 47396
rect 137139 47348 137145 47400
rect 137197 47372 141045 47400
rect 137197 47348 137203 47372
rect 136490 47260 136496 47284
rect 44895 47232 136496 47260
rect 136548 47232 136554 47284
rect 137333 47236 137339 47288
rect 137391 47260 140933 47288
rect 137391 47236 137397 47260
rect 137562 47204 137568 47228
rect 44839 47176 137568 47204
rect 137620 47176 137626 47228
rect 138335 47180 138341 47232
rect 138393 47204 140877 47232
rect 138393 47180 138399 47204
rect 137686 47092 137692 47116
rect 44671 47064 137692 47092
rect 137744 47064 137750 47116
rect 138529 47068 138535 47120
rect 138587 47092 140765 47120
rect 138587 47068 138593 47092
rect 138758 47036 138764 47060
rect 44615 47008 138764 47036
rect 138816 47008 138822 47060
rect 139531 47012 139537 47064
rect 139589 47036 140709 47064
rect 139589 47012 139595 47036
rect 138882 46924 138888 46948
rect 44447 46896 138888 46924
rect 138940 46896 138946 46948
rect 139725 46900 139731 46952
rect 139783 46924 140651 46952
rect 139783 46900 139789 46924
rect 139954 46868 139960 46892
rect 44391 46840 139960 46868
rect 140012 46840 140018 46892
rect 140078 46756 140084 46780
rect 44223 46728 140084 46756
rect 140136 46728 140142 46780
rect 44167 46672 140585 46700
rect 43999 46560 140526 46588
rect 43943 46504 140462 46532
rect 43775 46392 140403 46420
rect 43719 46336 140347 46364
rect 43551 46224 140287 46252
rect 43495 46168 140231 46196
rect 140203 46084 140231 46168
rect 140259 46140 140287 46224
rect 140319 46196 140347 46336
rect 140375 46252 140403 46392
rect 140434 46308 140462 46504
rect 140498 46364 140526 46560
rect 140557 46420 140585 46672
rect 140623 46616 140651 46924
rect 140681 46672 140709 47036
rect 140737 46728 140765 47092
rect 140849 46784 140877 47204
rect 140905 46840 140933 47260
rect 141017 46896 141045 47372
rect 141073 46952 141101 47428
rect 141185 47008 141213 47540
rect 141241 47064 141269 47596
rect 155603 47596 429504 47624
rect 429556 47596 429562 47648
rect 430341 47600 430347 47652
rect 430399 47624 487832 47652
rect 430399 47600 430405 47624
rect 155603 47064 155631 47596
rect 430570 47568 430576 47592
rect 141241 47036 155631 47064
rect 155659 47540 430576 47568
rect 430628 47540 430634 47592
rect 431343 47544 431349 47596
rect 431401 47568 487776 47596
rect 431401 47544 431407 47568
rect 155659 47008 155687 47540
rect 430694 47456 430700 47480
rect 141185 46980 155687 47008
rect 155771 47428 430700 47456
rect 430752 47428 430758 47480
rect 431537 47432 431543 47484
rect 431595 47456 487608 47484
rect 431595 47432 431601 47456
rect 155771 46952 155799 47428
rect 431766 47400 431772 47424
rect 141073 46924 155799 46952
rect 155827 47372 431772 47400
rect 431824 47372 431830 47424
rect 432539 47376 432545 47428
rect 432597 47400 487552 47428
rect 432597 47376 432603 47400
rect 155827 46896 155855 47372
rect 431890 47288 431896 47312
rect 141017 46868 155855 46896
rect 155939 47260 431896 47288
rect 431948 47260 431954 47312
rect 432733 47264 432739 47316
rect 432791 47288 487384 47316
rect 432791 47264 432797 47288
rect 155939 46840 155967 47260
rect 432962 47232 432968 47256
rect 140905 46812 155967 46840
rect 155995 47204 432968 47232
rect 433020 47204 433026 47256
rect 433735 47208 433741 47260
rect 433793 47232 487328 47260
rect 433793 47208 433799 47232
rect 155995 46784 156023 47204
rect 433086 47120 433092 47144
rect 140849 46756 156023 46784
rect 156107 47092 433092 47120
rect 433144 47092 433150 47144
rect 433929 47096 433935 47148
rect 433987 47120 487160 47148
rect 433987 47096 433993 47120
rect 156107 46728 156135 47092
rect 434158 47064 434164 47088
rect 140737 46700 156135 46728
rect 156163 47036 434164 47064
rect 434216 47036 434222 47088
rect 434931 47040 434937 47092
rect 434989 47064 487104 47092
rect 434989 47040 434995 47064
rect 156163 46672 156191 47036
rect 434282 46952 434288 46976
rect 140681 46644 156191 46672
rect 156275 46924 434288 46952
rect 434340 46924 434346 46976
rect 435125 46928 435131 46980
rect 435183 46952 486936 46980
rect 435183 46928 435189 46952
rect 156275 46616 156303 46924
rect 435354 46896 435360 46920
rect 140623 46588 156303 46616
rect 156331 46868 435360 46896
rect 435412 46868 435418 46920
rect 436127 46872 436133 46924
rect 436185 46896 486880 46924
rect 436185 46872 436191 46896
rect 156331 46560 156359 46868
rect 435478 46784 435484 46808
rect 140727 46508 140733 46560
rect 140785 46532 156359 46560
rect 156443 46756 435484 46784
rect 435536 46756 435542 46808
rect 436297 46760 436303 46812
rect 436355 46784 486712 46812
rect 436355 46760 436361 46784
rect 140785 46508 140791 46532
rect 156443 46504 156471 46756
rect 436550 46728 436556 46752
rect 140897 46452 140903 46504
rect 140955 46476 156471 46504
rect 156499 46700 436556 46728
rect 436608 46700 436614 46752
rect 437323 46704 437329 46756
rect 437381 46728 486656 46756
rect 437381 46704 437387 46728
rect 140955 46452 140961 46476
rect 156499 46448 156527 46700
rect 436674 46616 436680 46640
rect 141150 46420 141156 46444
rect 140557 46392 141156 46420
rect 141208 46392 141214 46444
rect 141923 46396 141929 46448
rect 141981 46420 156527 46448
rect 156611 46588 436680 46616
rect 436732 46588 436738 46640
rect 437517 46592 437523 46644
rect 437575 46616 486488 46644
rect 437575 46592 437581 46616
rect 141981 46396 141987 46420
rect 156611 46392 156639 46588
rect 437746 46560 437752 46584
rect 141274 46364 141280 46388
rect 140498 46336 141280 46364
rect 141332 46336 141338 46388
rect 142117 46340 142123 46392
rect 142175 46364 156639 46392
rect 156667 46532 437752 46560
rect 437804 46532 437810 46584
rect 438519 46536 438525 46588
rect 438577 46560 486432 46588
rect 438577 46536 438583 46560
rect 142175 46340 142181 46364
rect 156667 46336 156695 46532
rect 437870 46448 437876 46472
rect 142346 46308 142352 46332
rect 140434 46280 142352 46308
rect 142404 46280 142410 46332
rect 143119 46284 143125 46336
rect 143177 46308 156695 46336
rect 156779 46420 437876 46448
rect 437928 46420 437934 46472
rect 438689 46424 438695 46476
rect 438747 46448 486264 46476
rect 438747 46424 438753 46448
rect 143177 46284 143183 46308
rect 156779 46280 156807 46420
rect 438942 46392 438948 46416
rect 142470 46252 142476 46276
rect 140375 46224 142476 46252
rect 142528 46224 142534 46276
rect 143289 46228 143295 46280
rect 143347 46252 156807 46280
rect 156835 46364 438948 46392
rect 439000 46364 439006 46416
rect 439715 46368 439721 46420
rect 439773 46392 486208 46420
rect 439773 46368 439779 46392
rect 143347 46228 143353 46252
rect 156835 46224 156863 46364
rect 439066 46280 439072 46304
rect 143542 46196 143548 46220
rect 140319 46168 143548 46196
rect 143600 46168 143606 46220
rect 144315 46172 144321 46224
rect 144373 46196 156863 46224
rect 156947 46252 439072 46280
rect 439124 46252 439130 46304
rect 439909 46256 439915 46308
rect 439967 46280 486040 46308
rect 439967 46256 439973 46280
rect 144373 46172 144379 46196
rect 156947 46168 156975 46252
rect 440138 46224 440144 46248
rect 143666 46140 143672 46164
rect 140259 46112 143672 46140
rect 143724 46112 143730 46164
rect 144509 46116 144515 46168
rect 144567 46140 156975 46168
rect 157003 46196 440144 46224
rect 440196 46196 440202 46248
rect 440911 46200 440917 46252
rect 440969 46224 485984 46252
rect 440969 46200 440975 46224
rect 144567 46116 144573 46140
rect 157003 46112 157031 46196
rect 440262 46112 440268 46136
rect 144738 46084 144744 46108
rect 43327 46056 140168 46084
rect 140203 46056 144744 46084
rect 144796 46056 144802 46108
rect 145511 46060 145517 46112
rect 145569 46084 157031 46112
rect 157072 46084 440268 46112
rect 440320 46084 440326 46136
rect 441105 46088 441111 46140
rect 441163 46112 485816 46140
rect 441163 46088 441169 46112
rect 145569 46060 145575 46084
rect 157072 46056 157100 46084
rect 441334 46056 441340 46080
rect 140140 46028 140168 46056
rect 144862 46028 144868 46052
rect 43271 46000 140109 46028
rect 140140 46000 144868 46028
rect 144920 46000 144926 46052
rect 145705 46004 145711 46056
rect 145763 46028 157100 46056
rect 157173 46028 441340 46056
rect 441392 46028 441398 46080
rect 442107 46032 442113 46084
rect 442165 46056 485760 46084
rect 442165 46032 442171 46056
rect 145763 46004 145769 46028
rect 157173 46000 157201 46028
rect 140081 45972 140109 46000
rect 145934 45972 145940 45996
rect 140081 45944 145940 45972
rect 145992 45944 145998 45996
rect 146707 45948 146713 46000
rect 146765 45972 157201 46000
rect 146765 45948 146771 45972
rect 441458 45944 441464 45968
rect 146058 45916 146064 45940
rect 43103 45888 146064 45916
rect 146116 45888 146122 45940
rect 146901 45892 146907 45944
rect 146959 45916 441464 45944
rect 441516 45916 441522 45968
rect 442301 45920 442307 45972
rect 442359 45944 485592 45972
rect 442359 45920 442365 45944
rect 146959 45892 146965 45916
rect 442530 45888 442536 45912
rect 147130 45860 147136 45884
rect 43047 45832 147136 45860
rect 147188 45832 147194 45884
rect 147903 45836 147909 45888
rect 147961 45860 442536 45888
rect 442588 45860 442594 45912
rect 443303 45864 443309 45916
rect 443361 45888 485536 45916
rect 443361 45864 443367 45888
rect 147961 45836 147967 45860
rect 442654 45776 442660 45800
rect 147254 45748 147260 45772
rect 42879 45720 147260 45748
rect 147312 45720 147318 45772
rect 148097 45724 148103 45776
rect 148155 45748 442660 45776
rect 442712 45748 442718 45800
rect 443497 45752 443503 45804
rect 443555 45776 485368 45804
rect 443555 45752 443561 45776
rect 148155 45724 148161 45748
rect 443726 45720 443732 45744
rect 148326 45692 148332 45716
rect 42823 45664 148332 45692
rect 148384 45664 148390 45716
rect 149099 45668 149105 45720
rect 149157 45692 443732 45720
rect 443784 45692 443790 45744
rect 444499 45696 444505 45748
rect 444557 45720 485312 45748
rect 444557 45696 444563 45720
rect 149157 45668 149163 45692
rect 443850 45608 443856 45632
rect 148450 45580 148456 45604
rect 42655 45552 148456 45580
rect 148508 45552 148514 45604
rect 149293 45556 149299 45608
rect 149351 45580 443856 45608
rect 443908 45580 443914 45632
rect 444693 45584 444699 45636
rect 444751 45608 485144 45636
rect 444751 45584 444757 45608
rect 149351 45556 149357 45580
rect 444922 45552 444928 45576
rect 149522 45524 149528 45548
rect 42599 45496 149528 45524
rect 149580 45496 149586 45548
rect 150295 45500 150301 45552
rect 150353 45524 444928 45552
rect 444980 45524 444986 45576
rect 445695 45528 445701 45580
rect 445753 45552 485088 45580
rect 445753 45528 445759 45552
rect 150353 45500 150359 45524
rect 445046 45440 445052 45464
rect 149646 45412 149652 45436
rect 42431 45384 149652 45412
rect 149704 45384 149710 45436
rect 150489 45388 150495 45440
rect 150547 45412 445052 45440
rect 445104 45412 445110 45464
rect 445889 45416 445895 45468
rect 445947 45440 484920 45468
rect 445947 45416 445953 45440
rect 150547 45388 150553 45412
rect 446118 45384 446124 45408
rect 150718 45356 150724 45380
rect 42375 45328 150724 45356
rect 150776 45328 150782 45380
rect 151491 45332 151497 45384
rect 151549 45356 446124 45384
rect 446176 45356 446182 45408
rect 446891 45360 446897 45412
rect 446949 45384 484864 45412
rect 446949 45360 446955 45384
rect 151549 45332 151555 45356
rect 446242 45272 446248 45296
rect 150842 45244 150848 45268
rect 42207 45216 150848 45244
rect 150900 45216 150906 45268
rect 151685 45220 151691 45272
rect 151743 45244 446248 45272
rect 446300 45244 446306 45296
rect 447085 45248 447091 45300
rect 447143 45272 484696 45300
rect 447143 45248 447149 45272
rect 151743 45220 151749 45244
rect 447314 45216 447320 45240
rect 151914 45188 151920 45212
rect 42151 45160 151920 45188
rect 151972 45160 151978 45212
rect 152687 45164 152693 45216
rect 152745 45188 447320 45216
rect 447372 45188 447378 45240
rect 448087 45192 448093 45244
rect 448145 45216 484640 45244
rect 448145 45192 448151 45216
rect 152745 45164 152751 45188
rect 447438 45104 447444 45128
rect 152038 45076 152044 45100
rect 131123 45048 152044 45076
rect 152096 45048 152102 45100
rect 152881 45052 152887 45104
rect 152939 45076 447444 45104
rect 447496 45076 447502 45128
rect 448281 45080 448287 45132
rect 448339 45104 484472 45132
rect 448339 45080 448345 45104
rect 152939 45052 152945 45076
rect 448510 45048 448516 45072
rect 153110 45020 153116 45044
rect 132046 44992 153116 45020
rect 153168 44992 153174 45044
rect 153883 44996 153889 45048
rect 153941 45020 448516 45048
rect 448568 45020 448574 45072
rect 449283 45024 449289 45076
rect 449341 45048 484416 45076
rect 449341 45024 449347 45048
rect 153941 44996 153947 45020
rect 131351 44964 132074 44992
rect 448634 44936 448640 44960
rect 153234 44908 153240 44932
rect 131523 44880 153240 44908
rect 153292 44880 153298 44932
rect 154077 44884 154083 44936
rect 154135 44908 448640 44936
rect 448692 44908 448698 44960
rect 449477 44912 449483 44964
rect 449535 44936 484248 44964
rect 449535 44912 449541 44936
rect 154135 44884 154141 44908
rect 449706 44880 449712 44904
rect 154306 44852 154312 44876
rect 132447 44824 154312 44852
rect 154364 44824 154370 44876
rect 155079 44828 155085 44880
rect 155137 44852 449712 44880
rect 449764 44852 449770 44904
rect 450479 44856 450485 44908
rect 450537 44880 484192 44908
rect 450537 44856 450543 44880
rect 155137 44828 155143 44852
rect 131751 44796 132475 44824
rect 449830 44768 449836 44792
rect 154430 44740 154436 44764
rect 131923 44712 154436 44740
rect 154488 44712 154494 44764
rect 155249 44716 155255 44768
rect 155307 44740 449836 44768
rect 449888 44740 449894 44792
rect 450649 44744 450655 44796
rect 450707 44768 484024 44796
rect 450707 44744 450713 44768
rect 155307 44716 155313 44740
rect 450902 44712 450908 44736
rect 155502 44684 155508 44708
rect 132852 44656 155508 44684
rect 155560 44656 155566 44708
rect 156275 44660 156281 44712
rect 156333 44684 450908 44712
rect 450960 44684 450966 44736
rect 451675 44688 451681 44740
rect 451733 44712 483968 44740
rect 451733 44688 451739 44712
rect 156333 44660 156339 44684
rect 132151 44628 132880 44656
rect 451026 44600 451032 44624
rect 155626 44572 155632 44596
rect 132323 44544 155632 44572
rect 155684 44544 155690 44596
rect 156469 44548 156475 44600
rect 156527 44572 451032 44600
rect 451084 44572 451090 44624
rect 451869 44576 451875 44628
rect 451927 44600 483800 44628
rect 451927 44576 451933 44600
rect 156527 44548 156533 44572
rect 452098 44544 452104 44568
rect 156698 44516 156704 44540
rect 133260 44488 156704 44516
rect 156756 44488 156762 44540
rect 157471 44492 157477 44544
rect 157529 44516 452104 44544
rect 452156 44516 452162 44568
rect 452871 44520 452877 44572
rect 452929 44544 483744 44572
rect 452929 44520 452935 44544
rect 157529 44492 157535 44516
rect 132551 44460 133288 44488
rect 452222 44432 452228 44456
rect 156822 44404 156828 44428
rect 133443 44376 156828 44404
rect 156880 44376 156886 44428
rect 157641 44380 157647 44432
rect 157699 44404 452228 44432
rect 452280 44404 452286 44456
rect 453041 44408 453047 44460
rect 453099 44432 483576 44460
rect 453099 44408 453105 44432
rect 157699 44380 157705 44404
rect 132751 44348 133471 44376
rect 453294 44320 453300 44344
rect 157894 44292 157900 44316
rect 133649 44264 157900 44292
rect 157952 44264 157958 44316
rect 158667 44268 158673 44320
rect 158725 44292 453300 44320
rect 453352 44292 453358 44344
rect 454067 44296 454073 44348
rect 454125 44320 483408 44348
rect 454125 44296 454131 44320
rect 158725 44268 158731 44292
rect 132951 44236 133677 44264
rect 453418 44208 453424 44232
rect 158018 44180 158024 44204
rect 133838 44152 158024 44180
rect 158076 44152 158082 44204
rect 158861 44156 158867 44208
rect 158919 44180 453424 44208
rect 453476 44180 453482 44232
rect 454261 44184 454267 44236
rect 454319 44208 483240 44236
rect 454319 44184 454325 44208
rect 158919 44156 158925 44180
rect 133151 44124 133866 44152
rect 134094 43272 134146 43284
rect 135290 43272 135342 43284
rect 134836 43162 134848 43214
rect 135066 43162 135078 43214
rect 134094 43090 134146 43102
rect 136486 43272 136538 43284
rect 136032 43162 136044 43214
rect 136262 43162 136274 43214
rect 135290 43090 135342 43102
rect 137682 43272 137734 43284
rect 137228 43162 137240 43214
rect 137458 43162 137470 43214
rect 136486 43090 136538 43102
rect 138878 43272 138930 43284
rect 138424 43162 138436 43214
rect 138654 43162 138666 43214
rect 137682 43090 137734 43102
rect 140074 43272 140126 43284
rect 139620 43162 139632 43214
rect 139850 43162 139862 43214
rect 138878 43090 138930 43102
rect 141270 43272 141322 43284
rect 140816 43162 140828 43214
rect 141046 43162 141058 43214
rect 140074 43090 140126 43102
rect 142466 43272 142518 43284
rect 142012 43162 142024 43214
rect 142242 43162 142254 43214
rect 141270 43090 141322 43102
rect 143662 43272 143714 43284
rect 143208 43162 143220 43214
rect 143438 43162 143450 43214
rect 142466 43090 142518 43102
rect 144858 43272 144910 43284
rect 144404 43162 144416 43214
rect 144634 43162 144646 43214
rect 143662 43090 143714 43102
rect 146054 43272 146106 43284
rect 145600 43162 145612 43214
rect 145830 43162 145842 43214
rect 144858 43090 144910 43102
rect 147250 43272 147302 43284
rect 146796 43162 146808 43214
rect 147026 43162 147038 43214
rect 146054 43090 146106 43102
rect 148446 43272 148498 43284
rect 147992 43162 148004 43214
rect 148222 43162 148234 43214
rect 147250 43090 147302 43102
rect 149642 43272 149694 43284
rect 149188 43162 149200 43214
rect 149418 43162 149430 43214
rect 148446 43090 148498 43102
rect 150838 43272 150890 43284
rect 150384 43162 150396 43214
rect 150614 43162 150626 43214
rect 149642 43090 149694 43102
rect 152034 43272 152086 43284
rect 151580 43162 151592 43214
rect 151810 43162 151822 43214
rect 150838 43090 150890 43102
rect 153230 43272 153282 43284
rect 152776 43162 152788 43214
rect 153006 43162 153018 43214
rect 152034 43090 152086 43102
rect 154426 43272 154478 43284
rect 153972 43162 153984 43214
rect 154202 43162 154214 43214
rect 153230 43090 153282 43102
rect 155622 43272 155674 43284
rect 155168 43162 155180 43214
rect 155398 43162 155410 43214
rect 154426 43090 154478 43102
rect 156818 43272 156870 43284
rect 156364 43162 156376 43214
rect 156594 43162 156606 43214
rect 155622 43090 155674 43102
rect 158014 43272 158066 43284
rect 157560 43162 157572 43214
rect 157790 43162 157802 43214
rect 156818 43090 156870 43102
rect 429494 43272 429546 43284
rect 158756 43162 158768 43214
rect 158986 43162 158998 43214
rect 158014 43090 158066 43102
rect 430690 43272 430742 43284
rect 430236 43162 430248 43214
rect 430466 43162 430478 43214
rect 429494 43090 429546 43102
rect 431886 43272 431938 43284
rect 431432 43162 431444 43214
rect 431662 43162 431674 43214
rect 430690 43090 430742 43102
rect 433082 43272 433134 43284
rect 432628 43162 432640 43214
rect 432858 43162 432870 43214
rect 431886 43090 431938 43102
rect 434278 43272 434330 43284
rect 433824 43162 433836 43214
rect 434054 43162 434066 43214
rect 433082 43090 433134 43102
rect 435474 43272 435526 43284
rect 435020 43162 435032 43214
rect 435250 43162 435262 43214
rect 434278 43090 434330 43102
rect 436670 43272 436722 43284
rect 436216 43162 436228 43214
rect 436446 43162 436458 43214
rect 435474 43090 435526 43102
rect 437866 43272 437918 43284
rect 437412 43162 437424 43214
rect 437642 43162 437654 43214
rect 436670 43090 436722 43102
rect 439062 43272 439114 43284
rect 438608 43162 438620 43214
rect 438838 43162 438850 43214
rect 437866 43090 437918 43102
rect 440258 43272 440310 43284
rect 439804 43162 439816 43214
rect 440034 43162 440046 43214
rect 439062 43090 439114 43102
rect 441454 43272 441506 43284
rect 441000 43162 441012 43214
rect 441230 43162 441242 43214
rect 440258 43090 440310 43102
rect 442650 43272 442702 43284
rect 442196 43162 442208 43214
rect 442426 43162 442438 43214
rect 441454 43090 441506 43102
rect 443846 43272 443898 43284
rect 443392 43162 443404 43214
rect 443622 43162 443634 43214
rect 442650 43090 442702 43102
rect 445042 43272 445094 43284
rect 444588 43162 444600 43214
rect 444818 43162 444830 43214
rect 443846 43090 443898 43102
rect 446238 43272 446290 43284
rect 445784 43162 445796 43214
rect 446014 43162 446026 43214
rect 445042 43090 445094 43102
rect 447434 43272 447486 43284
rect 446980 43162 446992 43214
rect 447210 43162 447222 43214
rect 446238 43090 446290 43102
rect 448630 43272 448682 43284
rect 448176 43162 448188 43214
rect 448406 43162 448418 43214
rect 447434 43090 447486 43102
rect 449826 43272 449878 43284
rect 449372 43162 449384 43214
rect 449602 43162 449614 43214
rect 448630 43090 448682 43102
rect 451022 43272 451074 43284
rect 450568 43162 450580 43214
rect 450798 43162 450810 43214
rect 449826 43090 449878 43102
rect 452218 43272 452270 43284
rect 451764 43162 451776 43214
rect 451994 43162 452006 43214
rect 451022 43090 451074 43102
rect 453414 43272 453466 43284
rect 452960 43162 452972 43214
rect 453190 43162 453202 43214
rect 452218 43090 452270 43102
rect 454156 43162 454168 43214
rect 454386 43162 454398 43214
rect 453414 43090 453466 43102
rect 135936 42660 135988 42672
rect 135106 42550 135118 42602
rect 135336 42550 135348 42602
rect 137132 42660 137184 42672
rect 136302 42550 136314 42602
rect 136532 42550 136544 42602
rect 135936 42478 135988 42490
rect 138328 42660 138380 42672
rect 137498 42550 137510 42602
rect 137728 42550 137740 42602
rect 137132 42478 137184 42490
rect 139524 42660 139576 42672
rect 138694 42550 138706 42602
rect 138924 42550 138936 42602
rect 138328 42478 138380 42490
rect 140720 42660 140772 42672
rect 139890 42550 139902 42602
rect 140120 42550 140132 42602
rect 139524 42478 139576 42490
rect 141916 42660 141968 42672
rect 141086 42550 141098 42602
rect 141316 42550 141328 42602
rect 140720 42478 140772 42490
rect 143112 42660 143164 42672
rect 142282 42550 142294 42602
rect 142512 42550 142524 42602
rect 141916 42478 141968 42490
rect 144308 42660 144360 42672
rect 143478 42550 143490 42602
rect 143708 42550 143720 42602
rect 143112 42478 143164 42490
rect 145504 42660 145556 42672
rect 144674 42550 144686 42602
rect 144904 42550 144916 42602
rect 144308 42478 144360 42490
rect 146700 42660 146752 42672
rect 145870 42550 145882 42602
rect 146100 42550 146112 42602
rect 145504 42478 145556 42490
rect 147896 42660 147948 42672
rect 147066 42550 147078 42602
rect 147296 42550 147308 42602
rect 146700 42478 146752 42490
rect 149092 42660 149144 42672
rect 148262 42550 148274 42602
rect 148492 42550 148504 42602
rect 147896 42478 147948 42490
rect 150288 42660 150340 42672
rect 149458 42550 149470 42602
rect 149688 42550 149700 42602
rect 149092 42478 149144 42490
rect 151484 42660 151536 42672
rect 150654 42550 150666 42602
rect 150884 42550 150896 42602
rect 150288 42478 150340 42490
rect 152680 42660 152732 42672
rect 151850 42550 151862 42602
rect 152080 42550 152092 42602
rect 151484 42478 151536 42490
rect 153876 42660 153928 42672
rect 153046 42550 153058 42602
rect 153276 42550 153288 42602
rect 152680 42478 152732 42490
rect 155072 42660 155124 42672
rect 154242 42550 154254 42602
rect 154472 42550 154484 42602
rect 153876 42478 153928 42490
rect 156268 42660 156320 42672
rect 155438 42550 155450 42602
rect 155668 42550 155680 42602
rect 155072 42478 155124 42490
rect 157464 42660 157516 42672
rect 156634 42550 156646 42602
rect 156864 42550 156876 42602
rect 156268 42478 156320 42490
rect 157464 42478 157516 42490
rect 158016 42660 158068 42672
rect 431336 42660 431388 42672
rect 158656 42550 158668 42602
rect 158886 42550 158898 42602
rect 430506 42550 430518 42602
rect 430736 42550 430748 42602
rect 158016 42478 158068 42490
rect 432532 42660 432584 42672
rect 431702 42550 431714 42602
rect 431932 42550 431944 42602
rect 431336 42478 431388 42490
rect 433728 42660 433780 42672
rect 432898 42550 432910 42602
rect 433128 42550 433140 42602
rect 432532 42478 432584 42490
rect 434924 42660 434976 42672
rect 434094 42550 434106 42602
rect 434324 42550 434336 42602
rect 433728 42478 433780 42490
rect 436120 42660 436172 42672
rect 435290 42550 435302 42602
rect 435520 42550 435532 42602
rect 434924 42478 434976 42490
rect 437316 42660 437368 42672
rect 436486 42550 436498 42602
rect 436716 42550 436728 42602
rect 436120 42478 436172 42490
rect 438512 42660 438564 42672
rect 437682 42550 437694 42602
rect 437912 42550 437924 42602
rect 437316 42478 437368 42490
rect 439708 42660 439760 42672
rect 438878 42550 438890 42602
rect 439108 42550 439120 42602
rect 438512 42478 438564 42490
rect 440904 42660 440956 42672
rect 440074 42550 440086 42602
rect 440304 42550 440316 42602
rect 439708 42478 439760 42490
rect 442100 42660 442152 42672
rect 441270 42550 441282 42602
rect 441500 42550 441512 42602
rect 440904 42478 440956 42490
rect 443296 42660 443348 42672
rect 442466 42550 442478 42602
rect 442696 42550 442708 42602
rect 442100 42478 442152 42490
rect 444492 42660 444544 42672
rect 443662 42550 443674 42602
rect 443892 42550 443904 42602
rect 443296 42478 443348 42490
rect 445688 42660 445740 42672
rect 444858 42550 444870 42602
rect 445088 42550 445100 42602
rect 444492 42478 444544 42490
rect 446884 42660 446936 42672
rect 446054 42550 446066 42602
rect 446284 42550 446296 42602
rect 445688 42478 445740 42490
rect 448080 42660 448132 42672
rect 447250 42550 447262 42602
rect 447480 42550 447492 42602
rect 446884 42478 446936 42490
rect 449276 42660 449328 42672
rect 448446 42550 448458 42602
rect 448676 42550 448688 42602
rect 448080 42478 448132 42490
rect 450472 42660 450524 42672
rect 449642 42550 449654 42602
rect 449872 42550 449884 42602
rect 449276 42478 449328 42490
rect 451668 42660 451720 42672
rect 450838 42550 450850 42602
rect 451068 42550 451080 42602
rect 450472 42478 450524 42490
rect 452864 42660 452916 42672
rect 452034 42550 452046 42602
rect 452264 42550 452276 42602
rect 451668 42478 451720 42490
rect 452864 42478 452916 42490
rect 453416 42660 453468 42672
rect 454056 42550 454068 42602
rect 454286 42550 454298 42602
rect 453416 42478 453468 42490
rect 483212 42356 483240 44208
rect 483380 42412 483408 44320
rect 483548 42468 483576 44432
rect 483716 42524 483744 44544
rect 483772 42580 483800 44600
rect 483939 42636 483967 44712
rect 483996 42692 484024 44768
rect 484164 42748 484192 44880
rect 484220 42804 484248 44936
rect 484388 42860 484416 45048
rect 484444 42916 484472 45104
rect 484612 42972 484640 45216
rect 484668 43028 484696 45272
rect 484836 43084 484864 45384
rect 484892 43140 484920 45440
rect 485060 43196 485088 45552
rect 485116 43252 485144 45608
rect 485284 43308 485312 45720
rect 485340 43364 485368 45776
rect 485508 43420 485536 45888
rect 485564 43476 485592 45944
rect 485732 43532 485760 46056
rect 485788 43588 485816 46112
rect 485956 43644 485984 46224
rect 486012 43700 486040 46280
rect 486180 43756 486208 46392
rect 486236 43812 486264 46448
rect 486404 43868 486432 46560
rect 486460 43924 486488 46616
rect 486628 43980 486656 46728
rect 486684 44036 486712 46784
rect 486852 44092 486880 46896
rect 486908 44148 486936 46952
rect 487076 44204 487104 47064
rect 487132 44260 487160 47120
rect 487300 44316 487328 47232
rect 487356 44372 487384 47288
rect 487524 44428 487552 47400
rect 487580 44484 487608 47456
rect 487748 44540 487776 47568
rect 487804 44596 487832 47624
rect 670936 45852 670964 224350
rect 671048 223698 671076 224546
rect 502852 45824 670964 45852
rect 670992 223670 671076 223698
rect 502852 44596 502880 45824
rect 670992 45796 671020 223670
rect 487804 44568 502880 44596
rect 502908 45768 671020 45796
rect 502908 44540 502936 45768
rect 671160 45684 671188 224740
rect 671272 224218 671300 224938
rect 487748 44512 502936 44540
rect 503076 45656 671188 45684
rect 671216 224190 671300 224218
rect 503076 44484 503104 45656
rect 671216 45628 671244 224190
rect 487580 44456 503104 44484
rect 503132 45600 671244 45628
rect 503132 44428 503160 45600
rect 671384 45516 671412 225138
rect 671496 224630 671524 225348
rect 487524 44400 503160 44428
rect 503300 45488 671412 45516
rect 671440 224602 671524 224630
rect 503300 44372 503328 45488
rect 671440 45460 671468 224602
rect 487356 44344 503328 44372
rect 503356 45432 671468 45460
rect 503356 44316 503384 45432
rect 671608 45348 671636 225542
rect 671720 225006 671748 225744
rect 487300 44288 503384 44316
rect 503524 45320 671636 45348
rect 671664 224978 671748 225006
rect 503524 44260 503552 45320
rect 671664 45292 671692 224978
rect 487132 44232 503552 44260
rect 503580 45264 671692 45292
rect 503580 44204 503608 45264
rect 671832 45180 671860 225936
rect 671944 225402 671972 226140
rect 487076 44176 503608 44204
rect 503748 45152 671860 45180
rect 671888 225374 671972 225402
rect 503748 44148 503776 45152
rect 671888 45124 671916 225374
rect 486908 44120 503776 44148
rect 503804 45096 671916 45124
rect 503804 44092 503832 45096
rect 672056 45012 672084 226340
rect 672168 225782 672196 226536
rect 486852 44064 503832 44092
rect 503972 44984 672084 45012
rect 672112 225754 672196 225782
rect 503972 44036 504000 44984
rect 672112 44956 672140 225754
rect 486684 44008 504000 44036
rect 504028 44928 672140 44956
rect 504028 43980 504056 44928
rect 672280 44844 672308 226738
rect 672392 226186 672420 226942
rect 486628 43952 504056 43980
rect 504196 44816 672308 44844
rect 672336 226158 672420 226186
rect 504196 43924 504224 44816
rect 672336 44788 672364 226158
rect 486460 43896 504224 43924
rect 504252 44760 672364 44788
rect 504252 43868 504280 44760
rect 672504 44676 672532 227138
rect 672616 226622 672644 227336
rect 486404 43840 504280 43868
rect 504420 44648 672532 44676
rect 672560 226594 672644 226622
rect 504420 43812 504448 44648
rect 672560 44620 672588 226594
rect 486236 43784 504448 43812
rect 504476 44592 672588 44620
rect 504476 43756 504504 44592
rect 672728 44508 672756 227538
rect 672840 227012 672868 227736
rect 486180 43728 504504 43756
rect 504644 44480 672756 44508
rect 672784 226984 672868 227012
rect 504644 43700 504672 44480
rect 672784 44452 672812 226984
rect 486012 43672 504672 43700
rect 504700 44424 672812 44452
rect 504700 43644 504728 44424
rect 672952 44340 672980 227938
rect 673064 227468 673092 228138
rect 485956 43616 504728 43644
rect 504868 44312 672980 44340
rect 673008 227440 673092 227468
rect 504868 43588 504896 44312
rect 673008 44284 673036 227440
rect 485788 43560 504896 43588
rect 504924 44256 673036 44284
rect 504924 43532 504952 44256
rect 673176 44172 673204 228338
rect 673288 227758 673316 228540
rect 485732 43504 504952 43532
rect 505092 44144 673204 44172
rect 673232 227730 673316 227758
rect 505092 43476 505120 44144
rect 673232 44116 673260 227730
rect 485564 43448 505120 43476
rect 505148 44088 673260 44116
rect 505148 43420 505176 44088
rect 673400 44004 673428 228736
rect 673512 228168 673540 228938
rect 485508 43392 505176 43420
rect 505316 43976 673428 44004
rect 673456 228140 673540 228168
rect 505316 43364 505344 43976
rect 673456 43948 673484 228140
rect 485340 43336 505344 43364
rect 505372 43920 673484 43948
rect 505372 43308 505400 43920
rect 673624 43836 673652 229138
rect 673736 228514 673764 229334
rect 485284 43280 505400 43308
rect 505540 43808 673652 43836
rect 673680 228486 673764 228514
rect 505540 43252 505568 43808
rect 673680 43780 673708 228486
rect 485116 43224 505568 43252
rect 505596 43752 673708 43780
rect 505596 43196 505624 43752
rect 673848 43668 673876 229534
rect 673960 228940 673988 229736
rect 485060 43168 505624 43196
rect 505764 43640 673876 43668
rect 673904 228912 673988 228940
rect 505764 43140 505792 43640
rect 673904 43612 673932 228912
rect 484892 43112 505792 43140
rect 505820 43584 673932 43612
rect 505820 43084 505848 43584
rect 674072 43500 674100 229936
rect 674184 229294 674212 230136
rect 484836 43056 505848 43084
rect 505988 43472 674100 43500
rect 674128 229266 674212 229294
rect 505988 43028 506016 43472
rect 674128 43444 674156 229266
rect 484668 43000 506016 43028
rect 506044 43416 674156 43444
rect 506044 42972 506072 43416
rect 674296 43332 674324 230288
rect 674408 229710 674436 230488
rect 484612 42944 506072 42972
rect 506212 43304 674324 43332
rect 674352 229682 674436 229710
rect 506212 42916 506240 43304
rect 674352 43276 674380 229682
rect 484444 42888 506240 42916
rect 506268 43248 674380 43276
rect 506268 42860 506296 43248
rect 674520 43164 674548 230690
rect 674632 230118 674660 230888
rect 484388 42832 506296 42860
rect 506436 43136 674548 43164
rect 674576 230090 674660 230118
rect 506436 42804 506464 43136
rect 674576 43108 674604 230090
rect 484220 42776 506464 42804
rect 506492 43080 674604 43108
rect 506492 42748 506520 43080
rect 674744 42996 674772 231088
rect 674856 230502 674884 231290
rect 484164 42720 506520 42748
rect 506660 42968 674772 42996
rect 674800 230474 674884 230502
rect 506660 42692 506688 42968
rect 674800 42940 674828 230474
rect 483996 42664 506688 42692
rect 506716 42912 674828 42940
rect 506716 42636 506744 42912
rect 674968 42828 674996 231490
rect 675080 230914 675108 231690
rect 483939 42608 506744 42636
rect 506884 42800 674996 42828
rect 675024 230886 675108 230914
rect 506884 42580 506912 42800
rect 675024 42772 675052 230886
rect 483772 42552 506912 42580
rect 506940 42744 675052 42772
rect 506940 42524 506968 42744
rect 675192 42660 675220 231888
rect 483716 42496 506968 42524
rect 507108 42632 675220 42660
rect 507108 42468 507136 42632
rect 675360 42548 675388 232090
rect 483548 42440 507136 42468
rect 507276 42520 675388 42548
rect 507276 42412 507304 42520
rect 675528 42449 675556 232290
rect 483380 42384 507304 42412
rect 507444 42421 675556 42449
rect 507444 42356 507472 42421
rect 483212 42328 507472 42356
<< via1 >>
rect 417027 997507 417384 997567
rect 663637 997425 663994 997485
rect 168590 997178 168947 997238
rect 416862 997217 416870 997387
rect 416870 997217 416904 997387
rect 416904 997217 416914 997387
rect 417514 997319 417732 997327
rect 417514 997285 417732 997319
rect 417514 997275 417732 997285
rect 662263 997135 662271 997305
rect 662271 997135 662305 997305
rect 662305 997135 662315 997305
rect 662915 997237 663133 997245
rect 662915 997203 663133 997237
rect 662915 997193 663133 997203
rect 663459 997135 663467 997305
rect 663467 997135 663501 997305
rect 663501 997135 663511 997305
rect 664111 997237 664329 997245
rect 664111 997203 664329 997237
rect 664111 997193 664329 997203
rect 664655 997135 664663 997305
rect 664663 997135 664697 997305
rect 664697 997135 664707 997305
rect 665307 997237 665525 997245
rect 665307 997203 665525 997237
rect 665307 997193 665525 997203
rect 665851 997135 665859 997305
rect 665859 997135 665893 997305
rect 665893 997135 665903 997305
rect 666503 997237 666721 997245
rect 666503 997203 666721 997237
rect 666503 997193 666721 997203
rect 167052 996994 167270 997002
rect 167052 996960 167270 996994
rect 167052 996950 167270 996960
rect 167870 996892 167880 997062
rect 167880 996892 167914 997062
rect 167914 996892 167922 997062
rect 168248 996994 168466 997002
rect 168248 996960 168466 996994
rect 168248 996950 168466 996960
rect 169066 996892 169076 997062
rect 169076 996892 169110 997062
rect 169110 996892 169118 997062
rect 169444 996994 169662 997002
rect 169444 996960 169662 996994
rect 169444 996950 169662 996960
rect 170262 996892 170272 997062
rect 170272 996892 170306 997062
rect 170306 996892 170314 997062
rect 418223 996966 418580 997026
rect 664833 996884 665190 996944
rect 169786 996637 170143 996697
rect 416588 996707 416806 996715
rect 416588 996673 416806 996707
rect 416588 996663 416806 996673
rect 417508 996605 417516 996775
rect 417516 996605 417550 996775
rect 417550 996605 417560 996775
rect 661989 996625 662207 996633
rect 661989 996591 662207 996625
rect 661989 996581 662207 996591
rect 662909 996523 662917 996693
rect 662917 996523 662951 996693
rect 662951 996523 662961 996693
rect 663185 996625 663403 996633
rect 663185 996591 663403 996625
rect 663185 996581 663403 996591
rect 664105 996523 664113 996693
rect 664113 996523 664147 996693
rect 664147 996523 664157 996693
rect 664381 996625 664599 996633
rect 664381 996591 664599 996625
rect 664381 996581 664599 996591
rect 665301 996523 665309 996693
rect 665309 996523 665343 996693
rect 665343 996523 665353 996693
rect 665577 996625 665795 996633
rect 665577 996591 665795 996625
rect 665577 996581 665795 996591
rect 666497 996523 666505 996693
rect 666505 996523 666539 996693
rect 666539 996523 666549 996693
rect 167224 996280 167234 996450
rect 167234 996280 167268 996450
rect 167268 996280 167276 996450
rect 167978 996382 168196 996390
rect 167978 996348 168196 996382
rect 167978 996338 168196 996348
rect 168420 996280 168430 996450
rect 168430 996280 168464 996450
rect 168464 996280 168472 996450
rect 169174 996382 169392 996390
rect 169174 996348 169392 996382
rect 169174 996338 169392 996348
rect 169616 996280 169626 996450
rect 169626 996280 169660 996450
rect 169660 996280 169668 996450
rect 417027 996425 417384 996485
rect 170370 996382 170588 996390
rect 170370 996348 170588 996382
rect 170370 996338 170588 996348
rect 663637 996343 663994 996403
rect 168590 996096 168947 996156
rect 418223 995878 418580 995938
rect 664833 995796 665190 995856
rect 169786 995549 170143 995609
rect 41194 891200 41202 891418
rect 41202 891200 41236 891418
rect 41236 891200 41246 891418
rect 169626 995405 169678 995457
rect 170469 995401 170521 995453
rect 42211 891299 42263 891351
rect 169502 995349 169554 995401
rect 416655 995359 416707 995411
rect 170275 995289 170327 995341
rect 417498 995307 417550 995359
rect 662056 995331 662108 995383
rect 662899 995335 662951 995387
rect 416849 995247 416901 995299
rect 417622 995251 417674 995303
rect 662250 995275 662302 995327
rect 663023 995279 663075 995331
rect 40522 891136 40692 891144
rect 40522 891102 40692 891136
rect 40522 891092 40692 891102
rect 42267 891105 42319 891157
rect 40582 890274 40590 890492
rect 40590 890274 40624 890492
rect 40624 890274 40634 890492
rect 41134 890490 41304 890498
rect 41134 890456 41304 890490
rect 41134 890446 41304 890456
rect 42207 890456 42259 890508
rect 41194 890004 41202 890222
rect 41202 890004 41236 890222
rect 41236 890004 41246 890222
rect 40522 889940 40692 889948
rect 40522 889906 40692 889940
rect 40522 889896 40692 889906
rect 40340 889384 40400 889741
rect 41422 889384 41482 889741
rect 40582 889078 40590 889296
rect 40590 889078 40624 889296
rect 40624 889078 40634 889296
rect 41134 889294 41304 889302
rect 41134 889260 41304 889294
rect 41134 889250 41304 889260
rect 41194 888808 41202 889026
rect 41202 888808 41236 889026
rect 41236 888808 41246 889026
rect 40522 888744 40692 888752
rect 40522 888710 40692 888744
rect 40522 888700 40692 888710
rect 40881 888188 40941 888545
rect 41969 888188 42029 888545
rect 40582 887882 40590 888100
rect 40590 887882 40624 888100
rect 40624 887882 40634 888100
rect 41134 888098 41304 888106
rect 41134 888064 41304 888098
rect 41134 888054 41304 888064
rect 41194 887612 41202 887830
rect 41202 887612 41236 887830
rect 41236 887612 41246 887830
rect 40522 887548 40692 887556
rect 40522 887514 40692 887548
rect 40522 887504 40692 887514
rect 40582 886686 40590 886904
rect 40590 886686 40624 886904
rect 40624 886686 40634 886904
rect 41134 886902 41304 886910
rect 41134 886868 41304 886902
rect 41134 886858 41304 886868
rect 41194 886416 41202 886634
rect 41202 886416 41236 886634
rect 41236 886416 41246 886634
rect 40522 886352 40692 886360
rect 40522 886318 40692 886352
rect 40522 886308 40692 886318
rect 40582 885490 40590 885708
rect 40590 885490 40624 885708
rect 40624 885490 40634 885708
rect 41134 885706 41304 885714
rect 41134 885672 41304 885706
rect 41134 885662 41304 885672
rect 41219 609954 41227 610172
rect 41227 609954 41261 610172
rect 41261 609954 41271 610172
rect 42183 610053 42235 610105
rect 42263 890332 42315 890384
rect 168430 995181 168482 995233
rect 169249 995177 169301 995229
rect 42435 890079 42487 890131
rect 168306 995125 168358 995177
rect 169079 995121 169131 995173
rect 663252 995107 663304 995159
rect 664095 995111 664147 995163
rect 663446 995051 663498 995103
rect 664219 995055 664271 995107
rect 42491 889909 42543 889961
rect 40547 609890 40717 609898
rect 40547 609856 40717 609890
rect 40547 609846 40717 609856
rect 42239 609859 42291 609911
rect 42431 889260 42483 889312
rect 40607 609028 40615 609246
rect 40615 609028 40649 609246
rect 40649 609028 40659 609246
rect 41159 609244 41329 609252
rect 41159 609210 41329 609244
rect 41159 609200 41329 609210
rect 42179 609210 42231 609262
rect 41219 608758 41227 608976
rect 41227 608758 41261 608976
rect 41261 608758 41271 608976
rect 40547 608694 40717 608702
rect 40547 608660 40717 608694
rect 40547 608650 40717 608660
rect 40607 607832 40615 608050
rect 40615 607832 40649 608050
rect 40649 607832 40659 608050
rect 41159 608048 41329 608056
rect 41159 608014 41329 608048
rect 41159 608004 41329 608014
rect 41219 607562 41227 607780
rect 41227 607562 41261 607780
rect 41261 607562 41271 607780
rect 40547 607498 40717 607506
rect 40547 607464 40717 607498
rect 40547 607454 40717 607464
rect 40607 606636 40615 606854
rect 40615 606636 40649 606854
rect 40649 606636 40659 606854
rect 41159 606852 41329 606860
rect 41159 606818 41329 606852
rect 41159 606808 41329 606818
rect 41219 606366 41227 606584
rect 41227 606366 41261 606584
rect 41261 606366 41271 606584
rect 40547 606302 40717 606310
rect 40547 606268 40717 606302
rect 40547 606258 40717 606268
rect 40607 605440 40615 605658
rect 40615 605440 40649 605658
rect 40649 605440 40659 605658
rect 41159 605656 41329 605664
rect 41159 605622 41329 605656
rect 41159 605612 41329 605622
rect 41219 605170 41227 605388
rect 41227 605170 41261 605388
rect 41261 605170 41271 605388
rect 40547 605106 40717 605114
rect 40547 605072 40717 605106
rect 40547 605062 40717 605072
rect 40371 604610 40431 604967
rect 41453 604610 41513 604967
rect 40607 604244 40615 604462
rect 40615 604244 40649 604462
rect 40649 604244 40659 604462
rect 41159 604460 41329 604468
rect 41159 604426 41329 604460
rect 41159 604416 41329 604426
rect 41219 603974 41227 604192
rect 41227 603974 41261 604192
rect 41261 603974 41271 604192
rect 40547 603910 40717 603918
rect 40547 603876 40717 603910
rect 40547 603866 40717 603876
rect 40912 603414 40972 603771
rect 42000 603414 42060 603771
rect 40607 603048 40615 603266
rect 40615 603048 40649 603266
rect 40649 603048 40659 603266
rect 41159 603264 41329 603272
rect 41159 603230 41329 603264
rect 41159 603220 41329 603230
rect 41219 602778 41227 602996
rect 41227 602778 41261 602996
rect 41261 602778 41271 602996
rect 40547 602714 40717 602722
rect 40547 602680 40717 602714
rect 40547 602670 40717 602680
rect 40607 601852 40615 602070
rect 40615 601852 40649 602070
rect 40649 601852 40659 602070
rect 41159 602068 41329 602076
rect 41159 602034 41329 602068
rect 41159 602024 41329 602034
rect 41219 601582 41227 601800
rect 41227 601582 41261 601800
rect 41261 601582 41271 601800
rect 40547 601518 40717 601526
rect 40547 601484 40717 601518
rect 40547 601474 40717 601484
rect 40607 600656 40615 600874
rect 40615 600656 40649 600874
rect 40649 600656 40659 600874
rect 41159 600872 41329 600880
rect 41159 600838 41329 600872
rect 41159 600828 41329 600838
rect 41219 600386 41227 600604
rect 41227 600386 41261 600604
rect 41261 600386 41271 600604
rect 40547 600322 40717 600330
rect 40547 600288 40717 600322
rect 40547 600278 40717 600288
rect 40607 599460 40615 599678
rect 40615 599460 40649 599678
rect 40649 599460 40659 599678
rect 41159 599676 41329 599684
rect 41159 599642 41329 599676
rect 41159 599632 41329 599642
rect 41219 599190 41227 599408
rect 41227 599190 41261 599408
rect 41261 599190 41271 599408
rect 40547 599126 40717 599134
rect 40547 599092 40717 599126
rect 40547 599082 40717 599092
rect 40607 598264 40615 598482
rect 40615 598264 40649 598482
rect 40649 598264 40659 598482
rect 41159 598480 41329 598488
rect 41159 598446 41329 598480
rect 41159 598436 41329 598446
rect 41219 597994 41227 598212
rect 41227 597994 41261 598212
rect 41261 597994 41271 598212
rect 40547 597930 40717 597938
rect 40547 597896 40717 597930
rect 40547 597886 40717 597896
rect 40607 597068 40615 597286
rect 40615 597068 40649 597286
rect 40649 597068 40659 597286
rect 41159 597284 41329 597292
rect 41159 597250 41329 597284
rect 41159 597240 41329 597250
rect 41241 352373 41249 352591
rect 41249 352373 41283 352591
rect 41283 352373 41293 352591
rect 42155 352472 42207 352524
rect 42235 609086 42287 609138
rect 42407 608833 42459 608885
rect 42487 889136 42539 889188
rect 167234 994957 167286 995009
rect 168077 994953 168129 995005
rect 42659 888907 42711 888959
rect 167110 994901 167162 994953
rect 167883 994897 167935 994949
rect 664448 994883 664500 994935
rect 665291 994887 665343 994939
rect 664642 994827 664694 994879
rect 665415 994831 665467 994883
rect 665644 994659 665696 994711
rect 666487 994663 666539 994715
rect 665838 994603 665890 994655
rect 666611 994607 666663 994659
rect 42715 888713 42767 888765
rect 42463 608663 42515 608715
rect 42655 888064 42707 888116
rect 40569 352309 40739 352317
rect 40569 352275 40739 352309
rect 40569 352265 40739 352275
rect 42211 352278 42263 352330
rect 42403 608014 42455 608066
rect 40629 351447 40637 351665
rect 40637 351447 40671 351665
rect 40671 351447 40681 351665
rect 41181 351663 41351 351671
rect 41181 351629 41351 351663
rect 41181 351619 41351 351629
rect 42151 351629 42203 351681
rect 41241 351177 41249 351395
rect 41249 351177 41283 351395
rect 41283 351177 41293 351395
rect 40569 351113 40739 351121
rect 40569 351079 40739 351113
rect 40569 351069 40739 351079
rect 40629 350251 40637 350469
rect 40637 350251 40671 350469
rect 40671 350251 40681 350469
rect 41171 350467 41341 350475
rect 41171 350433 41341 350467
rect 41171 350423 41341 350433
rect 41241 349981 41249 350199
rect 41249 349981 41283 350199
rect 41283 349981 41293 350199
rect 40569 349917 40739 349925
rect 40569 349883 40739 349917
rect 40569 349873 40739 349883
rect 40629 349055 40637 349273
rect 40637 349055 40671 349273
rect 40671 349055 40681 349273
rect 41181 349271 41351 349279
rect 41181 349237 41351 349271
rect 41181 349227 41351 349237
rect 41241 348785 41249 349003
rect 41249 348785 41283 349003
rect 41283 348785 41293 349003
rect 40569 348721 40739 348729
rect 40569 348687 40739 348721
rect 40569 348677 40739 348687
rect 40629 347859 40637 348077
rect 40637 347859 40671 348077
rect 40671 347859 40681 348077
rect 41181 348075 41351 348083
rect 41181 348041 41351 348075
rect 41181 348031 41351 348041
rect 41241 347589 41249 347807
rect 41249 347589 41283 347807
rect 41283 347589 41293 347807
rect 40569 347525 40739 347533
rect 40569 347491 40739 347525
rect 40569 347481 40739 347491
rect 40390 346959 40450 347316
rect 41472 346959 41532 347316
rect 40629 346663 40637 346881
rect 40637 346663 40671 346881
rect 40671 346663 40681 346881
rect 41181 346879 41351 346887
rect 41181 346845 41351 346879
rect 41181 346835 41351 346845
rect 41241 346393 41249 346611
rect 41249 346393 41283 346611
rect 41283 346393 41293 346611
rect 40569 346329 40739 346337
rect 40569 346295 40739 346329
rect 40569 346285 40739 346295
rect 40931 345763 40991 346120
rect 42019 345763 42079 346120
rect 40629 345467 40637 345685
rect 40637 345467 40671 345685
rect 40671 345467 40681 345685
rect 41181 345683 41351 345691
rect 41181 345649 41351 345683
rect 41181 345639 41351 345649
rect 41241 345197 41249 345415
rect 41249 345197 41283 345415
rect 41283 345197 41293 345415
rect 40569 345133 40739 345141
rect 40569 345099 40739 345133
rect 40569 345089 40739 345099
rect 40629 344271 40637 344489
rect 40637 344271 40671 344489
rect 40671 344271 40681 344489
rect 41181 344487 41351 344495
rect 41181 344453 41351 344487
rect 41181 344443 41351 344453
rect 41241 344001 41249 344219
rect 41249 344001 41283 344219
rect 41283 344001 41293 344219
rect 40569 343937 40739 343945
rect 40569 343903 40739 343937
rect 40569 343893 40739 343903
rect 40629 343161 40637 343293
rect 40637 343161 40671 343293
rect 40671 343161 40681 343293
rect 41181 343291 41351 343299
rect 41181 343257 41351 343291
rect 41181 343247 41351 343257
rect 40629 343075 40637 343133
rect 40637 343075 40671 343133
rect 40671 343075 40681 343133
rect 41241 342805 41249 343023
rect 41249 342805 41283 343023
rect 41283 342805 41293 343023
rect 40569 342741 40739 342749
rect 40569 342707 40739 342741
rect 40569 342697 40739 342707
rect 40629 341879 40637 342097
rect 40637 341879 40671 342097
rect 40671 341879 40681 342097
rect 41181 342095 41351 342103
rect 41181 342061 41351 342095
rect 41181 342051 41351 342061
rect 41241 341609 41249 341827
rect 41249 341609 41283 341827
rect 41283 341609 41293 341827
rect 40569 341545 40739 341553
rect 40569 341511 40739 341545
rect 40569 341501 40739 341511
rect 40629 340683 40637 340901
rect 40637 340683 40671 340901
rect 40671 340683 40681 340901
rect 41181 340899 41351 340907
rect 41181 340865 41351 340899
rect 41181 340855 41351 340865
rect 41241 340413 41249 340631
rect 41249 340413 41283 340631
rect 41283 340413 41293 340631
rect 40569 340349 40739 340357
rect 40569 340315 40739 340349
rect 40569 340305 40739 340315
rect 40629 339487 40637 339705
rect 40637 339487 40671 339705
rect 40671 339487 40681 339705
rect 41181 339703 41351 339711
rect 41181 339669 41351 339703
rect 41181 339659 41351 339669
rect 41241 339217 41249 339435
rect 41249 339217 41283 339435
rect 41283 339217 41293 339435
rect 40569 339153 40739 339161
rect 40569 339119 40739 339153
rect 40569 339109 40739 339119
rect 40629 338291 40637 338509
rect 40637 338291 40671 338509
rect 40671 338291 40681 338509
rect 41181 338507 41351 338515
rect 41181 338473 41351 338507
rect 41181 338463 41351 338473
rect 41241 338021 41249 338239
rect 41249 338021 41283 338239
rect 41283 338021 41293 338239
rect 40569 337957 40739 337965
rect 40569 337923 40739 337957
rect 40569 337913 40739 337923
rect 40629 337095 40637 337313
rect 40637 337095 40671 337313
rect 40671 337095 40681 337313
rect 41181 337311 41351 337319
rect 41181 337277 41351 337311
rect 41181 337267 41351 337277
rect 41241 336825 41249 337043
rect 41249 336825 41283 337043
rect 41283 336825 41293 337043
rect 40569 336761 40739 336769
rect 40569 336727 40739 336761
rect 40569 336717 40739 336727
rect 40629 335899 40637 336117
rect 40637 335899 40671 336117
rect 40671 335899 40681 336117
rect 41181 336115 41351 336123
rect 41181 336081 41351 336115
rect 41181 336071 41351 336081
rect 41241 335629 41249 335847
rect 41249 335629 41283 335847
rect 41283 335629 41293 335847
rect 40569 335565 40739 335573
rect 40569 335531 40739 335565
rect 40569 335521 40739 335531
rect 40629 334703 40637 334921
rect 40637 334703 40671 334921
rect 40671 334703 40681 334921
rect 41181 334919 41351 334927
rect 41181 334885 41351 334919
rect 41181 334875 41351 334885
rect 42207 351505 42259 351557
rect 42379 351252 42431 351304
rect 42459 607890 42511 607942
rect 42631 607661 42683 607713
rect 42711 887940 42763 887992
rect 42883 887687 42935 887739
rect 42939 887517 42991 887569
rect 42687 607467 42739 607519
rect 42879 886868 42931 886920
rect 42435 351082 42487 351134
rect 42627 606818 42679 606870
rect 42375 350433 42427 350485
rect 42431 350309 42483 350361
rect 42603 350080 42655 350132
rect 42683 606694 42735 606746
rect 42855 606441 42907 606493
rect 42935 886744 42987 886796
rect 43107 886515 43159 886567
rect 43163 886321 43215 886373
rect 42911 606271 42963 606323
rect 43103 885672 43155 885724
rect 42659 349886 42711 349938
rect 42851 605622 42903 605674
rect 42599 349237 42651 349289
rect 42655 349113 42707 349165
rect 42827 348860 42879 348912
rect 42907 605498 42959 605550
rect 43079 605269 43131 605321
rect 43159 885548 43211 885600
rect 675304 727515 675356 727567
rect 676328 727440 676338 727658
rect 676338 727440 676372 727658
rect 676372 727440 676380 727658
rect 675248 727345 675300 727397
rect 676882 727376 677052 727384
rect 676882 727342 677052 727376
rect 676882 727332 677052 727342
rect 675308 726696 675360 726748
rect 675252 726572 675304 726624
rect 675052 726343 675104 726395
rect 674996 726149 675048 726201
rect 675056 725500 675108 725552
rect 675000 725376 675052 725428
rect 674828 725147 674880 725199
rect 674772 724953 674824 725005
rect 674832 724304 674884 724356
rect 674776 724180 674828 724232
rect 674604 723951 674656 724003
rect 674548 723757 674600 723809
rect 674608 723108 674660 723160
rect 674552 722984 674604 723036
rect 674380 722755 674432 722807
rect 674324 722561 674376 722613
rect 674384 721912 674436 721964
rect 674328 721788 674380 721840
rect 674156 721559 674208 721611
rect 674100 721365 674152 721417
rect 674160 720716 674212 720768
rect 674104 720592 674156 720644
rect 43135 605075 43187 605127
rect 42883 348690 42935 348742
rect 43075 604426 43127 604478
rect 42823 348041 42875 348093
rect 42879 347917 42931 347969
rect 43051 347688 43103 347740
rect 43131 604302 43183 604354
rect 43303 604073 43355 604125
rect 43359 603879 43411 603931
rect 43107 347494 43159 347546
rect 43299 603230 43351 603282
rect 43047 346845 43099 346897
rect 43103 346721 43155 346773
rect 43275 346492 43327 346544
rect 43355 603106 43407 603158
rect 43527 602877 43579 602929
rect 43583 602683 43635 602735
rect 43331 346298 43383 346350
rect 43523 602034 43575 602086
rect 43271 345649 43323 345701
rect 43327 345525 43379 345577
rect 43499 345296 43551 345348
rect 43579 601910 43631 601962
rect 43751 601681 43803 601733
rect 43807 601487 43859 601539
rect 43555 345102 43607 345154
rect 43747 600838 43799 600890
rect 43495 344453 43547 344505
rect 43551 344329 43603 344381
rect 43723 344100 43775 344152
rect 43803 600714 43855 600766
rect 43975 600485 44027 600537
rect 44031 600291 44083 600343
rect 43779 343906 43831 343958
rect 43971 599642 44023 599694
rect 43719 343257 43771 343309
rect 43775 343133 43827 343185
rect 43947 342904 43999 342956
rect 44027 599518 44079 599570
rect 44199 599289 44251 599341
rect 44255 599095 44307 599147
rect 44003 342710 44055 342762
rect 44195 598446 44247 598498
rect 43943 342061 43995 342113
rect 43999 341937 44051 341989
rect 44171 341708 44223 341760
rect 44251 598322 44303 598374
rect 44423 598093 44475 598145
rect 44479 597899 44531 597951
rect 44227 341514 44279 341566
rect 44419 597250 44471 597302
rect 44167 340865 44219 340917
rect 44223 340741 44275 340793
rect 44395 340512 44447 340564
rect 44475 597126 44527 597178
rect 676270 726730 676440 726738
rect 676270 726696 676440 726730
rect 676270 726686 676440 726696
rect 676940 726514 676950 726732
rect 676950 726514 676984 726732
rect 676984 726514 676992 726732
rect 676328 726244 676338 726462
rect 676338 726244 676372 726462
rect 676372 726244 676380 726462
rect 676882 726180 677052 726188
rect 676882 726146 677052 726180
rect 676882 726136 677052 726146
rect 676270 725534 676440 725542
rect 676270 725500 676440 725534
rect 676270 725490 676440 725500
rect 676940 725318 676950 725536
rect 676950 725318 676984 725536
rect 676984 725318 676992 725536
rect 676328 725048 676338 725266
rect 676338 725048 676372 725266
rect 676372 725048 676380 725266
rect 676882 724984 677052 724992
rect 676882 724950 677052 724984
rect 676882 724940 677052 724950
rect 676093 724496 676153 724853
rect 677175 724496 677235 724853
rect 676270 724338 676440 724346
rect 676270 724304 676440 724338
rect 676270 724294 676440 724304
rect 676940 724122 676950 724340
rect 676950 724122 676984 724340
rect 676984 724122 676992 724340
rect 676328 723852 676338 724070
rect 676338 723852 676372 724070
rect 676372 723852 676380 724070
rect 676882 723788 677052 723796
rect 676882 723754 677052 723788
rect 676882 723744 677052 723754
rect 675546 723300 675606 723657
rect 676634 723300 676694 723657
rect 676270 723142 676440 723150
rect 676270 723108 676440 723142
rect 676270 723098 676440 723108
rect 676940 722926 676950 723144
rect 676950 722926 676984 723144
rect 676984 722926 676992 723144
rect 676328 722656 676338 722874
rect 676338 722656 676372 722874
rect 676372 722656 676380 722874
rect 676882 722592 677052 722600
rect 676882 722558 677052 722592
rect 676882 722548 677052 722558
rect 676270 721946 676440 721954
rect 676270 721912 676440 721946
rect 676270 721902 676440 721912
rect 676940 721730 676950 721948
rect 676950 721730 676984 721948
rect 676984 721730 676992 721948
rect 676328 721460 676338 721678
rect 676338 721460 676372 721678
rect 676372 721460 676380 721678
rect 676882 721396 677052 721404
rect 676882 721362 677052 721396
rect 676882 721352 677052 721362
rect 676270 720750 676440 720758
rect 676270 720716 676440 720750
rect 676270 720706 676440 720716
rect 676940 720534 676950 720752
rect 676950 720534 676984 720752
rect 676984 720534 676992 720752
rect 675332 453515 675384 453567
rect 676328 453416 676338 453634
rect 676338 453416 676372 453634
rect 676372 453416 676380 453634
rect 675276 453321 675328 453373
rect 676882 453352 677052 453360
rect 676882 453318 677052 453352
rect 676882 453308 677052 453318
rect 675336 452672 675388 452724
rect 675280 452548 675332 452600
rect 675080 452295 675132 452347
rect 675024 452125 675076 452177
rect 675084 451476 675136 451528
rect 675028 451352 675080 451404
rect 674856 451123 674908 451175
rect 674800 450929 674852 450981
rect 674860 450280 674912 450332
rect 674804 450156 674856 450208
rect 674632 449903 674684 449955
rect 674576 449733 674628 449785
rect 674636 449084 674688 449136
rect 674580 448960 674632 449012
rect 674408 448731 674460 448783
rect 674352 448537 674404 448589
rect 674412 447888 674464 447940
rect 674356 447764 674408 447816
rect 674184 447535 674236 447587
rect 674128 447341 674180 447393
rect 674188 446692 674240 446744
rect 674132 446568 674184 446620
rect 673960 446339 674012 446391
rect 673904 446145 673956 446197
rect 673964 445496 674016 445548
rect 673908 445372 673960 445424
rect 673736 445143 673788 445195
rect 673680 444949 673732 445001
rect 673740 444300 673792 444352
rect 673684 444176 673736 444228
rect 673512 443947 673564 443999
rect 673456 443753 673508 443805
rect 673516 443104 673568 443156
rect 673460 442980 673512 443032
rect 673288 442751 673340 442803
rect 673232 442557 673284 442609
rect 673292 441908 673344 441960
rect 673236 441784 673288 441836
rect 673064 441555 673116 441607
rect 673008 441361 673060 441413
rect 673068 440712 673120 440764
rect 673012 440588 673064 440640
rect 672840 440359 672892 440411
rect 672784 440165 672836 440217
rect 672844 439516 672896 439568
rect 672788 439392 672840 439444
rect 44451 340318 44503 340370
rect 44391 339669 44443 339721
rect 44447 339545 44499 339597
rect 44619 339316 44671 339368
rect 44675 339122 44727 339174
rect 44615 338473 44667 338525
rect 44671 338349 44723 338401
rect 44843 338120 44895 338172
rect 44899 337926 44951 337978
rect 44839 337277 44891 337329
rect 44895 337153 44947 337205
rect 45067 336900 45119 336952
rect 45123 336730 45175 336782
rect 45063 336081 45115 336133
rect 45119 335957 45171 336009
rect 45291 335728 45343 335780
rect 45347 335534 45399 335586
rect 45287 334885 45339 334937
rect 45343 334761 45395 334813
rect 676270 452706 676440 452714
rect 676270 452672 676440 452706
rect 676270 452662 676440 452672
rect 676940 452490 676950 452708
rect 676950 452490 676984 452708
rect 676984 452490 676992 452708
rect 676328 452220 676338 452438
rect 676338 452220 676372 452438
rect 676372 452220 676380 452438
rect 676882 452156 677052 452164
rect 676882 452122 677052 452156
rect 676882 452112 677052 452122
rect 676270 451510 676440 451518
rect 676270 451476 676440 451510
rect 676270 451466 676440 451476
rect 676940 451294 676950 451512
rect 676950 451294 676984 451512
rect 676984 451294 676992 451512
rect 676328 451024 676338 451242
rect 676338 451024 676372 451242
rect 676372 451024 676380 451242
rect 676882 450960 677052 450968
rect 676882 450926 677052 450960
rect 676882 450916 677052 450926
rect 676270 450314 676440 450322
rect 676270 450280 676440 450314
rect 676270 450270 676440 450280
rect 676940 450098 676950 450316
rect 676950 450098 676984 450316
rect 676984 450098 676992 450316
rect 676328 449828 676338 450046
rect 676338 449828 676372 450046
rect 676372 449828 676380 450046
rect 676882 449764 677052 449772
rect 676882 449730 677052 449764
rect 676882 449720 677052 449730
rect 676270 449118 676440 449126
rect 676270 449084 676440 449118
rect 676270 449074 676440 449084
rect 676940 448902 676950 449120
rect 676950 448902 676984 449120
rect 676984 448902 676992 449120
rect 676328 448632 676338 448850
rect 676338 448632 676372 448850
rect 676372 448632 676380 448850
rect 676882 448568 677052 448576
rect 676882 448534 677052 448568
rect 676882 448524 677052 448534
rect 676085 448095 676145 448452
rect 677167 448095 677227 448452
rect 676270 447922 676440 447930
rect 676270 447888 676440 447922
rect 676270 447878 676440 447888
rect 676940 447706 676950 447924
rect 676950 447706 676984 447924
rect 676984 447706 676992 447924
rect 676328 447436 676338 447654
rect 676338 447436 676372 447654
rect 676372 447436 676380 447654
rect 676882 447372 677052 447380
rect 676882 447338 677052 447372
rect 676882 447328 677052 447338
rect 675538 446899 675598 447256
rect 676626 446899 676686 447256
rect 676270 446726 676440 446734
rect 676270 446692 676440 446726
rect 676270 446682 676440 446692
rect 676940 446510 676950 446728
rect 676950 446510 676984 446728
rect 676984 446510 676992 446728
rect 676328 446240 676338 446458
rect 676338 446240 676372 446458
rect 676372 446240 676380 446458
rect 676882 446176 677052 446184
rect 676882 446142 677052 446176
rect 676882 446132 677052 446142
rect 676270 445530 676440 445538
rect 676270 445496 676440 445530
rect 676270 445486 676440 445496
rect 676940 445314 676950 445532
rect 676950 445314 676984 445532
rect 676984 445314 676992 445532
rect 676328 445044 676338 445262
rect 676338 445044 676372 445262
rect 676372 445044 676380 445262
rect 676882 444980 677052 444988
rect 676882 444946 677052 444980
rect 676882 444936 677052 444946
rect 676270 444334 676440 444342
rect 676270 444300 676440 444334
rect 676270 444290 676440 444300
rect 676940 444118 676950 444336
rect 676950 444118 676984 444336
rect 676984 444118 676992 444336
rect 676328 443848 676338 444066
rect 676338 443848 676372 444066
rect 676372 443848 676380 444066
rect 676882 443784 677052 443792
rect 676882 443750 677052 443784
rect 676882 443740 677052 443750
rect 676270 443138 676440 443146
rect 676270 443104 676440 443138
rect 676270 443094 676440 443104
rect 676940 442922 676950 443140
rect 676950 442922 676984 443140
rect 676984 442922 676992 443140
rect 676328 442652 676338 442870
rect 676338 442652 676372 442870
rect 676372 442652 676380 442870
rect 676882 442588 677052 442596
rect 676882 442554 677052 442588
rect 676882 442544 677052 442554
rect 676270 441942 676440 441950
rect 676270 441908 676440 441942
rect 676270 441898 676440 441908
rect 676940 441726 676950 441944
rect 676950 441726 676984 441944
rect 676984 441726 676992 441944
rect 676328 441456 676338 441674
rect 676338 441456 676372 441674
rect 676372 441456 676380 441674
rect 676882 441392 677052 441400
rect 676882 441358 677052 441392
rect 676882 441348 677052 441358
rect 676270 440746 676440 440754
rect 676270 440712 676440 440746
rect 676270 440702 676440 440712
rect 676940 440530 676950 440748
rect 676950 440530 676984 440748
rect 676984 440530 676992 440748
rect 676328 440260 676338 440478
rect 676338 440260 676372 440478
rect 676372 440260 676380 440478
rect 676882 440196 677052 440204
rect 676882 440162 677052 440196
rect 676882 440152 677052 440162
rect 676270 439550 676440 439558
rect 676270 439516 676440 439550
rect 676270 439506 676440 439516
rect 676940 439334 676950 439552
rect 676950 439334 676984 439552
rect 676984 439334 676992 439552
rect 134104 47568 134156 47620
rect 134947 47572 134999 47624
rect 135176 47512 135228 47564
rect 135949 47516 136001 47568
rect 135300 47400 135352 47452
rect 136143 47404 136195 47456
rect 136372 47344 136424 47396
rect 137145 47348 137197 47400
rect 136496 47232 136548 47284
rect 137339 47236 137391 47288
rect 137568 47176 137620 47228
rect 138341 47180 138393 47232
rect 137692 47064 137744 47116
rect 138535 47068 138587 47120
rect 138764 47008 138816 47060
rect 139537 47012 139589 47064
rect 138888 46896 138940 46948
rect 139731 46900 139783 46952
rect 139960 46840 140012 46892
rect 140084 46728 140136 46780
rect 429504 47596 429556 47648
rect 430347 47600 430399 47652
rect 430576 47540 430628 47592
rect 431349 47544 431401 47596
rect 430700 47428 430752 47480
rect 431543 47432 431595 47484
rect 431772 47372 431824 47424
rect 432545 47376 432597 47428
rect 431896 47260 431948 47312
rect 432739 47264 432791 47316
rect 432968 47204 433020 47256
rect 433741 47208 433793 47260
rect 433092 47092 433144 47144
rect 433935 47096 433987 47148
rect 434164 47036 434216 47088
rect 434937 47040 434989 47092
rect 434288 46924 434340 46976
rect 435131 46928 435183 46980
rect 435360 46868 435412 46920
rect 436133 46872 436185 46924
rect 140733 46508 140785 46560
rect 435484 46756 435536 46808
rect 436303 46760 436355 46812
rect 140903 46452 140955 46504
rect 436556 46700 436608 46752
rect 437329 46704 437381 46756
rect 141156 46392 141208 46444
rect 141929 46396 141981 46448
rect 436680 46588 436732 46640
rect 437523 46592 437575 46644
rect 141280 46336 141332 46388
rect 142123 46340 142175 46392
rect 437752 46532 437804 46584
rect 438525 46536 438577 46588
rect 142352 46280 142404 46332
rect 143125 46284 143177 46336
rect 437876 46420 437928 46472
rect 438695 46424 438747 46476
rect 142476 46224 142528 46276
rect 143295 46228 143347 46280
rect 438948 46364 439000 46416
rect 439721 46368 439773 46420
rect 143548 46168 143600 46220
rect 144321 46172 144373 46224
rect 439072 46252 439124 46304
rect 439915 46256 439967 46308
rect 143672 46112 143724 46164
rect 144515 46116 144567 46168
rect 440144 46196 440196 46248
rect 440917 46200 440969 46252
rect 144744 46056 144796 46108
rect 145517 46060 145569 46112
rect 440268 46084 440320 46136
rect 441111 46088 441163 46140
rect 144868 46000 144920 46052
rect 145711 46004 145763 46056
rect 441340 46028 441392 46080
rect 442113 46032 442165 46084
rect 145940 45944 145992 45996
rect 146713 45948 146765 46000
rect 146064 45888 146116 45940
rect 146907 45892 146959 45944
rect 441464 45916 441516 45968
rect 442307 45920 442359 45972
rect 147136 45832 147188 45884
rect 147909 45836 147961 45888
rect 442536 45860 442588 45912
rect 443309 45864 443361 45916
rect 147260 45720 147312 45772
rect 148103 45724 148155 45776
rect 442660 45748 442712 45800
rect 443503 45752 443555 45804
rect 148332 45664 148384 45716
rect 149105 45668 149157 45720
rect 443732 45692 443784 45744
rect 444505 45696 444557 45748
rect 148456 45552 148508 45604
rect 149299 45556 149351 45608
rect 443856 45580 443908 45632
rect 444699 45584 444751 45636
rect 149528 45496 149580 45548
rect 150301 45500 150353 45552
rect 444928 45524 444980 45576
rect 445701 45528 445753 45580
rect 149652 45384 149704 45436
rect 150495 45388 150547 45440
rect 445052 45412 445104 45464
rect 445895 45416 445947 45468
rect 150724 45328 150776 45380
rect 151497 45332 151549 45384
rect 446124 45356 446176 45408
rect 446897 45360 446949 45412
rect 150848 45216 150900 45268
rect 151691 45220 151743 45272
rect 446248 45244 446300 45296
rect 447091 45248 447143 45300
rect 151920 45160 151972 45212
rect 152693 45164 152745 45216
rect 447320 45188 447372 45240
rect 448093 45192 448145 45244
rect 152044 45048 152096 45100
rect 152887 45052 152939 45104
rect 447444 45076 447496 45128
rect 448287 45080 448339 45132
rect 153116 44992 153168 45044
rect 153889 44996 153941 45048
rect 448516 45020 448568 45072
rect 449289 45024 449341 45076
rect 153240 44880 153292 44932
rect 154083 44884 154135 44936
rect 448640 44908 448692 44960
rect 449483 44912 449535 44964
rect 154312 44824 154364 44876
rect 155085 44828 155137 44880
rect 449712 44852 449764 44904
rect 450485 44856 450537 44908
rect 154436 44712 154488 44764
rect 155255 44716 155307 44768
rect 449836 44740 449888 44792
rect 450655 44744 450707 44796
rect 155508 44656 155560 44708
rect 156281 44660 156333 44712
rect 450908 44684 450960 44736
rect 451681 44688 451733 44740
rect 155632 44544 155684 44596
rect 156475 44548 156527 44600
rect 451032 44572 451084 44624
rect 451875 44576 451927 44628
rect 156704 44488 156756 44540
rect 157477 44492 157529 44544
rect 452104 44516 452156 44568
rect 452877 44520 452929 44572
rect 156828 44376 156880 44428
rect 157647 44380 157699 44432
rect 452228 44404 452280 44456
rect 453047 44408 453099 44460
rect 157900 44264 157952 44316
rect 158673 44268 158725 44320
rect 453300 44292 453352 44344
rect 454073 44296 454125 44348
rect 158024 44152 158076 44204
rect 158867 44156 158919 44208
rect 453424 44180 453476 44232
rect 454267 44184 454319 44236
rect 146199 43944 146556 44004
rect 440430 43937 440787 43997
rect 147395 43397 147752 43457
rect 441626 43390 441983 43450
rect 134094 43102 134104 43272
rect 134104 43102 134138 43272
rect 134138 43102 134146 43272
rect 134848 43204 135066 43214
rect 134848 43170 135066 43204
rect 134848 43162 135066 43170
rect 135290 43102 135300 43272
rect 135300 43102 135334 43272
rect 135334 43102 135342 43272
rect 136044 43204 136262 43214
rect 136044 43170 136262 43204
rect 136044 43162 136262 43170
rect 136486 43102 136496 43272
rect 136496 43102 136530 43272
rect 136530 43102 136538 43272
rect 137240 43204 137458 43214
rect 137240 43170 137458 43204
rect 137240 43162 137458 43170
rect 137682 43102 137692 43272
rect 137692 43102 137726 43272
rect 137726 43102 137734 43272
rect 138436 43204 138654 43214
rect 138436 43170 138654 43204
rect 138436 43162 138654 43170
rect 138878 43102 138888 43272
rect 138888 43102 138922 43272
rect 138922 43102 138930 43272
rect 139632 43204 139850 43214
rect 139632 43170 139850 43204
rect 139632 43162 139850 43170
rect 140074 43102 140084 43272
rect 140084 43102 140118 43272
rect 140118 43102 140126 43272
rect 140828 43204 141046 43214
rect 140828 43170 141046 43204
rect 140828 43162 141046 43170
rect 141270 43102 141280 43272
rect 141280 43102 141314 43272
rect 141314 43102 141322 43272
rect 142024 43204 142242 43214
rect 142024 43170 142242 43204
rect 142024 43162 142242 43170
rect 142466 43102 142476 43272
rect 142476 43102 142510 43272
rect 142510 43102 142518 43272
rect 143220 43204 143438 43214
rect 143220 43170 143438 43204
rect 143220 43162 143438 43170
rect 143662 43102 143672 43272
rect 143672 43102 143706 43272
rect 143706 43102 143714 43272
rect 144416 43204 144634 43214
rect 144416 43170 144634 43204
rect 144416 43162 144634 43170
rect 144858 43102 144868 43272
rect 144868 43102 144902 43272
rect 144902 43102 144910 43272
rect 145612 43204 145830 43214
rect 145612 43170 145830 43204
rect 145612 43162 145830 43170
rect 146054 43102 146064 43272
rect 146064 43102 146098 43272
rect 146098 43102 146106 43272
rect 146808 43204 147026 43214
rect 146808 43170 147026 43204
rect 146808 43162 147026 43170
rect 147250 43102 147260 43272
rect 147260 43102 147294 43272
rect 147294 43102 147302 43272
rect 148004 43204 148222 43214
rect 148004 43170 148222 43204
rect 148004 43162 148222 43170
rect 148446 43102 148456 43272
rect 148456 43102 148490 43272
rect 148490 43102 148498 43272
rect 149200 43204 149418 43214
rect 149200 43170 149418 43204
rect 149200 43162 149418 43170
rect 149642 43102 149652 43272
rect 149652 43102 149686 43272
rect 149686 43102 149694 43272
rect 150396 43204 150614 43214
rect 150396 43170 150614 43204
rect 150396 43162 150614 43170
rect 150838 43102 150848 43272
rect 150848 43102 150882 43272
rect 150882 43102 150890 43272
rect 151592 43204 151810 43214
rect 151592 43170 151810 43204
rect 151592 43162 151810 43170
rect 152034 43102 152044 43272
rect 152044 43102 152078 43272
rect 152078 43102 152086 43272
rect 152788 43204 153006 43214
rect 152788 43170 153006 43204
rect 152788 43162 153006 43170
rect 153230 43102 153240 43272
rect 153240 43102 153274 43272
rect 153274 43102 153282 43272
rect 153984 43204 154202 43214
rect 153984 43170 154202 43204
rect 153984 43162 154202 43170
rect 154426 43102 154436 43272
rect 154436 43102 154470 43272
rect 154470 43102 154478 43272
rect 155180 43204 155398 43214
rect 155180 43170 155398 43204
rect 155180 43162 155398 43170
rect 155622 43102 155632 43272
rect 155632 43102 155666 43272
rect 155666 43102 155674 43272
rect 156376 43204 156594 43214
rect 156376 43170 156594 43204
rect 156376 43162 156594 43170
rect 156818 43102 156828 43272
rect 156828 43102 156862 43272
rect 156862 43102 156870 43272
rect 157572 43204 157790 43214
rect 157572 43170 157790 43204
rect 157572 43162 157790 43170
rect 158014 43102 158024 43272
rect 158024 43102 158058 43272
rect 158058 43102 158066 43272
rect 158768 43204 158986 43214
rect 158768 43170 158986 43204
rect 158768 43162 158986 43170
rect 429494 43102 429504 43272
rect 429504 43102 429538 43272
rect 429538 43102 429546 43272
rect 430248 43204 430466 43214
rect 430248 43170 430466 43204
rect 430248 43162 430466 43170
rect 430690 43102 430700 43272
rect 430700 43102 430734 43272
rect 430734 43102 430742 43272
rect 431444 43204 431662 43214
rect 431444 43170 431662 43204
rect 431444 43162 431662 43170
rect 431886 43102 431896 43272
rect 431896 43102 431930 43272
rect 431930 43102 431938 43272
rect 432640 43204 432858 43214
rect 432640 43170 432858 43204
rect 432640 43162 432858 43170
rect 433082 43102 433092 43272
rect 433092 43102 433126 43272
rect 433126 43102 433134 43272
rect 433836 43204 434054 43214
rect 433836 43170 434054 43204
rect 433836 43162 434054 43170
rect 434278 43102 434288 43272
rect 434288 43102 434322 43272
rect 434322 43102 434330 43272
rect 435032 43204 435250 43214
rect 435032 43170 435250 43204
rect 435032 43162 435250 43170
rect 435474 43102 435484 43272
rect 435484 43102 435518 43272
rect 435518 43102 435526 43272
rect 436228 43204 436446 43214
rect 436228 43170 436446 43204
rect 436228 43162 436446 43170
rect 436670 43102 436680 43272
rect 436680 43102 436714 43272
rect 436714 43102 436722 43272
rect 437424 43204 437642 43214
rect 437424 43170 437642 43204
rect 437424 43162 437642 43170
rect 437866 43102 437876 43272
rect 437876 43102 437910 43272
rect 437910 43102 437918 43272
rect 438620 43204 438838 43214
rect 438620 43170 438838 43204
rect 438620 43162 438838 43170
rect 439062 43102 439072 43272
rect 439072 43102 439106 43272
rect 439106 43102 439114 43272
rect 439816 43204 440034 43214
rect 439816 43170 440034 43204
rect 439816 43162 440034 43170
rect 440258 43102 440268 43272
rect 440268 43102 440302 43272
rect 440302 43102 440310 43272
rect 441012 43204 441230 43214
rect 441012 43170 441230 43204
rect 441012 43162 441230 43170
rect 441454 43102 441464 43272
rect 441464 43102 441498 43272
rect 441498 43102 441506 43272
rect 442208 43204 442426 43214
rect 442208 43170 442426 43204
rect 442208 43162 442426 43170
rect 442650 43102 442660 43272
rect 442660 43102 442694 43272
rect 442694 43102 442702 43272
rect 443404 43204 443622 43214
rect 443404 43170 443622 43204
rect 443404 43162 443622 43170
rect 443846 43102 443856 43272
rect 443856 43102 443890 43272
rect 443890 43102 443898 43272
rect 444600 43204 444818 43214
rect 444600 43170 444818 43204
rect 444600 43162 444818 43170
rect 445042 43102 445052 43272
rect 445052 43102 445086 43272
rect 445086 43102 445094 43272
rect 445796 43204 446014 43214
rect 445796 43170 446014 43204
rect 445796 43162 446014 43170
rect 446238 43102 446248 43272
rect 446248 43102 446282 43272
rect 446282 43102 446290 43272
rect 446992 43204 447210 43214
rect 446992 43170 447210 43204
rect 446992 43162 447210 43170
rect 447434 43102 447444 43272
rect 447444 43102 447478 43272
rect 447478 43102 447486 43272
rect 448188 43204 448406 43214
rect 448188 43170 448406 43204
rect 448188 43162 448406 43170
rect 448630 43102 448640 43272
rect 448640 43102 448674 43272
rect 448674 43102 448682 43272
rect 449384 43204 449602 43214
rect 449384 43170 449602 43204
rect 449384 43162 449602 43170
rect 449826 43102 449836 43272
rect 449836 43102 449870 43272
rect 449870 43102 449878 43272
rect 450580 43204 450798 43214
rect 450580 43170 450798 43204
rect 450580 43162 450798 43170
rect 451022 43102 451032 43272
rect 451032 43102 451066 43272
rect 451066 43102 451074 43272
rect 451776 43204 451994 43214
rect 451776 43170 451994 43204
rect 451776 43162 451994 43170
rect 452218 43102 452228 43272
rect 452228 43102 452262 43272
rect 452262 43102 452270 43272
rect 452972 43204 453190 43214
rect 452972 43170 453190 43204
rect 452972 43162 453190 43170
rect 453414 43102 453424 43272
rect 453424 43102 453458 43272
rect 453458 43102 453466 43272
rect 454168 43204 454386 43214
rect 454168 43170 454386 43204
rect 454168 43162 454386 43170
rect 146199 42856 146556 42916
rect 440430 42849 440787 42909
rect 135118 42592 135336 42602
rect 135118 42558 135336 42592
rect 135118 42550 135336 42558
rect 135936 42490 135946 42660
rect 135946 42490 135980 42660
rect 135980 42490 135988 42660
rect 136314 42592 136532 42602
rect 136314 42558 136532 42592
rect 136314 42550 136532 42558
rect 137132 42490 137142 42660
rect 137142 42490 137176 42660
rect 137176 42490 137184 42660
rect 137510 42592 137728 42602
rect 137510 42558 137728 42592
rect 137510 42550 137728 42558
rect 138328 42490 138338 42660
rect 138338 42490 138372 42660
rect 138372 42490 138380 42660
rect 138706 42592 138924 42602
rect 138706 42558 138924 42592
rect 138706 42550 138924 42558
rect 139524 42490 139534 42660
rect 139534 42490 139568 42660
rect 139568 42490 139576 42660
rect 139902 42592 140120 42602
rect 139902 42558 140120 42592
rect 139902 42550 140120 42558
rect 140720 42490 140730 42660
rect 140730 42490 140764 42660
rect 140764 42490 140772 42660
rect 141098 42592 141316 42602
rect 141098 42558 141316 42592
rect 141098 42550 141316 42558
rect 141916 42490 141926 42660
rect 141926 42490 141960 42660
rect 141960 42490 141968 42660
rect 142294 42592 142512 42602
rect 142294 42558 142512 42592
rect 142294 42550 142512 42558
rect 143112 42490 143122 42660
rect 143122 42490 143156 42660
rect 143156 42490 143164 42660
rect 143490 42592 143708 42602
rect 143490 42558 143708 42592
rect 143490 42550 143708 42558
rect 144308 42490 144318 42660
rect 144318 42490 144352 42660
rect 144352 42490 144360 42660
rect 144686 42592 144904 42602
rect 144686 42558 144904 42592
rect 144686 42550 144904 42558
rect 145504 42490 145514 42660
rect 145514 42490 145548 42660
rect 145548 42490 145556 42660
rect 145882 42592 146100 42602
rect 145882 42558 146100 42592
rect 145882 42550 146100 42558
rect 146700 42490 146710 42660
rect 146710 42490 146744 42660
rect 146744 42490 146752 42660
rect 147078 42592 147296 42602
rect 147078 42558 147296 42592
rect 147078 42550 147296 42558
rect 147896 42490 147906 42660
rect 147906 42490 147940 42660
rect 147940 42490 147948 42660
rect 148274 42592 148492 42602
rect 148274 42558 148492 42592
rect 148274 42550 148492 42558
rect 149092 42490 149102 42660
rect 149102 42490 149136 42660
rect 149136 42490 149144 42660
rect 149470 42592 149688 42602
rect 149470 42558 149688 42592
rect 149470 42550 149688 42558
rect 150288 42490 150298 42660
rect 150298 42490 150332 42660
rect 150332 42490 150340 42660
rect 150666 42592 150884 42602
rect 150666 42558 150884 42592
rect 150666 42550 150884 42558
rect 151484 42490 151494 42660
rect 151494 42490 151528 42660
rect 151528 42490 151536 42660
rect 151862 42592 152080 42602
rect 151862 42558 152080 42592
rect 151862 42550 152080 42558
rect 152680 42490 152690 42660
rect 152690 42490 152724 42660
rect 152724 42490 152732 42660
rect 153058 42592 153276 42602
rect 153058 42558 153276 42592
rect 153058 42550 153276 42558
rect 153876 42490 153886 42660
rect 153886 42490 153920 42660
rect 153920 42490 153928 42660
rect 154254 42592 154472 42602
rect 154254 42558 154472 42592
rect 154254 42550 154472 42558
rect 155072 42490 155082 42660
rect 155082 42490 155116 42660
rect 155116 42490 155124 42660
rect 155450 42592 155668 42602
rect 155450 42558 155668 42592
rect 155450 42550 155668 42558
rect 156268 42490 156278 42660
rect 156278 42490 156312 42660
rect 156312 42490 156320 42660
rect 156646 42592 156864 42602
rect 156646 42558 156864 42592
rect 156646 42550 156864 42558
rect 157464 42490 157474 42660
rect 157474 42490 157508 42660
rect 157508 42490 157516 42660
rect 158016 42490 158024 42660
rect 158024 42490 158058 42660
rect 158058 42490 158068 42660
rect 158668 42592 158886 42602
rect 158668 42558 158886 42592
rect 158668 42550 158886 42558
rect 430518 42592 430736 42602
rect 430518 42558 430736 42592
rect 430518 42550 430736 42558
rect 431336 42490 431346 42660
rect 431346 42490 431380 42660
rect 431380 42490 431388 42660
rect 431714 42592 431932 42602
rect 431714 42558 431932 42592
rect 431714 42550 431932 42558
rect 432532 42490 432542 42660
rect 432542 42490 432576 42660
rect 432576 42490 432584 42660
rect 432910 42592 433128 42602
rect 432910 42558 433128 42592
rect 432910 42550 433128 42558
rect 433728 42490 433738 42660
rect 433738 42490 433772 42660
rect 433772 42490 433780 42660
rect 434106 42592 434324 42602
rect 434106 42558 434324 42592
rect 434106 42550 434324 42558
rect 434924 42490 434934 42660
rect 434934 42490 434968 42660
rect 434968 42490 434976 42660
rect 435302 42592 435520 42602
rect 435302 42558 435520 42592
rect 435302 42550 435520 42558
rect 436120 42490 436130 42660
rect 436130 42490 436164 42660
rect 436164 42490 436172 42660
rect 436498 42592 436716 42602
rect 436498 42558 436716 42592
rect 436498 42550 436716 42558
rect 437316 42490 437326 42660
rect 437326 42490 437360 42660
rect 437360 42490 437368 42660
rect 437694 42592 437912 42602
rect 437694 42558 437912 42592
rect 437694 42550 437912 42558
rect 438512 42490 438522 42660
rect 438522 42490 438556 42660
rect 438556 42490 438564 42660
rect 438890 42592 439108 42602
rect 438890 42558 439108 42592
rect 438890 42550 439108 42558
rect 439708 42490 439718 42660
rect 439718 42490 439752 42660
rect 439752 42490 439760 42660
rect 440086 42592 440304 42602
rect 440086 42558 440304 42592
rect 440086 42550 440304 42558
rect 440904 42490 440914 42660
rect 440914 42490 440948 42660
rect 440948 42490 440956 42660
rect 441282 42592 441500 42602
rect 441282 42558 441500 42592
rect 441282 42550 441500 42558
rect 442100 42490 442110 42660
rect 442110 42490 442144 42660
rect 442144 42490 442152 42660
rect 442478 42592 442696 42602
rect 442478 42558 442696 42592
rect 442478 42550 442696 42558
rect 443296 42490 443306 42660
rect 443306 42490 443340 42660
rect 443340 42490 443348 42660
rect 443674 42592 443892 42602
rect 443674 42558 443892 42592
rect 443674 42550 443892 42558
rect 444492 42490 444502 42660
rect 444502 42490 444536 42660
rect 444536 42490 444544 42660
rect 444870 42592 445088 42602
rect 444870 42558 445088 42592
rect 444870 42550 445088 42558
rect 445688 42490 445698 42660
rect 445698 42490 445732 42660
rect 445732 42490 445740 42660
rect 446066 42592 446284 42602
rect 446066 42558 446284 42592
rect 446066 42550 446284 42558
rect 446884 42490 446894 42660
rect 446894 42490 446928 42660
rect 446928 42490 446936 42660
rect 447262 42592 447480 42602
rect 447262 42558 447480 42592
rect 447262 42550 447480 42558
rect 448080 42490 448090 42660
rect 448090 42490 448124 42660
rect 448124 42490 448132 42660
rect 448458 42592 448676 42602
rect 448458 42558 448676 42592
rect 448458 42550 448676 42558
rect 449276 42490 449286 42660
rect 449286 42490 449320 42660
rect 449320 42490 449328 42660
rect 449654 42592 449872 42602
rect 449654 42558 449872 42592
rect 449654 42550 449872 42558
rect 450472 42490 450482 42660
rect 450482 42490 450516 42660
rect 450516 42490 450524 42660
rect 450850 42592 451068 42602
rect 450850 42558 451068 42592
rect 450850 42550 451068 42558
rect 451668 42490 451678 42660
rect 451678 42490 451712 42660
rect 451712 42490 451720 42660
rect 452046 42592 452264 42602
rect 452046 42558 452264 42592
rect 452046 42550 452264 42558
rect 452864 42490 452874 42660
rect 452874 42490 452908 42660
rect 452908 42490 452916 42660
rect 453416 42490 453424 42660
rect 453424 42490 453458 42660
rect 453458 42490 453468 42660
rect 454068 42592 454286 42602
rect 454068 42558 454286 42592
rect 454068 42550 454286 42558
rect 147395 42315 147752 42375
rect 441626 42308 441983 42368
<< metal2 >>
rect 417019 997567 417392 997584
rect 417019 997507 417027 997567
rect 417384 997507 417392 997567
rect 417019 997498 417392 997507
rect 663629 997485 664002 997502
rect 663629 997425 663637 997485
rect 663994 997425 664002 997485
rect 663629 997416 664002 997425
rect 168582 997238 168955 997255
rect 168582 997178 168590 997238
rect 168947 997178 168955 997238
rect 416856 997217 416862 997387
rect 416914 997217 416920 997387
rect 417514 997327 417732 997333
rect 417514 997269 417732 997275
rect 168582 997169 168955 997178
rect 167052 997002 167270 997008
rect 167052 996944 167270 996950
rect 167110 994959 167138 996944
rect 167864 996892 167870 997062
rect 167922 996892 167928 997062
rect 168248 997002 168466 997008
rect 168248 996944 168466 996950
rect 167218 996280 167224 996450
rect 167276 996280 167282 996450
rect 167234 995015 167262 996280
rect 167234 995009 167286 995015
rect 167110 994953 167162 994959
rect 167110 994895 167162 994901
rect 167234 994951 167286 994957
rect 167883 994955 167911 996892
rect 167978 996390 168196 996396
rect 167978 996332 168196 996338
rect 168077 995011 168105 996332
rect 168306 995183 168334 996944
rect 169060 996892 169066 997062
rect 169118 996892 169124 997062
rect 169444 997002 169662 997008
rect 169444 996944 169662 996950
rect 168414 996280 168420 996450
rect 168472 996280 168478 996450
rect 168430 995239 168458 996280
rect 168582 996156 168955 996170
rect 168582 996096 168590 996156
rect 168947 996096 168955 996156
rect 168582 996084 168955 996096
rect 168430 995233 168482 995239
rect 168306 995177 168358 995183
rect 168306 995119 168358 995125
rect 168430 995175 168482 995181
rect 169079 995179 169107 996892
rect 169174 996390 169392 996396
rect 169174 996332 169392 996338
rect 169273 995235 169301 996332
rect 169249 995229 169301 995235
rect 168077 995005 168129 995011
rect 167110 994880 167138 994895
rect 167234 994880 167262 994951
rect 167883 994949 167935 994955
rect 167883 994891 167935 994897
rect 168077 994947 168129 994953
rect 167883 994880 167911 994891
rect 168077 994880 168105 994947
rect 168306 994880 168334 995119
rect 168430 994880 168458 995175
rect 169079 995173 169131 995179
rect 169249 995171 169301 995177
rect 169079 995115 169131 995121
rect 169079 995055 169107 995115
rect 169273 995055 169301 995171
rect 169502 995407 169530 996944
rect 170256 996892 170262 997062
rect 170314 996892 170320 997062
rect 169778 996697 170151 996709
rect 169778 996637 169786 996697
rect 170143 996637 170151 996697
rect 169778 996623 170151 996637
rect 169610 996280 169616 996450
rect 169668 996280 169674 996450
rect 169626 995463 169654 996280
rect 169778 995609 170151 995621
rect 169778 995549 169786 995609
rect 170143 995549 170151 995609
rect 169778 995535 170151 995549
rect 169626 995457 169678 995463
rect 169502 995401 169554 995407
rect 169502 995343 169554 995349
rect 169626 995399 169678 995405
rect 169502 995055 169530 995343
rect 169626 995055 169654 995399
rect 170275 995347 170303 996892
rect 416588 996715 416806 996721
rect 416588 996657 416806 996663
rect 170370 996390 170588 996396
rect 170370 996332 170588 996338
rect 170469 995459 170497 996332
rect 170469 995453 170521 995459
rect 416679 995417 416707 996657
rect 170469 995395 170521 995401
rect 416655 995411 416707 995417
rect 170275 995341 170327 995347
rect 170275 995283 170327 995289
rect 170275 995098 170303 995283
rect 170469 995098 170497 995395
rect 416655 995353 416707 995359
rect 416679 995213 416707 995353
rect 416873 995305 416901 997217
rect 417502 996605 417508 996775
rect 417560 996605 417566 996775
rect 417019 996485 417392 996499
rect 417019 996425 417027 996485
rect 417384 996425 417392 996485
rect 417019 996413 417392 996425
rect 417522 995365 417550 996605
rect 416849 995299 416901 995305
rect 417498 995359 417550 995365
rect 417646 995309 417674 997269
rect 662257 997135 662263 997305
rect 662315 997135 662321 997305
rect 662915 997245 663133 997251
rect 662915 997187 663133 997193
rect 418215 997026 418588 997038
rect 418215 996966 418223 997026
rect 418580 996966 418588 997026
rect 418215 996952 418588 996966
rect 661989 996633 662207 996639
rect 661989 996575 662207 996581
rect 418215 995938 418588 995950
rect 418215 995878 418223 995938
rect 418580 995878 418588 995938
rect 418215 995864 418588 995878
rect 662080 995389 662108 996575
rect 662056 995383 662108 995389
rect 662274 995333 662302 997135
rect 662903 996523 662909 996693
rect 662961 996523 662967 996693
rect 662923 995393 662951 996523
rect 662056 995325 662108 995331
rect 417498 995301 417550 995307
rect 417522 995286 417550 995301
rect 417622 995303 417674 995309
rect 416849 995241 416901 995247
rect 417622 995245 417674 995251
rect 416873 995213 416901 995241
rect 417646 995213 417674 995245
rect 662080 994569 662108 995325
rect 662250 995327 662302 995333
rect 662899 995387 662951 995393
rect 663047 995337 663075 997187
rect 663453 997135 663459 997305
rect 663511 997135 663517 997305
rect 664111 997245 664329 997251
rect 664111 997187 664329 997193
rect 663185 996633 663403 996639
rect 663185 996575 663403 996581
rect 662899 995329 662951 995335
rect 662250 995269 662302 995275
rect 662274 994569 662302 995269
rect 662923 994569 662951 995329
rect 663023 995331 663075 995337
rect 663023 995273 663075 995279
rect 663047 994569 663075 995273
rect 663276 995165 663304 996575
rect 663252 995159 663304 995165
rect 663470 995109 663498 997135
rect 664099 996523 664105 996693
rect 664157 996523 664163 996693
rect 663629 996403 664002 996417
rect 663629 996343 663637 996403
rect 663994 996343 664002 996403
rect 663629 996331 664002 996343
rect 664119 995169 664147 996523
rect 663252 995101 663304 995107
rect 663276 994569 663304 995101
rect 663446 995103 663498 995109
rect 664095 995163 664147 995169
rect 664243 995113 664271 997187
rect 664649 997135 664655 997305
rect 664707 997135 664713 997305
rect 665307 997245 665525 997251
rect 665307 997187 665525 997193
rect 664381 996633 664599 996639
rect 664381 996575 664599 996581
rect 664095 995105 664147 995111
rect 663446 995045 663498 995051
rect 663470 994569 663498 995045
rect 664119 994569 664147 995105
rect 664219 995107 664271 995113
rect 664219 995049 664271 995055
rect 664243 994569 664271 995049
rect 664472 994941 664500 996575
rect 664448 994935 664500 994941
rect 664666 994885 664694 997135
rect 664825 996944 665198 996956
rect 664825 996884 664833 996944
rect 665190 996884 665198 996944
rect 664825 996870 665198 996884
rect 665295 996523 665301 996693
rect 665353 996523 665359 996693
rect 664825 995856 665198 995868
rect 664825 995796 664833 995856
rect 665190 995796 665198 995856
rect 664825 995782 665198 995796
rect 665315 994945 665343 996523
rect 664448 994877 664500 994883
rect 664472 994569 664500 994877
rect 664642 994879 664694 994885
rect 665291 994939 665343 994945
rect 665439 994889 665467 997187
rect 665845 997135 665851 997305
rect 665903 997135 665909 997305
rect 666503 997245 666721 997251
rect 666503 997187 666721 997193
rect 665577 996633 665795 996639
rect 665577 996575 665795 996581
rect 665291 994881 665343 994887
rect 664642 994821 664694 994827
rect 664666 994569 664694 994821
rect 665315 994569 665343 994881
rect 665415 994883 665467 994889
rect 665415 994825 665467 994831
rect 665439 994569 665467 994825
rect 665668 994717 665696 996575
rect 665644 994711 665696 994717
rect 665862 994661 665890 997135
rect 666491 996523 666497 996693
rect 666549 996523 666555 996693
rect 666511 994721 666539 996523
rect 665644 994653 665696 994659
rect 665668 994569 665696 994653
rect 665838 994655 665890 994661
rect 666487 994715 666539 994721
rect 666635 994665 666663 997187
rect 666487 994657 666539 994663
rect 665838 994597 665890 994603
rect 665862 994569 665890 994597
rect 666511 994569 666539 994657
rect 666611 994659 666663 994665
rect 666611 994601 666663 994607
rect 666635 994569 666663 994601
rect 41188 891200 41194 891418
rect 41246 891327 41252 891418
rect 42205 891327 42211 891351
rect 41246 891299 42211 891327
rect 42263 891327 42269 891351
rect 42263 891299 43227 891327
rect 41246 891200 41252 891299
rect 40522 891144 40692 891150
rect 42261 891133 42267 891157
rect 40692 891105 42267 891133
rect 42319 891133 42325 891157
rect 42319 891105 43227 891133
rect 40522 891086 40692 891092
rect 41134 890498 41304 890504
rect 40576 890274 40582 890492
rect 40634 890360 40640 890492
rect 42201 890484 42207 890508
rect 41304 890456 42207 890484
rect 42259 890484 42265 890508
rect 42259 890456 43227 890484
rect 41134 890440 41304 890446
rect 42257 890360 42263 890384
rect 40634 890332 42263 890360
rect 42315 890360 42321 890384
rect 42315 890332 43227 890360
rect 40634 890274 40640 890332
rect 41188 890004 41194 890222
rect 41246 890131 41252 890222
rect 41246 890103 42435 890131
rect 41246 890004 41252 890103
rect 42429 890079 42435 890103
rect 42487 890103 43227 890131
rect 42487 890079 42493 890103
rect 40522 889948 40692 889954
rect 42485 889937 42491 889961
rect 40692 889909 42491 889937
rect 42543 889937 42549 889961
rect 42543 889909 43227 889937
rect 40522 889890 40692 889896
rect 40323 889741 40409 889749
rect 40323 889384 40340 889741
rect 40400 889384 40409 889741
rect 40323 889376 40409 889384
rect 41408 889741 41494 889749
rect 41408 889384 41422 889741
rect 41482 889384 41494 889741
rect 41408 889376 41494 889384
rect 41134 889302 41304 889308
rect 40576 889078 40582 889296
rect 40634 889164 40640 889296
rect 42425 889288 42431 889312
rect 41304 889260 42431 889288
rect 42483 889288 42489 889312
rect 42483 889260 43227 889288
rect 41134 889244 41304 889250
rect 42481 889164 42487 889188
rect 40634 889136 42487 889164
rect 42539 889164 42545 889188
rect 42539 889136 43227 889164
rect 40634 889078 40640 889136
rect 41188 888808 41194 889026
rect 41246 888935 41252 889026
rect 42653 888935 42659 888959
rect 41246 888907 42659 888935
rect 42711 888935 42717 888959
rect 42711 888907 43227 888935
rect 41246 888808 41252 888907
rect 40522 888752 40692 888758
rect 42709 888741 42715 888765
rect 40692 888713 42715 888741
rect 42767 888741 42773 888765
rect 42767 888713 43227 888741
rect 40522 888694 40692 888700
rect 40869 888545 40955 888553
rect 40869 888188 40881 888545
rect 40941 888188 40955 888545
rect 40869 888180 40955 888188
rect 41957 888545 42043 888553
rect 41957 888188 41969 888545
rect 42029 888188 42043 888545
rect 41957 888180 42043 888188
rect 41134 888106 41304 888112
rect 40576 887882 40582 888100
rect 40634 887968 40640 888100
rect 42649 888092 42655 888116
rect 41304 888064 42655 888092
rect 42707 888092 42713 888116
rect 42707 888064 43227 888092
rect 41134 888048 41304 888054
rect 42705 887968 42711 887992
rect 40634 887940 42711 887968
rect 42763 887968 42769 887992
rect 42763 887940 43227 887968
rect 40634 887882 40640 887940
rect 41188 887612 41194 887830
rect 41246 887739 41252 887830
rect 41246 887711 42883 887739
rect 41246 887612 41252 887711
rect 42877 887687 42883 887711
rect 42935 887711 43227 887739
rect 42935 887687 42941 887711
rect 40522 887556 40692 887562
rect 42933 887545 42939 887569
rect 40692 887517 42939 887545
rect 42991 887545 42997 887569
rect 42991 887517 43227 887545
rect 40522 887498 40692 887504
rect 41134 886910 41304 886916
rect 40576 886686 40582 886904
rect 40634 886772 40640 886904
rect 42873 886896 42879 886920
rect 41304 886868 42879 886896
rect 42931 886896 42937 886920
rect 42931 886868 43227 886896
rect 41134 886852 41304 886858
rect 42929 886772 42935 886796
rect 40634 886744 42935 886772
rect 42987 886772 42993 886796
rect 42987 886744 43227 886772
rect 40634 886686 40640 886744
rect 41188 886416 41194 886634
rect 41246 886543 41252 886634
rect 43101 886543 43107 886567
rect 41246 886515 43107 886543
rect 43159 886543 43165 886567
rect 43159 886515 43227 886543
rect 41246 886416 41252 886515
rect 40522 886360 40692 886366
rect 43157 886349 43163 886373
rect 40692 886321 43163 886349
rect 43215 886349 43221 886373
rect 43215 886321 43227 886349
rect 40522 886302 40692 886308
rect 41134 885714 41304 885720
rect 40576 885490 40582 885708
rect 40634 885576 40640 885708
rect 43097 885700 43103 885724
rect 41304 885672 43103 885700
rect 43155 885700 43161 885724
rect 43155 885672 43227 885700
rect 41134 885656 41304 885662
rect 43153 885576 43159 885600
rect 40634 885548 43159 885576
rect 43211 885576 43217 885600
rect 43211 885548 43227 885576
rect 40634 885490 40640 885548
rect 676322 727567 676328 727658
rect 675230 727539 675304 727567
rect 675298 727515 675304 727539
rect 675356 727539 676328 727567
rect 675356 727515 675362 727539
rect 676322 727440 676328 727539
rect 676380 727440 676386 727658
rect 675242 727373 675248 727397
rect 675230 727345 675248 727373
rect 675300 727373 675306 727397
rect 676882 727384 677052 727390
rect 675300 727345 676882 727373
rect 676882 727326 677052 727332
rect 675302 726724 675308 726748
rect 675253 726696 675308 726724
rect 675360 726724 675366 726748
rect 676270 726738 676440 726744
rect 675360 726696 676270 726724
rect 676270 726680 676440 726686
rect 675246 726572 675252 726624
rect 675304 726600 675310 726624
rect 676934 726600 676940 726732
rect 675304 726572 676940 726600
rect 676934 726514 676940 726572
rect 676992 726514 676998 726732
rect 675046 726371 675052 726395
rect 673842 726343 675052 726371
rect 675104 726371 675110 726395
rect 676322 726371 676328 726462
rect 675104 726343 676328 726371
rect 676322 726244 676328 726343
rect 676380 726244 676386 726462
rect 674990 726177 674996 726201
rect 673842 726149 674996 726177
rect 675048 726177 675054 726201
rect 676882 726188 677052 726194
rect 675048 726149 676882 726177
rect 676882 726130 677052 726136
rect 675050 725528 675056 725552
rect 673842 725500 675056 725528
rect 675108 725528 675114 725552
rect 676270 725542 676440 725548
rect 675108 725500 676270 725528
rect 676270 725484 676440 725490
rect 674994 725404 675000 725428
rect 673842 725376 675000 725404
rect 675052 725404 675058 725428
rect 676934 725404 676940 725536
rect 675052 725376 676940 725404
rect 676934 725318 676940 725376
rect 676992 725318 676998 725536
rect 674822 725175 674828 725199
rect 673842 725147 674828 725175
rect 674880 725175 674886 725199
rect 676322 725175 676328 725266
rect 674880 725147 676328 725175
rect 676322 725048 676328 725147
rect 676380 725048 676386 725266
rect 674766 724981 674772 725005
rect 673842 724953 674772 724981
rect 674824 724981 674830 725005
rect 676882 724992 677052 724998
rect 674824 724953 676882 724981
rect 676882 724934 677052 724940
rect 676081 724853 676167 724861
rect 676081 724496 676093 724853
rect 676153 724496 676167 724853
rect 676081 724488 676167 724496
rect 677166 724853 677252 724861
rect 677166 724496 677175 724853
rect 677235 724496 677252 724853
rect 677166 724488 677252 724496
rect 674826 724332 674832 724356
rect 673842 724304 674832 724332
rect 674884 724332 674890 724356
rect 676270 724346 676440 724352
rect 674884 724304 676270 724332
rect 676270 724288 676440 724294
rect 674770 724208 674776 724232
rect 673842 724180 674776 724208
rect 674828 724208 674834 724232
rect 676934 724208 676940 724340
rect 674828 724180 676940 724208
rect 676934 724122 676940 724180
rect 676992 724122 676998 724340
rect 674598 723979 674604 724003
rect 673842 723951 674604 723979
rect 674656 723979 674662 724003
rect 676322 723979 676328 724070
rect 674656 723951 676328 723979
rect 676322 723852 676328 723951
rect 676380 723852 676386 724070
rect 674542 723785 674548 723809
rect 673842 723757 674548 723785
rect 674600 723785 674606 723809
rect 676882 723796 677052 723802
rect 674600 723757 676882 723785
rect 676882 723738 677052 723744
rect 675532 723657 675618 723665
rect 675532 723300 675546 723657
rect 675606 723300 675618 723657
rect 675532 723292 675618 723300
rect 676620 723657 676706 723665
rect 676620 723300 676634 723657
rect 676694 723300 676706 723657
rect 676620 723292 676706 723300
rect 674602 723136 674608 723160
rect 673842 723108 674608 723136
rect 674660 723136 674666 723160
rect 676270 723150 676440 723156
rect 674660 723108 676270 723136
rect 676270 723092 676440 723098
rect 674546 723012 674552 723036
rect 673842 722984 674552 723012
rect 674604 723012 674610 723036
rect 676934 723012 676940 723144
rect 674604 722984 676940 723012
rect 676934 722926 676940 722984
rect 676992 722926 676998 723144
rect 674374 722783 674380 722807
rect 673842 722755 674380 722783
rect 674432 722783 674438 722807
rect 676322 722783 676328 722874
rect 674432 722755 676328 722783
rect 676322 722656 676328 722755
rect 676380 722656 676386 722874
rect 674318 722589 674324 722613
rect 673842 722561 674324 722589
rect 674376 722589 674382 722613
rect 676882 722600 677052 722606
rect 674376 722561 676882 722589
rect 676882 722542 677052 722548
rect 674378 721940 674384 721964
rect 673842 721912 674384 721940
rect 674436 721940 674442 721964
rect 676270 721954 676440 721960
rect 674436 721912 676270 721940
rect 676270 721896 676440 721902
rect 674322 721816 674328 721840
rect 673842 721788 674328 721816
rect 674380 721816 674386 721840
rect 676934 721816 676940 721948
rect 674380 721788 676940 721816
rect 676934 721730 676940 721788
rect 676992 721730 676998 721948
rect 674150 721587 674156 721611
rect 674066 721559 674156 721587
rect 674208 721587 674214 721611
rect 676322 721587 676328 721678
rect 674208 721559 676328 721587
rect 676322 721460 676328 721559
rect 676380 721460 676386 721678
rect 674094 721393 674100 721417
rect 674066 721365 674100 721393
rect 674152 721393 674158 721417
rect 676882 721404 677052 721410
rect 674152 721365 676882 721393
rect 676882 721346 677052 721352
rect 674154 720744 674160 720768
rect 674066 720716 674160 720744
rect 674212 720744 674218 720768
rect 676270 720758 676440 720764
rect 674212 720716 676270 720744
rect 676270 720700 676440 720706
rect 674098 720620 674104 720644
rect 674066 720592 674104 720620
rect 674156 720620 674162 720644
rect 676934 720620 676940 720752
rect 674156 720592 676940 720620
rect 676934 720534 676940 720592
rect 676992 720534 676998 720752
rect 41213 609954 41219 610172
rect 41271 610081 41277 610172
rect 42177 610081 42183 610105
rect 41271 610053 42183 610081
rect 42235 610081 42241 610105
rect 42235 610053 44320 610081
rect 41271 609954 41277 610053
rect 40547 609898 40717 609904
rect 42233 609887 42239 609911
rect 40717 609859 42239 609887
rect 42291 609887 42297 609911
rect 42291 609859 44320 609887
rect 40547 609840 40717 609846
rect 41159 609252 41329 609258
rect 40601 609028 40607 609246
rect 40659 609114 40665 609246
rect 42173 609238 42179 609262
rect 41329 609210 42179 609238
rect 42231 609238 42237 609262
rect 42231 609210 44320 609238
rect 41159 609194 41329 609200
rect 42229 609114 42235 609138
rect 40659 609086 42235 609114
rect 42287 609114 42293 609138
rect 42287 609086 44320 609114
rect 40659 609028 40665 609086
rect 41213 608758 41219 608976
rect 41271 608885 41277 608976
rect 41271 608857 42407 608885
rect 41271 608758 41277 608857
rect 42401 608833 42407 608857
rect 42459 608857 44320 608885
rect 42459 608833 42465 608857
rect 40547 608702 40717 608708
rect 42457 608691 42463 608715
rect 40717 608663 42463 608691
rect 42515 608691 42521 608715
rect 42515 608663 44320 608691
rect 40547 608644 40717 608650
rect 41159 608056 41329 608062
rect 40601 607832 40607 608050
rect 40659 607918 40665 608050
rect 42397 608042 42403 608066
rect 41329 608014 42403 608042
rect 42455 608042 42461 608066
rect 42455 608014 44320 608042
rect 41159 607998 41329 608004
rect 42453 607918 42459 607942
rect 40659 607890 42459 607918
rect 42511 607918 42517 607942
rect 42511 607890 44320 607918
rect 40659 607832 40665 607890
rect 41213 607562 41219 607780
rect 41271 607689 41277 607780
rect 42625 607689 42631 607713
rect 41271 607661 42631 607689
rect 42683 607689 42689 607713
rect 42683 607661 44320 607689
rect 41271 607562 41277 607661
rect 40547 607506 40717 607512
rect 42681 607495 42687 607519
rect 40717 607467 42687 607495
rect 42739 607495 42745 607519
rect 42739 607467 44320 607495
rect 40547 607448 40717 607454
rect 41159 606860 41329 606866
rect 40601 606636 40607 606854
rect 40659 606722 40665 606854
rect 42621 606846 42627 606870
rect 41329 606818 42627 606846
rect 42679 606846 42685 606870
rect 42679 606818 44320 606846
rect 41159 606802 41329 606808
rect 42677 606722 42683 606746
rect 40659 606694 42683 606722
rect 42735 606722 42741 606746
rect 42735 606694 44320 606722
rect 40659 606636 40665 606694
rect 41213 606366 41219 606584
rect 41271 606493 41277 606584
rect 41271 606465 42855 606493
rect 41271 606366 41277 606465
rect 42849 606441 42855 606465
rect 42907 606465 44320 606493
rect 42907 606441 42913 606465
rect 40547 606310 40717 606316
rect 42905 606299 42911 606323
rect 40717 606271 42911 606299
rect 42963 606299 42969 606323
rect 42963 606271 44320 606299
rect 40547 606252 40717 606258
rect 41159 605664 41329 605670
rect 40601 605440 40607 605658
rect 40659 605526 40665 605658
rect 42845 605650 42851 605674
rect 41329 605622 42851 605650
rect 42903 605650 42909 605674
rect 42903 605622 44320 605650
rect 41159 605606 41329 605612
rect 42901 605526 42907 605550
rect 40659 605498 42907 605526
rect 42959 605526 42965 605550
rect 42959 605498 44320 605526
rect 40659 605440 40665 605498
rect 41213 605170 41219 605388
rect 41271 605297 41277 605388
rect 43073 605297 43079 605321
rect 41271 605269 43079 605297
rect 43131 605297 43137 605321
rect 43131 605269 44320 605297
rect 41271 605170 41277 605269
rect 40547 605114 40717 605120
rect 43129 605103 43135 605127
rect 40717 605075 43135 605103
rect 43187 605103 43193 605127
rect 43187 605075 44320 605103
rect 40547 605056 40717 605062
rect 40354 604967 40440 604975
rect 40354 604610 40371 604967
rect 40431 604610 40440 604967
rect 40354 604602 40440 604610
rect 41439 604967 41525 604975
rect 41439 604610 41453 604967
rect 41513 604610 41525 604967
rect 41439 604602 41525 604610
rect 41159 604468 41329 604474
rect 40601 604244 40607 604462
rect 40659 604330 40665 604462
rect 43069 604454 43075 604478
rect 41329 604426 43075 604454
rect 43127 604454 43133 604478
rect 43127 604426 44320 604454
rect 41159 604410 41329 604416
rect 43125 604330 43131 604354
rect 40659 604302 43131 604330
rect 43183 604330 43189 604354
rect 43183 604302 44320 604330
rect 40659 604244 40665 604302
rect 41213 603974 41219 604192
rect 41271 604101 41277 604192
rect 43297 604101 43303 604125
rect 41271 604073 43303 604101
rect 43355 604101 43361 604125
rect 43355 604073 44320 604101
rect 41271 603974 41277 604073
rect 40547 603918 40717 603924
rect 43353 603907 43359 603931
rect 40717 603879 43359 603907
rect 43411 603907 43417 603931
rect 43411 603879 44320 603907
rect 40547 603860 40717 603866
rect 40900 603771 40986 603779
rect 40900 603414 40912 603771
rect 40972 603414 40986 603771
rect 40900 603406 40986 603414
rect 41988 603771 42074 603779
rect 41988 603414 42000 603771
rect 42060 603414 42074 603771
rect 41988 603406 42074 603414
rect 41159 603272 41329 603278
rect 40601 603048 40607 603266
rect 40659 603134 40665 603266
rect 43293 603258 43299 603282
rect 41329 603230 43299 603258
rect 43351 603258 43357 603282
rect 43351 603230 44320 603258
rect 41159 603214 41329 603220
rect 43349 603134 43355 603158
rect 40659 603106 43355 603134
rect 43407 603134 43413 603158
rect 43407 603106 44320 603134
rect 40659 603048 40665 603106
rect 41213 602778 41219 602996
rect 41271 602905 41277 602996
rect 43521 602905 43527 602929
rect 41271 602877 43527 602905
rect 43579 602905 43585 602929
rect 43579 602877 44320 602905
rect 41271 602778 41277 602877
rect 40547 602722 40717 602728
rect 43577 602711 43583 602735
rect 40717 602683 43583 602711
rect 43635 602711 43641 602735
rect 43635 602683 44320 602711
rect 40547 602664 40717 602670
rect 41159 602076 41329 602082
rect 40601 601852 40607 602070
rect 40659 601938 40665 602070
rect 43517 602062 43523 602086
rect 41329 602034 43523 602062
rect 43575 602062 43581 602086
rect 43575 602034 44320 602062
rect 41159 602018 41329 602024
rect 43573 601938 43579 601962
rect 40659 601910 43579 601938
rect 43631 601938 43637 601962
rect 43631 601910 44320 601938
rect 40659 601852 40665 601910
rect 41213 601582 41219 601800
rect 41271 601709 41277 601800
rect 43745 601709 43751 601733
rect 41271 601681 43751 601709
rect 43803 601709 43809 601733
rect 43803 601681 44320 601709
rect 41271 601582 41277 601681
rect 40547 601526 40717 601532
rect 43801 601515 43807 601539
rect 40717 601487 43807 601515
rect 43859 601515 43865 601539
rect 43859 601487 44320 601515
rect 40547 601468 40717 601474
rect 41159 600880 41329 600886
rect 40601 600656 40607 600874
rect 40659 600742 40665 600874
rect 43741 600866 43747 600890
rect 41329 600838 43747 600866
rect 43799 600866 43805 600890
rect 43799 600838 44320 600866
rect 41159 600822 41329 600828
rect 43797 600742 43803 600766
rect 40659 600714 43803 600742
rect 43855 600742 43861 600766
rect 43855 600714 44320 600742
rect 40659 600656 40665 600714
rect 41213 600386 41219 600604
rect 41271 600513 41277 600604
rect 43969 600513 43975 600537
rect 41271 600485 43975 600513
rect 44027 600513 44033 600537
rect 44027 600485 44320 600513
rect 41271 600386 41277 600485
rect 40547 600330 40717 600336
rect 44025 600319 44031 600343
rect 40717 600291 44031 600319
rect 44083 600319 44089 600343
rect 44083 600291 44320 600319
rect 40547 600272 40717 600278
rect 41159 599684 41329 599690
rect 40601 599460 40607 599678
rect 40659 599546 40665 599678
rect 43965 599670 43971 599694
rect 41329 599642 43971 599670
rect 44023 599670 44029 599694
rect 44023 599642 44320 599670
rect 41159 599626 41329 599632
rect 44021 599546 44027 599570
rect 40659 599518 44027 599546
rect 44079 599546 44085 599570
rect 44079 599518 44320 599546
rect 40659 599460 40665 599518
rect 41213 599190 41219 599408
rect 41271 599317 41277 599408
rect 44193 599317 44199 599341
rect 41271 599289 44199 599317
rect 44251 599317 44257 599341
rect 44251 599289 44321 599317
rect 41271 599190 41277 599289
rect 40547 599134 40717 599140
rect 44249 599123 44255 599147
rect 40717 599095 44255 599123
rect 44307 599123 44313 599147
rect 44307 599095 44321 599123
rect 40547 599076 40717 599082
rect 41159 598488 41329 598494
rect 40601 598264 40607 598482
rect 40659 598350 40665 598482
rect 44189 598474 44195 598498
rect 41329 598446 44195 598474
rect 44247 598474 44253 598498
rect 44247 598446 44335 598474
rect 41159 598430 41329 598436
rect 44245 598350 44251 598374
rect 40659 598322 44251 598350
rect 44303 598350 44309 598374
rect 44303 598322 44335 598350
rect 40659 598264 40665 598322
rect 41213 597994 41219 598212
rect 41271 598121 41277 598212
rect 44417 598121 44423 598145
rect 41271 598093 44423 598121
rect 44475 598121 44481 598145
rect 44475 598093 44544 598121
rect 41271 597994 41277 598093
rect 40547 597938 40717 597944
rect 44473 597927 44479 597951
rect 40717 597899 44479 597927
rect 44531 597927 44537 597951
rect 44531 597899 44544 597927
rect 40547 597880 40717 597886
rect 41159 597292 41329 597298
rect 40601 597068 40607 597286
rect 40659 597154 40665 597286
rect 44413 597278 44419 597302
rect 41329 597250 44419 597278
rect 44471 597278 44477 597302
rect 44471 597250 44544 597278
rect 41159 597234 41329 597240
rect 44469 597154 44475 597178
rect 40659 597126 44475 597154
rect 44527 597154 44533 597178
rect 44527 597126 44544 597154
rect 40659 597068 40665 597126
rect 675326 453543 675332 453567
rect 673198 453515 675332 453543
rect 675384 453543 675390 453567
rect 676322 453543 676328 453634
rect 675384 453515 676328 453543
rect 676322 453416 676328 453515
rect 676380 453416 676386 453634
rect 675270 453349 675276 453373
rect 673198 453321 675276 453349
rect 675328 453349 675334 453373
rect 676882 453360 677052 453366
rect 675328 453321 676882 453349
rect 676882 453302 677052 453308
rect 675330 452700 675336 452724
rect 673198 452672 675336 452700
rect 675388 452700 675394 452724
rect 676270 452714 676440 452720
rect 675388 452672 676270 452700
rect 676270 452656 676440 452662
rect 675274 452576 675280 452600
rect 673198 452548 675149 452576
rect 675208 452548 675280 452576
rect 675332 452576 675338 452600
rect 676934 452576 676940 452708
rect 675332 452548 676940 452576
rect 676934 452490 676940 452548
rect 676992 452490 676998 452708
rect 676322 452347 676328 452438
rect 673198 452319 675080 452347
rect 675074 452295 675080 452319
rect 675132 452319 676328 452347
rect 675132 452295 675138 452319
rect 676322 452220 676328 452319
rect 676380 452220 676386 452438
rect 675018 452153 675024 452177
rect 673198 452125 675024 452153
rect 675076 452153 675082 452177
rect 676882 452164 677052 452170
rect 675076 452125 676882 452153
rect 676882 452106 677052 452112
rect 675078 451504 675084 451528
rect 673198 451476 675084 451504
rect 675136 451504 675142 451528
rect 676270 451518 676440 451524
rect 675136 451476 676270 451504
rect 676270 451460 676440 451466
rect 675022 451380 675028 451404
rect 673198 451352 675028 451380
rect 675080 451380 675086 451404
rect 676934 451380 676940 451512
rect 675080 451352 676940 451380
rect 676934 451294 676940 451352
rect 676992 451294 676998 451512
rect 674850 451151 674856 451175
rect 673198 451123 674856 451151
rect 674908 451151 674914 451175
rect 676322 451151 676328 451242
rect 674908 451123 676328 451151
rect 676322 451024 676328 451123
rect 676380 451024 676386 451242
rect 674794 450957 674800 450981
rect 673198 450929 674800 450957
rect 674852 450957 674858 450981
rect 676882 450968 677052 450974
rect 674852 450929 676882 450957
rect 676882 450910 677052 450916
rect 674854 450308 674860 450332
rect 673198 450280 674860 450308
rect 674912 450308 674918 450332
rect 676270 450322 676440 450328
rect 674912 450280 676270 450308
rect 676270 450264 676440 450270
rect 674798 450184 674804 450208
rect 673198 450156 674804 450184
rect 674856 450184 674862 450208
rect 676934 450184 676940 450316
rect 674856 450156 676940 450184
rect 676934 450098 676940 450156
rect 676992 450098 676998 450316
rect 676322 449955 676328 450046
rect 673198 449927 674632 449955
rect 674626 449903 674632 449927
rect 674684 449927 676328 449955
rect 674684 449903 674690 449927
rect 676322 449828 676328 449927
rect 676380 449828 676386 450046
rect 674570 449761 674576 449785
rect 673198 449733 674576 449761
rect 674628 449761 674634 449785
rect 676882 449772 677052 449778
rect 674628 449733 676882 449761
rect 676882 449714 677052 449720
rect 674630 449112 674636 449136
rect 673198 449084 674636 449112
rect 674688 449112 674694 449136
rect 676270 449126 676440 449132
rect 674688 449084 676270 449112
rect 676270 449068 676440 449074
rect 674574 448988 674580 449012
rect 673198 448960 674580 448988
rect 674632 448988 674638 449012
rect 676934 448988 676940 449120
rect 674632 448960 676940 448988
rect 676934 448902 676940 448960
rect 676992 448902 676998 449120
rect 674402 448759 674408 448783
rect 673198 448731 674408 448759
rect 674460 448759 674466 448783
rect 676322 448759 676328 448850
rect 674460 448731 676328 448759
rect 676322 448632 676328 448731
rect 676380 448632 676386 448850
rect 674346 448565 674352 448589
rect 673198 448537 674352 448565
rect 674404 448565 674410 448589
rect 676882 448576 677052 448582
rect 674404 448537 676882 448565
rect 676882 448518 677052 448524
rect 676073 448452 676159 448460
rect 676073 448095 676085 448452
rect 676145 448095 676159 448452
rect 676073 448087 676159 448095
rect 677158 448452 677244 448460
rect 677158 448095 677167 448452
rect 677227 448095 677244 448452
rect 677158 448087 677244 448095
rect 674406 447916 674412 447940
rect 673198 447888 674412 447916
rect 674464 447916 674470 447940
rect 676270 447930 676440 447936
rect 674464 447888 676270 447916
rect 676270 447872 676440 447878
rect 674350 447792 674356 447816
rect 673198 447764 674356 447792
rect 674408 447792 674414 447816
rect 676934 447792 676940 447924
rect 674408 447764 676940 447792
rect 676934 447706 676940 447764
rect 676992 447706 676998 447924
rect 674178 447563 674184 447587
rect 673198 447535 674184 447563
rect 674236 447563 674242 447587
rect 676322 447563 676328 447654
rect 674236 447535 676328 447563
rect 676322 447436 676328 447535
rect 676380 447436 676386 447654
rect 674122 447369 674128 447393
rect 673198 447341 674128 447369
rect 674180 447369 674186 447393
rect 676882 447380 677052 447386
rect 674180 447341 676882 447369
rect 676882 447322 677052 447328
rect 675524 447256 675610 447264
rect 675524 446899 675538 447256
rect 675598 446899 675610 447256
rect 675524 446891 675610 446899
rect 676612 447256 676698 447264
rect 676612 446899 676626 447256
rect 676686 446899 676698 447256
rect 676612 446891 676698 446899
rect 674182 446720 674188 446744
rect 673198 446692 674188 446720
rect 674240 446720 674246 446744
rect 676270 446734 676440 446740
rect 674240 446692 676270 446720
rect 676270 446676 676440 446682
rect 674126 446596 674132 446620
rect 673198 446568 674132 446596
rect 674184 446596 674190 446620
rect 676934 446596 676940 446728
rect 674184 446568 676940 446596
rect 676934 446510 676940 446568
rect 676992 446510 676998 446728
rect 673954 446367 673960 446391
rect 673198 446339 673960 446367
rect 674012 446367 674018 446391
rect 676322 446367 676328 446458
rect 674012 446339 676328 446367
rect 676322 446240 676328 446339
rect 676380 446240 676386 446458
rect 673898 446173 673904 446197
rect 673198 446145 673904 446173
rect 673956 446173 673962 446197
rect 676882 446184 677052 446190
rect 673956 446145 676882 446173
rect 676882 446126 677052 446132
rect 673958 445524 673964 445548
rect 673198 445496 673964 445524
rect 674016 445524 674022 445548
rect 676270 445538 676440 445544
rect 674016 445496 676270 445524
rect 676270 445480 676440 445486
rect 673902 445400 673908 445424
rect 673198 445372 673908 445400
rect 673960 445400 673966 445424
rect 676934 445400 676940 445532
rect 673960 445372 676940 445400
rect 676934 445314 676940 445372
rect 676992 445314 676998 445532
rect 673730 445171 673736 445195
rect 673198 445143 673736 445171
rect 673788 445171 673794 445195
rect 676322 445171 676328 445262
rect 673788 445143 676328 445171
rect 676322 445044 676328 445143
rect 676380 445044 676386 445262
rect 673674 444977 673680 445001
rect 673198 444949 673680 444977
rect 673732 444977 673738 445001
rect 676882 444988 677052 444994
rect 673732 444949 676882 444977
rect 676882 444930 677052 444936
rect 673734 444328 673740 444352
rect 673198 444300 673740 444328
rect 673792 444328 673798 444352
rect 676270 444342 676440 444348
rect 673792 444300 676270 444328
rect 676270 444284 676440 444290
rect 673678 444204 673684 444228
rect 673198 444176 673684 444204
rect 673736 444204 673742 444228
rect 676934 444204 676940 444336
rect 673736 444176 676940 444204
rect 676934 444118 676940 444176
rect 676992 444118 676998 444336
rect 673506 443975 673512 443999
rect 673198 443947 673512 443975
rect 673564 443975 673570 443999
rect 676322 443975 676328 444066
rect 673564 443947 676328 443975
rect 676322 443848 676328 443947
rect 676380 443848 676386 444066
rect 673450 443781 673456 443805
rect 673198 443753 673456 443781
rect 673508 443781 673514 443805
rect 676882 443792 677052 443798
rect 673508 443753 676882 443781
rect 676882 443734 677052 443740
rect 673510 443132 673516 443156
rect 673198 443104 673516 443132
rect 673568 443132 673574 443156
rect 676270 443146 676440 443152
rect 673568 443104 676270 443132
rect 676270 443088 676440 443094
rect 673454 443008 673460 443032
rect 673198 442980 673460 443008
rect 673512 443008 673518 443032
rect 676934 443008 676940 443140
rect 673512 442980 676940 443008
rect 676934 442922 676940 442980
rect 676992 442922 676998 443140
rect 673282 442779 673288 442803
rect 673198 442751 673288 442779
rect 673340 442779 673346 442803
rect 676322 442779 676328 442870
rect 673340 442751 676328 442779
rect 676322 442652 676328 442751
rect 676380 442652 676386 442870
rect 673226 442585 673232 442609
rect 673198 442557 673232 442585
rect 673284 442585 673290 442609
rect 676882 442596 677052 442602
rect 673284 442557 676882 442585
rect 676882 442538 677052 442544
rect 673286 441936 673292 441960
rect 673198 441908 673292 441936
rect 673344 441936 673350 441960
rect 676270 441950 676440 441956
rect 673344 441908 676270 441936
rect 676270 441892 676440 441898
rect 673230 441812 673236 441836
rect 673198 441784 673236 441812
rect 673288 441812 673294 441836
rect 676934 441812 676940 441944
rect 673288 441784 676940 441812
rect 676934 441726 676940 441784
rect 676992 441726 676998 441944
rect 673058 441583 673064 441607
rect 672973 441555 673064 441583
rect 673116 441583 673122 441607
rect 676322 441583 676328 441674
rect 673116 441555 676328 441583
rect 676322 441456 676328 441555
rect 676380 441456 676386 441674
rect 673002 441389 673008 441413
rect 672973 441361 673008 441389
rect 673060 441389 673066 441413
rect 676882 441400 677052 441406
rect 673060 441361 676882 441389
rect 676882 441342 677052 441348
rect 673062 440740 673068 440764
rect 672980 440712 673068 440740
rect 673120 440740 673126 440764
rect 676270 440754 676440 440760
rect 673120 440712 676270 440740
rect 676270 440696 676440 440702
rect 673006 440616 673012 440640
rect 672980 440588 673012 440616
rect 673064 440616 673070 440640
rect 676934 440616 676940 440748
rect 673064 440588 676940 440616
rect 676934 440530 676940 440588
rect 676992 440530 676998 440748
rect 672834 440387 672840 440411
rect 672750 440359 672840 440387
rect 672892 440387 672898 440411
rect 676322 440387 676328 440478
rect 672892 440359 676328 440387
rect 676322 440260 676328 440359
rect 676380 440260 676386 440478
rect 672778 440193 672784 440217
rect 672750 440165 672784 440193
rect 672836 440193 672842 440217
rect 676882 440204 677052 440210
rect 672836 440165 676882 440193
rect 676882 440146 677052 440152
rect 672838 439544 672844 439568
rect 672750 439516 672844 439544
rect 672896 439544 672902 439568
rect 676270 439558 676440 439564
rect 672896 439516 676270 439544
rect 676270 439500 676440 439506
rect 672782 439420 672788 439444
rect 672750 439392 672788 439420
rect 672840 439420 672846 439444
rect 676934 439420 676940 439552
rect 672840 439392 676940 439420
rect 676934 439334 676940 439392
rect 676992 439334 676998 439552
rect 41235 352373 41241 352591
rect 41293 352500 41299 352591
rect 42149 352500 42155 352524
rect 41293 352472 42155 352500
rect 42207 352500 42213 352524
rect 42207 352472 44748 352500
rect 41293 352373 41299 352472
rect 40569 352317 40739 352323
rect 42205 352306 42211 352330
rect 40739 352278 42211 352306
rect 42263 352306 42269 352330
rect 42263 352278 44748 352306
rect 40569 352259 40739 352265
rect 41181 351671 41351 351677
rect 40623 351447 40629 351665
rect 40681 351533 40687 351665
rect 42145 351657 42151 351681
rect 41351 351629 42151 351657
rect 42203 351657 42209 351681
rect 42203 351629 44748 351657
rect 41181 351613 41351 351619
rect 42201 351533 42207 351557
rect 40681 351505 42207 351533
rect 42259 351533 42266 351557
rect 42259 351505 44748 351533
rect 40681 351447 40687 351505
rect 41235 351177 41241 351395
rect 41293 351304 41299 351395
rect 41293 351276 42379 351304
rect 41293 351177 41299 351276
rect 42373 351252 42379 351276
rect 42431 351276 44748 351304
rect 42431 351252 42437 351276
rect 40569 351121 40739 351127
rect 42429 351110 42435 351134
rect 40739 351082 42435 351110
rect 42487 351110 42493 351134
rect 42487 351082 44748 351110
rect 40569 351063 40739 351069
rect 41171 350475 41341 350481
rect 40623 350251 40629 350469
rect 40681 350337 40687 350469
rect 42369 350461 42375 350485
rect 41341 350433 42375 350461
rect 42427 350461 42433 350485
rect 42427 350433 44748 350461
rect 41171 350417 41341 350423
rect 42425 350337 42431 350361
rect 40681 350309 42431 350337
rect 42483 350337 42489 350361
rect 42483 350309 44748 350337
rect 40681 350251 40687 350309
rect 41235 349981 41241 350199
rect 41293 350108 41299 350199
rect 42597 350108 42603 350132
rect 41293 350080 42603 350108
rect 42655 350108 42661 350132
rect 42655 350080 44748 350108
rect 41293 349981 41299 350080
rect 40569 349925 40739 349931
rect 42653 349914 42659 349938
rect 40739 349886 42659 349914
rect 42711 349914 42717 349938
rect 42711 349886 44748 349914
rect 40569 349867 40739 349873
rect 41181 349279 41351 349285
rect 40623 349055 40629 349273
rect 40681 349141 40687 349273
rect 42593 349265 42599 349289
rect 41351 349237 42599 349265
rect 42651 349265 42657 349289
rect 42651 349237 44748 349265
rect 41181 349221 41351 349227
rect 42649 349141 42655 349165
rect 40681 349113 42655 349141
rect 42707 349141 42713 349165
rect 42707 349113 44748 349141
rect 40681 349055 40687 349113
rect 41235 348785 41241 349003
rect 41293 348912 41299 349003
rect 41293 348884 42827 348912
rect 41293 348785 41299 348884
rect 42821 348860 42827 348884
rect 42879 348884 44748 348912
rect 42879 348860 42885 348884
rect 40569 348729 40739 348735
rect 42877 348718 42883 348742
rect 40739 348690 42883 348718
rect 42935 348718 42941 348742
rect 42935 348690 44748 348718
rect 40569 348671 40739 348677
rect 41181 348083 41351 348089
rect 40623 347859 40629 348077
rect 40681 347945 40687 348077
rect 42817 348069 42823 348093
rect 41351 348041 42823 348069
rect 42875 348069 42881 348093
rect 42875 348041 44748 348069
rect 41181 348025 41351 348031
rect 42873 347945 42879 347969
rect 40681 347917 42879 347945
rect 42931 347945 42937 347969
rect 42931 347917 44748 347945
rect 40681 347859 40687 347917
rect 41235 347589 41241 347807
rect 41293 347716 41299 347807
rect 43045 347716 43051 347740
rect 41293 347688 43051 347716
rect 43103 347716 43109 347740
rect 43103 347688 44748 347716
rect 41293 347589 41299 347688
rect 40569 347533 40739 347539
rect 43101 347522 43107 347546
rect 40739 347494 43107 347522
rect 43159 347522 43165 347546
rect 43159 347494 44748 347522
rect 40569 347475 40739 347481
rect 40373 347316 40459 347324
rect 40373 346959 40390 347316
rect 40450 346959 40459 347316
rect 40373 346951 40459 346959
rect 41458 347316 41544 347324
rect 41458 346959 41472 347316
rect 41532 346959 41544 347316
rect 41458 346951 41544 346959
rect 41181 346887 41351 346893
rect 40623 346663 40629 346881
rect 40681 346749 40687 346881
rect 43041 346873 43047 346897
rect 41351 346845 43047 346873
rect 43099 346873 43105 346897
rect 43099 346845 44748 346873
rect 41181 346829 41351 346835
rect 43097 346749 43103 346773
rect 40681 346721 43103 346749
rect 43155 346749 43161 346773
rect 43155 346721 44748 346749
rect 40681 346663 40687 346721
rect 41235 346393 41241 346611
rect 41293 346520 41299 346611
rect 43269 346520 43275 346544
rect 41293 346492 43275 346520
rect 43327 346520 43333 346544
rect 43327 346492 44748 346520
rect 41293 346393 41299 346492
rect 40569 346337 40739 346343
rect 43325 346326 43331 346350
rect 40739 346298 43331 346326
rect 43383 346326 43389 346350
rect 43383 346298 44748 346326
rect 40569 346279 40739 346285
rect 40919 346120 41005 346128
rect 40919 345763 40931 346120
rect 40991 345763 41005 346120
rect 40919 345755 41005 345763
rect 42007 346120 42093 346128
rect 42007 345763 42019 346120
rect 42079 345763 42093 346120
rect 42007 345755 42093 345763
rect 41181 345691 41351 345697
rect 40623 345467 40629 345685
rect 40681 345553 40687 345685
rect 43265 345677 43271 345701
rect 41351 345649 43271 345677
rect 43323 345677 43329 345701
rect 43323 345649 44748 345677
rect 41181 345633 41351 345639
rect 43321 345553 43327 345577
rect 40681 345525 43327 345553
rect 43379 345553 43385 345577
rect 43379 345525 44748 345553
rect 40681 345467 40687 345525
rect 41235 345197 41241 345415
rect 41293 345324 41299 345415
rect 43493 345324 43499 345348
rect 41293 345296 43499 345324
rect 43551 345324 43557 345348
rect 43551 345296 44748 345324
rect 41293 345197 41299 345296
rect 40569 345141 40739 345147
rect 43549 345130 43555 345154
rect 40739 345102 43555 345130
rect 43607 345130 43613 345154
rect 43607 345102 44748 345130
rect 40569 345083 40739 345089
rect 41181 344495 41351 344501
rect 40623 344271 40629 344489
rect 40681 344357 40687 344489
rect 43489 344481 43495 344505
rect 41351 344453 43495 344481
rect 43547 344481 43553 344505
rect 43547 344453 44748 344481
rect 41181 344437 41351 344443
rect 43545 344357 43551 344381
rect 40681 344329 43551 344357
rect 43603 344357 43609 344381
rect 43603 344329 44748 344357
rect 40681 344271 40687 344329
rect 41235 344001 41241 344219
rect 41293 344128 41299 344219
rect 43717 344128 43723 344152
rect 41293 344100 43723 344128
rect 43775 344128 43781 344152
rect 43775 344100 44748 344128
rect 41293 344001 41299 344100
rect 40569 343945 40739 343951
rect 43773 343934 43779 343958
rect 40739 343906 43779 343934
rect 43831 343934 43837 343958
rect 43831 343906 44748 343934
rect 40569 343887 40739 343893
rect 41181 343299 41351 343305
rect 40623 343161 40629 343293
rect 40681 343161 40687 343293
rect 43713 343285 43719 343309
rect 41351 343257 43719 343285
rect 43771 343285 43777 343309
rect 43771 343257 44748 343285
rect 41181 343241 41351 343247
rect 43769 343161 43775 343185
rect 40569 343133 43775 343161
rect 43827 343161 43833 343185
rect 43827 343133 44748 343161
rect 40623 343075 40629 343133
rect 40681 343075 40687 343133
rect 41235 342805 41241 343023
rect 41293 342932 41299 343023
rect 43941 342932 43947 342956
rect 41293 342904 43947 342932
rect 43999 342932 44005 342956
rect 43999 342904 44748 342932
rect 41293 342805 41299 342904
rect 40569 342749 40739 342755
rect 43997 342738 44003 342762
rect 40739 342710 44003 342738
rect 44055 342738 44061 342762
rect 44055 342710 44748 342738
rect 40569 342691 40739 342697
rect 41181 342103 41351 342109
rect 40623 341879 40629 342097
rect 40681 341965 40687 342097
rect 43937 342089 43943 342113
rect 41351 342061 43943 342089
rect 43995 342089 44001 342113
rect 43995 342061 44748 342089
rect 41181 342045 41351 342051
rect 43993 341965 43999 341989
rect 40681 341937 43999 341965
rect 44051 341965 44057 341989
rect 44051 341937 44748 341965
rect 40681 341879 40687 341937
rect 41235 341609 41241 341827
rect 41293 341736 41299 341827
rect 44165 341736 44171 341760
rect 41293 341708 44171 341736
rect 44223 341736 44229 341760
rect 44223 341708 44748 341736
rect 41293 341609 41299 341708
rect 40569 341553 40739 341559
rect 44221 341542 44227 341566
rect 40739 341514 44227 341542
rect 44279 341542 44285 341566
rect 44279 341514 44748 341542
rect 40569 341495 40739 341501
rect 41181 340907 41351 340913
rect 40623 340683 40629 340901
rect 40681 340769 40687 340901
rect 44161 340893 44167 340917
rect 41351 340865 44167 340893
rect 44219 340893 44225 340917
rect 44219 340865 44748 340893
rect 41181 340849 41351 340855
rect 44217 340769 44223 340793
rect 40681 340741 44223 340769
rect 44275 340769 44281 340793
rect 44275 340741 44748 340769
rect 40681 340683 40687 340741
rect 41235 340413 41241 340631
rect 41293 340540 41299 340631
rect 44389 340540 44395 340564
rect 41293 340512 44395 340540
rect 44447 340540 44453 340564
rect 44447 340512 44748 340540
rect 41293 340413 41299 340512
rect 40569 340357 40739 340363
rect 44445 340346 44451 340370
rect 40739 340318 44451 340346
rect 44503 340346 44509 340370
rect 44503 340318 44748 340346
rect 40569 340299 40739 340305
rect 41181 339711 41351 339717
rect 40623 339487 40629 339705
rect 40681 339573 40687 339705
rect 44385 339697 44391 339721
rect 41351 339669 44391 339697
rect 44443 339697 44449 339721
rect 44443 339669 44748 339697
rect 41181 339653 41351 339659
rect 44441 339573 44447 339597
rect 40681 339545 44447 339573
rect 44499 339573 44505 339597
rect 44499 339545 44748 339573
rect 40681 339487 40687 339545
rect 41235 339217 41241 339435
rect 41293 339344 41299 339435
rect 44613 339344 44619 339368
rect 41293 339316 44619 339344
rect 44671 339344 44677 339368
rect 44671 339316 44768 339344
rect 41293 339217 41299 339316
rect 40569 339161 40739 339167
rect 44669 339150 44675 339174
rect 40739 339122 44675 339150
rect 44727 339150 44733 339174
rect 44727 339122 44768 339150
rect 40569 339103 40739 339109
rect 41181 338515 41351 338521
rect 40623 338291 40629 338509
rect 40681 338377 40687 338509
rect 44609 338501 44615 338525
rect 41351 338473 44615 338501
rect 44667 338501 44673 338525
rect 44667 338473 44749 338501
rect 41181 338457 41351 338463
rect 44665 338377 44671 338401
rect 40681 338349 44671 338377
rect 44723 338377 44729 338401
rect 44723 338349 44749 338377
rect 40681 338291 40687 338349
rect 41235 338021 41241 338239
rect 41293 338148 41299 338239
rect 44837 338148 44843 338172
rect 41293 338120 44843 338148
rect 44895 338148 44901 338172
rect 44895 338120 44982 338148
rect 41293 338021 41299 338120
rect 40569 337965 40739 337971
rect 44893 337954 44899 337978
rect 40739 337926 44899 337954
rect 44951 337954 44957 337978
rect 44951 337926 44982 337954
rect 40569 337907 40739 337913
rect 41181 337319 41351 337325
rect 40623 337095 40629 337313
rect 40681 337181 40687 337313
rect 44833 337305 44839 337329
rect 41351 337277 44839 337305
rect 44891 337305 44897 337329
rect 44891 337277 44961 337305
rect 41181 337261 41351 337267
rect 44889 337181 44895 337205
rect 40681 337153 44895 337181
rect 44947 337181 44953 337205
rect 44947 337153 44961 337181
rect 40681 337095 40687 337153
rect 41235 336825 41241 337043
rect 41293 336952 41299 337043
rect 41293 336924 45067 336952
rect 41293 336825 41299 336924
rect 45061 336900 45067 336924
rect 45119 336924 45195 336952
rect 45119 336900 45125 336924
rect 40569 336769 40739 336775
rect 45117 336758 45123 336782
rect 40739 336730 45123 336758
rect 45175 336758 45181 336782
rect 45175 336730 45195 336758
rect 40569 336711 40739 336717
rect 41181 336123 41351 336129
rect 40623 335899 40629 336117
rect 40681 335985 40687 336117
rect 45057 336109 45063 336133
rect 41351 336081 45063 336109
rect 45115 336109 45121 336133
rect 45115 336081 45206 336109
rect 41181 336065 41351 336071
rect 45113 335985 45119 336009
rect 40681 335957 45119 335985
rect 45171 335985 45177 336009
rect 45171 335957 45206 335985
rect 40681 335899 40687 335957
rect 41235 335629 41241 335847
rect 41293 335756 41299 335847
rect 45285 335756 45291 335780
rect 41293 335728 45291 335756
rect 45343 335756 45349 335780
rect 45343 335728 45420 335756
rect 41293 335629 41299 335728
rect 40569 335573 40739 335579
rect 45341 335562 45347 335586
rect 40739 335534 45347 335562
rect 45399 335562 45405 335586
rect 45399 335534 45420 335562
rect 40569 335515 40739 335521
rect 41181 334927 41351 334933
rect 40623 334703 40629 334921
rect 40681 334789 40687 334921
rect 45281 334913 45287 334937
rect 41351 334885 45287 334913
rect 45339 334913 45345 334937
rect 45339 334885 45420 334913
rect 41181 334869 41351 334875
rect 45337 334789 45343 334813
rect 40681 334761 45343 334789
rect 45395 334789 45401 334813
rect 45395 334761 45420 334789
rect 40681 334703 40687 334761
rect 429504 47654 429532 47673
rect 430347 47658 430375 47673
rect 429504 47648 429556 47654
rect 134104 47626 134132 47645
rect 134947 47630 134975 47645
rect 134104 47620 134156 47626
rect 134104 47562 134156 47568
rect 134947 47624 134999 47630
rect 429504 47590 429556 47596
rect 430347 47652 430399 47658
rect 430347 47594 430399 47600
rect 430576 47598 430604 47610
rect 431349 47602 431377 47617
rect 134947 47566 134999 47572
rect 135176 47570 135204 47580
rect 135949 47574 135977 47585
rect 134104 43272 134132 47562
rect 134088 43102 134094 43272
rect 134146 43102 134152 43272
rect 134947 43220 134975 47566
rect 135176 47564 135228 47570
rect 135176 47506 135228 47512
rect 135949 47568 136001 47574
rect 135949 47510 136001 47516
rect 134848 43214 135066 43220
rect 134848 43156 135066 43162
rect 135176 42608 135204 47506
rect 135300 47458 135328 47480
rect 135300 47452 135352 47458
rect 135300 47394 135352 47400
rect 135300 43272 135328 47394
rect 135284 43102 135290 43272
rect 135342 43102 135348 43272
rect 135949 42660 135977 47510
rect 136143 47462 136171 47480
rect 136143 47456 136195 47462
rect 136143 47398 136195 47404
rect 136372 47402 136400 47410
rect 137145 47406 137173 47417
rect 136143 43220 136171 47398
rect 136372 47396 136424 47402
rect 136372 47338 136424 47344
rect 137145 47400 137197 47406
rect 137145 47342 137197 47348
rect 136044 43214 136262 43220
rect 136044 43156 136262 43162
rect 135118 42602 135336 42608
rect 135118 42544 135336 42550
rect 135930 42490 135936 42660
rect 135988 42490 135994 42660
rect 136372 42608 136400 47338
rect 136496 47290 136524 47309
rect 136496 47284 136548 47290
rect 136496 47226 136548 47232
rect 136496 43272 136524 47226
rect 136480 43102 136486 43272
rect 136538 43102 136544 43272
rect 137145 42660 137173 47342
rect 137339 47294 137367 47304
rect 137339 47288 137391 47294
rect 137339 47230 137391 47236
rect 137568 47234 137596 47247
rect 138341 47238 138369 47252
rect 137339 43220 137367 47230
rect 137568 47228 137620 47234
rect 137568 47170 137620 47176
rect 138341 47232 138393 47238
rect 138341 47174 138393 47180
rect 137240 43214 137458 43220
rect 137240 43156 137458 43162
rect 136314 42602 136532 42608
rect 136314 42544 136532 42550
rect 137126 42490 137132 42660
rect 137184 42490 137190 42660
rect 137568 42608 137596 47170
rect 137692 47122 137720 47163
rect 137692 47116 137744 47122
rect 137692 47058 137744 47064
rect 137692 43272 137720 47058
rect 137676 43102 137682 43272
rect 137734 43102 137740 43272
rect 138341 42660 138369 47174
rect 138535 47126 138563 47139
rect 138535 47120 138587 47126
rect 138535 47062 138587 47068
rect 138764 47066 138792 47090
rect 139537 47070 139565 47094
rect 138535 43220 138563 47062
rect 138764 47060 138816 47066
rect 138764 47002 138816 47008
rect 139537 47064 139589 47070
rect 139537 47006 139589 47012
rect 138436 43214 138654 43220
rect 138436 43156 138654 43162
rect 137510 42602 137728 42608
rect 137510 42544 137728 42550
rect 138322 42490 138328 42660
rect 138380 42490 138386 42660
rect 138764 42608 138792 47002
rect 138888 46954 138916 46974
rect 138888 46948 138940 46954
rect 138888 46890 138940 46896
rect 138888 43272 138916 46890
rect 138872 43102 138878 43272
rect 138930 43102 138936 43272
rect 139537 42660 139565 47006
rect 139731 46958 139759 46981
rect 139731 46952 139783 46958
rect 139731 46894 139783 46900
rect 139960 46898 139988 46903
rect 139731 43220 139759 46894
rect 139960 46892 140012 46898
rect 139960 46834 140012 46840
rect 139632 43214 139850 43220
rect 139632 43156 139850 43162
rect 138706 42602 138924 42608
rect 138706 42544 138924 42550
rect 139518 42490 139524 42660
rect 139576 42490 139582 42660
rect 139960 42608 139988 46834
rect 140084 46786 140112 46812
rect 140084 46780 140136 46786
rect 140084 46722 140136 46728
rect 140084 43272 140112 46722
rect 140733 46566 140761 46578
rect 140733 46560 140785 46566
rect 140927 46510 140955 46536
rect 140733 46502 140785 46508
rect 140903 46504 140955 46510
rect 140068 43102 140074 43272
rect 140126 43102 140132 43272
rect 140733 42660 140761 46502
rect 140903 46446 140955 46452
rect 140927 43220 140955 46446
rect 141156 46450 141184 46463
rect 141929 46454 141957 46462
rect 141156 46444 141208 46450
rect 141929 46448 141981 46454
rect 141156 46386 141208 46392
rect 141280 46394 141308 46430
rect 141280 46388 141332 46394
rect 140828 43214 141046 43220
rect 140828 43156 141046 43162
rect 139902 42602 140120 42608
rect 139902 42544 140120 42550
rect 140714 42490 140720 42660
rect 140772 42490 140778 42660
rect 141156 42608 141184 46386
rect 141280 46330 141332 46336
rect 141929 46390 141981 46396
rect 142123 46398 142151 46438
rect 142123 46392 142175 46398
rect 141280 43272 141308 46330
rect 141264 43102 141270 43272
rect 141322 43102 141328 43272
rect 141929 42660 141957 46390
rect 142123 46334 142175 46340
rect 142352 46338 142380 46350
rect 143125 46342 143153 46356
rect 142123 43220 142151 46334
rect 142352 46332 142404 46338
rect 143125 46336 143177 46342
rect 142352 46274 142404 46280
rect 142476 46282 142504 46301
rect 143319 46286 143347 46305
rect 142476 46276 142528 46282
rect 142024 43214 142242 43220
rect 142024 43156 142242 43162
rect 141098 42602 141316 42608
rect 141098 42544 141316 42550
rect 141910 42490 141916 42660
rect 141968 42490 141974 42660
rect 142352 42608 142380 46274
rect 142476 46218 142528 46224
rect 143125 46278 143177 46284
rect 143295 46280 143347 46286
rect 142476 43272 142504 46218
rect 142460 43102 142466 43272
rect 142518 43102 142524 43272
rect 143125 42660 143153 46278
rect 143295 46222 143347 46228
rect 143319 43220 143347 46222
rect 143548 46226 143576 46469
rect 143548 46220 143600 46226
rect 143548 46162 143600 46168
rect 143672 46170 143700 46469
rect 144321 46230 144349 46469
rect 144321 46224 144373 46230
rect 143672 46164 143724 46170
rect 143220 43214 143438 43220
rect 143220 43156 143438 43162
rect 142294 42602 142512 42608
rect 142294 42544 142512 42550
rect 143106 42490 143112 42660
rect 143164 42490 143170 42660
rect 143548 42608 143576 46162
rect 143672 46106 143724 46112
rect 144321 46166 144373 46172
rect 144515 46174 144543 46469
rect 144515 46168 144567 46174
rect 143672 43272 143700 46106
rect 143656 43102 143662 43272
rect 143714 43102 143720 43272
rect 144321 42660 144349 46166
rect 144515 46110 144567 46116
rect 144744 46114 144772 46469
rect 144515 43220 144543 46110
rect 144744 46108 144796 46114
rect 144744 46050 144796 46056
rect 144868 46058 144896 46469
rect 145517 46118 145545 46469
rect 145517 46112 145569 46118
rect 144868 46052 144920 46058
rect 144416 43214 144634 43220
rect 144416 43156 144634 43162
rect 143490 42602 143708 42608
rect 143490 42544 143708 42550
rect 144302 42490 144308 42660
rect 144360 42490 144366 42660
rect 144744 42608 144772 46050
rect 144868 45994 144920 46000
rect 145517 46054 145569 46060
rect 145711 46062 145739 46469
rect 145711 46056 145763 46062
rect 144868 43272 144896 45994
rect 144852 43102 144858 43272
rect 144910 43102 144916 43272
rect 145517 42660 145545 46054
rect 145711 45998 145763 46004
rect 145940 46002 145968 46469
rect 145711 43220 145739 45998
rect 145940 45996 145992 46002
rect 145940 45938 145992 45944
rect 146064 45946 146092 46469
rect 146713 46006 146741 46469
rect 146713 46000 146765 46006
rect 146064 45940 146116 45946
rect 145612 43214 145830 43220
rect 145612 43156 145830 43162
rect 144686 42602 144904 42608
rect 144686 42544 144904 42550
rect 145498 42490 145504 42660
rect 145556 42490 145562 42660
rect 145940 42608 145968 45938
rect 146064 45882 146116 45888
rect 146713 45942 146765 45948
rect 146907 45950 146935 46469
rect 146907 45944 146959 45950
rect 146064 43272 146092 45882
rect 146191 44004 146564 44018
rect 146191 43944 146199 44004
rect 146556 43944 146564 44004
rect 146191 43932 146564 43944
rect 146048 43102 146054 43272
rect 146106 43102 146112 43272
rect 146191 42916 146564 42930
rect 146191 42856 146199 42916
rect 146556 42856 146564 42916
rect 146191 42844 146564 42856
rect 146713 42660 146741 45942
rect 146907 45886 146959 45892
rect 147136 45890 147164 46469
rect 146907 43220 146935 45886
rect 147136 45884 147188 45890
rect 147136 45826 147188 45832
rect 146808 43214 147026 43220
rect 146808 43156 147026 43162
rect 145882 42602 146100 42608
rect 145882 42544 146100 42550
rect 146694 42490 146700 42660
rect 146752 42490 146758 42660
rect 147136 42608 147164 45826
rect 147260 45778 147288 46469
rect 147909 45894 147937 46469
rect 147909 45888 147961 45894
rect 147909 45830 147961 45836
rect 147260 45772 147312 45778
rect 147260 45714 147312 45720
rect 147260 43272 147288 45714
rect 147387 43457 147760 43469
rect 147387 43397 147395 43457
rect 147752 43397 147760 43457
rect 147387 43383 147760 43397
rect 147244 43102 147250 43272
rect 147302 43102 147308 43272
rect 147909 42660 147937 45830
rect 148103 45782 148131 46469
rect 148103 45776 148155 45782
rect 148103 45718 148155 45724
rect 148332 45722 148360 46469
rect 148103 43220 148131 45718
rect 148332 45716 148384 45722
rect 148332 45658 148384 45664
rect 148004 43214 148222 43220
rect 148004 43156 148222 43162
rect 147078 42602 147296 42608
rect 147078 42544 147296 42550
rect 147890 42490 147896 42660
rect 147948 42490 147954 42660
rect 148332 42608 148360 45658
rect 148456 45610 148484 46469
rect 149105 45726 149133 46469
rect 149105 45720 149157 45726
rect 149105 45662 149157 45668
rect 148456 45604 148508 45610
rect 148456 45546 148508 45552
rect 148456 43272 148484 45546
rect 148440 43102 148446 43272
rect 148498 43102 148504 43272
rect 149105 42660 149133 45662
rect 149299 45614 149327 46469
rect 149299 45608 149351 45614
rect 149299 45550 149351 45556
rect 149528 45554 149556 46469
rect 149299 43220 149327 45550
rect 149528 45548 149580 45554
rect 149528 45490 149580 45496
rect 149200 43214 149418 43220
rect 149200 43156 149418 43162
rect 148274 42602 148492 42608
rect 148274 42544 148492 42550
rect 149086 42490 149092 42660
rect 149144 42490 149150 42660
rect 149528 42608 149556 45490
rect 149652 45442 149680 46469
rect 150301 45558 150329 46469
rect 150301 45552 150353 45558
rect 150301 45494 150353 45500
rect 149652 45436 149704 45442
rect 149652 45378 149704 45384
rect 149652 43272 149680 45378
rect 149636 43102 149642 43272
rect 149694 43102 149700 43272
rect 150301 42660 150329 45494
rect 150495 45446 150523 46469
rect 150495 45440 150547 45446
rect 150495 45382 150547 45388
rect 150724 45386 150752 46469
rect 150495 43220 150523 45382
rect 150724 45380 150776 45386
rect 150724 45322 150776 45328
rect 150396 43214 150614 43220
rect 150396 43156 150614 43162
rect 149470 42602 149688 42608
rect 149470 42544 149688 42550
rect 150282 42490 150288 42660
rect 150340 42490 150346 42660
rect 150724 42608 150752 45322
rect 150848 45274 150876 46469
rect 151497 45390 151525 46469
rect 151497 45384 151549 45390
rect 151497 45326 151549 45332
rect 150848 45268 150900 45274
rect 150848 45210 150900 45216
rect 150848 43272 150876 45210
rect 150832 43102 150838 43272
rect 150890 43102 150896 43272
rect 151497 42660 151525 45326
rect 151691 45278 151719 46469
rect 151691 45272 151743 45278
rect 151691 45214 151743 45220
rect 151920 45218 151948 46469
rect 151691 43220 151719 45214
rect 151920 45212 151972 45218
rect 151920 45154 151972 45160
rect 151592 43214 151810 43220
rect 151592 43156 151810 43162
rect 150666 42602 150884 42608
rect 150666 42544 150884 42550
rect 151478 42490 151484 42660
rect 151536 42490 151542 42660
rect 151920 42608 151948 45154
rect 152044 45106 152072 46469
rect 152693 45222 152721 46469
rect 152693 45216 152745 45222
rect 152693 45158 152745 45164
rect 152044 45100 152096 45106
rect 152044 45042 152096 45048
rect 152044 43272 152072 45042
rect 152028 43102 152034 43272
rect 152086 43102 152092 43272
rect 152693 42660 152721 45158
rect 152887 45110 152915 46469
rect 152887 45104 152939 45110
rect 152887 45046 152939 45052
rect 153116 45050 153144 46469
rect 152887 43220 152915 45046
rect 153116 45044 153168 45050
rect 153116 44986 153168 44992
rect 152788 43214 153006 43220
rect 152788 43156 153006 43162
rect 151862 42602 152080 42608
rect 151862 42544 152080 42550
rect 152674 42490 152680 42660
rect 152732 42490 152738 42660
rect 153116 42608 153144 44986
rect 153240 44938 153268 46469
rect 153889 45054 153917 46469
rect 153889 45048 153941 45054
rect 153889 44990 153941 44996
rect 153240 44932 153292 44938
rect 153240 44874 153292 44880
rect 153240 43272 153268 44874
rect 153224 43102 153230 43272
rect 153282 43102 153288 43272
rect 153889 42660 153917 44990
rect 154083 44942 154111 46469
rect 154083 44936 154135 44942
rect 154083 44878 154135 44884
rect 154312 44882 154340 46469
rect 154083 43220 154111 44878
rect 154312 44876 154364 44882
rect 154312 44818 154364 44824
rect 153984 43214 154202 43220
rect 153984 43156 154202 43162
rect 153058 42602 153276 42608
rect 153058 42544 153276 42550
rect 153870 42490 153876 42660
rect 153928 42490 153934 42660
rect 154312 42608 154340 44818
rect 154436 44770 154464 46469
rect 155085 44886 155113 46469
rect 155085 44880 155137 44886
rect 155085 44822 155137 44828
rect 154436 44764 154488 44770
rect 154436 44706 154488 44712
rect 154436 43272 154464 44706
rect 154420 43102 154426 43272
rect 154478 43102 154484 43272
rect 155085 42660 155113 44822
rect 155279 44774 155307 46469
rect 155255 44768 155307 44774
rect 155255 44710 155307 44716
rect 155279 43220 155307 44710
rect 155508 44714 155536 46469
rect 155508 44708 155560 44714
rect 155508 44650 155560 44656
rect 155180 43214 155398 43220
rect 155180 43156 155398 43162
rect 154254 42602 154472 42608
rect 154254 42544 154472 42550
rect 155066 42490 155072 42660
rect 155124 42490 155130 42660
rect 155508 42608 155536 44650
rect 155632 44602 155660 46469
rect 156281 44718 156309 46469
rect 156281 44712 156333 44718
rect 156281 44654 156333 44660
rect 155632 44596 155684 44602
rect 155632 44538 155684 44544
rect 155632 43272 155660 44538
rect 155616 43102 155622 43272
rect 155674 43102 155680 43272
rect 156281 42660 156309 44654
rect 156475 44606 156503 46469
rect 156475 44600 156527 44606
rect 156475 44542 156527 44548
rect 156704 44546 156732 46469
rect 156475 43220 156503 44542
rect 156704 44540 156756 44546
rect 156704 44482 156756 44488
rect 156376 43214 156594 43220
rect 156376 43156 156594 43162
rect 155450 42602 155668 42608
rect 155450 42544 155668 42550
rect 156262 42490 156268 42660
rect 156320 42490 156326 42660
rect 156704 42608 156732 44482
rect 156828 44434 156856 46469
rect 157477 44550 157505 46469
rect 157477 44544 157529 44550
rect 157477 44486 157529 44492
rect 156828 44428 156880 44434
rect 156828 44370 156880 44376
rect 156828 43272 156856 44370
rect 156812 43102 156818 43272
rect 156870 43102 156876 43272
rect 157477 42660 157505 44486
rect 157671 44438 157699 46469
rect 157647 44432 157699 44438
rect 157647 44374 157699 44380
rect 157671 43220 157699 44374
rect 157900 44322 157928 46469
rect 157900 44316 157952 44322
rect 157900 44258 157952 44264
rect 157572 43214 157790 43220
rect 157572 43156 157790 43162
rect 157900 42848 157928 44258
rect 158024 44210 158052 46469
rect 158673 44326 158701 46469
rect 158673 44320 158725 44326
rect 158673 44262 158725 44268
rect 158024 44204 158076 44210
rect 158024 44146 158076 44152
rect 158024 43272 158052 44146
rect 158008 43102 158014 43272
rect 158066 43102 158072 43272
rect 158673 42848 158701 44262
rect 158867 44214 158895 46469
rect 158867 44208 158919 44214
rect 158867 44150 158919 44156
rect 158867 43220 158895 44150
rect 429504 43272 429532 47590
rect 158768 43214 158986 43220
rect 158768 43156 158986 43162
rect 429488 43102 429494 43272
rect 429546 43102 429552 43272
rect 430347 43220 430375 47594
rect 430576 47592 430628 47598
rect 430576 47534 430628 47540
rect 431349 47596 431401 47602
rect 431349 47538 431401 47544
rect 430248 43214 430466 43220
rect 430248 43156 430466 43162
rect 157900 42820 158055 42848
rect 158673 42820 158828 42848
rect 158027 42660 158055 42820
rect 156646 42602 156864 42608
rect 156646 42544 156864 42550
rect 157458 42490 157464 42660
rect 157516 42490 157522 42660
rect 158010 42490 158016 42660
rect 158068 42490 158074 42660
rect 158800 42608 158828 42820
rect 430576 42608 430604 47534
rect 430700 47486 430728 47505
rect 430700 47480 430752 47486
rect 430700 47422 430752 47428
rect 430700 43272 430728 47422
rect 430684 43102 430690 43272
rect 430742 43102 430748 43272
rect 431349 42660 431377 47538
rect 431543 47490 431571 47515
rect 431543 47484 431595 47490
rect 431543 47426 431595 47432
rect 431772 47430 431800 47447
rect 432545 47434 432573 47445
rect 431543 43220 431571 47426
rect 431772 47424 431824 47430
rect 431772 47366 431824 47372
rect 432545 47428 432597 47434
rect 432545 47370 432597 47376
rect 431444 43214 431662 43220
rect 431444 43156 431662 43162
rect 158668 42602 158886 42608
rect 158668 42544 158886 42550
rect 430518 42602 430736 42608
rect 430518 42544 430736 42550
rect 431330 42490 431336 42660
rect 431388 42490 431394 42660
rect 431772 42608 431800 47366
rect 431896 47318 431924 47341
rect 431896 47312 431948 47318
rect 431896 47254 431948 47260
rect 431896 43272 431924 47254
rect 431880 43102 431886 43272
rect 431938 43102 431944 43272
rect 432545 42660 432573 47370
rect 432739 47322 432767 47344
rect 432739 47316 432791 47322
rect 432739 47258 432791 47264
rect 432968 47262 432996 47279
rect 433741 47266 433769 47280
rect 432739 43220 432767 47258
rect 432968 47256 433020 47262
rect 432968 47198 433020 47204
rect 433741 47260 433793 47266
rect 433741 47202 433793 47208
rect 432640 43214 432858 43220
rect 432640 43156 432858 43162
rect 431714 42602 431932 42608
rect 431714 42544 431932 42550
rect 432526 42490 432532 42660
rect 432584 42490 432590 42660
rect 432968 42608 432996 47198
rect 433092 47150 433120 47163
rect 433092 47144 433144 47150
rect 433092 47086 433144 47092
rect 433092 43272 433120 47086
rect 433076 43102 433082 43272
rect 433134 43102 433140 43272
rect 433741 42660 433769 47202
rect 433935 47154 433963 47186
rect 433935 47148 433987 47154
rect 433935 47090 433987 47096
rect 434164 47094 434192 47108
rect 434937 47098 434965 47106
rect 433935 43220 433963 47090
rect 434164 47088 434216 47094
rect 434164 47030 434216 47036
rect 434937 47092 434989 47098
rect 434937 47034 434989 47040
rect 433836 43214 434054 43220
rect 433836 43156 434054 43162
rect 432910 42602 433128 42608
rect 432910 42544 433128 42550
rect 433722 42490 433728 42660
rect 433780 42490 433786 42660
rect 434164 42608 434192 47030
rect 434288 46982 434316 46998
rect 434288 46976 434340 46982
rect 434288 46918 434340 46924
rect 434288 43272 434316 46918
rect 434272 43102 434278 43272
rect 434330 43102 434336 43272
rect 434937 42660 434965 47034
rect 435131 46986 435159 47002
rect 435131 46980 435183 46986
rect 435131 46922 435183 46928
rect 435360 46926 435388 46935
rect 436133 46930 436161 46941
rect 435131 43220 435159 46922
rect 435360 46920 435412 46926
rect 435360 46862 435412 46868
rect 436133 46924 436185 46930
rect 436133 46866 436185 46872
rect 435032 43214 435250 43220
rect 435032 43156 435250 43162
rect 434106 42602 434324 42608
rect 434106 42544 434324 42550
rect 434918 42490 434924 42660
rect 434976 42490 434982 42660
rect 435360 42608 435388 46862
rect 435484 46814 435512 46836
rect 435484 46808 435536 46814
rect 435484 46750 435536 46756
rect 435484 43272 435512 46750
rect 435468 43102 435474 43272
rect 435526 43102 435532 43272
rect 436133 42660 436161 46866
rect 436327 46818 436355 46840
rect 436303 46812 436355 46818
rect 436303 46754 436355 46760
rect 436327 43220 436355 46754
rect 436556 46758 436584 46769
rect 437329 46762 437357 46774
rect 436556 46752 436608 46758
rect 436556 46694 436608 46700
rect 437329 46756 437381 46762
rect 437329 46698 437381 46704
rect 436228 43214 436446 43220
rect 436228 43156 436446 43162
rect 435302 42602 435520 42608
rect 435302 42544 435520 42550
rect 436114 42490 436120 42660
rect 436172 42490 436178 42660
rect 436556 42608 436584 46694
rect 436680 46646 436708 46662
rect 436680 46640 436732 46646
rect 436680 46582 436732 46588
rect 436680 43272 436708 46582
rect 436664 43102 436670 43272
rect 436722 43102 436728 43272
rect 437329 42660 437357 46698
rect 437523 46650 437551 46673
rect 437523 46644 437575 46650
rect 437523 46586 437575 46592
rect 437752 46590 437780 46600
rect 438525 46594 438553 46602
rect 437523 43220 437551 46586
rect 437752 46584 437804 46590
rect 437752 46526 437804 46532
rect 438525 46588 438577 46594
rect 438525 46530 438577 46536
rect 437424 43214 437642 43220
rect 437424 43156 437642 43162
rect 436498 42602 436716 42608
rect 436498 42544 436716 42550
rect 437310 42490 437316 42660
rect 437368 42490 437374 42660
rect 437752 42608 437780 46526
rect 437876 46478 437904 46497
rect 437876 46472 437928 46478
rect 437876 46414 437928 46420
rect 437876 43272 437904 46414
rect 437860 43102 437866 43272
rect 437918 43102 437924 43272
rect 438525 42660 438553 46530
rect 438719 46482 438747 46497
rect 438695 46476 438747 46482
rect 438695 46418 438747 46424
rect 438719 43220 438747 46418
rect 438948 46422 438976 46497
rect 438948 46416 439000 46422
rect 438948 46358 439000 46364
rect 438620 43214 438838 43220
rect 438620 43156 438838 43162
rect 437694 42602 437912 42608
rect 437694 42544 437912 42550
rect 438506 42490 438512 42660
rect 438564 42490 438570 42660
rect 438948 42608 438976 46358
rect 439072 46310 439100 46497
rect 439721 46426 439749 46497
rect 439721 46420 439773 46426
rect 439721 46362 439773 46368
rect 439072 46304 439124 46310
rect 439072 46246 439124 46252
rect 439072 43272 439100 46246
rect 439056 43102 439062 43272
rect 439114 43102 439120 43272
rect 439721 42660 439749 46362
rect 439915 46314 439943 46497
rect 439915 46308 439967 46314
rect 439915 46250 439967 46256
rect 440144 46254 440172 46497
rect 439915 43220 439943 46250
rect 440144 46248 440196 46254
rect 440144 46190 440196 46196
rect 439816 43214 440034 43220
rect 439816 43156 440034 43162
rect 438890 42602 439108 42608
rect 438890 42544 439108 42550
rect 439702 42490 439708 42660
rect 439760 42490 439766 42660
rect 440144 42608 440172 46190
rect 440268 46142 440296 46497
rect 440917 46258 440945 46497
rect 440917 46252 440969 46258
rect 440917 46194 440969 46200
rect 440268 46136 440320 46142
rect 440268 46078 440320 46084
rect 440268 43272 440296 46078
rect 440422 43997 440795 44011
rect 440422 43937 440430 43997
rect 440787 43937 440795 43997
rect 440422 43925 440795 43937
rect 440252 43102 440258 43272
rect 440310 43102 440316 43272
rect 440422 42909 440795 42923
rect 440422 42849 440430 42909
rect 440787 42849 440795 42909
rect 440422 42837 440795 42849
rect 440917 42660 440945 46194
rect 441111 46146 441139 46497
rect 441111 46140 441163 46146
rect 441111 46082 441163 46088
rect 441340 46086 441368 46497
rect 441111 43220 441139 46082
rect 441340 46080 441392 46086
rect 441340 46022 441392 46028
rect 441012 43214 441230 43220
rect 441012 43156 441230 43162
rect 440086 42602 440304 42608
rect 440086 42544 440304 42550
rect 440898 42490 440904 42660
rect 440956 42490 440962 42660
rect 441340 42608 441368 46022
rect 441464 45974 441492 46497
rect 442113 46090 442141 46497
rect 442113 46084 442165 46090
rect 442113 46026 442165 46032
rect 441464 45968 441516 45974
rect 441464 45910 441516 45916
rect 441464 43272 441492 45910
rect 441618 43450 441991 43462
rect 441618 43390 441626 43450
rect 441983 43390 441991 43450
rect 441618 43376 441991 43390
rect 441448 43102 441454 43272
rect 441506 43102 441512 43272
rect 442113 42660 442141 46026
rect 442307 45978 442335 46497
rect 442307 45972 442359 45978
rect 442307 45914 442359 45920
rect 442536 45918 442564 46497
rect 442307 43220 442335 45914
rect 442536 45912 442588 45918
rect 442536 45854 442588 45860
rect 442208 43214 442426 43220
rect 442208 43156 442426 43162
rect 441282 42602 441500 42608
rect 441282 42544 441500 42550
rect 442094 42490 442100 42660
rect 442152 42490 442158 42660
rect 442536 42608 442564 45854
rect 442660 45806 442688 46497
rect 443309 45922 443337 46497
rect 443309 45916 443361 45922
rect 443309 45858 443361 45864
rect 442660 45800 442712 45806
rect 442660 45742 442712 45748
rect 442660 43272 442688 45742
rect 442644 43102 442650 43272
rect 442702 43102 442708 43272
rect 443309 42660 443337 45858
rect 443503 45810 443531 46497
rect 443503 45804 443555 45810
rect 443503 45746 443555 45752
rect 443732 45750 443760 46497
rect 443503 43220 443531 45746
rect 443732 45744 443784 45750
rect 443732 45686 443784 45692
rect 443404 43214 443622 43220
rect 443404 43156 443622 43162
rect 442478 42602 442696 42608
rect 442478 42544 442696 42550
rect 443290 42490 443296 42660
rect 443348 42490 443354 42660
rect 443732 42608 443760 45686
rect 443856 45638 443884 46497
rect 444505 45754 444533 46497
rect 444505 45748 444557 45754
rect 444505 45690 444557 45696
rect 443856 45632 443908 45638
rect 443856 45574 443908 45580
rect 443856 43272 443884 45574
rect 443840 43102 443846 43272
rect 443898 43102 443904 43272
rect 444505 42660 444533 45690
rect 444699 45642 444727 46497
rect 444699 45636 444751 45642
rect 444699 45578 444751 45584
rect 444928 45582 444956 46497
rect 444699 43220 444727 45578
rect 444928 45576 444980 45582
rect 444928 45518 444980 45524
rect 444600 43214 444818 43220
rect 444600 43156 444818 43162
rect 443674 42602 443892 42608
rect 443674 42544 443892 42550
rect 444486 42490 444492 42660
rect 444544 42490 444550 42660
rect 444928 42608 444956 45518
rect 445052 45470 445080 46497
rect 445701 45586 445729 46497
rect 445701 45580 445753 45586
rect 445701 45522 445753 45528
rect 445052 45464 445104 45470
rect 445052 45406 445104 45412
rect 445052 43272 445080 45406
rect 445036 43102 445042 43272
rect 445094 43102 445100 43272
rect 445701 42660 445729 45522
rect 445895 45474 445923 46497
rect 445895 45468 445947 45474
rect 445895 45410 445947 45416
rect 446124 45414 446152 46497
rect 445895 43220 445923 45410
rect 446124 45408 446176 45414
rect 446124 45350 446176 45356
rect 445796 43214 446014 43220
rect 445796 43156 446014 43162
rect 444870 42602 445088 42608
rect 444870 42544 445088 42550
rect 445682 42490 445688 42660
rect 445740 42490 445746 42660
rect 446124 42608 446152 45350
rect 446248 45302 446276 46497
rect 446897 45418 446925 46497
rect 446897 45412 446949 45418
rect 446897 45354 446949 45360
rect 446248 45296 446300 45302
rect 446248 45238 446300 45244
rect 446248 43272 446276 45238
rect 446232 43102 446238 43272
rect 446290 43102 446296 43272
rect 446897 42660 446925 45354
rect 447091 45306 447119 46497
rect 447091 45300 447143 45306
rect 447091 45242 447143 45248
rect 447320 45246 447348 46497
rect 447091 43220 447119 45242
rect 447320 45240 447372 45246
rect 447320 45182 447372 45188
rect 446992 43214 447210 43220
rect 446992 43156 447210 43162
rect 446066 42602 446284 42608
rect 446066 42544 446284 42550
rect 446878 42490 446884 42660
rect 446936 42490 446942 42660
rect 447320 42608 447348 45182
rect 447444 45134 447472 46497
rect 448093 45250 448121 46497
rect 448093 45244 448145 45250
rect 448093 45186 448145 45192
rect 447444 45128 447496 45134
rect 447444 45070 447496 45076
rect 447444 43272 447472 45070
rect 447428 43102 447434 43272
rect 447486 43102 447492 43272
rect 448093 42660 448121 45186
rect 448287 45138 448315 46497
rect 448287 45132 448339 45138
rect 448287 45074 448339 45080
rect 448516 45078 448544 46497
rect 448287 43220 448315 45074
rect 448516 45072 448568 45078
rect 448516 45014 448568 45020
rect 448188 43214 448406 43220
rect 448188 43156 448406 43162
rect 447262 42602 447480 42608
rect 447262 42544 447480 42550
rect 448074 42490 448080 42660
rect 448132 42490 448138 42660
rect 448516 42608 448544 45014
rect 448640 44966 448668 46497
rect 449289 45082 449317 46497
rect 449289 45076 449341 45082
rect 449289 45018 449341 45024
rect 448640 44960 448692 44966
rect 448640 44902 448692 44908
rect 448640 43272 448668 44902
rect 448624 43102 448630 43272
rect 448682 43102 448688 43272
rect 449289 42660 449317 45018
rect 449483 44970 449511 46497
rect 449483 44964 449535 44970
rect 449483 44906 449535 44912
rect 449712 44910 449740 46497
rect 449483 43220 449511 44906
rect 449712 44904 449764 44910
rect 449712 44846 449764 44852
rect 449384 43214 449602 43220
rect 449384 43156 449602 43162
rect 448458 42602 448676 42608
rect 448458 42544 448676 42550
rect 449270 42490 449276 42660
rect 449328 42490 449334 42660
rect 449712 42608 449740 44846
rect 449836 44798 449864 46497
rect 450485 44914 450513 46497
rect 450485 44908 450537 44914
rect 450485 44850 450537 44856
rect 449836 44792 449888 44798
rect 449836 44734 449888 44740
rect 449836 43272 449864 44734
rect 449820 43102 449826 43272
rect 449878 43102 449884 43272
rect 450485 42660 450513 44850
rect 450679 44802 450707 46497
rect 450655 44796 450707 44802
rect 450655 44738 450707 44744
rect 450679 43220 450707 44738
rect 450908 44742 450936 46497
rect 450908 44736 450960 44742
rect 450908 44678 450960 44684
rect 450580 43214 450798 43220
rect 450580 43156 450798 43162
rect 449654 42602 449872 42608
rect 449654 42544 449872 42550
rect 450466 42490 450472 42660
rect 450524 42490 450530 42660
rect 450908 42608 450936 44678
rect 451032 44630 451060 46497
rect 451681 44746 451709 46497
rect 451681 44740 451733 44746
rect 451681 44682 451733 44688
rect 451032 44624 451084 44630
rect 451032 44566 451084 44572
rect 451032 43272 451060 44566
rect 451016 43102 451022 43272
rect 451074 43102 451080 43272
rect 451681 42660 451709 44682
rect 451875 44634 451903 46497
rect 451875 44628 451927 44634
rect 451875 44570 451927 44576
rect 452104 44574 452132 46497
rect 451875 43220 451903 44570
rect 452104 44568 452156 44574
rect 452104 44510 452156 44516
rect 451776 43214 451994 43220
rect 451776 43156 451994 43162
rect 450850 42602 451068 42608
rect 450850 42544 451068 42550
rect 451662 42490 451668 42660
rect 451720 42490 451726 42660
rect 452104 42608 452132 44510
rect 452228 44462 452256 46497
rect 452877 44578 452905 46497
rect 452877 44572 452929 44578
rect 452877 44514 452929 44520
rect 452228 44456 452280 44462
rect 452228 44398 452280 44404
rect 452228 43272 452256 44398
rect 452212 43102 452218 43272
rect 452270 43102 452276 43272
rect 452877 42660 452905 44514
rect 453071 44466 453099 46497
rect 453047 44460 453099 44466
rect 453047 44402 453099 44408
rect 453071 43220 453099 44402
rect 453300 44350 453328 46497
rect 453300 44344 453352 44350
rect 453300 44286 453352 44292
rect 452972 43214 453190 43220
rect 452972 43156 453190 43162
rect 453300 42834 453328 44286
rect 453424 44238 453452 46497
rect 454073 44354 454101 46497
rect 454073 44348 454125 44354
rect 454073 44290 454125 44296
rect 453424 44232 453476 44238
rect 453424 44174 453476 44180
rect 453424 43272 453452 44174
rect 453408 43102 453414 43272
rect 453466 43102 453472 43272
rect 454073 42834 454101 44290
rect 454267 44242 454295 46497
rect 454267 44236 454319 44242
rect 454267 44178 454319 44184
rect 454267 43220 454295 44178
rect 454168 43214 454386 43220
rect 454168 43156 454386 43162
rect 453300 42806 453455 42834
rect 454073 42806 454228 42834
rect 453427 42660 453455 42806
rect 452046 42602 452264 42608
rect 452046 42544 452264 42550
rect 452858 42490 452864 42660
rect 452916 42490 452922 42660
rect 453410 42490 453416 42660
rect 453468 42490 453474 42660
rect 454200 42608 454228 42806
rect 454068 42602 454286 42608
rect 454068 42544 454286 42550
rect 147387 42375 147760 42384
rect 147387 42315 147395 42375
rect 147752 42315 147760 42375
rect 147387 42298 147760 42315
rect 441618 42368 441991 42377
rect 441618 42308 441626 42368
rect 441983 42308 441991 42368
rect 441618 42291 441991 42308
<< via2 >>
rect 417027 997507 417384 997567
rect 663637 997425 663994 997485
rect 168590 997178 168947 997238
rect 168590 996096 168947 996156
rect 169786 996637 170143 996697
rect 169786 995549 170143 995609
rect 417027 996425 417384 996485
rect 418223 996966 418580 997026
rect 418223 995878 418580 995938
rect 663637 996343 663994 996403
rect 664833 996884 665190 996944
rect 664833 995796 665190 995856
rect 40340 889384 40400 889741
rect 41422 889384 41482 889741
rect 40881 888188 40941 888545
rect 41969 888188 42029 888545
rect 676093 724496 676153 724853
rect 677175 724496 677235 724853
rect 675546 723300 675606 723657
rect 676634 723300 676694 723657
rect 40371 604610 40431 604967
rect 41453 604610 41513 604967
rect 40912 603414 40972 603771
rect 42000 603414 42060 603771
rect 676085 448095 676145 448452
rect 677167 448095 677227 448452
rect 675538 446899 675598 447256
rect 676626 446899 676686 447256
rect 40390 346959 40450 347316
rect 41472 346959 41532 347316
rect 40931 345763 40991 346120
rect 42019 345763 42079 346120
rect 146199 43944 146556 44004
rect 146199 42856 146556 42916
rect 147395 43397 147752 43457
rect 440430 43937 440787 43997
rect 440430 42849 440787 42909
rect 441626 43390 441983 43450
rect 147395 42315 147752 42375
rect 441626 42308 441983 42368
<< metal3 >>
rect 168581 997238 168954 997586
rect 168581 997178 168590 997238
rect 168947 997178 168954 997238
rect 168581 996156 168954 997178
rect 168581 996096 168590 996156
rect 168947 996096 168954 996156
rect 168581 996081 168954 996096
rect 169779 996697 170149 997586
rect 169779 996637 169786 996697
rect 170143 996637 170149 996697
rect 169779 995609 170149 996637
rect 417018 997567 417391 997915
rect 417018 997507 417027 997567
rect 417384 997507 417391 997567
rect 417018 996485 417391 997507
rect 417018 996425 417027 996485
rect 417384 996425 417391 996485
rect 417018 996410 417391 996425
rect 418216 997026 418586 997915
rect 418216 996966 418223 997026
rect 418580 996966 418586 997026
rect 418216 995938 418586 996966
rect 663628 997485 664001 997833
rect 663628 997425 663637 997485
rect 663994 997425 664001 997485
rect 663628 996403 664001 997425
rect 663628 996343 663637 996403
rect 663994 996343 664001 996403
rect 663628 996328 664001 996343
rect 664826 996944 665196 997833
rect 664826 996884 664833 996944
rect 665190 996884 665196 996944
rect 418216 995878 418223 995938
rect 418580 995878 418586 995938
rect 418216 995864 418586 995878
rect 664826 995856 665196 996884
rect 664826 995796 664833 995856
rect 665190 995796 665196 995856
rect 664826 995782 665196 995796
rect 169779 995549 169786 995609
rect 170143 995549 170149 995609
rect 169779 995535 170149 995549
rect 39992 889741 41497 889748
rect 39992 889384 40340 889741
rect 40400 889384 41422 889741
rect 41482 889384 41497 889741
rect 39992 889375 41497 889384
rect 39992 888545 42043 888551
rect 39992 888188 40881 888545
rect 40941 888188 41969 888545
rect 42029 888188 42043 888545
rect 39992 888181 42043 888188
rect 676078 724853 677583 724862
rect 676078 724496 676093 724853
rect 676153 724496 677175 724853
rect 677235 724496 677583 724853
rect 676078 724489 677583 724496
rect 675532 723657 677583 723664
rect 675532 723300 675546 723657
rect 675606 723300 676634 723657
rect 676694 723300 677583 723657
rect 675532 723294 677583 723300
rect 40023 604967 41528 604974
rect 40023 604610 40371 604967
rect 40431 604610 41453 604967
rect 41513 604610 41528 604967
rect 40023 604601 41528 604610
rect 40023 603771 42074 603777
rect 40023 603414 40912 603771
rect 40972 603414 42000 603771
rect 42060 603414 42074 603771
rect 40023 603407 42074 603414
rect 676070 448452 677575 448461
rect 676070 448095 676085 448452
rect 676145 448095 677167 448452
rect 677227 448095 677575 448452
rect 676070 448088 677575 448095
rect 675524 447256 677575 447263
rect 675524 446899 675538 447256
rect 675598 446899 676626 447256
rect 676686 446899 677575 447256
rect 675524 446893 677575 446899
rect 40042 347316 41547 347323
rect 40042 346959 40390 347316
rect 40450 346959 41472 347316
rect 41532 346959 41547 347316
rect 40042 346950 41547 346959
rect 40042 346120 42093 346126
rect 40042 345763 40931 346120
rect 40991 345763 42019 346120
rect 42079 345763 42093 346120
rect 40042 345756 42093 345763
rect 146193 44004 146563 44018
rect 146193 43944 146199 44004
rect 146556 43944 146563 44004
rect 146193 42916 146563 43944
rect 440424 43997 440794 44011
rect 440424 43937 440430 43997
rect 440787 43937 440794 43997
rect 146193 42856 146199 42916
rect 146556 42856 146563 42916
rect 146193 41967 146563 42856
rect 147388 43457 147761 43472
rect 147388 43397 147395 43457
rect 147752 43397 147761 43457
rect 147388 42375 147761 43397
rect 147388 42315 147395 42375
rect 147752 42315 147761 42375
rect 147388 41967 147761 42315
rect 440424 42909 440794 43937
rect 440424 42849 440430 42909
rect 440787 42849 440794 42909
rect 440424 41960 440794 42849
rect 441619 43450 441992 43465
rect 441619 43390 441626 43450
rect 441983 43390 441992 43450
rect 441619 42368 441992 43390
rect 441619 42308 441626 42368
rect 441983 42308 441992 42368
rect 441619 41960 441992 42308
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 434076 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_1
timestamp 1663859327
transform 1 0 429292 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_2
timestamp 1663859327
transform 1 0 430488 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_3
timestamp 1663859327
transform 1 0 431684 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_4
timestamp 1663859327
transform 1 0 432880 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_5
timestamp 1663859327
transform 1 0 441252 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_6
timestamp 1663859327
transform 1 0 435272 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_7
timestamp 1663859327
transform 1 0 436468 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_8
timestamp 1663859327
transform 1 0 437664 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_9
timestamp 1663859327
transform 1 0 438860 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_10
timestamp 1663859327
transform 1 0 440056 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_11
timestamp 1663859327
transform 1 0 442448 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_12
timestamp 1663859327
transform 1 0 444840 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_13
timestamp 1663859327
transform 1 0 443644 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_14
timestamp 1663859327
transform 1 0 446036 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_15
timestamp 1663859327
transform 1 0 447232 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_16
timestamp 1663859327
transform 1 0 448428 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_17
timestamp 1663859327
transform 1 0 450820 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_18
timestamp 1663859327
transform 1 0 449624 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_19
timestamp 1663859327
transform 1 0 452016 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_20
timestamp 1663859327
transform 1 0 453212 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_21
timestamp 1663859327
transform 1 0 133892 0 1 42337
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_22
timestamp 1663859327
transform 1 0 429292 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_23
timestamp 1663859327
transform 1 0 135088 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_24
timestamp 1663859327
transform 1 0 133892 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_25
timestamp 1663859327
transform 1 0 137480 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_26
timestamp 1663859327
transform 1 0 136284 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_27
timestamp 1663859327
transform 1 0 138676 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_28
timestamp 1663859327
transform 1 0 141068 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_29
timestamp 1663859327
transform 1 0 139872 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_30
timestamp 1663859327
transform 1 0 142264 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_31
timestamp 1663859327
transform 1 0 144656 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_32
timestamp 1663859327
transform 1 0 143460 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_33
timestamp 1663859327
transform 1 0 147048 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_34
timestamp 1663859327
transform 1 0 145852 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_35
timestamp 1663859327
transform 1 0 149440 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_36
timestamp 1663859327
transform 1 0 148244 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_37
timestamp 1663859327
transform 1 0 150636 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_38
timestamp 1663859327
transform 1 0 154224 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_39
timestamp 1663859327
transform 1 0 151832 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_40
timestamp 1663859327
transform 1 0 153028 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_41
timestamp 1663859327
transform 1 0 156616 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_42
timestamp 1663859327
transform 1 0 155420 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_43
timestamp 1663859327
transform 1 0 157812 0 1 43425
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_44
timestamp 1663859327
transform 0 1 41504 -1 0 338169
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_45
timestamp 1663859327
transform 0 1 41504 -1 0 340561
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_46
timestamp 1663859327
transform 0 1 41504 -1 0 339365
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_47
timestamp 1663859327
transform 0 1 41504 -1 0 341757
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_48
timestamp 1663859327
transform 0 1 41504 -1 0 344149
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_49
timestamp 1663859327
transform 0 1 41504 -1 0 342953
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_50
timestamp 1663859327
transform 0 1 41504 -1 0 345345
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_51
timestamp 1663859327
transform 0 1 41504 -1 0 346541
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_52
timestamp 1663859327
transform 0 1 41504 -1 0 348933
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_53
timestamp 1663859327
transform 0 1 41504 -1 0 347737
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_54
timestamp 1663859327
transform 0 1 41504 -1 0 351325
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_55
timestamp 1663859327
transform 0 1 41504 -1 0 352521
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_56
timestamp 1663859327
transform 0 1 41504 -1 0 336973
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_57
timestamp 1663859327
transform 0 1 41504 -1 0 335777
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_58
timestamp 1663859327
transform 0 1 41482 -1 0 610102
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_59
timestamp 1663859327
transform 0 1 41482 -1 0 607710
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_60
timestamp 1663859327
transform 0 1 41482 -1 0 608906
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_61
timestamp 1663859327
transform 0 1 41482 -1 0 605318
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_62
timestamp 1663859327
transform 0 1 41482 -1 0 606514
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_63
timestamp 1663859327
transform 0 1 41482 -1 0 602926
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_64
timestamp 1663859327
transform 0 1 41482 -1 0 604122
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_65
timestamp 1663859327
transform 0 1 41482 -1 0 600534
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_66
timestamp 1663859327
transform 0 1 41482 -1 0 601730
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_67
timestamp 1663859327
transform 0 1 41482 -1 0 599338
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_68
timestamp 1663859327
transform 0 1 41482 -1 0 598142
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_69
timestamp 1663859327
transform 0 1 41457 -1 0 891348
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_70
timestamp 1663859327
transform 0 1 41457 -1 0 890152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_71
timestamp 1663859327
transform 0 1 41457 -1 0 888956
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_72
timestamp 1663859327
transform 0 1 41457 -1 0 887760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_73
timestamp 1663859327
transform 0 1 41457 -1 0 886564
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_74
timestamp 1663859327
transform -1 0 170518 0 -1 996127
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_75
timestamp 1663859327
transform -1 0 168126 0 -1 996127
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_76
timestamp 1663859327
transform -1 0 169322 0 -1 996127
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_77
timestamp 1663859327
transform -1 0 417762 0 -1 996452
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_78
timestamp 1663859327
transform -1 0 665555 0 -1 996370
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_79
timestamp 1663859327
transform -1 0 666751 0 -1 996370
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_80
timestamp 1663859327
transform -1 0 664359 0 -1 996370
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_81
timestamp 1663859327
transform -1 0 663163 0 -1 996370
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_82
timestamp 1663859327
transform 0 -1 676117 -1 0 726392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_83
timestamp 1663859327
transform 0 -1 676117 -1 0 725196
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_84
timestamp 1663859327
transform 0 -1 676117 -1 0 727588
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_85
timestamp 1663859327
transform 0 -1 676117 -1 0 722804
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_86
timestamp 1663859327
transform 0 -1 676117 -1 0 721608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_87
timestamp 1663859327
transform 0 -1 676117 -1 0 724000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_88
timestamp 1663859327
transform 0 -1 676117 -1 0 453564
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_89
timestamp 1663859327
transform 0 -1 676117 -1 0 451172
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_90
timestamp 1663859327
transform 0 -1 676117 -1 0 452368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_91
timestamp 1663859327
transform 0 -1 676117 -1 0 448780
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_92
timestamp 1663859327
transform 0 -1 676117 -1 0 449976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_93
timestamp 1663859327
transform 0 -1 676117 -1 0 446388
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_94
timestamp 1663859327
transform 0 -1 676117 -1 0 447584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_95
timestamp 1663859327
transform 0 -1 676117 -1 0 445192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_96
timestamp 1663859327
transform 0 -1 676117 -1 0 442800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_97
timestamp 1663859327
transform 0 -1 676117 -1 0 443996
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_98
timestamp 1663859327
transform 0 -1 676117 -1 0 440408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_99
timestamp 1663859327
transform 0 -1 676117 -1 0 441604
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_100
timestamp 1663859327
transform 0 1 41504 -1 0 350129
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 0 -1 41504 -1 0 351325
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_1
timestamp 1663859327
transform -1 0 134996 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_2
timestamp 1663859327
transform 1 0 153028 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_3
timestamp 1663859327
transform -1 0 154132 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_4
timestamp 1663859327
transform 1 0 155420 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_5
timestamp 1663859327
transform -1 0 156524 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_6
timestamp 1663859327
transform 1 0 156616 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_7
timestamp 1663859327
transform -1 0 157720 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_8
timestamp 1663859327
transform -1 0 158916 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_9
timestamp 1663859327
transform -1 0 158916 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_10
timestamp 1663859327
transform -1 0 417762 0 -1 997540
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_11
timestamp 1663859327
transform 1 0 416658 0 1 996452
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_12
timestamp 1663859327
transform 0 -1 677205 1 0 439304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_13
timestamp 1663859327
transform 0 1 676117 -1 0 440408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_14
timestamp 1663859327
transform 0 1 676117 -1 0 448780
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_15
timestamp 1663859327
transform 0 -1 677205 1 0 447676
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_16
timestamp 1663859327
transform 0 1 676117 -1 0 452368
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_17
timestamp 1663859327
transform 0 -1 677205 1 0 451264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_18
timestamp 1663859327
transform 0 1 676117 -1 0 449976
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_19
timestamp 1663859327
transform 0 -1 677205 1 0 448872
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_20
timestamp 1663859327
transform 0 1 676117 -1 0 451172
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_21
timestamp 1663859327
transform 0 -1 677205 1 0 450068
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_22
timestamp 1663859327
transform 0 1 676117 -1 0 453564
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_23
timestamp 1663859327
transform 0 -1 677205 1 0 452460
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_24
timestamp 1663859327
transform 0 -1 677205 1 0 720504
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_25
timestamp 1663859327
transform 0 1 676117 -1 0 721608
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_26
timestamp 1663859327
transform 0 1 676117 -1 0 722804
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_27
timestamp 1663859327
transform 0 -1 677205 1 0 721700
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_28
timestamp 1663859327
transform 0 1 676117 -1 0 724000
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_29
timestamp 1663859327
transform 0 -1 677205 1 0 722896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_30
timestamp 1663859327
transform 0 1 676117 -1 0 725196
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_31
timestamp 1663859327
transform 0 -1 677205 1 0 724092
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_32
timestamp 1663859327
transform 0 1 676117 -1 0 727588
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_33
timestamp 1663859327
transform 0 -1 677205 1 0 726484
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_34
timestamp 1663859327
transform 0 1 676117 -1 0 446388
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_35
timestamp 1663859327
transform 0 -1 677205 1 0 445284
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_36
timestamp 1663859327
transform 0 1 676117 -1 0 447584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_37
timestamp 1663859327
transform 0 -1 677205 1 0 446480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_38
timestamp 1663859327
transform -1 0 169322 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_39
timestamp 1663859327
transform -1 0 168126 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_40
timestamp 1663859327
transform 0 -1 677205 1 0 725288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_41
timestamp 1663859327
transform 0 1 676117 -1 0 726392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_42
timestamp 1663859327
transform -1 0 170518 0 1 996127
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_43
timestamp 1663859327
transform 1 0 169414 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_44
timestamp 1663859327
transform 1 0 168218 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_45
timestamp 1663859327
transform 1 0 167022 0 -1 997215
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_46
timestamp 1663859327
transform 0 1 676117 -1 0 441604
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_47
timestamp 1663859327
transform 0 -1 677205 1 0 440500
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_48
timestamp 1663859327
transform 0 -1 677205 1 0 441696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_49
timestamp 1663859327
transform 0 1 676117 -1 0 442800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_50
timestamp 1663859327
transform 0 -1 677205 1 0 442892
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_51
timestamp 1663859327
transform 0 1 676117 -1 0 443996
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_52
timestamp 1663859327
transform 0 -1 677205 1 0 444088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_53
timestamp 1663859327
transform 0 1 676117 -1 0 445192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_54
timestamp 1663859327
transform 1 0 151832 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_55
timestamp 1663859327
transform -1 0 152936 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_56
timestamp 1663859327
transform 1 0 150636 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_57
timestamp 1663859327
transform -1 0 151740 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_58
timestamp 1663859327
transform 1 0 149440 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_59
timestamp 1663859327
transform -1 0 150544 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_60
timestamp 1663859327
transform 1 0 148244 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_61
timestamp 1663859327
transform -1 0 149348 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_62
timestamp 1663859327
transform 1 0 147048 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_63
timestamp 1663859327
transform -1 0 148152 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_64
timestamp 1663859327
transform 1 0 145852 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_65
timestamp 1663859327
transform -1 0 146956 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_66
timestamp 1663859327
transform -1 0 145760 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_67
timestamp 1663859327
transform 1 0 144656 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_68
timestamp 1663859327
transform 1 0 143460 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_69
timestamp 1663859327
transform -1 0 144564 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_70
timestamp 1663859327
transform 1 0 142264 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_71
timestamp 1663859327
transform -1 0 143368 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_72
timestamp 1663859327
transform 1 0 141068 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_73
timestamp 1663859327
transform -1 0 142172 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_74
timestamp 1663859327
transform 1 0 139872 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_75
timestamp 1663859327
transform -1 0 140976 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_76
timestamp 1663859327
transform 1 0 138676 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_77
timestamp 1663859327
transform -1 0 139780 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_78
timestamp 1663859327
transform -1 0 138584 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_79
timestamp 1663859327
transform 1 0 137480 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_80
timestamp 1663859327
transform 1 0 136284 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_81
timestamp 1663859327
transform -1 0 137388 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_82
timestamp 1663859327
transform 1 0 135088 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_83
timestamp 1663859327
transform -1 0 136192 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_84
timestamp 1663859327
transform -1 0 155328 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_85
timestamp 1663859327
transform 1 0 154224 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_86
timestamp 1663859327
transform -1 0 430396 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_88
timestamp 1663859327
transform -1 0 431592 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_89
timestamp 1663859327
transform 1 0 430488 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_90
timestamp 1663859327
transform 1 0 431684 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_91
timestamp 1663859327
transform -1 0 432788 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_92
timestamp 1663859327
transform -1 0 433984 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_93
timestamp 1663859327
transform 1 0 432880 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_94
timestamp 1663859327
transform -1 0 435180 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_95
timestamp 1663859327
transform 1 0 434076 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_96
timestamp 1663859327
transform 1 0 435272 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_97
timestamp 1663859327
transform 1 0 436468 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_98
timestamp 1663859327
transform -1 0 436376 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_99
timestamp 1663859327
transform -1 0 437572 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_100
timestamp 1663859327
transform 1 0 437664 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_101
timestamp 1663859327
transform 1 0 438860 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_102
timestamp 1663859327
transform 1 0 440056 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_103
timestamp 1663859327
transform -1 0 438768 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_104
timestamp 1663859327
transform -1 0 439964 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_105
timestamp 1663859327
transform -1 0 441160 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_106
timestamp 1663859327
transform -1 0 442356 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_107
timestamp 1663859327
transform 1 0 441252 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_108
timestamp 1663859327
transform -1 0 443552 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_109
timestamp 1663859327
transform 1 0 442448 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_110
timestamp 1663859327
transform 1 0 443644 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_111
timestamp 1663859327
transform -1 0 444748 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_112
timestamp 1663859327
transform 1 0 444840 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_113
timestamp 1663859327
transform -1 0 445944 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_114
timestamp 1663859327
transform 1 0 446036 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_115
timestamp 1663859327
transform -1 0 447140 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_116
timestamp 1663859327
transform 1 0 447232 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_117
timestamp 1663859327
transform -1 0 448336 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_118
timestamp 1663859327
transform -1 0 449532 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_119
timestamp 1663859327
transform 1 0 448428 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_120
timestamp 1663859327
transform -1 0 450728 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_121
timestamp 1663859327
transform 1 0 449624 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_122
timestamp 1663859327
transform 1 0 450820 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_123
timestamp 1663859327
transform -1 0 451924 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_124
timestamp 1663859327
transform 1 0 452016 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_125
timestamp 1663859327
transform -1 0 454316 0 1 42337
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_126
timestamp 1663859327
transform -1 0 453120 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_127
timestamp 1663859327
transform -1 0 454316 0 -1 43425
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_128
timestamp 1663859327
transform 0 -1 41504 -1 0 335777
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_129
timestamp 1663859327
transform 0 1 40416 1 0 334673
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_130
timestamp 1663859327
transform 0 -1 41504 -1 0 336973
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_131
timestamp 1663859327
transform 0 1 40416 1 0 335869
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_132
timestamp 1663859327
transform 0 -1 41504 -1 0 338169
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_133
timestamp 1663859327
transform 0 1 40416 1 0 337065
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_134
timestamp 1663859327
transform 0 -1 41504 -1 0 341757
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_135
timestamp 1663859327
transform 0 1 40416 1 0 340653
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_136
timestamp 1663859327
transform 0 -1 41504 -1 0 340561
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_137
timestamp 1663859327
transform 0 1 40416 1 0 339457
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_138
timestamp 1663859327
transform 0 1 40416 1 0 338261
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_139
timestamp 1663859327
transform 0 -1 41504 -1 0 339365
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_140
timestamp 1663859327
transform 0 1 40416 1 0 343045
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_141
timestamp 1663859327
transform 0 -1 41504 -1 0 344149
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_142
timestamp 1663859327
transform 0 1 40416 1 0 341849
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_143
timestamp 1663859327
transform 0 -1 41504 -1 0 342953
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_144
timestamp 1663859327
transform 0 -1 41504 -1 0 347737
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_145
timestamp 1663859327
transform 0 1 40416 1 0 346633
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_146
timestamp 1663859327
transform 0 1 40416 1 0 345437
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_147
timestamp 1663859327
transform 0 -1 41504 -1 0 346541
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_148
timestamp 1663859327
transform 0 1 40416 1 0 344241
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_149
timestamp 1663859327
transform 0 -1 41504 -1 0 345345
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_151
timestamp 1663859327
transform 0 1 40416 1 0 350221
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_152
timestamp 1663859327
transform 0 -1 41504 -1 0 350129
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_153
timestamp 1663859327
transform 0 1 40416 1 0 349025
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_154
timestamp 1663859327
transform 0 1 40416 1 0 347829
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_155
timestamp 1663859327
transform 0 -1 41504 -1 0 348933
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_156
timestamp 1663859327
transform 0 -1 41504 -1 0 352521
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_157
timestamp 1663859327
transform 0 1 40416 1 0 351417
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_158
timestamp 1663859327
transform 0 1 40394 1 0 608998
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_159
timestamp 1663859327
transform 0 -1 41482 -1 0 610102
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_160
timestamp 1663859327
transform 0 1 40394 1 0 607802
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_161
timestamp 1663859327
transform 0 -1 41482 -1 0 608906
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_162
timestamp 1663859327
transform 0 1 40394 1 0 606606
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_163
timestamp 1663859327
transform 0 -1 41482 -1 0 607710
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_164
timestamp 1663859327
transform 0 1 40394 1 0 605410
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_165
timestamp 1663859327
transform 0 -1 41482 -1 0 606514
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_166
timestamp 1663859327
transform 0 1 40394 1 0 604214
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_167
timestamp 1663859327
transform 0 -1 41482 -1 0 605318
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_168
timestamp 1663859327
transform 0 1 40394 1 0 603018
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_169
timestamp 1663859327
transform 0 -1 41482 -1 0 604122
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_170
timestamp 1663859327
transform 0 1 40394 1 0 601822
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_171
timestamp 1663859327
transform 0 -1 41482 -1 0 602926
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_172
timestamp 1663859327
transform 0 -1 41482 -1 0 601730
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_173
timestamp 1663859327
transform 0 1 40394 1 0 600626
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_174
timestamp 1663859327
transform 0 1 40394 1 0 599430
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_175
timestamp 1663859327
transform 0 -1 41482 -1 0 600534
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_176
timestamp 1663859327
transform 0 1 40394 1 0 598234
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_177
timestamp 1663859327
transform 0 -1 41482 -1 0 599338
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_178
timestamp 1663859327
transform 0 1 40394 1 0 597038
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_179
timestamp 1663859327
transform 0 -1 41482 -1 0 598142
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_180
timestamp 1663859327
transform 1 0 662059 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_181
timestamp 1663859327
transform 0 -1 41457 -1 0 890152
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_182
timestamp 1663859327
transform 0 1 40369 1 0 889048
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_183
timestamp 1663859327
transform 0 -1 41457 -1 0 891348
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_184
timestamp 1663859327
transform 0 1 40369 1 0 890244
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_185
timestamp 1663859327
transform 0 1 40369 1 0 885460
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_186
timestamp 1663859327
transform 0 -1 41457 -1 0 886564
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_187
timestamp 1663859327
transform 0 1 40369 1 0 886656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_188
timestamp 1663859327
transform 0 -1 41457 -1 0 887760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_189
timestamp 1663859327
transform 0 -1 41457 -1 0 888956
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_190
timestamp 1663859327
transform 0 1 40369 1 0 887852
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_191
timestamp 1663859327
transform 1 0 663255 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_192
timestamp 1663859327
transform 1 0 664451 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_193
timestamp 1663859327
transform 1 0 665647 0 1 996370
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_194
timestamp 1663859327
transform -1 0 663163 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_195
timestamp 1663859327
transform -1 0 664359 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_196
timestamp 1663859327
transform -1 0 665555 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_197
timestamp 1663859327
transform -1 0 666751 0 -1 997458
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 0 -1 676117 -1 0 722896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1663859327
transform 0 -1 677205 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1663859327
transform -1 0 434076 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1663859327
transform -1 0 133892 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1663859327
transform -1 0 155420 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1663859327
transform -1 0 155420 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1663859327
transform -1 0 153028 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1663859327
transform -1 0 153028 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1663859327
transform -1 0 156616 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1663859327
transform -1 0 156616 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1663859327
transform -1 0 157812 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1663859327
transform -1 0 157812 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1663859327
transform -1 0 159008 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1663859327
transform -1 0 159008 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1663859327
transform 1 0 417762 0 1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1663859327
transform 1 0 417762 0 -1 997540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1663859327
transform 0 1 676117 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1663859327
transform 0 -1 677205 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1663859327
transform 0 1 676117 -1 0 451264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1663859327
transform 0 -1 677205 -1 0 451264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1663859327
transform 0 1 676117 -1 0 448872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1663859327
transform 0 -1 677205 -1 0 448872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1663859327
transform 0 1 676117 -1 0 450068
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1663859327
transform 0 -1 677205 -1 0 450068
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1663859327
transform 0 1 676117 -1 0 452460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1663859327
transform 0 -1 677205 -1 0 452460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1663859327
transform 0 -1 677205 -1 0 453656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1663859327
transform 0 1 676117 -1 0 453656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1663859327
transform 0 1 676117 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1663859327
transform 0 1 676117 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1663859327
transform 0 1 676117 -1 0 722896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1663859327
transform 0 -1 677205 -1 0 722896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1663859327
transform 0 1 676117 -1 0 724092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1663859327
transform 0 -1 677205 -1 0 724092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1663859327
transform 0 1 676117 -1 0 725288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1663859327
transform 0 -1 677205 -1 0 725288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1663859327
transform 0 1 676117 -1 0 727680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1663859327
transform 0 -1 677205 -1 0 727680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1663859327
transform 0 1 676117 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1663859327
transform 0 -1 677205 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1663859327
transform 1 0 416566 0 1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1663859327
transform 1 0 417762 0 -1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1663859327
transform -1 0 169414 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1663859327
transform -1 0 169414 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1663859327
transform 0 -1 677205 -1 0 726484
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1663859327
transform 0 1 676117 -1 0 726484
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1663859327
transform -1 0 170610 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1663859327
transform -1 0 170610 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1663859327
transform -1 0 168218 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1663859327
transform -1 0 168218 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1663859327
transform -1 0 167022 0 1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1663859327
transform -1 0 168218 0 -1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1663859327
transform 0 -1 676117 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1663859327
transform 0 1 676117 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1663859327
transform 0 -1 677205 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1663859327
transform 0 1 676117 -1 0 440500
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1663859327
transform 0 -1 677205 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1663859327
transform 0 1 676117 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1663859327
transform 0 -1 677205 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1663859327
transform 0 1 676117 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1663859327
transform 0 -1 677205 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1663859327
transform 0 1 676117 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1663859327
transform 0 -1 677205 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1663859327
transform 0 1 676117 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1663859327
transform -1 0 151832 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1663859327
transform -1 0 151832 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1663859327
transform -1 0 150636 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1663859327
transform -1 0 150636 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1663859327
transform -1 0 149440 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1663859327
transform -1 0 149440 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1663859327
transform -1 0 148244 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1663859327
transform -1 0 148244 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1663859327
transform -1 0 147048 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1663859327
transform -1 0 147048 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1663859327
transform -1 0 145852 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1663859327
transform -1 0 145852 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1663859327
transform -1 0 144656 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1663859327
transform -1 0 144656 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1663859327
transform -1 0 143460 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1663859327
transform -1 0 143460 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1663859327
transform -1 0 142264 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1663859327
transform -1 0 142264 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1663859327
transform -1 0 141068 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1663859327
transform -1 0 141068 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1663859327
transform -1 0 139872 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1663859327
transform -1 0 139872 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1663859327
transform -1 0 138676 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1663859327
transform -1 0 138676 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1663859327
transform -1 0 137480 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1663859327
transform -1 0 137480 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1663859327
transform -1 0 136284 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1663859327
transform -1 0 136284 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1663859327
transform -1 0 135088 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1663859327
transform -1 0 135088 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1663859327
transform -1 0 154224 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1663859327
transform -1 0 154224 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1663859327
transform -1 0 429292 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1663859327
transform -1 0 429292 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1663859327
transform -1 0 430488 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1663859327
transform -1 0 430488 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1663859327
transform -1 0 431684 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1663859327
transform -1 0 431684 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1663859327
transform -1 0 434076 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1663859327
transform -1 0 434076 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1663859327
transform -1 0 432880 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1663859327
transform -1 0 432880 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1663859327
transform -1 0 435272 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1663859327
transform -1 0 436468 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1663859327
transform -1 0 437664 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1663859327
transform -1 0 435272 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1663859327
transform -1 0 436468 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1663859327
transform -1 0 437664 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1663859327
transform -1 0 438860 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1663859327
transform -1 0 440056 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1663859327
transform -1 0 438860 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1663859327
transform -1 0 440056 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1663859327
transform -1 0 441252 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1663859327
transform -1 0 441252 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1663859327
transform -1 0 442448 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1663859327
transform -1 0 442448 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1663859327
transform -1 0 443644 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1663859327
transform -1 0 443644 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1663859327
transform -1 0 444840 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1663859327
transform -1 0 444840 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1663859327
transform -1 0 446036 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1663859327
transform -1 0 446036 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1663859327
transform -1 0 447232 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1663859327
transform -1 0 447232 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1663859327
transform -1 0 448428 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1663859327
transform -1 0 448428 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1663859327
transform -1 0 449624 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1663859327
transform -1 0 449624 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1663859327
transform -1 0 450820 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1663859327
transform -1 0 450820 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1663859327
transform -1 0 452016 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1663859327
transform -1 0 453212 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1663859327
transform -1 0 454408 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1663859327
transform -1 0 452016 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1663859327
transform -1 0 453212 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1663859327
transform -1 0 454408 0 -1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1663859327
transform 0 -1 41504 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1663859327
transform 0 1 41504 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1663859327
transform 0 -1 41504 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1663859327
transform 0 1 40416 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1663859327
transform 0 -1 41504 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1663859327
transform 0 1 40416 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1663859327
transform 0 1 40416 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1663859327
transform 0 -1 41504 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1663859327
transform 0 1 40416 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1663859327
transform 0 -1 41504 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1663859327
transform 0 1 40416 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1663859327
transform 0 -1 41504 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1663859327
transform 0 -1 41504 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1663859327
transform 0 1 40416 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1663859327
transform 0 -1 41504 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1663859327
transform 0 1 40416 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1663859327
transform 0 -1 41504 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1663859327
transform 0 1 40416 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1663859327
transform 0 -1 41504 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1663859327
transform 0 1 40416 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1663859327
transform 0 -1 41504 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1663859327
transform 0 1 40416 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1663859327
transform 0 1 41504 -1 0 349025
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1663859327
transform 0 1 40416 -1 0 350221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1663859327
transform 0 -1 41504 -1 0 349025
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1663859327
transform 0 1 40416 -1 0 349025
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1663859327
transform 0 1 40416 -1 0 347829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1663859327
transform 0 -1 41504 -1 0 347829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1663859327
transform 0 1 40416 -1 0 352613
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1663859327
transform 0 -1 41504 -1 0 352613
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1663859327
transform 0 -1 41504 -1 0 351417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1663859327
transform 0 1 40416 -1 0 351417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1663859327
transform 0 1 40394 -1 0 610194
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1663859327
transform 0 -1 41482 -1 0 610194
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1663859327
transform 0 1 40394 -1 0 608998
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1663859327
transform 0 -1 41482 -1 0 608998
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1663859327
transform 0 1 40394 -1 0 607802
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1663859327
transform 0 -1 41482 -1 0 607802
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1663859327
transform 0 1 40394 -1 0 606606
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1663859327
transform 0 -1 41482 -1 0 606606
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1663859327
transform 0 1 40394 -1 0 605410
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1663859327
transform 0 -1 41482 -1 0 605410
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1663859327
transform 0 1 40394 -1 0 604214
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1663859327
transform 0 -1 41482 -1 0 604214
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1663859327
transform 0 1 40394 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1663859327
transform 0 -1 41482 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1663859327
transform 0 -1 41482 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1663859327
transform 0 1 40394 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1663859327
transform 0 1 40394 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1663859327
transform 0 -1 41482 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1663859327
transform 0 1 40394 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1663859327
transform 0 1 40394 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1663859327
transform 0 -1 41482 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1663859327
transform 0 -1 41482 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1663859327
transform 0 1 40394 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1663859327
transform 0 -1 41482 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1663859327
transform 0 1 40369 -1 0 890244
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1663859327
transform 0 -1 41457 -1 0 890244
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1663859327
transform 0 -1 41457 -1 0 891440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1663859327
transform 0 1 40369 -1 0 891440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1663859327
transform 0 -1 41457 -1 0 885460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1663859327
transform 0 1 40369 -1 0 885460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1663859327
transform 0 -1 41457 -1 0 886656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1663859327
transform 0 1 40369 -1 0 886656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1663859327
transform 0 1 40369 -1 0 887852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1663859327
transform 0 -1 41457 -1 0 887852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1663859327
transform 0 1 40369 -1 0 889048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1663859327
transform 0 -1 41457 -1 0 889048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1663859327
transform 1 0 661967 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1663859327
transform 1 0 663163 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1663859327
transform 1 0 664359 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1663859327
transform 1 0 665555 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1663859327
transform 1 0 661967 0 -1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1663859327
transform 1 0 663163 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1663859327
transform 1 0 664359 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1663859327
transform 1 0 665555 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1663859327
transform 1 0 666751 0 1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1663859327
transform 1 0 666751 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1663859327
transform -1 0 430488 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1663859327
transform -1 0 431684 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1663859327
transform -1 0 432880 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1663859327
transform -1 0 441252 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1663859327
transform -1 0 435272 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1663859327
transform -1 0 436468 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_224
timestamp 1663859327
transform -1 0 437664 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_225
timestamp 1663859327
transform -1 0 438860 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_226
timestamp 1663859327
transform -1 0 440056 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_227
timestamp 1663859327
transform -1 0 442448 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_228
timestamp 1663859327
transform -1 0 444840 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_229
timestamp 1663859327
transform -1 0 443644 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_230
timestamp 1663859327
transform -1 0 446036 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_231
timestamp 1663859327
transform -1 0 447232 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_232
timestamp 1663859327
transform -1 0 448428 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_233
timestamp 1663859327
transform -1 0 450820 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_234
timestamp 1663859327
transform -1 0 449624 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_235
timestamp 1663859327
transform -1 0 453212 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_236
timestamp 1663859327
transform -1 0 452016 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_237
timestamp 1663859327
transform -1 0 454408 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_238
timestamp 1663859327
transform -1 0 133892 0 1 42337
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_239
timestamp 1663859327
transform -1 0 429292 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_240
timestamp 1663859327
transform -1 0 135088 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_241
timestamp 1663859327
transform -1 0 133892 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_242
timestamp 1663859327
transform -1 0 136284 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_243
timestamp 1663859327
transform -1 0 137480 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_244
timestamp 1663859327
transform -1 0 138676 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_245
timestamp 1663859327
transform -1 0 141068 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_246
timestamp 1663859327
transform -1 0 139872 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_247
timestamp 1663859327
transform -1 0 142264 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_248
timestamp 1663859327
transform -1 0 144656 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_249
timestamp 1663859327
transform -1 0 143460 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_250
timestamp 1663859327
transform -1 0 145852 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_251
timestamp 1663859327
transform -1 0 147048 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_252
timestamp 1663859327
transform -1 0 149440 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_253
timestamp 1663859327
transform -1 0 148244 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_254
timestamp 1663859327
transform -1 0 150636 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_255
timestamp 1663859327
transform -1 0 154224 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_256
timestamp 1663859327
transform -1 0 151832 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_257
timestamp 1663859327
transform -1 0 153028 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_258
timestamp 1663859327
transform -1 0 156616 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_259
timestamp 1663859327
transform -1 0 155420 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_260
timestamp 1663859327
transform -1 0 157812 0 1 43425
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_261
timestamp 1663859327
transform 0 -1 677205 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_262
timestamp 1663859327
transform 0 -1 676117 -1 0 439304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_263
timestamp 1663859327
transform 0 -1 676117 -1 0 442892
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_264
timestamp 1663859327
transform 0 -1 676117 -1 0 441696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_265
timestamp 1663859327
transform 0 -1 676117 -1 0 444088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_266
timestamp 1663859327
transform 0 -1 676117 -1 0 446480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_267
timestamp 1663859327
transform 0 -1 676117 -1 0 445284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_268
timestamp 1663859327
transform 0 -1 676117 -1 0 448872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_269
timestamp 1663859327
transform 0 -1 676117 -1 0 447676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_270
timestamp 1663859327
transform 0 -1 676117 -1 0 451264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_271
timestamp 1663859327
transform 0 -1 676117 -1 0 450068
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_272
timestamp 1663859327
transform 0 -1 677205 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_273
timestamp 1663859327
transform 0 -1 676117 -1 0 453656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_274
timestamp 1663859327
transform 0 -1 676117 -1 0 720504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_275
timestamp 1663859327
transform 0 -1 676117 -1 0 721700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_276
timestamp 1663859327
transform 0 -1 676117 -1 0 726484
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_277
timestamp 1663859327
transform 0 -1 676117 -1 0 724092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_278
timestamp 1663859327
transform 0 -1 676117 -1 0 725288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_279
timestamp 1663859327
transform 0 -1 676117 -1 0 727680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_280
timestamp 1663859327
transform 1 0 661967 0 -1 997458
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_281
timestamp 1663859327
transform 1 0 663163 0 -1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_282
timestamp 1663859327
transform 1 0 665555 0 -1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_283
timestamp 1663859327
transform 1 0 664359 0 -1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_284
timestamp 1663859327
transform 1 0 666751 0 -1 996370
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_285
timestamp 1663859327
transform 1 0 416566 0 -1 997540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_286
timestamp 1663859327
transform 1 0 416566 0 -1 996452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_287
timestamp 1663859327
transform -1 0 167022 0 -1 997215
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_288
timestamp 1663859327
transform -1 0 167022 0 -1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_289
timestamp 1663859327
transform -1 0 169414 0 -1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_290
timestamp 1663859327
transform -1 0 170610 0 -1 996127
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_291
timestamp 1663859327
transform 0 1 41457 -1 0 885460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_292
timestamp 1663859327
transform 0 1 41457 -1 0 886656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_293
timestamp 1663859327
transform 0 1 41457 -1 0 887852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_294
timestamp 1663859327
transform 0 1 41457 -1 0 889048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_295
timestamp 1663859327
transform 0 1 41457 -1 0 891440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_296
timestamp 1663859327
transform 0 1 41457 -1 0 890244
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_297
timestamp 1663859327
transform 0 1 41482 -1 0 597038
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_298
timestamp 1663859327
transform 0 1 41482 -1 0 599430
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_299
timestamp 1663859327
transform 0 1 41482 -1 0 598234
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_300
timestamp 1663859327
transform 0 1 41482 -1 0 600626
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_301
timestamp 1663859327
transform 0 1 41482 -1 0 603018
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_302
timestamp 1663859327
transform 0 1 41482 -1 0 601822
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_303
timestamp 1663859327
transform 0 1 41482 -1 0 605410
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_304
timestamp 1663859327
transform 0 1 41482 -1 0 604214
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_305
timestamp 1663859327
transform 0 1 41482 -1 0 607802
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_306
timestamp 1663859327
transform 0 1 41482 -1 0 606606
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_307
timestamp 1663859327
transform 0 1 41482 -1 0 610194
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_308
timestamp 1663859327
transform 0 1 41482 -1 0 608998
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_309
timestamp 1663859327
transform 0 1 40416 -1 0 334673
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_310
timestamp 1663859327
transform 0 1 41504 -1 0 335869
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_311
timestamp 1663859327
transform 0 1 41504 -1 0 338261
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_312
timestamp 1663859327
transform 0 1 41504 -1 0 337065
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_313
timestamp 1663859327
transform 0 1 41504 -1 0 339457
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_314
timestamp 1663859327
transform 0 1 41504 -1 0 340653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_315
timestamp 1663859327
transform 0 1 41504 -1 0 343045
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_316
timestamp 1663859327
transform 0 1 41504 -1 0 341849
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_317
timestamp 1663859327
transform 0 1 41504 -1 0 344241
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_318
timestamp 1663859327
transform 0 1 41504 -1 0 345437
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_319
timestamp 1663859327
transform 0 1 41504 -1 0 347829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_320
timestamp 1663859327
transform 0 1 41504 -1 0 346633
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_321
timestamp 1663859327
transform 0 1 41504 -1 0 350221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_322
timestamp 1663859327
transform 0 1 41504 -1 0 351417
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_323
timestamp 1663859327
transform 0 -1 41504 -1 0 350221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_324
timestamp 1663859327
transform 0 1 41504 -1 0 352613
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_325
timestamp 1663859327
transform 0 -1 676117 -1 0 452460
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_326
timestamp 1663859327
transform -1 0 159008 0 1 43425
box -38 -48 130 592
<< labels >>
flabel metal3 418245 997803 418551 997897 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 417057 997799 417363 997893 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 169809 997465 170115 997559 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 168616 997465 168922 997559 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal1 171829 995401 172109 995429 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[12]
port 50 nsew signal input
flabel metal1 171030 994953 171310 994981 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[14]
port 53 nsew signal input
flabel metal1 171431 995177 171711 995205 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[13]
port 52 nsew signal input
flabel metal3 663663 997712 663969 997806 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 664858 997701 665164 997795 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 677462 446931 677552 447228 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 677464 448130 677554 448427 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal1 660323 995107 660632 995135 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[10]
port 4 nsew signal input
flabel metal3 677461 723330 677551 723627 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 677470 724527 677560 724824 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal1 660723 994883 661032 994911 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[9]
port 5 nsew signal input
flabel metal1 661123 994659 661432 994687 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[8]
port 6 nsew signal input
flabel metal1 673736 455568 673764 455855 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[4]
port 14 nsew signal input
flabel metal1 674380 728434 674408 728721 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[7]
port 9 nsew signal input
flabel metal1 674156 728034 674184 728321 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[6]
port 10 nsew signal input
flabel metal1 673960 455968 673988 456255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[5]
port 13 nsew signal input
flabel metal1 672840 453968 672868 454255 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[0]
port 18 nsew signal input
flabel metal1 673064 454368 673092 454655 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[1]
port 17 nsew signal input
flabel metal1 673288 454768 673316 455055 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[2]
port 16 nsew signal input
flabel metal1 673512 455168 673540 455455 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[3]
port 15 nsew signal input
flabel metal3 147432 41997 147738 42091 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 146226 41997 146532 42091 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal3 441644 41978 441950 42072 0 FreeSans 400 0 0 0 vssd
port 135 nsew ground input
flabel metal3 440451 41984 440757 42078 0 FreeSans 400 0 0 0 vccd
port 136 nsew power input
flabel metal1 131123 45048 131374 45076 0 FreeSans 288 0 0 0 mgmt_io_out_buf[27]
port 83 nsew signal output
flabel metal1 131523 44880 131774 44908 0 FreeSans 288 0 0 0 mgmt_io_out_buf[28]
port 84 nsew signal output
flabel metal1 131923 44712 132174 44740 0 FreeSans 288 0 0 0 mgmt_io_out_buf[29]
port 85 nsew signal output
flabel metal1 132323 44544 132574 44572 0 FreeSans 288 0 0 0 mgmt_io_out_buf[30]
port 86 nsew signal output
flabel metal1 44055 611295 44083 611556 0 FreeSans 288 90 0 0 mgmt_io_out_buf[20]
port 65 nsew signal output
flabel metal3 40074 346985 40164 347282 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 40076 345792 40166 346089 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 40053 604641 40143 604938 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 40053 603440 40143 603737 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal3 40025 889407 40115 889704 0 FreeSans 400 90 0 0 vssd
port 135 nsew ground input
flabel metal3 40022 888213 40112 888510 0 FreeSans 400 90 0 0 vccd
port 136 nsew power input
flabel metal1 42963 892082 42991 892317 0 FreeSans 288 90 0 0 mgmt_io_out_buf[15]
port 58 nsew signal output
flabel metal1 43187 891682 43215 891917 0 FreeSans 288 90 0 0 mgmt_io_out_buf[16]
port 59 nsew signal output
flabel metal1 43383 612495 43411 612756 0 FreeSans 288 90 0 0 mgmt_io_out_buf[17]
port 62 nsew signal output
flabel metal1 43607 612095 43635 612356 0 FreeSans 288 90 0 0 mgmt_io_out_buf[18]
port 63 nsew signal output
flabel metal1 43831 611695 43859 611956 0 FreeSans 288 90 0 0 mgmt_io_out_buf[19]
port 64 nsew signal output
flabel metal1 45371 353036 45399 353330 0 FreeSans 288 90 0 0 mgmt_io_out_buf[26]
port 77 nsew signal output
flabel metal1 45147 353436 45175 353730 0 FreeSans 288 90 0 0 mgmt_io_out_buf[25]
port 76 nsew signal output
flabel metal1 44923 353836 44951 354130 0 FreeSans 288 90 0 0 mgmt_io_out_buf[24]
port 75 nsew signal output
flabel metal1 44699 354236 44727 354530 0 FreeSans 288 90 0 0 mgmt_io_out_buf[23]
port 74 nsew signal output
flabel metal1 44503 610495 44531 610756 0 FreeSans 288 90 0 0 mgmt_io_out_buf[22]
port 67 nsew signal output
flabel metal1 44279 610895 44307 611156 0 FreeSans 288 90 0 0 mgmt_io_out_buf[21]
port 66 nsew signal output
flabel metal1 673624 228850 673652 229133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[14]
port 117 nsew signal input
flabel metal1 673764 236250 673792 236537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[4]
port 44 nsew signal output
flabel metal1 675360 233450 675388 233737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[11]
port 37 nsew signal output
flabel metal1 675108 233850 675136 234137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[10]
port 38 nsew signal output
flabel metal1 674884 234250 674912 234537 0 FreeSans 288 90 0 0 mgmt_io_in_buf[9]
port 39 nsew signal output
flabel metal1 674660 234650 674688 234937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[8]
port 40 nsew signal output
flabel metal1 674436 235050 674464 235337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[7]
port 41 nsew signal output
flabel metal1 674212 235450 674240 235737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[6]
port 42 nsew signal output
flabel metal1 673988 235850 674016 236137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[5]
port 43 nsew signal output
flabel metal1 672868 237850 672896 238137 0 FreeSans 288 90 0 0 mgmt_io_in_buf[0]
port 48 nsew signal output
flabel metal1 673092 237450 673120 237737 0 FreeSans 288 90 0 0 mgmt_io_in_buf[1]
port 47 nsew signal output
flabel metal1 673316 237050 673344 237337 0 FreeSans 288 90 0 0 mgmt_io_in_buf[2]
port 46 nsew signal output
flabel metal1 673540 236650 673568 236937 0 FreeSans 288 90 0 0 mgmt_io_in_buf[3]
port 45 nsew signal output
flabel metal1 670936 224050 670964 224333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[26]
port 105 nsew signal input
flabel metal1 671160 224450 671188 224733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[25]
port 106 nsew signal input
flabel metal1 671384 224850 671412 225133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[24]
port 107 nsew signal input
flabel metal1 671608 225250 671636 225533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[23]
port 108 nsew signal input
flabel metal1 671832 225650 671860 225933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[22]
port 109 nsew signal input
flabel metal1 672056 226050 672084 226333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[21]
port 110 nsew signal input
flabel metal1 672280 226450 672308 226733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[20]
port 111 nsew signal input
flabel metal1 672504 226850 672532 227133 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[19]
port 112 nsew signal input
flabel metal1 672728 227250 672756 227533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[18]
port 113 nsew signal input
flabel metal1 672952 227650 672980 227933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[17]
port 114 nsew signal input
flabel metal1 673176 228050 673204 228333 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[16]
port 115 nsew signal input
flabel metal1 673400 228450 673428 228733 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[15]
port 116 nsew signal input
flabel metal1 674296 230050 674324 230287 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[27]
port 101 nsew signal input
flabel metal1 674520 230450 674548 230687 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[28]
port 102 nsew signal input
flabel metal1 674744 230850 674772 231087 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[29]
port 103 nsew signal input
flabel metal1 674968 231250 674996 231487 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[30]
port 104 nsew signal input
flabel metal1 675192 231650 675220 231887 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[0]
port 96 nsew signal input
flabel metal1 675528 232050 675556 232287 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[2]
port 94 nsew signal input
flabel metal1 675360 231850 675388 232087 0 FreeSans 288 90 0 0 mgmt_io_oeb_unbuf[1]
port 95 nsew signal input
flabel metal1 673848 229250 673876 229533 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[13]
port 118 nsew signal input
flabel metal1 674072 229650 674100 229933 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[12]
port 119 nsew signal input
flabel metal1 416107 995247 416416 995275 0 FreeSans 288 0 0 0 mgmt_io_out_buf[11]
port 1 nsew signal output
flabel metal1 675080 231450 675108 231687 0 FreeSans 288 90 0 0 mgmt_io_in_buf[30]
port 97 nsew signal output
flabel metal1 674856 231050 674884 231287 0 FreeSans 288 90 0 0 mgmt_io_in_buf[29]
port 98 nsew signal output
flabel metal1 674632 230650 674660 230887 0 FreeSans 288 90 0 0 mgmt_io_in_buf[28]
port 99 nsew signal output
flabel metal1 674408 230250 674436 230487 0 FreeSans 288 90 0 0 mgmt_io_in_buf[27]
port 100 nsew signal output
flabel metal1 674184 229850 674212 230133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[12]
port 120 nsew signal output
flabel metal1 673960 229450 673988 229733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[13]
port 121 nsew signal output
flabel metal1 673736 229050 673764 229333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[14]
port 122 nsew signal output
flabel metal1 673512 228650 673540 228933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[15]
port 123 nsew signal output
flabel metal1 673288 228250 673316 228533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[16]
port 124 nsew signal output
flabel metal1 673064 227850 673092 228133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[17]
port 125 nsew signal output
flabel metal1 672840 227450 672868 227733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[18]
port 126 nsew signal output
flabel metal1 672616 227050 672644 227333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[19]
port 127 nsew signal output
flabel metal1 672392 226650 672420 226933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[20]
port 128 nsew signal output
flabel metal1 672168 226250 672196 226533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[21]
port 129 nsew signal output
flabel metal1 671944 225850 671972 226133 0 FreeSans 288 90 0 0 mgmt_io_in_buf[22]
port 130 nsew signal output
flabel metal1 671720 225450 671748 225733 0 FreeSans 288 90 0 0 mgmt_io_in_buf[23]
port 131 nsew signal output
flabel metal1 671496 225050 671524 225333 0 FreeSans 288 90 0 0 mgmt_io_in_buf[24]
port 132 nsew signal output
flabel metal1 671272 224650 671300 224933 0 FreeSans 288 90 0 0 mgmt_io_in_buf[25]
port 133 nsew signal output
flabel metal1 671048 224250 671076 224533 0 FreeSans 288 90 0 0 mgmt_io_in_buf[26]
port 134 nsew signal output
flabel metal1 672980 237650 673008 237937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[1]
port 26 nsew signal input
flabel metal1 673204 237250 673232 237537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[2]
port 27 nsew signal input
flabel metal1 672756 238050 672784 238337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[0]
port 25 nsew signal input
flabel metal1 673428 236850 673456 237137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[3]
port 28 nsew signal input
flabel metal1 673652 236450 673680 236737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[4]
port 29 nsew signal input
flabel metal1 673876 236050 673904 236337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[5]
port 30 nsew signal input
flabel metal1 674100 235650 674128 235937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[6]
port 31 nsew signal input
flabel metal1 674324 235250 674352 235537 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[7]
port 32 nsew signal input
flabel metal1 674548 234850 674576 235137 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[8]
port 33 nsew signal input
flabel metal1 674772 234450 674800 234737 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[9]
port 34 nsew signal input
flabel metal1 674996 234050 675024 234337 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[10]
port 35 nsew signal input
flabel metal1 675248 233650 675276 233937 0 FreeSans 288 90 0 0 mgmt_io_out_unbuf[11]
port 36 nsew signal input
flabel metal1 672728 453768 672756 454055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[0]
port 19 nsew signal output
flabel metal1 672952 454168 672980 454455 0 FreeSans 288 90 0 0 mgmt_io_out_buf[1]
port 20 nsew signal output
flabel metal1 673176 454568 673204 454855 0 FreeSans 288 90 0 0 mgmt_io_out_buf[2]
port 21 nsew signal output
flabel metal1 673400 454968 673428 455255 0 FreeSans 288 90 0 0 mgmt_io_out_buf[3]
port 22 nsew signal output
flabel metal1 673624 455368 673652 455655 0 FreeSans 288 90 0 0 mgmt_io_out_buf[4]
port 23 nsew signal output
flabel metal1 673848 455768 673876 456055 0 FreeSans 288 90 0 0 mgmt_io_out_buf[5]
port 24 nsew signal output
flabel metal1 674044 727834 674072 728121 0 FreeSans 288 90 0 0 mgmt_io_out_buf[6]
port 12 nsew signal output
flabel metal1 674268 728234 674296 728521 0 FreeSans 288 90 0 0 mgmt_io_out_buf[7]
port 11 nsew signal output
flabel metal1 660523 994995 660832 995023 0 FreeSans 288 0 0 0 mgmt_io_out_buf[10]
port 2 nsew signal output
flabel metal1 660923 994771 661232 994799 0 FreeSans 288 0 0 0 mgmt_io_out_buf[9]
port 3 nsew signal output
flabel metal1 661323 994547 661632 994575 0 FreeSans 288 0 0 0 mgmt_io_out_buf[8]
port 7 nsew signal output
flabel metal1 415907 995359 416216 995387 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[11]
port 0 nsew signal input
flabel metal1 171629 995289 171909 995317 0 FreeSans 288 0 0 0 mgmt_io_out_buf[12]
port 56 nsew signal output
flabel metal1 171231 995065 171511 995093 0 FreeSans 288 0 0 0 mgmt_io_out_buf[13]
port 55 nsew signal output
flabel metal1 170830 994841 171110 994869 0 FreeSans 288 0 0 0 mgmt_io_out_buf[14]
port 54 nsew signal output
flabel metal1 42851 892282 42879 892517 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[15]
port 61 nsew signal input
flabel metal1 43075 891882 43103 892117 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[16]
port 60 nsew signal input
flabel metal1 43271 612695 43299 612956 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[17]
port 73 nsew signal input
flabel metal1 43495 612295 43523 612556 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[18]
port 72 nsew signal input
flabel metal1 43719 611895 43747 612156 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[19]
port 71 nsew signal input
flabel metal1 43943 611495 43971 611756 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[20]
port 70 nsew signal input
flabel metal1 44167 611095 44195 611356 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[21]
port 69 nsew signal input
flabel metal1 44391 610695 44419 610956 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[22]
port 68 nsew signal input
flabel metal1 44587 354436 44615 354730 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[23]
port 81 nsew signal input
flabel metal1 44811 354036 44839 354330 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[24]
port 80 nsew signal input
flabel metal1 45035 353636 45063 353930 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[25]
port 79 nsew signal input
flabel metal1 45259 353236 45287 353530 0 FreeSans 288 90 0 0 mgmt_io_in_unbuf[26]
port 78 nsew signal input
flabel metal1 133151 44124 133402 44152 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[2]
port 93 nsew signal output
flabel metal1 132951 44236 133202 44264 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[1]
port 92 nsew signal output
flabel metal1 132751 44348 133002 44376 0 FreeSans 288 0 0 0 mgmt_io_oeb_buf[0]
port 91 nsew signal output
flabel metal1 132551 44460 132802 44488 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[30]
port 87 nsew signal input
flabel metal1 132151 44628 132402 44656 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[29]
port 88 nsew signal input
flabel metal1 131751 44796 132002 44824 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[28]
port 89 nsew signal input
flabel metal1 131351 44964 131602 44992 0 FreeSans 288 0 0 0 mgmt_io_in_unbuf[27]
port 90 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
