VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3165.000 BY 4767.000 ;
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.135 -2.000 725.415 4.000 ;
    END
  END clock_core
  PIN flash_clk_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.335 -2.000 1597.615 4.000 ;
    END
  END flash_clk_frame
  PIN flash_clk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.975 -2.000 1613.255 4.000 ;
    END
  END flash_clk_oeb
  PIN flash_csb_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.335 -2.000 1323.615 4.000 ;
    END
  END flash_csb_frame
  PIN flash_csb_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.975 -2.000 1339.255 4.000 ;
    END
  END flash_csb_oeb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.135 -2.000 1816.415 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.335 -2.000 1871.615 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.715 -2.000 1849.995 4.000 ;
    END
  END flash_io0_ieb
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.975 -2.000 1887.255 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.135 -2.000 2090.415 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.335 -2.000 2145.615 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ieb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2123.715 -2.000 2123.995 4.000 ;
    END
  END flash_io1_ieb
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.975 -2.000 2161.255 4.000 ;
    END
  END flash_io1_oeb
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.135 -2.000 2364.415 4.000 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2397.715 -2.000 2397.995 4.000 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2391.735 -2.000 2392.015 4.000 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.355 -2.000 2413.635 4.000 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.335 -2.000 2419.615 4.000 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.975 -2.000 2435.255 4.000 ;
    END
  END gpio_outenb_core
  PIN mprj_analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2545.395 3167.185 2545.995 ;
    END
  END mprj_analog_io[0]
  PIN mprj_analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.165 4763.000 2215.445 4768.935 ;
    END
  END mprj_analog_io[10]
  PIN mprj_analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.165 4763.000 1770.445 4768.935 ;
    END
  END mprj_analog_io[11]
  PIN mprj_analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.165 4763.000 1261.445 4768.935 ;
    END
  END mprj_analog_io[12]
  PIN mprj_analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.165 4763.000 1003.445 4768.935 ;
    END
  END mprj_analog_io[13]
  PIN mprj_analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.165 4763.000 746.445 4768.935 ;
    END
  END mprj_analog_io[14]
  PIN mprj_analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.165 4763.000 489.445 4768.935 ;
    END
  END mprj_analog_io[15]
  PIN mprj_analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.165 4763.000 232.445 4768.935 ;
    END
  END mprj_analog_io[16]
  PIN mprj_analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4623.005 4.000 4623.605 ;
    END
  END mprj_analog_io[17]
  PIN mprj_analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3774.005 4.000 3774.605 ;
    END
  END mprj_analog_io[18]
  PIN mprj_analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3558.005 4.000 3558.605 ;
    END
  END mprj_analog_io[19]
  PIN mprj_analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2771.395 3167.185 2771.995 ;
    END
  END mprj_analog_io[1]
  PIN mprj_analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3342.005 4.000 3342.605 ;
    END
  END mprj_analog_io[20]
  PIN mprj_analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3126.005 4.000 3126.605 ;
    END
  END mprj_analog_io[21]
  PIN mprj_analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2910.005 4.000 2910.605 ;
    END
  END mprj_analog_io[22]
  PIN mprj_analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2694.005 4.000 2694.605 ;
    END
  END mprj_analog_io[23]
  PIN mprj_analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2478.005 4.000 2478.605 ;
    END
  END mprj_analog_io[24]
  PIN mprj_analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1840.005 4.000 1840.605 ;
    END
  END mprj_analog_io[25]
  PIN mprj_analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1624.005 4.000 1624.605 ;
    END
  END mprj_analog_io[26]
  PIN mprj_analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1408.005 4.000 1408.605 ;
    END
  END mprj_analog_io[27]
  PIN mprj_analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1192.005 4.000 1192.605 ;
    END
  END mprj_analog_io[28]
  PIN mprj_analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2996.395 3167.185 2996.995 ;
    END
  END mprj_analog_io[2]
  PIN mprj_analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3222.395 3167.185 3222.995 ;
    END
  END mprj_analog_io[3]
  PIN mprj_analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3447.395 3167.185 3447.995 ;
    END
  END mprj_analog_io[4]
  PIN mprj_analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3672.395 3167.185 3672.995 ;
    END
  END mprj_analog_io[5]
  PIN mprj_analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4118.395 3167.185 4118.995 ;
    END
  END mprj_analog_io[6]
  PIN mprj_analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4564.395 3167.185 4564.995 ;
    END
  END mprj_analog_io[7]
  PIN mprj_analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2981.165 4763.000 2981.445 4768.935 ;
    END
  END mprj_analog_io[8]
  PIN mprj_analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.165 4763.000 2472.445 4768.935 ;
    END
  END mprj_analog_io[9]
  PIN mprj_io_analog_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 318.355 3167.185 318.955 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_en[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3234.355 3167.185 3234.955 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_en[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3459.355 3167.185 3459.955 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_en[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3684.355 3167.185 3684.955 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_en[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4130.355 3167.185 4130.955 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_en[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4576.355 3167.185 4576.955 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_en[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2969.205 4763.000 2969.485 4768.935 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_en[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.205 4763.000 2460.485 4768.935 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_en[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.205 4763.000 2203.485 4768.935 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_en[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.205 4763.000 1758.485 4768.935 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_en[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.205 4763.000 1249.485 4768.935 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 544.355 3167.185 544.955 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_en[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.205 4763.000 991.485 4768.935 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_en[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.205 4763.000 734.485 4768.935 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_en[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.205 4763.000 477.485 4768.935 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_en[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.205 4763.000 220.485 4768.935 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_en[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4611.045 4.000 4611.645 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_en[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3762.045 4.000 3762.645 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_en[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3546.045 4.000 3546.645 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_en[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3330.045 4.000 3330.645 ;
    END
  END mprj_io_analog_en[27]
  PIN mprj_io_analog_en[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3114.045 4.000 3114.645 ;
    END
  END mprj_io_analog_en[28]
  PIN mprj_io_analog_en[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2898.045 4.000 2898.645 ;
    END
  END mprj_io_analog_en[29]
  PIN mprj_io_analog_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 769.355 3167.185 769.955 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_en[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2682.045 4.000 2682.645 ;
    END
  END mprj_io_analog_en[30]
  PIN mprj_io_analog_en[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2466.045 4.000 2466.645 ;
    END
  END mprj_io_analog_en[31]
  PIN mprj_io_analog_en[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1828.045 4.000 1828.645 ;
    END
  END mprj_io_analog_en[32]
  PIN mprj_io_analog_en[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1612.045 4.000 1612.645 ;
    END
  END mprj_io_analog_en[33]
  PIN mprj_io_analog_en[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1396.045 4.000 1396.645 ;
    END
  END mprj_io_analog_en[34]
  PIN mprj_io_analog_en[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1180.045 4.000 1180.645 ;
    END
  END mprj_io_analog_en[35]
  PIN mprj_io_analog_en[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 964.045 4.000 964.645 ;
    END
  END mprj_io_analog_en[36]
  PIN mprj_io_analog_en[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 748.045 4.000 748.645 ;
    END
  END mprj_io_analog_en[37]
  PIN mprj_io_analog_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 995.355 3167.185 995.955 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_en[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1220.355 3167.185 1220.955 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_en[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1445.355 3167.185 1445.955 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_en[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1671.355 3167.185 1671.955 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_en[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2557.355 3167.185 2557.955 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_en[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2783.355 3167.185 2783.955 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_en[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3008.355 3167.185 3008.955 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 324.795 3167.185 325.395 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_pol[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3240.795 3167.185 3241.395 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_pol[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3465.795 3167.185 3466.395 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_pol[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3690.795 3167.185 3691.395 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_pol[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4136.795 3167.185 4137.395 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_pol[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4582.795 3167.185 4583.395 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_pol[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2962.765 4763.000 2963.045 4768.935 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_pol[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.765 4763.000 2454.045 4768.935 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_pol[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.765 4763.000 2197.045 4768.935 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_pol[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.765 4763.000 1752.045 4768.935 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_pol[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.765 4763.000 1243.045 4768.935 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_pol[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 550.795 3167.185 551.395 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_pol[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.765 4763.000 985.045 4768.935 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_pol[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.765 4763.000 728.045 4768.935 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_pol[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.765 4763.000 471.045 4768.935 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_pol[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.765 4763.000 214.045 4768.935 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_pol[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4604.605 4.000 4605.205 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_pol[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3755.605 4.000 3756.205 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_pol[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3539.605 4.000 3540.205 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_pol[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3323.605 4.000 3324.205 ;
    END
  END mprj_io_analog_pol[27]
  PIN mprj_io_analog_pol[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3107.605 4.000 3108.205 ;
    END
  END mprj_io_analog_pol[28]
  PIN mprj_io_analog_pol[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2891.605 4.000 2892.205 ;
    END
  END mprj_io_analog_pol[29]
  PIN mprj_io_analog_pol[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 775.795 3167.185 776.395 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_pol[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2675.605 4.000 2676.205 ;
    END
  END mprj_io_analog_pol[30]
  PIN mprj_io_analog_pol[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2459.605 4.000 2460.205 ;
    END
  END mprj_io_analog_pol[31]
  PIN mprj_io_analog_pol[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1821.605 4.000 1822.205 ;
    END
  END mprj_io_analog_pol[32]
  PIN mprj_io_analog_pol[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1605.605 4.000 1606.205 ;
    END
  END mprj_io_analog_pol[33]
  PIN mprj_io_analog_pol[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1389.605 4.000 1390.205 ;
    END
  END mprj_io_analog_pol[34]
  PIN mprj_io_analog_pol[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1173.605 4.000 1174.205 ;
    END
  END mprj_io_analog_pol[35]
  PIN mprj_io_analog_pol[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 957.605 4.000 958.205 ;
    END
  END mprj_io_analog_pol[36]
  PIN mprj_io_analog_pol[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 741.605 4.000 742.205 ;
    END
  END mprj_io_analog_pol[37]
  PIN mprj_io_analog_pol[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1001.795 3167.185 1002.395 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_pol[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1226.795 3167.185 1227.395 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_pol[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1451.795 3167.185 1452.395 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_pol[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1677.795 3167.185 1678.395 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_pol[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2563.795 3167.185 2564.395 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_pol[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2789.795 3167.185 2790.395 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_pol[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3014.795 3167.185 3015.395 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 339.975 3167.185 340.575 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_analog_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3255.975 3167.185 3256.575 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_analog_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3480.975 3167.185 3481.575 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_analog_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3705.975 3167.185 3706.575 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_analog_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4151.975 3167.185 4152.575 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_analog_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4597.975 3167.185 4598.575 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_analog_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2947.585 4763.000 2947.865 4768.935 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_analog_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.585 4763.000 2438.865 4768.935 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_analog_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2181.585 4763.000 2181.865 4768.935 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_analog_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.585 4763.000 1736.865 4768.935 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_analog_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.585 4763.000 1227.865 4768.935 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_analog_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 565.975 3167.185 566.575 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_analog_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.585 4763.000 969.865 4768.935 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_analog_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.585 4763.000 712.865 4768.935 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_analog_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.585 4763.000 455.865 4768.935 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_analog_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.585 4763.000 198.865 4768.935 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_analog_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4589.425 4.000 4590.025 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_analog_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3740.425 4.000 3741.025 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_analog_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3524.425 4.000 3525.025 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_analog_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3308.425 4.000 3309.025 ;
    END
  END mprj_io_analog_sel[27]
  PIN mprj_io_analog_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3092.425 4.000 3093.025 ;
    END
  END mprj_io_analog_sel[28]
  PIN mprj_io_analog_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2876.425 4.000 2877.025 ;
    END
  END mprj_io_analog_sel[29]
  PIN mprj_io_analog_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 790.975 3167.185 791.575 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_analog_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2660.425 4.000 2661.025 ;
    END
  END mprj_io_analog_sel[30]
  PIN mprj_io_analog_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2444.425 4.000 2445.025 ;
    END
  END mprj_io_analog_sel[31]
  PIN mprj_io_analog_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1806.425 4.000 1807.025 ;
    END
  END mprj_io_analog_sel[32]
  PIN mprj_io_analog_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1590.425 4.000 1591.025 ;
    END
  END mprj_io_analog_sel[33]
  PIN mprj_io_analog_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1374.425 4.000 1375.025 ;
    END
  END mprj_io_analog_sel[34]
  PIN mprj_io_analog_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1158.425 4.000 1159.025 ;
    END
  END mprj_io_analog_sel[35]
  PIN mprj_io_analog_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 942.425 4.000 943.025 ;
    END
  END mprj_io_analog_sel[36]
  PIN mprj_io_analog_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 726.425 4.000 727.025 ;
    END
  END mprj_io_analog_sel[37]
  PIN mprj_io_analog_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1016.975 3167.185 1017.575 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_analog_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1241.975 3167.185 1242.575 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_analog_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1466.975 3167.185 1467.575 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_analog_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1692.975 3167.185 1693.575 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_analog_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2578.975 3167.185 2579.575 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_analog_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2804.975 3167.185 2805.575 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_analog_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3029.975 3167.185 3030.575 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 321.575 3167.185 322.175 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1618.025 4.000 1618.625 ;
    END
  END mprj_io_dm[100]
  PIN mprj_io_dm[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1587.205 4.000 1587.805 ;
    END
  END mprj_io_dm[101]
  PIN mprj_io_dm[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1392.825 4.000 1393.425 ;
    END
  END mprj_io_dm[102]
  PIN mprj_io_dm[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1402.025 4.000 1402.625 ;
    END
  END mprj_io_dm[103]
  PIN mprj_io_dm[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1371.205 4.000 1371.805 ;
    END
  END mprj_io_dm[104]
  PIN mprj_io_dm[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1176.825 4.000 1177.425 ;
    END
  END mprj_io_dm[105]
  PIN mprj_io_dm[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1186.025 4.000 1186.625 ;
    END
  END mprj_io_dm[106]
  PIN mprj_io_dm[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1155.205 4.000 1155.805 ;
    END
  END mprj_io_dm[107]
  PIN mprj_io_dm[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 960.825 4.000 961.425 ;
    END
  END mprj_io_dm[108]
  PIN mprj_io_dm[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 970.025 4.000 970.625 ;
    END
  END mprj_io_dm[109]
  PIN mprj_io_dm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 989.375 3167.185 989.975 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 939.205 4.000 939.805 ;
    END
  END mprj_io_dm[110]
  PIN mprj_io_dm[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 744.825 4.000 745.425 ;
    END
  END mprj_io_dm[111]
  PIN mprj_io_dm[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 754.025 4.000 754.625 ;
    END
  END mprj_io_dm[112]
  PIN mprj_io_dm[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 723.205 4.000 723.805 ;
    END
  END mprj_io_dm[113]
  PIN mprj_io_dm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1020.195 3167.185 1020.795 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1223.575 3167.185 1224.175 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1214.375 3167.185 1214.975 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1245.195 3167.185 1245.795 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_dm[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1448.575 3167.185 1449.175 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1439.375 3167.185 1439.975 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1470.195 3167.185 1470.795 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_dm[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1674.575 3167.185 1675.175 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1665.375 3167.185 1665.975 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 312.375 3167.185 312.975 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1696.195 3167.185 1696.795 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_dm[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2560.575 3167.185 2561.175 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2551.375 3167.185 2551.975 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2582.195 3167.185 2582.795 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_dm[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2786.575 3167.185 2787.175 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2777.375 3167.185 2777.975 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2808.195 3167.185 2808.795 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_dm[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3011.575 3167.185 3012.175 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3002.375 3167.185 3002.975 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3033.195 3167.185 3033.795 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 343.195 3167.185 343.795 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_dm[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3237.575 3167.185 3238.175 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3228.375 3167.185 3228.975 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3259.195 3167.185 3259.795 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_dm[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3462.575 3167.185 3463.175 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3453.375 3167.185 3453.975 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3484.195 3167.185 3484.795 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_dm[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3687.575 3167.185 3688.175 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3678.375 3167.185 3678.975 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3709.195 3167.185 3709.795 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_dm[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4133.575 3167.185 4134.175 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 547.575 3167.185 548.175 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4124.375 3167.185 4124.975 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4155.195 3167.185 4155.795 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_dm[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4579.575 3167.185 4580.175 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4570.375 3167.185 4570.975 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4601.195 3167.185 4601.795 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_dm[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2965.985 4763.000 2966.265 4768.935 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2975.185 4763.000 2975.465 4768.935 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2944.365 4763.000 2944.645 4768.935 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_dm[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.985 4763.000 2457.265 4768.935 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.185 4763.000 2466.465 4768.935 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 538.375 3167.185 538.975 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2435.365 4763.000 2435.645 4768.935 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_dm[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.985 4763.000 2200.265 4768.935 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.185 4763.000 2209.465 4768.935 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.365 4763.000 2178.645 4768.935 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_dm[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.985 4763.000 1755.265 4768.935 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.185 4763.000 1764.465 4768.935 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.365 4763.000 1733.645 4768.935 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_dm[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.985 4763.000 1246.265 4768.935 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.185 4763.000 1255.465 4768.935 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.365 4763.000 1224.645 4768.935 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_dm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 569.195 3167.185 569.795 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_dm[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.985 4763.000 988.265 4768.935 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.185 4763.000 997.465 4768.935 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.365 4763.000 966.645 4768.935 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_dm[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.985 4763.000 731.265 4768.935 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.185 4763.000 740.465 4768.935 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.365 4763.000 709.645 4768.935 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_dm[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.985 4763.000 474.265 4768.935 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.185 4763.000 483.465 4768.935 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.365 4763.000 452.645 4768.935 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_dm[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.985 4763.000 217.265 4768.935 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 772.575 3167.185 773.175 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.185 4763.000 226.465 4768.935 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.365 4763.000 195.645 4768.935 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_dm[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4607.825 4.000 4608.425 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4617.025 4.000 4617.625 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4586.205 4.000 4586.805 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_dm[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3758.825 4.000 3759.425 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3768.025 4.000 3768.625 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3737.205 4.000 3737.805 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_dm[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3542.825 4.000 3543.425 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3552.025 4.000 3552.625 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 763.375 3167.185 763.975 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3521.205 4.000 3521.805 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_dm[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3326.825 4.000 3327.425 ;
    END
  END mprj_io_dm[81]
  PIN mprj_io_dm[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3336.025 4.000 3336.625 ;
    END
  END mprj_io_dm[82]
  PIN mprj_io_dm[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3305.205 4.000 3305.805 ;
    END
  END mprj_io_dm[83]
  PIN mprj_io_dm[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3110.825 4.000 3111.425 ;
    END
  END mprj_io_dm[84]
  PIN mprj_io_dm[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3120.025 4.000 3120.625 ;
    END
  END mprj_io_dm[85]
  PIN mprj_io_dm[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3089.205 4.000 3089.805 ;
    END
  END mprj_io_dm[86]
  PIN mprj_io_dm[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2894.825 4.000 2895.425 ;
    END
  END mprj_io_dm[87]
  PIN mprj_io_dm[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2904.025 4.000 2904.625 ;
    END
  END mprj_io_dm[88]
  PIN mprj_io_dm[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2873.205 4.000 2873.805 ;
    END
  END mprj_io_dm[89]
  PIN mprj_io_dm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 794.195 3167.185 794.795 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_dm[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2678.825 4.000 2679.425 ;
    END
  END mprj_io_dm[90]
  PIN mprj_io_dm[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2688.025 4.000 2688.625 ;
    END
  END mprj_io_dm[91]
  PIN mprj_io_dm[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2657.205 4.000 2657.805 ;
    END
  END mprj_io_dm[92]
  PIN mprj_io_dm[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2462.825 4.000 2463.425 ;
    END
  END mprj_io_dm[93]
  PIN mprj_io_dm[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2472.025 4.000 2472.625 ;
    END
  END mprj_io_dm[94]
  PIN mprj_io_dm[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2441.205 4.000 2441.805 ;
    END
  END mprj_io_dm[95]
  PIN mprj_io_dm[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1824.825 4.000 1825.425 ;
    END
  END mprj_io_dm[96]
  PIN mprj_io_dm[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1834.025 4.000 1834.625 ;
    END
  END mprj_io_dm[97]
  PIN mprj_io_dm[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1803.205 4.000 1803.805 ;
    END
  END mprj_io_dm[98]
  PIN mprj_io_dm[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1608.825 4.000 1609.425 ;
    END
  END mprj_io_dm[99]
  PIN mprj_io_dm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 998.575 3167.185 999.175 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 346.415 3167.185 347.015 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_holdover[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3262.415 3167.185 3263.015 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_holdover[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3487.415 3167.185 3488.015 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_holdover[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3712.415 3167.185 3713.015 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_holdover[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4158.415 3167.185 4159.015 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_holdover[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4604.415 3167.185 4605.015 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_holdover[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2941.145 4763.000 2941.425 4768.935 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_holdover[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2432.145 4763.000 2432.425 4768.935 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_holdover[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.145 4763.000 2175.425 4768.935 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_holdover[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.145 4763.000 1730.425 4768.935 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_holdover[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.145 4763.000 1221.425 4768.935 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_holdover[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 572.415 3167.185 573.015 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_holdover[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.145 4763.000 963.425 4768.935 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_holdover[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.145 4763.000 706.425 4768.935 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_holdover[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.145 4763.000 449.425 4768.935 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_holdover[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.145 4763.000 192.425 4768.935 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_holdover[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4582.985 4.000 4583.585 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_holdover[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3733.985 4.000 3734.585 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_holdover[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3517.985 4.000 3518.585 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_holdover[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3301.985 4.000 3302.585 ;
    END
  END mprj_io_holdover[27]
  PIN mprj_io_holdover[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3085.985 4.000 3086.585 ;
    END
  END mprj_io_holdover[28]
  PIN mprj_io_holdover[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2869.985 4.000 2870.585 ;
    END
  END mprj_io_holdover[29]
  PIN mprj_io_holdover[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 797.415 3167.185 798.015 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_holdover[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2653.985 4.000 2654.585 ;
    END
  END mprj_io_holdover[30]
  PIN mprj_io_holdover[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2437.985 4.000 2438.585 ;
    END
  END mprj_io_holdover[31]
  PIN mprj_io_holdover[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1799.985 4.000 1800.585 ;
    END
  END mprj_io_holdover[32]
  PIN mprj_io_holdover[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1583.985 4.000 1584.585 ;
    END
  END mprj_io_holdover[33]
  PIN mprj_io_holdover[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1367.985 4.000 1368.585 ;
    END
  END mprj_io_holdover[34]
  PIN mprj_io_holdover[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1151.985 4.000 1152.585 ;
    END
  END mprj_io_holdover[35]
  PIN mprj_io_holdover[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 935.985 4.000 936.585 ;
    END
  END mprj_io_holdover[36]
  PIN mprj_io_holdover[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 719.985 4.000 720.585 ;
    END
  END mprj_io_holdover[37]
  PIN mprj_io_holdover[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1023.415 3167.185 1024.015 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_holdover[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1248.415 3167.185 1249.015 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_holdover[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1473.415 3167.185 1474.015 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_holdover[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1699.415 3167.185 1700.015 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_holdover[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2585.415 3167.185 2586.015 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_holdover[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2811.415 3167.185 2812.015 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_holdover[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3036.415 3167.185 3037.015 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 361.595 3167.185 362.195 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3277.595 3167.185 3278.195 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3502.595 3167.185 3503.195 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3727.595 3167.185 3728.195 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4173.595 3167.185 4174.195 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4619.595 3167.185 4620.195 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2925.965 4763.000 2926.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.965 4763.000 2417.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.965 4763.000 2160.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.965 4763.000 1715.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.965 4763.000 1206.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 587.595 3167.185 588.195 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.965 4763.000 948.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.965 4763.000 691.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.965 4763.000 434.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.965 4763.000 177.245 4768.935 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4567.805 4.000 4568.405 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3718.805 4.000 3719.405 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3502.805 4.000 3503.405 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3286.805 4.000 3287.405 ;
    END
  END mprj_io_ib_mode_sel[27]
  PIN mprj_io_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3070.805 4.000 3071.405 ;
    END
  END mprj_io_ib_mode_sel[28]
  PIN mprj_io_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2854.805 4.000 2855.405 ;
    END
  END mprj_io_ib_mode_sel[29]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 812.595 3167.185 813.195 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2638.805 4.000 2639.405 ;
    END
  END mprj_io_ib_mode_sel[30]
  PIN mprj_io_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2422.805 4.000 2423.405 ;
    END
  END mprj_io_ib_mode_sel[31]
  PIN mprj_io_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1784.805 4.000 1785.405 ;
    END
  END mprj_io_ib_mode_sel[32]
  PIN mprj_io_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1568.805 4.000 1569.405 ;
    END
  END mprj_io_ib_mode_sel[33]
  PIN mprj_io_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1352.805 4.000 1353.405 ;
    END
  END mprj_io_ib_mode_sel[34]
  PIN mprj_io_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1136.805 4.000 1137.405 ;
    END
  END mprj_io_ib_mode_sel[35]
  PIN mprj_io_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 920.805 4.000 921.405 ;
    END
  END mprj_io_ib_mode_sel[36]
  PIN mprj_io_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 704.805 4.000 705.405 ;
    END
  END mprj_io_ib_mode_sel[37]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1038.595 3167.185 1039.195 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1263.595 3167.185 1264.195 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1488.595 3167.185 1489.195 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1714.595 3167.185 1715.195 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2600.595 3167.185 2601.195 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2826.595 3167.185 2827.195 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3051.595 3167.185 3052.195 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 293.975 3167.185 294.575 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3209.975 3167.185 3210.575 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3434.975 3167.185 3435.575 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3659.975 3167.185 3660.575 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4105.975 3167.185 4106.575 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4551.975 3167.185 4552.575 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2993.585 4763.000 2993.865 4768.935 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2484.585 4763.000 2484.865 4768.935 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.585 4763.000 2227.865 4768.935 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.585 4763.000 1782.865 4768.935 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.585 4763.000 1273.865 4768.935 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 519.975 3167.185 520.575 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.585 4763.000 1015.865 4768.935 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.585 4763.000 758.865 4768.935 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.585 4763.000 501.865 4768.935 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.585 4763.000 244.865 4768.935 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4635.425 4.000 4636.025 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3786.425 4.000 3787.025 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3570.425 4.000 3571.025 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3354.425 4.000 3355.025 ;
    END
  END mprj_io_in[27]
  PIN mprj_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3138.425 4.000 3139.025 ;
    END
  END mprj_io_in[28]
  PIN mprj_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2922.425 4.000 2923.025 ;
    END
  END mprj_io_in[29]
  PIN mprj_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 744.975 3167.185 745.575 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2706.425 4.000 2707.025 ;
    END
  END mprj_io_in[30]
  PIN mprj_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2490.425 4.000 2491.025 ;
    END
  END mprj_io_in[31]
  PIN mprj_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1852.425 4.000 1853.025 ;
    END
  END mprj_io_in[32]
  PIN mprj_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1636.425 4.000 1637.025 ;
    END
  END mprj_io_in[33]
  PIN mprj_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1420.425 4.000 1421.025 ;
    END
  END mprj_io_in[34]
  PIN mprj_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1204.425 4.000 1205.025 ;
    END
  END mprj_io_in[35]
  PIN mprj_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 988.425 4.000 989.025 ;
    END
  END mprj_io_in[36]
  PIN mprj_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 772.425 4.000 773.025 ;
    END
  END mprj_io_in[37]
  PIN mprj_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 970.975 3167.185 971.575 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1195.975 3167.185 1196.575 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1420.975 3167.185 1421.575 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1646.975 3167.185 1647.575 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2532.975 3167.185 2533.575 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2758.975 3167.185 2759.575 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2983.975 3167.185 2984.575 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_inp_dis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 327.555 3167.185 328.155 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_inp_dis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3243.555 3167.185 3244.155 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_inp_dis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3468.555 3167.185 3469.155 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_inp_dis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3693.555 3167.185 3694.155 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_inp_dis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4139.555 3167.185 4140.155 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_inp_dis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4585.555 3167.185 4586.155 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_inp_dis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2960.005 4763.000 2960.285 4768.935 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_inp_dis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.005 4763.000 2451.285 4768.935 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_inp_dis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.005 4763.000 2194.285 4768.935 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_inp_dis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.005 4763.000 1749.285 4768.935 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_inp_dis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.005 4763.000 1240.285 4768.935 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_inp_dis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 553.555 3167.185 554.155 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_inp_dis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.005 4763.000 982.285 4768.935 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_inp_dis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.005 4763.000 725.285 4768.935 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_inp_dis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.005 4763.000 468.285 4768.935 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_inp_dis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.005 4763.000 211.285 4768.935 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_inp_dis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4601.845 4.000 4602.445 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_inp_dis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3752.845 4.000 3753.445 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_inp_dis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3536.845 4.000 3537.445 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_inp_dis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3320.845 4.000 3321.445 ;
    END
  END mprj_io_inp_dis[27]
  PIN mprj_io_inp_dis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3104.845 4.000 3105.445 ;
    END
  END mprj_io_inp_dis[28]
  PIN mprj_io_inp_dis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2888.845 4.000 2889.445 ;
    END
  END mprj_io_inp_dis[29]
  PIN mprj_io_inp_dis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 778.555 3167.185 779.155 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_inp_dis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2672.845 4.000 2673.445 ;
    END
  END mprj_io_inp_dis[30]
  PIN mprj_io_inp_dis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2456.845 4.000 2457.445 ;
    END
  END mprj_io_inp_dis[31]
  PIN mprj_io_inp_dis[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1818.845 4.000 1819.445 ;
    END
  END mprj_io_inp_dis[32]
  PIN mprj_io_inp_dis[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1602.845 4.000 1603.445 ;
    END
  END mprj_io_inp_dis[33]
  PIN mprj_io_inp_dis[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1386.845 4.000 1387.445 ;
    END
  END mprj_io_inp_dis[34]
  PIN mprj_io_inp_dis[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1170.845 4.000 1171.445 ;
    END
  END mprj_io_inp_dis[35]
  PIN mprj_io_inp_dis[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 954.845 4.000 955.445 ;
    END
  END mprj_io_inp_dis[36]
  PIN mprj_io_inp_dis[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 738.845 4.000 739.445 ;
    END
  END mprj_io_inp_dis[37]
  PIN mprj_io_inp_dis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1004.555 3167.185 1005.155 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_inp_dis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1229.555 3167.185 1230.155 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_inp_dis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1454.555 3167.185 1455.155 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_inp_dis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1680.555 3167.185 1681.155 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_inp_dis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2566.555 3167.185 2567.155 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_inp_dis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2792.555 3167.185 2793.155 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_inp_dis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3017.555 3167.185 3018.155 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 364.815 3167.185 365.415 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3280.815 3167.185 3281.415 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3505.815 3167.185 3506.415 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3730.815 3167.185 3731.415 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4176.815 3167.185 4177.415 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4622.815 3167.185 4623.415 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2922.745 4763.000 2923.025 4768.935 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.745 4763.000 2414.025 4768.935 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.745 4763.000 2157.025 4768.935 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.745 4763.000 1712.025 4768.935 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.745 4763.000 1203.025 4768.935 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 590.815 3167.185 591.415 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.745 4763.000 945.025 4768.935 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.745 4763.000 688.025 4768.935 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.745 4763.000 431.025 4768.935 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.745 4763.000 174.025 4768.935 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4564.585 4.000 4565.185 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3715.585 4.000 3716.185 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3499.585 4.000 3500.185 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3283.585 4.000 3284.185 ;
    END
  END mprj_io_oeb[27]
  PIN mprj_io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3067.585 4.000 3068.185 ;
    END
  END mprj_io_oeb[28]
  PIN mprj_io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2851.585 4.000 2852.185 ;
    END
  END mprj_io_oeb[29]
  PIN mprj_io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 815.815 3167.185 816.415 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2635.585 4.000 2636.185 ;
    END
  END mprj_io_oeb[30]
  PIN mprj_io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2419.585 4.000 2420.185 ;
    END
  END mprj_io_oeb[31]
  PIN mprj_io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1781.585 4.000 1782.185 ;
    END
  END mprj_io_oeb[32]
  PIN mprj_io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1565.585 4.000 1566.185 ;
    END
  END mprj_io_oeb[33]
  PIN mprj_io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1349.585 4.290 1350.185 ;
    END
  END mprj_io_oeb[34]
  PIN mprj_io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1133.585 4.000 1134.185 ;
    END
  END mprj_io_oeb[35]
  PIN mprj_io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 917.585 4.000 918.185 ;
    END
  END mprj_io_oeb[36]
  PIN mprj_io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 701.585 4.000 702.185 ;
    END
  END mprj_io_oeb[37]
  PIN mprj_io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1041.815 3167.185 1042.415 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1266.815 3167.185 1267.415 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1491.815 3167.185 1492.415 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1717.815 3167.185 1718.415 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2603.815 3167.185 2604.415 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2829.815 3167.185 2830.415 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3054.815 3167.185 3055.415 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_one[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 299.955 3167.185 300.555 ;
    END
  END mprj_io_one[0]
  PIN mprj_io_one[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3215.955 3167.185 3216.555 ;
    END
  END mprj_io_one[10]
  PIN mprj_io_one[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3440.955 3167.185 3441.555 ;
    END
  END mprj_io_one[11]
  PIN mprj_io_one[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3665.955 3167.185 3666.555 ;
    END
  END mprj_io_one[12]
  PIN mprj_io_one[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4111.955 3167.185 4112.555 ;
    END
  END mprj_io_one[13]
  PIN mprj_io_one[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4557.955 3167.185 4558.555 ;
    END
  END mprj_io_one[14]
  PIN mprj_io_one[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2987.605 4763.000 2987.885 4768.935 ;
    END
  END mprj_io_one[15]
  PIN mprj_io_one[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2478.605 4763.000 2478.885 4768.935 ;
    END
  END mprj_io_one[16]
  PIN mprj_io_one[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.605 4763.000 2221.885 4768.935 ;
    END
  END mprj_io_one[17]
  PIN mprj_io_one[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.605 4763.000 1776.885 4768.935 ;
    END
  END mprj_io_one[18]
  PIN mprj_io_one[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.605 4763.000 1267.885 4768.935 ;
    END
  END mprj_io_one[19]
  PIN mprj_io_one[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 525.955 3167.185 526.555 ;
    END
  END mprj_io_one[1]
  PIN mprj_io_one[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.605 4763.000 1009.885 4768.935 ;
    END
  END mprj_io_one[20]
  PIN mprj_io_one[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.605 4763.000 752.885 4768.935 ;
    END
  END mprj_io_one[21]
  PIN mprj_io_one[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.605 4763.000 495.885 4768.935 ;
    END
  END mprj_io_one[22]
  PIN mprj_io_one[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.605 4763.000 238.885 4768.935 ;
    END
  END mprj_io_one[23]
  PIN mprj_io_one[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4629.445 4.000 4630.045 ;
    END
  END mprj_io_one[24]
  PIN mprj_io_one[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3780.445 4.000 3781.045 ;
    END
  END mprj_io_one[25]
  PIN mprj_io_one[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3564.445 4.000 3565.045 ;
    END
  END mprj_io_one[26]
  PIN mprj_io_one[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3348.445 4.000 3349.045 ;
    END
  END mprj_io_one[27]
  PIN mprj_io_one[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3132.445 4.000 3133.045 ;
    END
  END mprj_io_one[28]
  PIN mprj_io_one[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2916.445 4.000 2917.045 ;
    END
  END mprj_io_one[29]
  PIN mprj_io_one[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 750.955 3167.185 751.555 ;
    END
  END mprj_io_one[2]
  PIN mprj_io_one[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2700.445 4.000 2701.045 ;
    END
  END mprj_io_one[30]
  PIN mprj_io_one[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2484.445 4.000 2485.045 ;
    END
  END mprj_io_one[31]
  PIN mprj_io_one[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1846.445 4.000 1847.045 ;
    END
  END mprj_io_one[32]
  PIN mprj_io_one[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1630.445 4.000 1631.045 ;
    END
  END mprj_io_one[33]
  PIN mprj_io_one[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1414.445 4.000 1415.045 ;
    END
  END mprj_io_one[34]
  PIN mprj_io_one[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1198.445 4.290 1199.045 ;
    END
  END mprj_io_one[35]
  PIN mprj_io_one[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 982.445 4.000 983.045 ;
    END
  END mprj_io_one[36]
  PIN mprj_io_one[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 766.445 4.000 767.045 ;
    END
  END mprj_io_one[37]
  PIN mprj_io_one[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 976.955 3167.185 977.555 ;
    END
  END mprj_io_one[3]
  PIN mprj_io_one[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1201.955 3167.185 1202.555 ;
    END
  END mprj_io_one[4]
  PIN mprj_io_one[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1426.955 3167.185 1427.555 ;
    END
  END mprj_io_one[5]
  PIN mprj_io_one[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1652.955 3167.185 1653.555 ;
    END
  END mprj_io_one[6]
  PIN mprj_io_one[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2538.955 3167.185 2539.555 ;
    END
  END mprj_io_one[7]
  PIN mprj_io_one[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2764.955 3167.185 2765.555 ;
    END
  END mprj_io_one[8]
  PIN mprj_io_one[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2989.955 3167.185 2990.555 ;
    END
  END mprj_io_one[9]
  PIN mprj_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 349.175 3167.185 349.775 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3265.175 3167.185 3265.775 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3490.175 3167.185 3490.775 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3715.175 3167.185 3715.775 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4161.175 3167.185 4161.775 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4607.175 3167.185 4607.775 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2938.385 4763.000 2938.665 4768.935 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.385 4763.000 2429.665 4768.935 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.385 4763.000 2172.665 4768.935 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.385 4763.000 1727.665 4768.935 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.385 4763.000 1218.665 4768.935 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 575.175 3167.185 575.775 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.385 4763.000 960.665 4768.935 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.385 4763.000 703.665 4768.935 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.385 4763.000 446.665 4768.935 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.385 4763.000 189.665 4768.935 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4580.225 4.000 4580.825 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3731.225 4.000 3731.825 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3515.225 4.000 3515.825 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3299.225 4.000 3299.825 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3083.225 4.000 3083.825 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2867.225 4.000 2867.825 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 800.175 3167.185 800.775 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2651.225 4.000 2651.825 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2435.225 4.000 2435.825 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1797.225 4.000 1797.825 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1581.225 4.000 1581.825 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1365.225 4.000 1365.825 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1149.225 4.000 1149.825 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 933.225 4.000 933.825 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 717.225 4.000 717.825 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1026.175 3167.185 1026.775 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1251.175 3167.185 1251.775 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1476.175 3167.185 1476.775 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1702.175 3167.185 1702.775 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2588.175 3167.185 2588.775 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2814.175 3167.185 2814.775 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3039.175 3167.185 3039.775 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 303.175 3167.185 303.775 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3219.175 3167.185 3219.775 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3444.175 3167.185 3444.775 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3669.175 3167.185 3669.775 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4115.175 3167.185 4115.775 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4561.175 3167.185 4561.775 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2984.385 4763.000 2984.665 4768.935 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.385 4763.000 2475.665 4768.935 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.385 4763.000 2218.665 4768.935 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.385 4763.000 1773.665 4768.935 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.385 4763.000 1264.665 4768.935 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 529.175 3167.185 529.775 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.385 4763.000 1006.665 4768.935 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.385 4763.000 749.665 4768.935 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.385 4763.000 492.665 4768.935 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.385 4763.000 235.665 4768.935 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4626.225 4.000 4626.825 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3777.225 4.000 3777.825 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3561.225 4.000 3561.825 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3345.225 4.000 3345.825 ;
    END
  END mprj_io_slow_sel[27]
  PIN mprj_io_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3129.225 4.000 3129.825 ;
    END
  END mprj_io_slow_sel[28]
  PIN mprj_io_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2913.225 4.000 2913.825 ;
    END
  END mprj_io_slow_sel[29]
  PIN mprj_io_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 754.175 3167.185 754.775 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2697.225 4.000 2697.825 ;
    END
  END mprj_io_slow_sel[30]
  PIN mprj_io_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2481.225 4.000 2481.825 ;
    END
  END mprj_io_slow_sel[31]
  PIN mprj_io_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1843.225 4.000 1843.825 ;
    END
  END mprj_io_slow_sel[32]
  PIN mprj_io_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1627.225 4.000 1627.825 ;
    END
  END mprj_io_slow_sel[33]
  PIN mprj_io_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1411.225 4.000 1411.825 ;
    END
  END mprj_io_slow_sel[34]
  PIN mprj_io_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1195.225 4.000 1195.825 ;
    END
  END mprj_io_slow_sel[35]
  PIN mprj_io_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 979.225 4.000 979.825 ;
    END
  END mprj_io_slow_sel[36]
  PIN mprj_io_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 763.225 4.000 763.825 ;
    END
  END mprj_io_slow_sel[37]
  PIN mprj_io_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 980.175 3167.185 980.775 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1205.175 3167.185 1205.775 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1430.175 3167.185 1430.775 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1656.175 3167.185 1656.775 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2542.175 3167.185 2542.775 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2768.175 3167.185 2768.775 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2993.175 3167.185 2993.775 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 358.375 3167.185 358.975 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3274.375 3167.185 3274.975 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3499.375 3167.185 3499.975 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3724.375 3167.185 3724.975 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4170.375 3167.185 4170.975 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 4616.375 3167.185 4616.975 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2929.185 4763.000 2929.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.185 4763.000 2420.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.185 4763.000 2163.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.185 4763.000 1718.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.185 4763.000 1209.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 584.375 3167.185 584.975 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.185 4763.000 951.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.185 4763.000 694.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.185 4763.000 437.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.185 4763.000 180.465 4768.935 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 4571.025 4.000 4571.625 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3722.025 4.000 3722.625 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3506.025 4.000 3506.625 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3290.025 4.000 3290.625 ;
    END
  END mprj_io_vtrip_sel[27]
  PIN mprj_io_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 3074.025 4.000 3074.625 ;
    END
  END mprj_io_vtrip_sel[28]
  PIN mprj_io_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2858.025 4.000 2858.625 ;
    END
  END mprj_io_vtrip_sel[29]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 809.375 3167.185 809.975 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2642.025 4.000 2642.625 ;
    END
  END mprj_io_vtrip_sel[30]
  PIN mprj_io_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 2426.025 4.000 2426.625 ;
    END
  END mprj_io_vtrip_sel[31]
  PIN mprj_io_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1788.025 4.000 1788.625 ;
    END
  END mprj_io_vtrip_sel[32]
  PIN mprj_io_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1572.025 4.000 1572.625 ;
    END
  END mprj_io_vtrip_sel[33]
  PIN mprj_io_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1356.025 4.000 1356.625 ;
    END
  END mprj_io_vtrip_sel[34]
  PIN mprj_io_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 1140.025 4.000 1140.625 ;
    END
  END mprj_io_vtrip_sel[35]
  PIN mprj_io_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 924.025 4.000 924.625 ;
    END
  END mprj_io_vtrip_sel[36]
  PIN mprj_io_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.185 708.025 4.000 708.625 ;
    END
  END mprj_io_vtrip_sel[37]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1035.375 3167.185 1035.975 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1260.375 3167.185 1260.975 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1485.375 3167.185 1485.975 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 1711.375 3167.185 1711.975 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2597.375 3167.185 2597.975 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 2823.375 3167.185 2823.975 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3161.000 3048.375 3167.185 3048.975 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN por_l
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.715 -2.000 758.995 4.000 ;
    END
  END por_l
  PIN porb_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.775 -2.000 1330.055 4.000 ;
    END
  END porb_h
  PIN rstb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.835 -10.525 497.115 4.000 ;
    END
  END rstb_h
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.920 0.000 15.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3147.180 0.000 3152.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 10.880 3165.000 20.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4739.560 3165.000 4749.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.515 10.640 73.515 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3086.585 10.640 3088.585 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.520 10.640 128.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.520 669.885 128.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.520 4596.300 128.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.520 10.640 228.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.520 669.885 228.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.520 4596.300 228.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.520 10.640 328.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.520 669.885 328.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.520 4596.300 328.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.520 10.640 428.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.520 669.885 428.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.520 4596.300 428.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.520 10.640 528.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.520 669.885 528.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.520 4596.300 528.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.520 10.640 628.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.520 669.885 628.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.520 4596.300 628.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.520 10.640 728.720 132.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.520 677.100 728.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.520 4603.350 728.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.520 10.640 828.720 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.520 669.885 828.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.520 4596.300 828.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.520 10.640 928.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.520 936.205 928.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.520 4596.300 928.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.520 10.640 1028.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.520 936.205 1028.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.520 4596.300 1028.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.520 10.640 1128.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.520 936.205 1128.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.520 4596.300 1128.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.520 10.640 1228.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.520 936.205 1228.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.520 4596.300 1228.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.520 10.640 1328.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.520 936.205 1328.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.520 4596.300 1328.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.520 10.640 1428.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.520 936.205 1428.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.520 4596.300 1428.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.520 10.640 1528.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.520 936.205 1528.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.520 4596.300 1528.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.520 10.640 1628.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.520 936.205 1628.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.520 4603.350 1628.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.520 10.640 1728.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.520 936.205 1728.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.520 4596.300 1728.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.520 10.640 1828.720 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.520 582.645 1828.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.520 936.205 1828.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.520 4596.300 1828.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.520 10.640 1928.720 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.520 582.645 1928.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.520 936.205 1928.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.520 4596.300 1928.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.520 10.640 2028.720 142.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.520 586.460 2028.720 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.520 936.205 2028.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.520 4596.300 2028.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2125.520 10.640 2128.720 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2125.520 582.645 2128.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2125.520 4596.300 2128.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.520 10.640 2228.720 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.520 582.645 2228.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.520 4596.300 2228.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.520 10.640 2328.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.520 4596.300 2328.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.520 10.640 2428.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.520 4596.300 2428.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.520 10.640 2528.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.520 4603.350 2528.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2625.520 10.640 2628.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2625.520 4596.300 2628.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2725.520 10.640 2728.720 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2725.520 735.325 2728.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2725.520 4596.300 2728.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2825.520 10.640 2828.720 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2825.520 735.325 2828.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2825.520 4596.300 2828.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2925.520 10.640 2928.720 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2925.520 735.325 2928.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2925.520 4596.300 2928.720 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3025.520 10.640 3028.720 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 3025.520 735.325 3028.720 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3025.520 4596.300 3028.720 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 190.280 3154.920 193.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 310.280 3154.920 313.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 430.280 3154.920 433.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 550.280 3154.920 553.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 670.280 3154.920 673.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 790.280 3154.920 793.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 910.280 3154.920 913.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1030.280 76.000 1033.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1150.280 76.000 1153.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1270.280 76.000 1273.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1390.280 76.000 1393.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1510.280 76.000 1513.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1630.280 76.000 1633.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1750.280 76.000 1753.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1870.280 76.000 1873.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1990.280 76.000 1993.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2110.280 76.000 2113.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2230.280 76.000 2233.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2350.280 76.000 2353.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2470.280 76.000 2473.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2590.280 76.000 2593.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2710.280 76.000 2713.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2830.280 76.000 2833.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2950.280 76.000 2953.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3070.280 76.000 3073.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3190.280 76.000 3193.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3310.280 76.000 3313.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3430.280 76.000 3433.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3550.280 76.000 3553.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3670.280 76.000 3673.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3790.280 76.000 3793.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3910.280 76.000 3913.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4030.280 76.000 4033.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4150.280 76.000 4153.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4270.280 76.000 4273.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4390.280 76.000 4393.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4510.280 76.000 4513.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4630.280 3154.920 4633.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1030.280 3154.920 1033.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1150.280 3154.920 1153.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1270.280 3154.920 1273.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1390.280 3154.920 1393.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1510.280 3154.920 1513.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1630.280 3154.920 1633.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1750.280 3154.920 1753.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1870.280 3154.920 1873.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1990.280 3154.920 1993.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2110.280 3154.920 2113.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2230.280 3154.920 2233.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2350.280 3154.920 2353.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2470.280 3154.920 2473.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2590.280 3154.920 2593.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2710.280 3154.920 2713.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2830.280 3154.920 2833.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2950.280 3154.920 2953.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3070.280 3154.920 3073.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3190.280 3154.920 3193.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3310.280 3154.920 3313.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3430.280 3154.920 3433.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3550.280 3154.920 3553.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3670.280 3154.920 3673.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3790.280 3154.920 3793.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3910.280 3154.920 3913.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4030.280 3154.920 4033.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4150.280 3154.920 4153.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4270.280 3154.920 4273.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4390.280 3154.920 4393.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4510.280 3154.920 4513.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 247.480 3154.920 252.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 367.480 3154.920 372.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 487.480 3154.920 492.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 607.480 3154.920 612.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 825.520 948.700 2238.320 958.700 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.920 0.000 27.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3135.180 0.000 3140.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.080 3165.000 44.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4716.360 3165.000 4726.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 815.480 3154.920 820.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 262.240 4596.300 263.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 562.240 4596.300 563.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.240 669.885 863.840 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.240 4596.300 863.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1162.240 4596.300 1163.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1462.240 4596.300 1463.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1762.240 4596.300 1763.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2062.240 4596.300 2063.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2362.240 10.640 2363.840 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2362.240 4596.300 2363.840 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2662.240 10.640 2663.840 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2662.240 4596.300 2663.840 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4609.480 3154.920 4612.680 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 34.920 0.000 39.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3123.180 0.000 3128.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 57.280 3165.000 67.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4693.160 3165.000 4703.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 831.480 3154.920 836.280 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 46.920 0.000 51.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3111.180 0.000 3116.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 80.480 3165.000 90.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4669.960 3165.000 4679.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 847.480 3154.920 852.280 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 58.920 0.000 63.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3099.180 0.000 3104.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 103.680 3165.000 113.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4646.760 3165.000 4656.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 863.480 3154.920 868.280 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 52.920 0.000 57.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3105.180 0.000 3110.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 92.080 3165.000 102.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4658.360 3165.000 4668.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 855.480 3154.920 860.280 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 64.920 0.000 69.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3093.180 0.000 3098.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 115.280 3165.000 125.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4635.160 3165.000 4645.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 871.480 3154.920 876.280 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.920 0.000 21.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3141.180 0.000 3146.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 22.480 3165.000 32.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4727.960 3165.000 4737.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.515 10.640 76.515 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3089.585 10.640 3091.585 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.120 10.640 138.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.120 669.885 138.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.120 4596.300 138.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 235.120 10.640 238.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 235.120 669.885 238.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 235.120 4596.300 238.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.120 10.640 338.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.120 669.885 338.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.120 4596.300 338.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.120 10.640 438.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.120 669.885 438.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.120 4596.300 438.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.120 10.640 538.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.120 669.885 538.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.120 4596.300 538.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.120 10.640 638.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.120 669.885 638.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.120 4603.350 638.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.120 10.640 738.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.120 669.885 738.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.120 4596.300 738.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 835.120 10.640 838.320 169.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 835.120 669.885 838.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 835.120 4596.300 838.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.120 10.640 938.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.120 936.205 938.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 935.120 4596.300 938.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.120 10.640 1038.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.120 936.205 1038.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.120 4596.300 1038.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.120 10.640 1138.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.120 936.205 1138.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1135.120 4596.300 1138.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.120 10.640 1238.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.120 936.205 1238.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.120 4596.300 1238.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.120 10.640 1338.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.120 936.205 1338.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.120 4596.300 1338.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.120 10.640 1438.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.120 936.205 1438.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1435.120 4596.300 1438.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.120 10.640 1538.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.120 936.205 1538.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.120 4603.350 1538.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1635.120 10.640 1638.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1635.120 936.205 1638.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1635.120 4596.300 1638.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.120 10.640 1738.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.120 936.205 1738.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1735.120 4596.300 1738.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1835.120 10.640 1838.320 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 1835.120 582.645 1838.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1835.120 936.205 1838.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1835.120 4596.300 1838.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.120 10.640 1938.320 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.120 582.645 1938.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.120 936.205 1938.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.120 4596.300 1938.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.120 10.640 2038.320 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.120 582.645 2038.320 779.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.120 936.205 2038.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.120 4596.300 2038.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.120 10.640 2138.320 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.120 582.645 2138.320 784.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.120 929.820 2138.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2135.120 4596.300 2138.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2235.120 10.640 2238.320 151.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2235.120 582.645 2238.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2235.120 4596.300 2238.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2335.120 10.640 2338.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2335.120 4596.300 2338.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2435.120 10.640 2438.320 784.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2435.120 929.820 2438.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2435.120 4603.350 2438.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2535.120 10.640 2538.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2535.120 4596.300 2538.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2635.120 10.640 2638.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2635.120 4596.300 2638.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.120 10.640 2738.320 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.120 735.325 2738.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.120 4596.300 2738.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.120 10.640 2838.320 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.120 735.325 2838.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.120 4596.300 2838.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2935.120 10.640 2938.320 192.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2935.120 735.325 2938.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2935.120 4596.300 2938.320 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 3035.120 10.640 3038.320 192.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 3035.120 737.100 3038.320 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3035.120 4596.300 3038.320 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 199.880 3154.920 203.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 319.880 3154.920 323.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 439.880 3154.920 443.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 559.880 3154.920 563.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 679.880 3154.920 683.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 799.880 3154.920 803.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 919.880 3154.920 923.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1039.880 76.000 1043.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1159.880 76.000 1163.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1279.880 76.000 1283.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1399.880 76.000 1403.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1519.880 76.000 1523.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1639.880 76.000 1643.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1759.880 76.000 1763.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1879.880 76.000 1883.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 1999.880 76.000 2003.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2119.880 76.000 2123.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2239.880 76.000 2243.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2359.880 76.000 2363.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2479.880 76.000 2483.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2599.880 76.000 2603.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2719.880 76.000 2723.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2839.880 76.000 2843.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 2959.880 76.000 2963.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3079.880 76.000 3083.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3199.880 76.000 3203.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3319.880 76.000 3323.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3439.880 76.000 3443.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3559.880 76.000 3563.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3679.880 76.000 3683.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3799.880 76.000 3803.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 3919.880 76.000 3923.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4039.880 76.000 4043.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4159.880 76.000 4163.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4279.880 76.000 4283.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4399.880 76.000 4403.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4519.880 76.000 4523.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1039.880 3154.920 1043.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1159.880 3154.920 1163.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1279.880 3154.920 1283.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1399.880 3154.920 1403.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1519.880 3154.920 1523.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1639.880 3154.920 1643.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1759.880 3154.920 1763.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1879.880 3154.920 1883.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 1999.880 3154.920 2003.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2119.880 3154.920 2123.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2239.880 3154.920 2243.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2359.880 3154.920 2363.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2479.880 3154.920 2483.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2599.880 3154.920 2603.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2719.880 3154.920 2723.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2839.880 3154.920 2843.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 2959.880 3154.920 2963.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3079.880 3154.920 3083.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3199.880 3154.920 3203.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3319.880 3154.920 3323.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3439.880 3154.920 3443.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3559.880 3154.920 3563.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3679.880 3154.920 3683.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3799.880 3154.920 3803.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 3919.880 3154.920 3923.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4039.880 3154.920 4043.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4159.880 3154.920 4163.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4279.880 3154.920 4283.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4399.880 3154.920 4403.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 3087.000 4519.880 3154.920 4523.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 258.680 3154.920 263.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 378.680 3154.920 383.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 498.680 3154.920 503.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 618.680 3154.920 623.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 825.520 962.300 2238.320 972.300 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.920 0.000 33.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3129.180 0.000 3134.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.680 3165.000 55.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4704.760 3165.000 4714.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 823.480 3154.920 828.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.440 4596.300 260.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.440 4596.300 560.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.440 669.885 860.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.440 4596.300 860.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.440 4596.300 1160.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.440 4596.300 1460.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.440 4596.300 1760.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.440 4596.300 2060.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.440 10.640 2360.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.440 4596.300 2360.040 4754.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.440 10.640 2660.040 989.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.440 4596.300 2660.040 4754.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 4604.040 3154.920 4607.240 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 40.920 0.000 45.920 4767.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 3117.180 0.000 3122.180 4767.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.880 3165.000 78.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 4681.560 3165.000 4691.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 839.480 3154.920 844.280 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 3154.680 4754.645 ;
      LAYER met1 ;
        RECT 5.590 10.640 3159.210 4754.800 ;
      LAYER met2 ;
        RECT 5.610 4762.720 173.465 4764.490 ;
        RECT 174.305 4762.720 176.685 4764.490 ;
        RECT 177.525 4762.720 179.905 4764.490 ;
        RECT 180.745 4762.720 189.105 4764.490 ;
        RECT 189.945 4762.720 191.865 4764.490 ;
        RECT 192.705 4762.720 195.085 4764.490 ;
        RECT 195.925 4762.720 198.305 4764.490 ;
        RECT 199.145 4762.720 210.725 4764.490 ;
        RECT 211.565 4762.720 213.485 4764.490 ;
        RECT 214.325 4762.720 216.705 4764.490 ;
        RECT 217.545 4762.720 219.925 4764.490 ;
        RECT 220.765 4762.720 225.905 4764.490 ;
        RECT 226.745 4762.720 231.885 4764.490 ;
        RECT 232.725 4762.720 235.105 4764.490 ;
        RECT 235.945 4762.720 238.325 4764.490 ;
        RECT 239.165 4762.720 244.305 4764.490 ;
        RECT 245.145 4762.720 430.465 4764.490 ;
        RECT 431.305 4762.720 433.685 4764.490 ;
        RECT 434.525 4762.720 436.905 4764.490 ;
        RECT 437.745 4762.720 446.105 4764.490 ;
        RECT 446.945 4762.720 448.865 4764.490 ;
        RECT 449.705 4762.720 452.085 4764.490 ;
        RECT 452.925 4762.720 455.305 4764.490 ;
        RECT 456.145 4762.720 467.725 4764.490 ;
        RECT 468.565 4762.720 470.485 4764.490 ;
        RECT 471.325 4762.720 473.705 4764.490 ;
        RECT 474.545 4762.720 476.925 4764.490 ;
        RECT 477.765 4762.720 482.905 4764.490 ;
        RECT 483.745 4762.720 488.885 4764.490 ;
        RECT 489.725 4762.720 492.105 4764.490 ;
        RECT 492.945 4762.720 495.325 4764.490 ;
        RECT 496.165 4762.720 501.305 4764.490 ;
        RECT 502.145 4762.720 687.465 4764.490 ;
        RECT 688.305 4762.720 690.685 4764.490 ;
        RECT 691.525 4762.720 693.905 4764.490 ;
        RECT 694.745 4762.720 703.105 4764.490 ;
        RECT 703.945 4762.720 705.865 4764.490 ;
        RECT 706.705 4762.720 709.085 4764.490 ;
        RECT 709.925 4762.720 712.305 4764.490 ;
        RECT 713.145 4762.720 724.725 4764.490 ;
        RECT 725.565 4762.720 727.485 4764.490 ;
        RECT 728.325 4762.720 730.705 4764.490 ;
        RECT 731.545 4762.720 733.925 4764.490 ;
        RECT 734.765 4762.720 739.905 4764.490 ;
        RECT 740.745 4762.720 745.885 4764.490 ;
        RECT 746.725 4762.720 749.105 4764.490 ;
        RECT 749.945 4762.720 752.325 4764.490 ;
        RECT 753.165 4762.720 758.305 4764.490 ;
        RECT 759.145 4762.720 944.465 4764.490 ;
        RECT 945.305 4762.720 947.685 4764.490 ;
        RECT 948.525 4762.720 950.905 4764.490 ;
        RECT 951.745 4762.720 960.105 4764.490 ;
        RECT 960.945 4762.720 962.865 4764.490 ;
        RECT 963.705 4762.720 966.085 4764.490 ;
        RECT 966.925 4762.720 969.305 4764.490 ;
        RECT 970.145 4762.720 981.725 4764.490 ;
        RECT 982.565 4762.720 984.485 4764.490 ;
        RECT 985.325 4762.720 987.705 4764.490 ;
        RECT 988.545 4762.720 990.925 4764.490 ;
        RECT 991.765 4762.720 996.905 4764.490 ;
        RECT 997.745 4762.720 1002.885 4764.490 ;
        RECT 1003.725 4762.720 1006.105 4764.490 ;
        RECT 1006.945 4762.720 1009.325 4764.490 ;
        RECT 1010.165 4762.720 1015.305 4764.490 ;
        RECT 1016.145 4762.720 1202.465 4764.490 ;
        RECT 1203.305 4762.720 1205.685 4764.490 ;
        RECT 1206.525 4762.720 1208.905 4764.490 ;
        RECT 1209.745 4762.720 1218.105 4764.490 ;
        RECT 1218.945 4762.720 1220.865 4764.490 ;
        RECT 1221.705 4762.720 1224.085 4764.490 ;
        RECT 1224.925 4762.720 1227.305 4764.490 ;
        RECT 1228.145 4762.720 1239.725 4764.490 ;
        RECT 1240.565 4762.720 1242.485 4764.490 ;
        RECT 1243.325 4762.720 1245.705 4764.490 ;
        RECT 1246.545 4762.720 1248.925 4764.490 ;
        RECT 1249.765 4762.720 1254.905 4764.490 ;
        RECT 1255.745 4762.720 1260.885 4764.490 ;
        RECT 1261.725 4762.720 1264.105 4764.490 ;
        RECT 1264.945 4762.720 1267.325 4764.490 ;
        RECT 1268.165 4762.720 1273.305 4764.490 ;
        RECT 1274.145 4762.720 1711.465 4764.490 ;
        RECT 1712.305 4762.720 1714.685 4764.490 ;
        RECT 1715.525 4762.720 1717.905 4764.490 ;
        RECT 1718.745 4762.720 1727.105 4764.490 ;
        RECT 1727.945 4762.720 1729.865 4764.490 ;
        RECT 1730.705 4762.720 1733.085 4764.490 ;
        RECT 1733.925 4762.720 1736.305 4764.490 ;
        RECT 1737.145 4762.720 1748.725 4764.490 ;
        RECT 1749.565 4762.720 1751.485 4764.490 ;
        RECT 1752.325 4762.720 1754.705 4764.490 ;
        RECT 1755.545 4762.720 1757.925 4764.490 ;
        RECT 1758.765 4762.720 1763.905 4764.490 ;
        RECT 1764.745 4762.720 1769.885 4764.490 ;
        RECT 1770.725 4762.720 1773.105 4764.490 ;
        RECT 1773.945 4762.720 1776.325 4764.490 ;
        RECT 1777.165 4762.720 1782.305 4764.490 ;
        RECT 1783.145 4762.720 2156.465 4764.490 ;
        RECT 2157.305 4762.720 2159.685 4764.490 ;
        RECT 2160.525 4762.720 2162.905 4764.490 ;
        RECT 2163.745 4762.720 2172.105 4764.490 ;
        RECT 2172.945 4762.720 2174.865 4764.490 ;
        RECT 2175.705 4762.720 2178.085 4764.490 ;
        RECT 2178.925 4762.720 2181.305 4764.490 ;
        RECT 2182.145 4762.720 2193.725 4764.490 ;
        RECT 2194.565 4762.720 2196.485 4764.490 ;
        RECT 2197.325 4762.720 2199.705 4764.490 ;
        RECT 2200.545 4762.720 2202.925 4764.490 ;
        RECT 2203.765 4762.720 2208.905 4764.490 ;
        RECT 2209.745 4762.720 2214.885 4764.490 ;
        RECT 2215.725 4762.720 2218.105 4764.490 ;
        RECT 2218.945 4762.720 2221.325 4764.490 ;
        RECT 2222.165 4762.720 2227.305 4764.490 ;
        RECT 2228.145 4762.720 2413.465 4764.490 ;
        RECT 2414.305 4762.720 2416.685 4764.490 ;
        RECT 2417.525 4762.720 2419.905 4764.490 ;
        RECT 2420.745 4762.720 2429.105 4764.490 ;
        RECT 2429.945 4762.720 2431.865 4764.490 ;
        RECT 2432.705 4762.720 2435.085 4764.490 ;
        RECT 2435.925 4762.720 2438.305 4764.490 ;
        RECT 2439.145 4762.720 2450.725 4764.490 ;
        RECT 2451.565 4762.720 2453.485 4764.490 ;
        RECT 2454.325 4762.720 2456.705 4764.490 ;
        RECT 2457.545 4762.720 2459.925 4764.490 ;
        RECT 2460.765 4762.720 2465.905 4764.490 ;
        RECT 2466.745 4762.720 2471.885 4764.490 ;
        RECT 2472.725 4762.720 2475.105 4764.490 ;
        RECT 2475.945 4762.720 2478.325 4764.490 ;
        RECT 2479.165 4762.720 2484.305 4764.490 ;
        RECT 2485.145 4762.720 2922.465 4764.490 ;
        RECT 2923.305 4762.720 2925.685 4764.490 ;
        RECT 2926.525 4762.720 2928.905 4764.490 ;
        RECT 2929.745 4762.720 2938.105 4764.490 ;
        RECT 2938.945 4762.720 2940.865 4764.490 ;
        RECT 2941.705 4762.720 2944.085 4764.490 ;
        RECT 2944.925 4762.720 2947.305 4764.490 ;
        RECT 2948.145 4762.720 2959.725 4764.490 ;
        RECT 2960.565 4762.720 2962.485 4764.490 ;
        RECT 2963.325 4762.720 2965.705 4764.490 ;
        RECT 2966.545 4762.720 2968.925 4764.490 ;
        RECT 2969.765 4762.720 2974.905 4764.490 ;
        RECT 2975.745 4762.720 2980.885 4764.490 ;
        RECT 2981.725 4762.720 2984.105 4764.490 ;
        RECT 2984.945 4762.720 2987.325 4764.490 ;
        RECT 2988.165 4762.720 2993.305 4764.490 ;
        RECT 2994.145 4762.720 3159.190 4764.490 ;
        RECT 5.610 4.280 3159.190 4762.720 ;
        RECT 5.610 3.670 496.555 4.280 ;
        RECT 497.395 3.670 724.855 4.280 ;
        RECT 725.695 3.670 758.435 4.280 ;
        RECT 759.275 3.670 1323.055 4.280 ;
        RECT 1323.895 3.670 1329.495 4.280 ;
        RECT 1330.335 3.670 1338.695 4.280 ;
        RECT 1339.535 3.670 1597.055 4.280 ;
        RECT 1597.895 3.670 1612.695 4.280 ;
        RECT 1613.535 3.670 1815.855 4.280 ;
        RECT 1816.695 3.670 1849.435 4.280 ;
        RECT 1850.275 3.670 1871.055 4.280 ;
        RECT 1871.895 3.670 1886.695 4.280 ;
        RECT 1887.535 3.670 2089.855 4.280 ;
        RECT 2090.695 3.670 2123.435 4.280 ;
        RECT 2124.275 3.670 2145.055 4.280 ;
        RECT 2145.895 3.670 2160.695 4.280 ;
        RECT 2161.535 3.670 2363.855 4.280 ;
        RECT 2364.695 3.670 2391.455 4.280 ;
        RECT 2392.295 3.670 2397.435 4.280 ;
        RECT 2398.275 3.670 2413.075 4.280 ;
        RECT 2413.915 3.670 2419.055 4.280 ;
        RECT 2419.895 3.670 2434.695 4.280 ;
        RECT 2435.535 3.670 3159.190 4.280 ;
      LAYER met3 ;
        RECT 3.070 4636.425 3161.730 4754.725 ;
        RECT 4.400 4635.025 3161.730 4636.425 ;
        RECT 3.070 4630.445 3161.730 4635.025 ;
        RECT 4.400 4629.045 3161.730 4630.445 ;
        RECT 3.070 4627.225 3161.730 4629.045 ;
        RECT 4.400 4625.825 3161.730 4627.225 ;
        RECT 3.070 4624.005 3161.730 4625.825 ;
        RECT 4.400 4623.815 3161.730 4624.005 ;
        RECT 4.400 4622.605 3160.600 4623.815 ;
        RECT 3.070 4622.415 3160.600 4622.605 ;
        RECT 3.070 4620.595 3161.730 4622.415 ;
        RECT 3.070 4619.195 3160.600 4620.595 ;
        RECT 3.070 4618.025 3161.730 4619.195 ;
        RECT 4.400 4617.375 3161.730 4618.025 ;
        RECT 4.400 4616.625 3160.600 4617.375 ;
        RECT 3.070 4615.975 3160.600 4616.625 ;
        RECT 3.070 4612.045 3161.730 4615.975 ;
        RECT 4.400 4610.645 3161.730 4612.045 ;
        RECT 3.070 4608.825 3161.730 4610.645 ;
        RECT 4.400 4608.175 3161.730 4608.825 ;
        RECT 4.400 4607.425 3160.600 4608.175 ;
        RECT 3.070 4606.775 3160.600 4607.425 ;
        RECT 3.070 4605.605 3161.730 4606.775 ;
        RECT 4.400 4605.415 3161.730 4605.605 ;
        RECT 4.400 4604.205 3160.600 4605.415 ;
        RECT 3.070 4604.015 3160.600 4604.205 ;
        RECT 3.070 4602.845 3161.730 4604.015 ;
        RECT 4.400 4602.195 3161.730 4602.845 ;
        RECT 4.400 4601.445 3160.600 4602.195 ;
        RECT 3.070 4600.795 3160.600 4601.445 ;
        RECT 3.070 4598.975 3161.730 4600.795 ;
        RECT 3.070 4597.575 3160.600 4598.975 ;
        RECT 3.070 4590.425 3161.730 4597.575 ;
        RECT 4.400 4589.025 3161.730 4590.425 ;
        RECT 3.070 4587.205 3161.730 4589.025 ;
        RECT 4.400 4586.555 3161.730 4587.205 ;
        RECT 4.400 4585.805 3160.600 4586.555 ;
        RECT 3.070 4585.155 3160.600 4585.805 ;
        RECT 3.070 4583.985 3161.730 4585.155 ;
        RECT 4.400 4583.795 3161.730 4583.985 ;
        RECT 4.400 4582.585 3160.600 4583.795 ;
        RECT 3.070 4582.395 3160.600 4582.585 ;
        RECT 3.070 4581.225 3161.730 4582.395 ;
        RECT 4.400 4580.575 3161.730 4581.225 ;
        RECT 4.400 4579.825 3160.600 4580.575 ;
        RECT 3.070 4579.175 3160.600 4579.825 ;
        RECT 3.070 4577.355 3161.730 4579.175 ;
        RECT 3.070 4575.955 3160.600 4577.355 ;
        RECT 3.070 4572.025 3161.730 4575.955 ;
        RECT 4.400 4571.375 3161.730 4572.025 ;
        RECT 4.400 4570.625 3160.600 4571.375 ;
        RECT 3.070 4569.975 3160.600 4570.625 ;
        RECT 3.070 4568.805 3161.730 4569.975 ;
        RECT 4.400 4567.405 3161.730 4568.805 ;
        RECT 3.070 4565.585 3161.730 4567.405 ;
        RECT 4.400 4565.395 3161.730 4565.585 ;
        RECT 4.400 4564.185 3160.600 4565.395 ;
        RECT 3.070 4563.995 3160.600 4564.185 ;
        RECT 3.070 4562.175 3161.730 4563.995 ;
        RECT 3.070 4560.775 3160.600 4562.175 ;
        RECT 3.070 4558.955 3161.730 4560.775 ;
        RECT 3.070 4557.555 3160.600 4558.955 ;
        RECT 3.070 4552.975 3161.730 4557.555 ;
        RECT 3.070 4551.575 3160.600 4552.975 ;
        RECT 3.070 4177.815 3161.730 4551.575 ;
        RECT 3.070 4176.415 3160.600 4177.815 ;
        RECT 3.070 4174.595 3161.730 4176.415 ;
        RECT 3.070 4173.195 3160.600 4174.595 ;
        RECT 3.070 4171.375 3161.730 4173.195 ;
        RECT 3.070 4169.975 3160.600 4171.375 ;
        RECT 3.070 4162.175 3161.730 4169.975 ;
        RECT 3.070 4160.775 3160.600 4162.175 ;
        RECT 3.070 4159.415 3161.730 4160.775 ;
        RECT 3.070 4158.015 3160.600 4159.415 ;
        RECT 3.070 4156.195 3161.730 4158.015 ;
        RECT 3.070 4154.795 3160.600 4156.195 ;
        RECT 3.070 4152.975 3161.730 4154.795 ;
        RECT 3.070 4151.575 3160.600 4152.975 ;
        RECT 3.070 4140.555 3161.730 4151.575 ;
        RECT 3.070 4139.155 3160.600 4140.555 ;
        RECT 3.070 4137.795 3161.730 4139.155 ;
        RECT 3.070 4136.395 3160.600 4137.795 ;
        RECT 3.070 4134.575 3161.730 4136.395 ;
        RECT 3.070 4133.175 3160.600 4134.575 ;
        RECT 3.070 4131.355 3161.730 4133.175 ;
        RECT 3.070 4129.955 3160.600 4131.355 ;
        RECT 3.070 4125.375 3161.730 4129.955 ;
        RECT 3.070 4123.975 3160.600 4125.375 ;
        RECT 3.070 4119.395 3161.730 4123.975 ;
        RECT 3.070 4117.995 3160.600 4119.395 ;
        RECT 3.070 4116.175 3161.730 4117.995 ;
        RECT 3.070 4114.775 3160.600 4116.175 ;
        RECT 3.070 4112.955 3161.730 4114.775 ;
        RECT 3.070 4111.555 3160.600 4112.955 ;
        RECT 3.070 4106.975 3161.730 4111.555 ;
        RECT 3.070 4105.575 3160.600 4106.975 ;
        RECT 3.070 3787.425 3161.730 4105.575 ;
        RECT 4.400 3786.025 3161.730 3787.425 ;
        RECT 3.070 3781.445 3161.730 3786.025 ;
        RECT 4.400 3780.045 3161.730 3781.445 ;
        RECT 3.070 3778.225 3161.730 3780.045 ;
        RECT 4.400 3776.825 3161.730 3778.225 ;
        RECT 3.070 3775.005 3161.730 3776.825 ;
        RECT 4.400 3773.605 3161.730 3775.005 ;
        RECT 3.070 3769.025 3161.730 3773.605 ;
        RECT 4.400 3767.625 3161.730 3769.025 ;
        RECT 3.070 3763.045 3161.730 3767.625 ;
        RECT 4.400 3761.645 3161.730 3763.045 ;
        RECT 3.070 3759.825 3161.730 3761.645 ;
        RECT 4.400 3758.425 3161.730 3759.825 ;
        RECT 3.070 3756.605 3161.730 3758.425 ;
        RECT 4.400 3755.205 3161.730 3756.605 ;
        RECT 3.070 3753.845 3161.730 3755.205 ;
        RECT 4.400 3752.445 3161.730 3753.845 ;
        RECT 3.070 3741.425 3161.730 3752.445 ;
        RECT 4.400 3740.025 3161.730 3741.425 ;
        RECT 3.070 3738.205 3161.730 3740.025 ;
        RECT 4.400 3736.805 3161.730 3738.205 ;
        RECT 3.070 3734.985 3161.730 3736.805 ;
        RECT 4.400 3733.585 3161.730 3734.985 ;
        RECT 3.070 3732.225 3161.730 3733.585 ;
        RECT 4.400 3731.815 3161.730 3732.225 ;
        RECT 4.400 3730.825 3160.600 3731.815 ;
        RECT 3.070 3730.415 3160.600 3730.825 ;
        RECT 3.070 3728.595 3161.730 3730.415 ;
        RECT 3.070 3727.195 3160.600 3728.595 ;
        RECT 3.070 3725.375 3161.730 3727.195 ;
        RECT 3.070 3723.975 3160.600 3725.375 ;
        RECT 3.070 3723.025 3161.730 3723.975 ;
        RECT 4.400 3721.625 3161.730 3723.025 ;
        RECT 3.070 3719.805 3161.730 3721.625 ;
        RECT 4.400 3718.405 3161.730 3719.805 ;
        RECT 3.070 3716.585 3161.730 3718.405 ;
        RECT 4.400 3716.175 3161.730 3716.585 ;
        RECT 4.400 3715.185 3160.600 3716.175 ;
        RECT 3.070 3714.775 3160.600 3715.185 ;
        RECT 3.070 3713.415 3161.730 3714.775 ;
        RECT 3.070 3712.015 3160.600 3713.415 ;
        RECT 3.070 3710.195 3161.730 3712.015 ;
        RECT 3.070 3708.795 3160.600 3710.195 ;
        RECT 3.070 3706.975 3161.730 3708.795 ;
        RECT 3.070 3705.575 3160.600 3706.975 ;
        RECT 3.070 3694.555 3161.730 3705.575 ;
        RECT 3.070 3693.155 3160.600 3694.555 ;
        RECT 3.070 3691.795 3161.730 3693.155 ;
        RECT 3.070 3690.395 3160.600 3691.795 ;
        RECT 3.070 3688.575 3161.730 3690.395 ;
        RECT 3.070 3687.175 3160.600 3688.575 ;
        RECT 3.070 3685.355 3161.730 3687.175 ;
        RECT 3.070 3683.955 3160.600 3685.355 ;
        RECT 3.070 3679.375 3161.730 3683.955 ;
        RECT 3.070 3677.975 3160.600 3679.375 ;
        RECT 3.070 3673.395 3161.730 3677.975 ;
        RECT 3.070 3671.995 3160.600 3673.395 ;
        RECT 3.070 3670.175 3161.730 3671.995 ;
        RECT 3.070 3668.775 3160.600 3670.175 ;
        RECT 3.070 3666.955 3161.730 3668.775 ;
        RECT 3.070 3665.555 3160.600 3666.955 ;
        RECT 3.070 3660.975 3161.730 3665.555 ;
        RECT 3.070 3659.575 3160.600 3660.975 ;
        RECT 3.070 3571.425 3161.730 3659.575 ;
        RECT 4.400 3570.025 3161.730 3571.425 ;
        RECT 3.070 3565.445 3161.730 3570.025 ;
        RECT 4.400 3564.045 3161.730 3565.445 ;
        RECT 3.070 3562.225 3161.730 3564.045 ;
        RECT 4.400 3560.825 3161.730 3562.225 ;
        RECT 3.070 3559.005 3161.730 3560.825 ;
        RECT 4.400 3557.605 3161.730 3559.005 ;
        RECT 3.070 3553.025 3161.730 3557.605 ;
        RECT 4.400 3551.625 3161.730 3553.025 ;
        RECT 3.070 3547.045 3161.730 3551.625 ;
        RECT 4.400 3545.645 3161.730 3547.045 ;
        RECT 3.070 3543.825 3161.730 3545.645 ;
        RECT 4.400 3542.425 3161.730 3543.825 ;
        RECT 3.070 3540.605 3161.730 3542.425 ;
        RECT 4.400 3539.205 3161.730 3540.605 ;
        RECT 3.070 3537.845 3161.730 3539.205 ;
        RECT 4.400 3536.445 3161.730 3537.845 ;
        RECT 3.070 3525.425 3161.730 3536.445 ;
        RECT 4.400 3524.025 3161.730 3525.425 ;
        RECT 3.070 3522.205 3161.730 3524.025 ;
        RECT 4.400 3520.805 3161.730 3522.205 ;
        RECT 3.070 3518.985 3161.730 3520.805 ;
        RECT 4.400 3517.585 3161.730 3518.985 ;
        RECT 3.070 3516.225 3161.730 3517.585 ;
        RECT 4.400 3514.825 3161.730 3516.225 ;
        RECT 3.070 3507.025 3161.730 3514.825 ;
        RECT 4.400 3506.815 3161.730 3507.025 ;
        RECT 4.400 3505.625 3160.600 3506.815 ;
        RECT 3.070 3505.415 3160.600 3505.625 ;
        RECT 3.070 3503.805 3161.730 3505.415 ;
        RECT 4.400 3503.595 3161.730 3503.805 ;
        RECT 4.400 3502.405 3160.600 3503.595 ;
        RECT 3.070 3502.195 3160.600 3502.405 ;
        RECT 3.070 3500.585 3161.730 3502.195 ;
        RECT 4.400 3500.375 3161.730 3500.585 ;
        RECT 4.400 3499.185 3160.600 3500.375 ;
        RECT 3.070 3498.975 3160.600 3499.185 ;
        RECT 3.070 3491.175 3161.730 3498.975 ;
        RECT 3.070 3489.775 3160.600 3491.175 ;
        RECT 3.070 3488.415 3161.730 3489.775 ;
        RECT 3.070 3487.015 3160.600 3488.415 ;
        RECT 3.070 3485.195 3161.730 3487.015 ;
        RECT 3.070 3483.795 3160.600 3485.195 ;
        RECT 3.070 3481.975 3161.730 3483.795 ;
        RECT 3.070 3480.575 3160.600 3481.975 ;
        RECT 3.070 3469.555 3161.730 3480.575 ;
        RECT 3.070 3468.155 3160.600 3469.555 ;
        RECT 3.070 3466.795 3161.730 3468.155 ;
        RECT 3.070 3465.395 3160.600 3466.795 ;
        RECT 3.070 3463.575 3161.730 3465.395 ;
        RECT 3.070 3462.175 3160.600 3463.575 ;
        RECT 3.070 3460.355 3161.730 3462.175 ;
        RECT 3.070 3458.955 3160.600 3460.355 ;
        RECT 3.070 3454.375 3161.730 3458.955 ;
        RECT 3.070 3452.975 3160.600 3454.375 ;
        RECT 3.070 3448.395 3161.730 3452.975 ;
        RECT 3.070 3446.995 3160.600 3448.395 ;
        RECT 3.070 3445.175 3161.730 3446.995 ;
        RECT 3.070 3443.775 3160.600 3445.175 ;
        RECT 3.070 3441.955 3161.730 3443.775 ;
        RECT 3.070 3440.555 3160.600 3441.955 ;
        RECT 3.070 3435.975 3161.730 3440.555 ;
        RECT 3.070 3434.575 3160.600 3435.975 ;
        RECT 3.070 3355.425 3161.730 3434.575 ;
        RECT 4.400 3354.025 3161.730 3355.425 ;
        RECT 3.070 3349.445 3161.730 3354.025 ;
        RECT 4.400 3348.045 3161.730 3349.445 ;
        RECT 3.070 3346.225 3161.730 3348.045 ;
        RECT 4.400 3344.825 3161.730 3346.225 ;
        RECT 3.070 3343.005 3161.730 3344.825 ;
        RECT 4.400 3341.605 3161.730 3343.005 ;
        RECT 3.070 3337.025 3161.730 3341.605 ;
        RECT 4.400 3335.625 3161.730 3337.025 ;
        RECT 3.070 3331.045 3161.730 3335.625 ;
        RECT 4.400 3329.645 3161.730 3331.045 ;
        RECT 3.070 3327.825 3161.730 3329.645 ;
        RECT 4.400 3326.425 3161.730 3327.825 ;
        RECT 3.070 3324.605 3161.730 3326.425 ;
        RECT 4.400 3323.205 3161.730 3324.605 ;
        RECT 3.070 3321.845 3161.730 3323.205 ;
        RECT 4.400 3320.445 3161.730 3321.845 ;
        RECT 3.070 3309.425 3161.730 3320.445 ;
        RECT 4.400 3308.025 3161.730 3309.425 ;
        RECT 3.070 3306.205 3161.730 3308.025 ;
        RECT 4.400 3304.805 3161.730 3306.205 ;
        RECT 3.070 3302.985 3161.730 3304.805 ;
        RECT 4.400 3301.585 3161.730 3302.985 ;
        RECT 3.070 3300.225 3161.730 3301.585 ;
        RECT 4.400 3298.825 3161.730 3300.225 ;
        RECT 3.070 3291.025 3161.730 3298.825 ;
        RECT 4.400 3289.625 3161.730 3291.025 ;
        RECT 3.070 3287.805 3161.730 3289.625 ;
        RECT 4.400 3286.405 3161.730 3287.805 ;
        RECT 3.070 3284.585 3161.730 3286.405 ;
        RECT 4.400 3283.185 3161.730 3284.585 ;
        RECT 3.070 3281.815 3161.730 3283.185 ;
        RECT 3.070 3280.415 3160.600 3281.815 ;
        RECT 3.070 3278.595 3161.730 3280.415 ;
        RECT 3.070 3277.195 3160.600 3278.595 ;
        RECT 3.070 3275.375 3161.730 3277.195 ;
        RECT 3.070 3273.975 3160.600 3275.375 ;
        RECT 3.070 3266.175 3161.730 3273.975 ;
        RECT 3.070 3264.775 3160.600 3266.175 ;
        RECT 3.070 3263.415 3161.730 3264.775 ;
        RECT 3.070 3262.015 3160.600 3263.415 ;
        RECT 3.070 3260.195 3161.730 3262.015 ;
        RECT 3.070 3258.795 3160.600 3260.195 ;
        RECT 3.070 3256.975 3161.730 3258.795 ;
        RECT 3.070 3255.575 3160.600 3256.975 ;
        RECT 3.070 3244.555 3161.730 3255.575 ;
        RECT 3.070 3243.155 3160.600 3244.555 ;
        RECT 3.070 3241.795 3161.730 3243.155 ;
        RECT 3.070 3240.395 3160.600 3241.795 ;
        RECT 3.070 3238.575 3161.730 3240.395 ;
        RECT 3.070 3237.175 3160.600 3238.575 ;
        RECT 3.070 3235.355 3161.730 3237.175 ;
        RECT 3.070 3233.955 3160.600 3235.355 ;
        RECT 3.070 3229.375 3161.730 3233.955 ;
        RECT 3.070 3227.975 3160.600 3229.375 ;
        RECT 3.070 3223.395 3161.730 3227.975 ;
        RECT 3.070 3221.995 3160.600 3223.395 ;
        RECT 3.070 3220.175 3161.730 3221.995 ;
        RECT 3.070 3218.775 3160.600 3220.175 ;
        RECT 3.070 3216.955 3161.730 3218.775 ;
        RECT 3.070 3215.555 3160.600 3216.955 ;
        RECT 3.070 3210.975 3161.730 3215.555 ;
        RECT 3.070 3209.575 3160.600 3210.975 ;
        RECT 3.070 3139.425 3161.730 3209.575 ;
        RECT 4.400 3138.025 3161.730 3139.425 ;
        RECT 3.070 3133.445 3161.730 3138.025 ;
        RECT 4.400 3132.045 3161.730 3133.445 ;
        RECT 3.070 3130.225 3161.730 3132.045 ;
        RECT 4.400 3128.825 3161.730 3130.225 ;
        RECT 3.070 3127.005 3161.730 3128.825 ;
        RECT 4.400 3125.605 3161.730 3127.005 ;
        RECT 3.070 3121.025 3161.730 3125.605 ;
        RECT 4.400 3119.625 3161.730 3121.025 ;
        RECT 3.070 3115.045 3161.730 3119.625 ;
        RECT 4.400 3113.645 3161.730 3115.045 ;
        RECT 3.070 3111.825 3161.730 3113.645 ;
        RECT 4.400 3110.425 3161.730 3111.825 ;
        RECT 3.070 3108.605 3161.730 3110.425 ;
        RECT 4.400 3107.205 3161.730 3108.605 ;
        RECT 3.070 3105.845 3161.730 3107.205 ;
        RECT 4.400 3104.445 3161.730 3105.845 ;
        RECT 3.070 3093.425 3161.730 3104.445 ;
        RECT 4.400 3092.025 3161.730 3093.425 ;
        RECT 3.070 3090.205 3161.730 3092.025 ;
        RECT 4.400 3088.805 3161.730 3090.205 ;
        RECT 3.070 3086.985 3161.730 3088.805 ;
        RECT 4.400 3085.585 3161.730 3086.985 ;
        RECT 3.070 3084.225 3161.730 3085.585 ;
        RECT 4.400 3082.825 3161.730 3084.225 ;
        RECT 3.070 3075.025 3161.730 3082.825 ;
        RECT 4.400 3073.625 3161.730 3075.025 ;
        RECT 3.070 3071.805 3161.730 3073.625 ;
        RECT 4.400 3070.405 3161.730 3071.805 ;
        RECT 3.070 3068.585 3161.730 3070.405 ;
        RECT 4.400 3067.185 3161.730 3068.585 ;
        RECT 3.070 3055.815 3161.730 3067.185 ;
        RECT 3.070 3054.415 3160.600 3055.815 ;
        RECT 3.070 3052.595 3161.730 3054.415 ;
        RECT 3.070 3051.195 3160.600 3052.595 ;
        RECT 3.070 3049.375 3161.730 3051.195 ;
        RECT 3.070 3047.975 3160.600 3049.375 ;
        RECT 3.070 3040.175 3161.730 3047.975 ;
        RECT 3.070 3038.775 3160.600 3040.175 ;
        RECT 3.070 3037.415 3161.730 3038.775 ;
        RECT 3.070 3036.015 3160.600 3037.415 ;
        RECT 3.070 3034.195 3161.730 3036.015 ;
        RECT 3.070 3032.795 3160.600 3034.195 ;
        RECT 3.070 3030.975 3161.730 3032.795 ;
        RECT 3.070 3029.575 3160.600 3030.975 ;
        RECT 3.070 3018.555 3161.730 3029.575 ;
        RECT 3.070 3017.155 3160.600 3018.555 ;
        RECT 3.070 3015.795 3161.730 3017.155 ;
        RECT 3.070 3014.395 3160.600 3015.795 ;
        RECT 3.070 3012.575 3161.730 3014.395 ;
        RECT 3.070 3011.175 3160.600 3012.575 ;
        RECT 3.070 3009.355 3161.730 3011.175 ;
        RECT 3.070 3007.955 3160.600 3009.355 ;
        RECT 3.070 3003.375 3161.730 3007.955 ;
        RECT 3.070 3001.975 3160.600 3003.375 ;
        RECT 3.070 2997.395 3161.730 3001.975 ;
        RECT 3.070 2995.995 3160.600 2997.395 ;
        RECT 3.070 2994.175 3161.730 2995.995 ;
        RECT 3.070 2992.775 3160.600 2994.175 ;
        RECT 3.070 2990.955 3161.730 2992.775 ;
        RECT 3.070 2989.555 3160.600 2990.955 ;
        RECT 3.070 2984.975 3161.730 2989.555 ;
        RECT 3.070 2983.575 3160.600 2984.975 ;
        RECT 3.070 2923.425 3161.730 2983.575 ;
        RECT 4.400 2922.025 3161.730 2923.425 ;
        RECT 3.070 2917.445 3161.730 2922.025 ;
        RECT 4.400 2916.045 3161.730 2917.445 ;
        RECT 3.070 2914.225 3161.730 2916.045 ;
        RECT 4.400 2912.825 3161.730 2914.225 ;
        RECT 3.070 2911.005 3161.730 2912.825 ;
        RECT 4.400 2909.605 3161.730 2911.005 ;
        RECT 3.070 2905.025 3161.730 2909.605 ;
        RECT 4.400 2903.625 3161.730 2905.025 ;
        RECT 3.070 2899.045 3161.730 2903.625 ;
        RECT 4.400 2897.645 3161.730 2899.045 ;
        RECT 3.070 2895.825 3161.730 2897.645 ;
        RECT 4.400 2894.425 3161.730 2895.825 ;
        RECT 3.070 2892.605 3161.730 2894.425 ;
        RECT 4.400 2891.205 3161.730 2892.605 ;
        RECT 3.070 2889.845 3161.730 2891.205 ;
        RECT 4.400 2888.445 3161.730 2889.845 ;
        RECT 3.070 2877.425 3161.730 2888.445 ;
        RECT 4.400 2876.025 3161.730 2877.425 ;
        RECT 3.070 2874.205 3161.730 2876.025 ;
        RECT 4.400 2872.805 3161.730 2874.205 ;
        RECT 3.070 2870.985 3161.730 2872.805 ;
        RECT 4.400 2869.585 3161.730 2870.985 ;
        RECT 3.070 2868.225 3161.730 2869.585 ;
        RECT 4.400 2866.825 3161.730 2868.225 ;
        RECT 3.070 2859.025 3161.730 2866.825 ;
        RECT 4.400 2857.625 3161.730 2859.025 ;
        RECT 3.070 2855.805 3161.730 2857.625 ;
        RECT 4.400 2854.405 3161.730 2855.805 ;
        RECT 3.070 2852.585 3161.730 2854.405 ;
        RECT 4.400 2851.185 3161.730 2852.585 ;
        RECT 3.070 2830.815 3161.730 2851.185 ;
        RECT 3.070 2829.415 3160.600 2830.815 ;
        RECT 3.070 2827.595 3161.730 2829.415 ;
        RECT 3.070 2826.195 3160.600 2827.595 ;
        RECT 3.070 2824.375 3161.730 2826.195 ;
        RECT 3.070 2822.975 3160.600 2824.375 ;
        RECT 3.070 2815.175 3161.730 2822.975 ;
        RECT 3.070 2813.775 3160.600 2815.175 ;
        RECT 3.070 2812.415 3161.730 2813.775 ;
        RECT 3.070 2811.015 3160.600 2812.415 ;
        RECT 3.070 2809.195 3161.730 2811.015 ;
        RECT 3.070 2807.795 3160.600 2809.195 ;
        RECT 3.070 2805.975 3161.730 2807.795 ;
        RECT 3.070 2804.575 3160.600 2805.975 ;
        RECT 3.070 2793.555 3161.730 2804.575 ;
        RECT 3.070 2792.155 3160.600 2793.555 ;
        RECT 3.070 2790.795 3161.730 2792.155 ;
        RECT 3.070 2789.395 3160.600 2790.795 ;
        RECT 3.070 2787.575 3161.730 2789.395 ;
        RECT 3.070 2786.175 3160.600 2787.575 ;
        RECT 3.070 2784.355 3161.730 2786.175 ;
        RECT 3.070 2782.955 3160.600 2784.355 ;
        RECT 3.070 2778.375 3161.730 2782.955 ;
        RECT 3.070 2776.975 3160.600 2778.375 ;
        RECT 3.070 2772.395 3161.730 2776.975 ;
        RECT 3.070 2770.995 3160.600 2772.395 ;
        RECT 3.070 2769.175 3161.730 2770.995 ;
        RECT 3.070 2767.775 3160.600 2769.175 ;
        RECT 3.070 2765.955 3161.730 2767.775 ;
        RECT 3.070 2764.555 3160.600 2765.955 ;
        RECT 3.070 2759.975 3161.730 2764.555 ;
        RECT 3.070 2758.575 3160.600 2759.975 ;
        RECT 3.070 2707.425 3161.730 2758.575 ;
        RECT 4.400 2706.025 3161.730 2707.425 ;
        RECT 3.070 2701.445 3161.730 2706.025 ;
        RECT 4.400 2700.045 3161.730 2701.445 ;
        RECT 3.070 2698.225 3161.730 2700.045 ;
        RECT 4.400 2696.825 3161.730 2698.225 ;
        RECT 3.070 2695.005 3161.730 2696.825 ;
        RECT 4.400 2693.605 3161.730 2695.005 ;
        RECT 3.070 2689.025 3161.730 2693.605 ;
        RECT 4.400 2687.625 3161.730 2689.025 ;
        RECT 3.070 2683.045 3161.730 2687.625 ;
        RECT 4.400 2681.645 3161.730 2683.045 ;
        RECT 3.070 2679.825 3161.730 2681.645 ;
        RECT 4.400 2678.425 3161.730 2679.825 ;
        RECT 3.070 2676.605 3161.730 2678.425 ;
        RECT 4.400 2675.205 3161.730 2676.605 ;
        RECT 3.070 2673.845 3161.730 2675.205 ;
        RECT 4.400 2672.445 3161.730 2673.845 ;
        RECT 3.070 2661.425 3161.730 2672.445 ;
        RECT 4.400 2660.025 3161.730 2661.425 ;
        RECT 3.070 2658.205 3161.730 2660.025 ;
        RECT 4.400 2656.805 3161.730 2658.205 ;
        RECT 3.070 2654.985 3161.730 2656.805 ;
        RECT 4.400 2653.585 3161.730 2654.985 ;
        RECT 3.070 2652.225 3161.730 2653.585 ;
        RECT 4.400 2650.825 3161.730 2652.225 ;
        RECT 3.070 2643.025 3161.730 2650.825 ;
        RECT 4.400 2641.625 3161.730 2643.025 ;
        RECT 3.070 2639.805 3161.730 2641.625 ;
        RECT 4.400 2638.405 3161.730 2639.805 ;
        RECT 3.070 2636.585 3161.730 2638.405 ;
        RECT 4.400 2635.185 3161.730 2636.585 ;
        RECT 3.070 2604.815 3161.730 2635.185 ;
        RECT 3.070 2603.415 3160.600 2604.815 ;
        RECT 3.070 2601.595 3161.730 2603.415 ;
        RECT 3.070 2600.195 3160.600 2601.595 ;
        RECT 3.070 2598.375 3161.730 2600.195 ;
        RECT 3.070 2596.975 3160.600 2598.375 ;
        RECT 3.070 2589.175 3161.730 2596.975 ;
        RECT 3.070 2587.775 3160.600 2589.175 ;
        RECT 3.070 2586.415 3161.730 2587.775 ;
        RECT 3.070 2585.015 3160.600 2586.415 ;
        RECT 3.070 2583.195 3161.730 2585.015 ;
        RECT 3.070 2581.795 3160.600 2583.195 ;
        RECT 3.070 2579.975 3161.730 2581.795 ;
        RECT 3.070 2578.575 3160.600 2579.975 ;
        RECT 3.070 2567.555 3161.730 2578.575 ;
        RECT 3.070 2566.155 3160.600 2567.555 ;
        RECT 3.070 2564.795 3161.730 2566.155 ;
        RECT 3.070 2563.395 3160.600 2564.795 ;
        RECT 3.070 2561.575 3161.730 2563.395 ;
        RECT 3.070 2560.175 3160.600 2561.575 ;
        RECT 3.070 2558.355 3161.730 2560.175 ;
        RECT 3.070 2556.955 3160.600 2558.355 ;
        RECT 3.070 2552.375 3161.730 2556.955 ;
        RECT 3.070 2550.975 3160.600 2552.375 ;
        RECT 3.070 2546.395 3161.730 2550.975 ;
        RECT 3.070 2544.995 3160.600 2546.395 ;
        RECT 3.070 2543.175 3161.730 2544.995 ;
        RECT 3.070 2541.775 3160.600 2543.175 ;
        RECT 3.070 2539.955 3161.730 2541.775 ;
        RECT 3.070 2538.555 3160.600 2539.955 ;
        RECT 3.070 2533.975 3161.730 2538.555 ;
        RECT 3.070 2532.575 3160.600 2533.975 ;
        RECT 3.070 2491.425 3161.730 2532.575 ;
        RECT 4.400 2490.025 3161.730 2491.425 ;
        RECT 3.070 2485.445 3161.730 2490.025 ;
        RECT 4.400 2484.045 3161.730 2485.445 ;
        RECT 3.070 2482.225 3161.730 2484.045 ;
        RECT 4.400 2480.825 3161.730 2482.225 ;
        RECT 3.070 2479.005 3161.730 2480.825 ;
        RECT 4.400 2477.605 3161.730 2479.005 ;
        RECT 3.070 2473.025 3161.730 2477.605 ;
        RECT 4.400 2471.625 3161.730 2473.025 ;
        RECT 3.070 2467.045 3161.730 2471.625 ;
        RECT 4.400 2465.645 3161.730 2467.045 ;
        RECT 3.070 2463.825 3161.730 2465.645 ;
        RECT 4.400 2462.425 3161.730 2463.825 ;
        RECT 3.070 2460.605 3161.730 2462.425 ;
        RECT 4.400 2459.205 3161.730 2460.605 ;
        RECT 3.070 2457.845 3161.730 2459.205 ;
        RECT 4.400 2456.445 3161.730 2457.845 ;
        RECT 3.070 2445.425 3161.730 2456.445 ;
        RECT 4.400 2444.025 3161.730 2445.425 ;
        RECT 3.070 2442.205 3161.730 2444.025 ;
        RECT 4.400 2440.805 3161.730 2442.205 ;
        RECT 3.070 2438.985 3161.730 2440.805 ;
        RECT 4.400 2437.585 3161.730 2438.985 ;
        RECT 3.070 2436.225 3161.730 2437.585 ;
        RECT 4.400 2434.825 3161.730 2436.225 ;
        RECT 3.070 2427.025 3161.730 2434.825 ;
        RECT 4.400 2425.625 3161.730 2427.025 ;
        RECT 3.070 2423.805 3161.730 2425.625 ;
        RECT 4.400 2422.405 3161.730 2423.805 ;
        RECT 3.070 2420.585 3161.730 2422.405 ;
        RECT 4.400 2419.185 3161.730 2420.585 ;
        RECT 3.070 1853.425 3161.730 2419.185 ;
        RECT 4.400 1852.025 3161.730 1853.425 ;
        RECT 3.070 1847.445 3161.730 1852.025 ;
        RECT 4.400 1846.045 3161.730 1847.445 ;
        RECT 3.070 1844.225 3161.730 1846.045 ;
        RECT 4.400 1842.825 3161.730 1844.225 ;
        RECT 3.070 1841.005 3161.730 1842.825 ;
        RECT 4.400 1839.605 3161.730 1841.005 ;
        RECT 3.070 1835.025 3161.730 1839.605 ;
        RECT 4.400 1833.625 3161.730 1835.025 ;
        RECT 3.070 1829.045 3161.730 1833.625 ;
        RECT 4.400 1827.645 3161.730 1829.045 ;
        RECT 3.070 1825.825 3161.730 1827.645 ;
        RECT 4.400 1824.425 3161.730 1825.825 ;
        RECT 3.070 1822.605 3161.730 1824.425 ;
        RECT 4.400 1821.205 3161.730 1822.605 ;
        RECT 3.070 1819.845 3161.730 1821.205 ;
        RECT 4.400 1818.445 3161.730 1819.845 ;
        RECT 3.070 1807.425 3161.730 1818.445 ;
        RECT 4.400 1806.025 3161.730 1807.425 ;
        RECT 3.070 1804.205 3161.730 1806.025 ;
        RECT 4.400 1802.805 3161.730 1804.205 ;
        RECT 3.070 1800.985 3161.730 1802.805 ;
        RECT 4.400 1799.585 3161.730 1800.985 ;
        RECT 3.070 1798.225 3161.730 1799.585 ;
        RECT 4.400 1796.825 3161.730 1798.225 ;
        RECT 3.070 1789.025 3161.730 1796.825 ;
        RECT 4.400 1787.625 3161.730 1789.025 ;
        RECT 3.070 1785.805 3161.730 1787.625 ;
        RECT 4.400 1784.405 3161.730 1785.805 ;
        RECT 3.070 1782.585 3161.730 1784.405 ;
        RECT 4.400 1781.185 3161.730 1782.585 ;
        RECT 3.070 1718.815 3161.730 1781.185 ;
        RECT 3.070 1717.415 3160.600 1718.815 ;
        RECT 3.070 1715.595 3161.730 1717.415 ;
        RECT 3.070 1714.195 3160.600 1715.595 ;
        RECT 3.070 1712.375 3161.730 1714.195 ;
        RECT 3.070 1710.975 3160.600 1712.375 ;
        RECT 3.070 1703.175 3161.730 1710.975 ;
        RECT 3.070 1701.775 3160.600 1703.175 ;
        RECT 3.070 1700.415 3161.730 1701.775 ;
        RECT 3.070 1699.015 3160.600 1700.415 ;
        RECT 3.070 1697.195 3161.730 1699.015 ;
        RECT 3.070 1695.795 3160.600 1697.195 ;
        RECT 3.070 1693.975 3161.730 1695.795 ;
        RECT 3.070 1692.575 3160.600 1693.975 ;
        RECT 3.070 1681.555 3161.730 1692.575 ;
        RECT 3.070 1680.155 3160.600 1681.555 ;
        RECT 3.070 1678.795 3161.730 1680.155 ;
        RECT 3.070 1677.395 3160.600 1678.795 ;
        RECT 3.070 1675.575 3161.730 1677.395 ;
        RECT 3.070 1674.175 3160.600 1675.575 ;
        RECT 3.070 1672.355 3161.730 1674.175 ;
        RECT 3.070 1670.955 3160.600 1672.355 ;
        RECT 3.070 1666.375 3161.730 1670.955 ;
        RECT 3.070 1664.975 3160.600 1666.375 ;
        RECT 3.070 1657.175 3161.730 1664.975 ;
        RECT 3.070 1655.775 3160.600 1657.175 ;
        RECT 3.070 1653.955 3161.730 1655.775 ;
        RECT 3.070 1652.555 3160.600 1653.955 ;
        RECT 3.070 1647.975 3161.730 1652.555 ;
        RECT 3.070 1646.575 3160.600 1647.975 ;
        RECT 3.070 1637.425 3161.730 1646.575 ;
        RECT 4.400 1636.025 3161.730 1637.425 ;
        RECT 3.070 1631.445 3161.730 1636.025 ;
        RECT 4.400 1630.045 3161.730 1631.445 ;
        RECT 3.070 1628.225 3161.730 1630.045 ;
        RECT 4.400 1626.825 3161.730 1628.225 ;
        RECT 3.070 1625.005 3161.730 1626.825 ;
        RECT 4.400 1623.605 3161.730 1625.005 ;
        RECT 3.070 1619.025 3161.730 1623.605 ;
        RECT 4.400 1617.625 3161.730 1619.025 ;
        RECT 3.070 1613.045 3161.730 1617.625 ;
        RECT 4.400 1611.645 3161.730 1613.045 ;
        RECT 3.070 1609.825 3161.730 1611.645 ;
        RECT 4.400 1608.425 3161.730 1609.825 ;
        RECT 3.070 1606.605 3161.730 1608.425 ;
        RECT 4.400 1605.205 3161.730 1606.605 ;
        RECT 3.070 1603.845 3161.730 1605.205 ;
        RECT 4.400 1602.445 3161.730 1603.845 ;
        RECT 3.070 1591.425 3161.730 1602.445 ;
        RECT 4.400 1590.025 3161.730 1591.425 ;
        RECT 3.070 1588.205 3161.730 1590.025 ;
        RECT 4.400 1586.805 3161.730 1588.205 ;
        RECT 3.070 1584.985 3161.730 1586.805 ;
        RECT 4.400 1583.585 3161.730 1584.985 ;
        RECT 3.070 1582.225 3161.730 1583.585 ;
        RECT 4.400 1580.825 3161.730 1582.225 ;
        RECT 3.070 1573.025 3161.730 1580.825 ;
        RECT 4.400 1571.625 3161.730 1573.025 ;
        RECT 3.070 1569.805 3161.730 1571.625 ;
        RECT 4.400 1568.405 3161.730 1569.805 ;
        RECT 3.070 1566.585 3161.730 1568.405 ;
        RECT 4.400 1565.185 3161.730 1566.585 ;
        RECT 3.070 1492.815 3161.730 1565.185 ;
        RECT 3.070 1491.415 3160.600 1492.815 ;
        RECT 3.070 1489.595 3161.730 1491.415 ;
        RECT 3.070 1488.195 3160.600 1489.595 ;
        RECT 3.070 1486.375 3161.730 1488.195 ;
        RECT 3.070 1484.975 3160.600 1486.375 ;
        RECT 3.070 1477.175 3161.730 1484.975 ;
        RECT 3.070 1475.775 3160.600 1477.175 ;
        RECT 3.070 1474.415 3161.730 1475.775 ;
        RECT 3.070 1473.015 3160.600 1474.415 ;
        RECT 3.070 1471.195 3161.730 1473.015 ;
        RECT 3.070 1469.795 3160.600 1471.195 ;
        RECT 3.070 1467.975 3161.730 1469.795 ;
        RECT 3.070 1466.575 3160.600 1467.975 ;
        RECT 3.070 1455.555 3161.730 1466.575 ;
        RECT 3.070 1454.155 3160.600 1455.555 ;
        RECT 3.070 1452.795 3161.730 1454.155 ;
        RECT 3.070 1451.395 3160.600 1452.795 ;
        RECT 3.070 1449.575 3161.730 1451.395 ;
        RECT 3.070 1448.175 3160.600 1449.575 ;
        RECT 3.070 1446.355 3161.730 1448.175 ;
        RECT 3.070 1444.955 3160.600 1446.355 ;
        RECT 3.070 1440.375 3161.730 1444.955 ;
        RECT 3.070 1438.975 3160.600 1440.375 ;
        RECT 3.070 1431.175 3161.730 1438.975 ;
        RECT 3.070 1429.775 3160.600 1431.175 ;
        RECT 3.070 1427.955 3161.730 1429.775 ;
        RECT 3.070 1426.555 3160.600 1427.955 ;
        RECT 3.070 1421.975 3161.730 1426.555 ;
        RECT 3.070 1421.425 3160.600 1421.975 ;
        RECT 4.400 1420.575 3160.600 1421.425 ;
        RECT 4.400 1420.025 3161.730 1420.575 ;
        RECT 3.070 1415.445 3161.730 1420.025 ;
        RECT 4.400 1414.045 3161.730 1415.445 ;
        RECT 3.070 1412.225 3161.730 1414.045 ;
        RECT 4.400 1410.825 3161.730 1412.225 ;
        RECT 3.070 1409.005 3161.730 1410.825 ;
        RECT 4.400 1407.605 3161.730 1409.005 ;
        RECT 3.070 1403.025 3161.730 1407.605 ;
        RECT 4.400 1401.625 3161.730 1403.025 ;
        RECT 3.070 1397.045 3161.730 1401.625 ;
        RECT 4.400 1395.645 3161.730 1397.045 ;
        RECT 3.070 1393.825 3161.730 1395.645 ;
        RECT 4.400 1392.425 3161.730 1393.825 ;
        RECT 3.070 1390.605 3161.730 1392.425 ;
        RECT 4.400 1389.205 3161.730 1390.605 ;
        RECT 3.070 1387.845 3161.730 1389.205 ;
        RECT 4.400 1386.445 3161.730 1387.845 ;
        RECT 3.070 1375.425 3161.730 1386.445 ;
        RECT 4.400 1374.025 3161.730 1375.425 ;
        RECT 3.070 1372.205 3161.730 1374.025 ;
        RECT 4.400 1370.805 3161.730 1372.205 ;
        RECT 3.070 1368.985 3161.730 1370.805 ;
        RECT 4.400 1367.585 3161.730 1368.985 ;
        RECT 3.070 1366.225 3161.730 1367.585 ;
        RECT 4.400 1364.825 3161.730 1366.225 ;
        RECT 3.070 1357.025 3161.730 1364.825 ;
        RECT 4.400 1355.625 3161.730 1357.025 ;
        RECT 3.070 1353.805 3161.730 1355.625 ;
        RECT 4.400 1352.405 3161.730 1353.805 ;
        RECT 3.070 1350.585 3161.730 1352.405 ;
        RECT 4.690 1349.185 3161.730 1350.585 ;
        RECT 3.070 1267.815 3161.730 1349.185 ;
        RECT 3.070 1266.415 3160.600 1267.815 ;
        RECT 3.070 1264.595 3161.730 1266.415 ;
        RECT 3.070 1263.195 3160.600 1264.595 ;
        RECT 3.070 1261.375 3161.730 1263.195 ;
        RECT 3.070 1259.975 3160.600 1261.375 ;
        RECT 3.070 1252.175 3161.730 1259.975 ;
        RECT 3.070 1250.775 3160.600 1252.175 ;
        RECT 3.070 1249.415 3161.730 1250.775 ;
        RECT 3.070 1248.015 3160.600 1249.415 ;
        RECT 3.070 1246.195 3161.730 1248.015 ;
        RECT 3.070 1244.795 3160.600 1246.195 ;
        RECT 3.070 1242.975 3161.730 1244.795 ;
        RECT 3.070 1241.575 3160.600 1242.975 ;
        RECT 3.070 1230.555 3161.730 1241.575 ;
        RECT 3.070 1229.155 3160.600 1230.555 ;
        RECT 3.070 1227.795 3161.730 1229.155 ;
        RECT 3.070 1226.395 3160.600 1227.795 ;
        RECT 3.070 1224.575 3161.730 1226.395 ;
        RECT 3.070 1223.175 3160.600 1224.575 ;
        RECT 3.070 1221.355 3161.730 1223.175 ;
        RECT 3.070 1219.955 3160.600 1221.355 ;
        RECT 3.070 1215.375 3161.730 1219.955 ;
        RECT 3.070 1213.975 3160.600 1215.375 ;
        RECT 3.070 1206.175 3161.730 1213.975 ;
        RECT 3.070 1205.425 3160.600 1206.175 ;
        RECT 4.400 1204.775 3160.600 1205.425 ;
        RECT 4.400 1204.025 3161.730 1204.775 ;
        RECT 3.070 1202.955 3161.730 1204.025 ;
        RECT 3.070 1201.555 3160.600 1202.955 ;
        RECT 3.070 1199.445 3161.730 1201.555 ;
        RECT 4.690 1198.045 3161.730 1199.445 ;
        RECT 3.070 1196.975 3161.730 1198.045 ;
        RECT 3.070 1196.225 3160.600 1196.975 ;
        RECT 4.400 1195.575 3160.600 1196.225 ;
        RECT 4.400 1194.825 3161.730 1195.575 ;
        RECT 3.070 1193.005 3161.730 1194.825 ;
        RECT 4.400 1191.605 3161.730 1193.005 ;
        RECT 3.070 1187.025 3161.730 1191.605 ;
        RECT 4.400 1185.625 3161.730 1187.025 ;
        RECT 3.070 1181.045 3161.730 1185.625 ;
        RECT 4.400 1179.645 3161.730 1181.045 ;
        RECT 3.070 1177.825 3161.730 1179.645 ;
        RECT 4.400 1176.425 3161.730 1177.825 ;
        RECT 3.070 1174.605 3161.730 1176.425 ;
        RECT 4.400 1173.205 3161.730 1174.605 ;
        RECT 3.070 1171.845 3161.730 1173.205 ;
        RECT 4.400 1170.445 3161.730 1171.845 ;
        RECT 3.070 1159.425 3161.730 1170.445 ;
        RECT 4.400 1158.025 3161.730 1159.425 ;
        RECT 3.070 1156.205 3161.730 1158.025 ;
        RECT 4.400 1154.805 3161.730 1156.205 ;
        RECT 3.070 1152.985 3161.730 1154.805 ;
        RECT 4.400 1151.585 3161.730 1152.985 ;
        RECT 3.070 1150.225 3161.730 1151.585 ;
        RECT 4.400 1148.825 3161.730 1150.225 ;
        RECT 3.070 1141.025 3161.730 1148.825 ;
        RECT 4.400 1139.625 3161.730 1141.025 ;
        RECT 3.070 1137.805 3161.730 1139.625 ;
        RECT 4.400 1136.405 3161.730 1137.805 ;
        RECT 3.070 1134.585 3161.730 1136.405 ;
        RECT 4.400 1133.185 3161.730 1134.585 ;
        RECT 3.070 1042.815 3161.730 1133.185 ;
        RECT 3.070 1041.415 3160.600 1042.815 ;
        RECT 3.070 1039.595 3161.730 1041.415 ;
        RECT 3.070 1038.195 3160.600 1039.595 ;
        RECT 3.070 1036.375 3161.730 1038.195 ;
        RECT 3.070 1034.975 3160.600 1036.375 ;
        RECT 3.070 1027.175 3161.730 1034.975 ;
        RECT 3.070 1025.775 3160.600 1027.175 ;
        RECT 3.070 1024.415 3161.730 1025.775 ;
        RECT 3.070 1023.015 3160.600 1024.415 ;
        RECT 3.070 1021.195 3161.730 1023.015 ;
        RECT 3.070 1019.795 3160.600 1021.195 ;
        RECT 3.070 1017.975 3161.730 1019.795 ;
        RECT 3.070 1016.575 3160.600 1017.975 ;
        RECT 3.070 1005.555 3161.730 1016.575 ;
        RECT 3.070 1004.155 3160.600 1005.555 ;
        RECT 3.070 1002.795 3161.730 1004.155 ;
        RECT 3.070 1001.395 3160.600 1002.795 ;
        RECT 3.070 999.575 3161.730 1001.395 ;
        RECT 3.070 998.175 3160.600 999.575 ;
        RECT 3.070 996.355 3161.730 998.175 ;
        RECT 3.070 994.955 3160.600 996.355 ;
        RECT 3.070 990.375 3161.730 994.955 ;
        RECT 3.070 989.425 3160.600 990.375 ;
        RECT 4.400 988.975 3160.600 989.425 ;
        RECT 4.400 988.025 3161.730 988.975 ;
        RECT 3.070 983.445 3161.730 988.025 ;
        RECT 4.400 982.045 3161.730 983.445 ;
        RECT 3.070 981.175 3161.730 982.045 ;
        RECT 3.070 980.225 3160.600 981.175 ;
        RECT 4.400 979.775 3160.600 980.225 ;
        RECT 4.400 978.825 3161.730 979.775 ;
        RECT 3.070 977.955 3161.730 978.825 ;
        RECT 3.070 976.555 3160.600 977.955 ;
        RECT 3.070 971.975 3161.730 976.555 ;
        RECT 3.070 971.025 3160.600 971.975 ;
        RECT 4.400 970.575 3160.600 971.025 ;
        RECT 4.400 969.625 3161.730 970.575 ;
        RECT 3.070 965.045 3161.730 969.625 ;
        RECT 4.400 963.645 3161.730 965.045 ;
        RECT 3.070 961.825 3161.730 963.645 ;
        RECT 4.400 960.425 3161.730 961.825 ;
        RECT 3.070 958.605 3161.730 960.425 ;
        RECT 4.400 957.205 3161.730 958.605 ;
        RECT 3.070 955.845 3161.730 957.205 ;
        RECT 4.400 954.445 3161.730 955.845 ;
        RECT 3.070 943.425 3161.730 954.445 ;
        RECT 4.400 942.025 3161.730 943.425 ;
        RECT 3.070 940.205 3161.730 942.025 ;
        RECT 4.400 938.805 3161.730 940.205 ;
        RECT 3.070 936.985 3161.730 938.805 ;
        RECT 4.400 935.585 3161.730 936.985 ;
        RECT 3.070 934.225 3161.730 935.585 ;
        RECT 4.400 932.825 3161.730 934.225 ;
        RECT 3.070 925.025 3161.730 932.825 ;
        RECT 4.400 923.625 3161.730 925.025 ;
        RECT 3.070 921.805 3161.730 923.625 ;
        RECT 4.400 920.405 3161.730 921.805 ;
        RECT 3.070 918.585 3161.730 920.405 ;
        RECT 4.400 917.185 3161.730 918.585 ;
        RECT 3.070 816.815 3161.730 917.185 ;
        RECT 3.070 815.415 3160.600 816.815 ;
        RECT 3.070 813.595 3161.730 815.415 ;
        RECT 3.070 812.195 3160.600 813.595 ;
        RECT 3.070 810.375 3161.730 812.195 ;
        RECT 3.070 808.975 3160.600 810.375 ;
        RECT 3.070 801.175 3161.730 808.975 ;
        RECT 3.070 799.775 3160.600 801.175 ;
        RECT 3.070 798.415 3161.730 799.775 ;
        RECT 3.070 797.015 3160.600 798.415 ;
        RECT 3.070 795.195 3161.730 797.015 ;
        RECT 3.070 793.795 3160.600 795.195 ;
        RECT 3.070 791.975 3161.730 793.795 ;
        RECT 3.070 790.575 3160.600 791.975 ;
        RECT 3.070 779.555 3161.730 790.575 ;
        RECT 3.070 778.155 3160.600 779.555 ;
        RECT 3.070 776.795 3161.730 778.155 ;
        RECT 3.070 775.395 3160.600 776.795 ;
        RECT 3.070 773.575 3161.730 775.395 ;
        RECT 3.070 773.425 3160.600 773.575 ;
        RECT 4.400 772.175 3160.600 773.425 ;
        RECT 4.400 772.025 3161.730 772.175 ;
        RECT 3.070 770.355 3161.730 772.025 ;
        RECT 3.070 768.955 3160.600 770.355 ;
        RECT 3.070 767.445 3161.730 768.955 ;
        RECT 4.400 766.045 3161.730 767.445 ;
        RECT 3.070 764.375 3161.730 766.045 ;
        RECT 3.070 764.225 3160.600 764.375 ;
        RECT 4.400 762.975 3160.600 764.225 ;
        RECT 4.400 762.825 3161.730 762.975 ;
        RECT 3.070 755.175 3161.730 762.825 ;
        RECT 3.070 755.025 3160.600 755.175 ;
        RECT 4.400 753.775 3160.600 755.025 ;
        RECT 4.400 753.625 3161.730 753.775 ;
        RECT 3.070 751.955 3161.730 753.625 ;
        RECT 3.070 750.555 3160.600 751.955 ;
        RECT 3.070 749.045 3161.730 750.555 ;
        RECT 4.400 747.645 3161.730 749.045 ;
        RECT 3.070 745.975 3161.730 747.645 ;
        RECT 3.070 745.825 3160.600 745.975 ;
        RECT 4.400 744.575 3160.600 745.825 ;
        RECT 4.400 744.425 3161.730 744.575 ;
        RECT 3.070 742.605 3161.730 744.425 ;
        RECT 4.400 741.205 3161.730 742.605 ;
        RECT 3.070 739.845 3161.730 741.205 ;
        RECT 4.400 738.445 3161.730 739.845 ;
        RECT 3.070 727.425 3161.730 738.445 ;
        RECT 4.400 726.025 3161.730 727.425 ;
        RECT 3.070 724.205 3161.730 726.025 ;
        RECT 4.400 722.805 3161.730 724.205 ;
        RECT 3.070 720.985 3161.730 722.805 ;
        RECT 4.400 719.585 3161.730 720.985 ;
        RECT 3.070 718.225 3161.730 719.585 ;
        RECT 4.400 716.825 3161.730 718.225 ;
        RECT 3.070 709.025 3161.730 716.825 ;
        RECT 4.400 707.625 3161.730 709.025 ;
        RECT 3.070 705.805 3161.730 707.625 ;
        RECT 4.400 704.405 3161.730 705.805 ;
        RECT 3.070 702.585 3161.730 704.405 ;
        RECT 4.400 701.185 3161.730 702.585 ;
        RECT 3.070 591.815 3161.730 701.185 ;
        RECT 3.070 590.415 3160.600 591.815 ;
        RECT 3.070 588.595 3161.730 590.415 ;
        RECT 3.070 587.195 3160.600 588.595 ;
        RECT 3.070 585.375 3161.730 587.195 ;
        RECT 3.070 583.975 3160.600 585.375 ;
        RECT 3.070 576.175 3161.730 583.975 ;
        RECT 3.070 574.775 3160.600 576.175 ;
        RECT 3.070 573.415 3161.730 574.775 ;
        RECT 3.070 572.015 3160.600 573.415 ;
        RECT 3.070 570.195 3161.730 572.015 ;
        RECT 3.070 568.795 3160.600 570.195 ;
        RECT 3.070 566.975 3161.730 568.795 ;
        RECT 3.070 565.575 3160.600 566.975 ;
        RECT 3.070 554.555 3161.730 565.575 ;
        RECT 3.070 553.155 3160.600 554.555 ;
        RECT 3.070 551.795 3161.730 553.155 ;
        RECT 3.070 550.395 3160.600 551.795 ;
        RECT 3.070 548.575 3161.730 550.395 ;
        RECT 3.070 547.175 3160.600 548.575 ;
        RECT 3.070 545.355 3161.730 547.175 ;
        RECT 3.070 543.955 3160.600 545.355 ;
        RECT 3.070 539.375 3161.730 543.955 ;
        RECT 3.070 537.975 3160.600 539.375 ;
        RECT 3.070 530.175 3161.730 537.975 ;
        RECT 3.070 528.775 3160.600 530.175 ;
        RECT 3.070 526.955 3161.730 528.775 ;
        RECT 3.070 525.555 3160.600 526.955 ;
        RECT 3.070 520.975 3161.730 525.555 ;
        RECT 3.070 519.575 3160.600 520.975 ;
        RECT 3.070 365.815 3161.730 519.575 ;
        RECT 3.070 364.415 3160.600 365.815 ;
        RECT 3.070 362.595 3161.730 364.415 ;
        RECT 3.070 361.195 3160.600 362.595 ;
        RECT 3.070 359.375 3161.730 361.195 ;
        RECT 3.070 357.975 3160.600 359.375 ;
        RECT 3.070 350.175 3161.730 357.975 ;
        RECT 3.070 348.775 3160.600 350.175 ;
        RECT 3.070 347.415 3161.730 348.775 ;
        RECT 3.070 346.015 3160.600 347.415 ;
        RECT 3.070 344.195 3161.730 346.015 ;
        RECT 3.070 342.795 3160.600 344.195 ;
        RECT 3.070 340.975 3161.730 342.795 ;
        RECT 3.070 339.575 3160.600 340.975 ;
        RECT 3.070 328.555 3161.730 339.575 ;
        RECT 3.070 327.155 3160.600 328.555 ;
        RECT 3.070 325.795 3161.730 327.155 ;
        RECT 3.070 324.395 3160.600 325.795 ;
        RECT 3.070 322.575 3161.730 324.395 ;
        RECT 3.070 321.175 3160.600 322.575 ;
        RECT 3.070 319.355 3161.730 321.175 ;
        RECT 3.070 317.955 3160.600 319.355 ;
        RECT 3.070 313.375 3161.730 317.955 ;
        RECT 3.070 311.975 3160.600 313.375 ;
        RECT 3.070 304.175 3161.730 311.975 ;
        RECT 3.070 302.775 3160.600 304.175 ;
        RECT 3.070 300.955 3161.730 302.775 ;
        RECT 3.070 299.555 3160.600 300.955 ;
        RECT 3.070 294.975 3161.730 299.555 ;
        RECT 3.070 293.575 3160.600 294.975 ;
        RECT 3.070 10.715 3161.730 293.575 ;
      LAYER met4 ;
        RECT 78.110 4595.900 125.120 4678.225 ;
        RECT 129.120 4595.900 134.720 4678.225 ;
        RECT 138.720 4595.900 225.120 4678.225 ;
        RECT 229.120 4595.900 234.720 4678.225 ;
        RECT 238.720 4595.900 258.040 4678.225 ;
        RECT 260.440 4595.900 261.840 4678.225 ;
        RECT 264.240 4595.900 325.120 4678.225 ;
        RECT 329.120 4595.900 334.720 4678.225 ;
        RECT 338.720 4595.900 425.120 4678.225 ;
        RECT 429.120 4595.900 434.720 4678.225 ;
        RECT 438.720 4595.900 525.120 4678.225 ;
        RECT 529.120 4595.900 534.720 4678.225 ;
        RECT 538.720 4595.900 558.040 4678.225 ;
        RECT 560.440 4595.900 561.840 4678.225 ;
        RECT 564.240 4595.900 625.120 4678.225 ;
        RECT 629.120 4602.950 634.720 4678.225 ;
        RECT 638.720 4602.950 725.120 4678.225 ;
        RECT 729.120 4602.950 734.720 4678.225 ;
        RECT 629.120 4595.900 734.720 4602.950 ;
        RECT 738.720 4595.900 825.120 4678.225 ;
        RECT 829.120 4595.900 834.720 4678.225 ;
        RECT 838.720 4595.900 858.040 4678.225 ;
        RECT 860.440 4595.900 861.840 4678.225 ;
        RECT 864.240 4595.900 925.120 4678.225 ;
        RECT 929.120 4595.900 934.720 4678.225 ;
        RECT 938.720 4595.900 1025.120 4678.225 ;
        RECT 1029.120 4595.900 1034.720 4678.225 ;
        RECT 1038.720 4595.900 1125.120 4678.225 ;
        RECT 1129.120 4595.900 1134.720 4678.225 ;
        RECT 1138.720 4595.900 1158.040 4678.225 ;
        RECT 1160.440 4595.900 1161.840 4678.225 ;
        RECT 1164.240 4595.900 1225.120 4678.225 ;
        RECT 1229.120 4595.900 1234.720 4678.225 ;
        RECT 1238.720 4595.900 1325.120 4678.225 ;
        RECT 1329.120 4595.900 1334.720 4678.225 ;
        RECT 1338.720 4595.900 1425.120 4678.225 ;
        RECT 1429.120 4595.900 1434.720 4678.225 ;
        RECT 1438.720 4595.900 1458.040 4678.225 ;
        RECT 1460.440 4595.900 1461.840 4678.225 ;
        RECT 1464.240 4595.900 1525.120 4678.225 ;
        RECT 1529.120 4602.950 1534.720 4678.225 ;
        RECT 1538.720 4602.950 1625.120 4678.225 ;
        RECT 1629.120 4602.950 1634.720 4678.225 ;
        RECT 1529.120 4595.900 1634.720 4602.950 ;
        RECT 1638.720 4595.900 1725.120 4678.225 ;
        RECT 1729.120 4595.900 1734.720 4678.225 ;
        RECT 1738.720 4595.900 1758.040 4678.225 ;
        RECT 1760.440 4595.900 1761.840 4678.225 ;
        RECT 1764.240 4595.900 1825.120 4678.225 ;
        RECT 1829.120 4595.900 1834.720 4678.225 ;
        RECT 1838.720 4595.900 1925.120 4678.225 ;
        RECT 1929.120 4595.900 1934.720 4678.225 ;
        RECT 1938.720 4595.900 2025.120 4678.225 ;
        RECT 2029.120 4595.900 2034.720 4678.225 ;
        RECT 2038.720 4595.900 2058.040 4678.225 ;
        RECT 2060.440 4595.900 2061.840 4678.225 ;
        RECT 2064.240 4595.900 2125.120 4678.225 ;
        RECT 2129.120 4595.900 2134.720 4678.225 ;
        RECT 2138.720 4595.900 2225.120 4678.225 ;
        RECT 2229.120 4595.900 2234.720 4678.225 ;
        RECT 2238.720 4595.900 2325.120 4678.225 ;
        RECT 2329.120 4595.900 2334.720 4678.225 ;
        RECT 2338.720 4595.900 2358.040 4678.225 ;
        RECT 2360.440 4595.900 2361.840 4678.225 ;
        RECT 2364.240 4595.900 2425.120 4678.225 ;
        RECT 2429.120 4602.950 2434.720 4678.225 ;
        RECT 2438.720 4602.950 2525.120 4678.225 ;
        RECT 2529.120 4602.950 2534.720 4678.225 ;
        RECT 2429.120 4595.900 2534.720 4602.950 ;
        RECT 2538.720 4595.900 2625.120 4678.225 ;
        RECT 2629.120 4595.900 2634.720 4678.225 ;
        RECT 2638.720 4595.900 2658.040 4678.225 ;
        RECT 2660.440 4595.900 2661.840 4678.225 ;
        RECT 2664.240 4595.900 2725.120 4678.225 ;
        RECT 2729.120 4595.900 2734.720 4678.225 ;
        RECT 2738.720 4595.900 2825.120 4678.225 ;
        RECT 2829.120 4595.900 2834.720 4678.225 ;
        RECT 2838.720 4595.900 2925.120 4678.225 ;
        RECT 2929.120 4595.900 2934.720 4678.225 ;
        RECT 2938.720 4595.900 3025.120 4678.225 ;
        RECT 3029.120 4595.900 3034.720 4678.225 ;
        RECT 3038.720 4595.900 3084.990 4678.225 ;
        RECT 78.110 989.400 3084.990 4595.900 ;
        RECT 78.110 669.485 125.120 989.400 ;
        RECT 129.120 669.485 134.720 989.400 ;
        RECT 138.720 669.485 225.120 989.400 ;
        RECT 229.120 669.485 234.720 989.400 ;
        RECT 238.720 669.485 325.120 989.400 ;
        RECT 329.120 669.485 334.720 989.400 ;
        RECT 338.720 669.485 425.120 989.400 ;
        RECT 429.120 669.485 434.720 989.400 ;
        RECT 438.720 669.485 525.120 989.400 ;
        RECT 529.120 669.485 534.720 989.400 ;
        RECT 538.720 669.485 625.120 989.400 ;
        RECT 629.120 669.485 634.720 989.400 ;
        RECT 638.720 676.700 725.120 989.400 ;
        RECT 729.120 676.700 734.720 989.400 ;
        RECT 638.720 669.485 734.720 676.700 ;
        RECT 738.720 669.485 825.120 989.400 ;
        RECT 829.120 669.485 834.720 989.400 ;
        RECT 838.720 669.485 858.040 989.400 ;
        RECT 860.440 669.485 861.840 989.400 ;
        RECT 864.240 935.805 925.120 989.400 ;
        RECT 929.120 935.805 934.720 989.400 ;
        RECT 938.720 935.805 1025.120 989.400 ;
        RECT 1029.120 935.805 1034.720 989.400 ;
        RECT 1038.720 935.805 1125.120 989.400 ;
        RECT 1129.120 935.805 1134.720 989.400 ;
        RECT 1138.720 935.805 1225.120 989.400 ;
        RECT 1229.120 935.805 1234.720 989.400 ;
        RECT 1238.720 935.805 1325.120 989.400 ;
        RECT 1329.120 935.805 1334.720 989.400 ;
        RECT 1338.720 935.805 1425.120 989.400 ;
        RECT 1429.120 935.805 1434.720 989.400 ;
        RECT 1438.720 935.805 1525.120 989.400 ;
        RECT 1529.120 935.805 1534.720 989.400 ;
        RECT 1538.720 935.805 1625.120 989.400 ;
        RECT 1629.120 935.805 1634.720 989.400 ;
        RECT 1638.720 935.805 1725.120 989.400 ;
        RECT 1729.120 935.805 1734.720 989.400 ;
        RECT 1738.720 935.805 1825.120 989.400 ;
        RECT 1829.120 935.805 1834.720 989.400 ;
        RECT 1838.720 935.805 1925.120 989.400 ;
        RECT 1929.120 935.805 1934.720 989.400 ;
        RECT 1938.720 935.805 2025.120 989.400 ;
        RECT 2029.120 935.805 2034.720 989.400 ;
        RECT 2038.720 935.805 2125.120 989.400 ;
        RECT 864.240 780.275 2125.120 935.805 ;
        RECT 864.240 669.485 925.120 780.275 ;
        RECT 78.110 169.875 925.120 669.485 ;
        RECT 78.110 25.335 125.120 169.875 ;
        RECT 129.120 25.335 134.720 169.875 ;
        RECT 138.720 25.335 225.120 169.875 ;
        RECT 229.120 25.335 234.720 169.875 ;
        RECT 238.720 25.335 325.120 169.875 ;
        RECT 329.120 25.335 334.720 169.875 ;
        RECT 338.720 25.335 425.120 169.875 ;
        RECT 429.120 25.335 434.720 169.875 ;
        RECT 438.720 25.335 525.120 169.875 ;
        RECT 529.120 25.335 534.720 169.875 ;
        RECT 538.720 25.335 625.120 169.875 ;
        RECT 629.120 25.335 634.720 169.875 ;
        RECT 638.720 132.740 734.720 169.875 ;
        RECT 638.720 25.335 725.120 132.740 ;
        RECT 729.120 25.335 734.720 132.740 ;
        RECT 738.720 25.335 825.120 169.875 ;
        RECT 829.120 25.335 834.720 169.875 ;
        RECT 838.720 25.335 925.120 169.875 ;
        RECT 929.120 25.335 934.720 780.275 ;
        RECT 938.720 25.335 1025.120 780.275 ;
        RECT 1029.120 25.335 1034.720 780.275 ;
        RECT 1038.720 25.335 1125.120 780.275 ;
        RECT 1129.120 25.335 1134.720 780.275 ;
        RECT 1138.720 25.335 1225.120 780.275 ;
        RECT 1229.120 25.335 1234.720 780.275 ;
        RECT 1238.720 25.335 1325.120 780.275 ;
        RECT 1329.120 25.335 1334.720 780.275 ;
        RECT 1338.720 25.335 1425.120 780.275 ;
        RECT 1429.120 25.335 1434.720 780.275 ;
        RECT 1438.720 25.335 1525.120 780.275 ;
        RECT 1529.120 25.335 1534.720 780.275 ;
        RECT 1538.720 25.335 1625.120 780.275 ;
        RECT 1629.120 25.335 1634.720 780.275 ;
        RECT 1638.720 25.335 1725.120 780.275 ;
        RECT 1729.120 25.335 1734.720 780.275 ;
        RECT 1738.720 582.245 1825.120 780.275 ;
        RECT 1829.120 582.245 1834.720 780.275 ;
        RECT 1838.720 582.245 1925.120 780.275 ;
        RECT 1929.120 582.245 1934.720 780.275 ;
        RECT 1938.720 586.060 2025.120 780.275 ;
        RECT 2029.120 586.060 2034.720 780.275 ;
        RECT 1938.720 582.245 2034.720 586.060 ;
        RECT 2038.720 582.245 2125.120 780.275 ;
        RECT 2129.120 929.420 2134.720 989.400 ;
        RECT 2138.720 929.420 2225.120 989.400 ;
        RECT 2129.120 785.300 2225.120 929.420 ;
        RECT 2129.120 582.245 2134.720 785.300 ;
        RECT 2138.720 582.245 2225.120 785.300 ;
        RECT 2229.120 582.245 2234.720 989.400 ;
        RECT 2238.720 582.245 2325.120 989.400 ;
        RECT 1738.720 151.995 2325.120 582.245 ;
        RECT 1738.720 25.335 1825.120 151.995 ;
        RECT 1829.120 25.335 1834.720 151.995 ;
        RECT 1838.720 25.335 1925.120 151.995 ;
        RECT 1929.120 25.335 1934.720 151.995 ;
        RECT 1938.720 142.740 2034.720 151.995 ;
        RECT 1938.720 25.335 2025.120 142.740 ;
        RECT 2029.120 25.335 2034.720 142.740 ;
        RECT 2038.720 25.335 2125.120 151.995 ;
        RECT 2129.120 25.335 2134.720 151.995 ;
        RECT 2138.720 25.335 2225.120 151.995 ;
        RECT 2229.120 25.335 2234.720 151.995 ;
        RECT 2238.720 25.335 2325.120 151.995 ;
        RECT 2329.120 25.335 2334.720 989.400 ;
        RECT 2338.720 25.335 2358.040 989.400 ;
        RECT 2360.440 25.335 2361.840 989.400 ;
        RECT 2364.240 25.335 2425.120 989.400 ;
        RECT 2429.120 929.420 2434.720 989.400 ;
        RECT 2438.720 929.420 2525.120 989.400 ;
        RECT 2429.120 785.300 2525.120 929.420 ;
        RECT 2429.120 25.335 2434.720 785.300 ;
        RECT 2438.720 25.335 2525.120 785.300 ;
        RECT 2529.120 25.335 2534.720 989.400 ;
        RECT 2538.720 25.335 2625.120 989.400 ;
        RECT 2629.120 25.335 2634.720 989.400 ;
        RECT 2638.720 25.335 2658.040 989.400 ;
        RECT 2660.440 25.335 2661.840 989.400 ;
        RECT 2664.240 734.925 2725.120 989.400 ;
        RECT 2729.120 734.925 2734.720 989.400 ;
        RECT 2738.720 734.925 2825.120 989.400 ;
        RECT 2829.120 734.925 2834.720 989.400 ;
        RECT 2838.720 734.925 2925.120 989.400 ;
        RECT 2929.120 734.925 2934.720 989.400 ;
        RECT 2938.720 734.925 3025.120 989.400 ;
        RECT 3029.120 736.700 3034.720 989.400 ;
        RECT 3038.720 736.700 3084.990 989.400 ;
        RECT 3029.120 734.925 3084.990 736.700 ;
        RECT 2664.240 193.155 3084.990 734.925 ;
        RECT 2664.240 25.335 2725.120 193.155 ;
        RECT 2729.120 25.335 2734.720 193.155 ;
        RECT 2738.720 25.335 2825.120 193.155 ;
        RECT 2829.120 25.335 2834.720 193.155 ;
        RECT 2838.720 25.335 2925.120 193.155 ;
        RECT 2929.120 25.335 2934.720 193.155 ;
        RECT 2938.720 25.335 3025.120 193.155 ;
        RECT 3029.120 192.740 3084.990 193.155 ;
        RECT 3029.120 25.335 3034.720 192.740 ;
        RECT 3038.720 25.335 3084.990 192.740 ;
      LAYER met5 ;
        RECT 78.110 973.900 3084.990 4594.950 ;
        RECT 78.110 960.700 823.920 973.900 ;
        RECT 2239.920 960.700 3084.990 973.900 ;
        RECT 78.110 960.300 3084.990 960.700 ;
        RECT 78.110 947.100 823.920 960.300 ;
        RECT 2239.920 947.100 3084.990 960.300 ;
        RECT 78.110 924.680 3084.990 947.100 ;
        RECT 78.110 915.080 3084.990 918.280 ;
        RECT 78.110 877.880 3084.990 908.680 ;
        RECT 78.110 804.680 3084.990 813.880 ;
        RECT 78.110 795.080 3084.990 798.280 ;
        RECT 78.110 684.680 3084.990 788.680 ;
        RECT 78.110 675.080 3084.990 678.280 ;
        RECT 78.110 625.080 3084.990 668.680 ;
        RECT 78.110 613.880 3084.990 617.080 ;
        RECT 78.110 564.680 3084.990 605.880 ;
        RECT 78.110 555.080 3084.990 558.280 ;
        RECT 78.110 505.080 3084.990 548.680 ;
        RECT 78.110 493.880 3084.990 497.080 ;
        RECT 78.110 444.680 3084.990 485.880 ;
        RECT 78.110 435.080 3084.990 438.280 ;
        RECT 78.110 385.080 3084.990 428.680 ;
        RECT 78.110 373.880 3084.990 377.080 ;
        RECT 78.110 324.680 3084.990 365.880 ;
        RECT 78.110 315.080 3084.990 318.280 ;
        RECT 78.110 265.080 3084.990 308.680 ;
        RECT 78.110 253.880 3084.990 257.080 ;
        RECT 78.110 204.680 3084.990 245.880 ;
        RECT 78.110 195.080 3084.990 198.280 ;
        RECT 78.110 133.500 3084.990 188.680 ;
  END
END caravel_core
END LIBRARY

