magic
tech sky130A
magscale 1 2
timestamp 1677507470
<< viali >>
rect 3617 18377 3651 18411
rect 4629 18377 4663 18411
rect 18429 18377 18463 18411
rect 17785 18309 17819 18343
rect 4261 18241 4295 18275
rect 6653 18241 6687 18275
rect 7205 18241 7239 18275
rect 10517 18241 10551 18275
rect 14841 18241 14875 18275
rect 1593 18173 1627 18207
rect 2053 18173 2087 18207
rect 5273 18173 5307 18207
rect 6009 18173 6043 18207
rect 6837 18173 6871 18207
rect 8217 18173 8251 18207
rect 9321 18173 9355 18207
rect 11253 18173 11287 18207
rect 11713 18173 11747 18207
rect 14232 18173 14266 18207
rect 16221 18173 16255 18207
rect 17969 18173 18003 18207
rect 5733 18105 5767 18139
rect 7849 18105 7883 18139
rect 10425 18105 10459 18139
rect 1777 18037 1811 18071
rect 4629 18037 4663 18071
rect 4813 18037 4847 18071
rect 8769 18037 8803 18071
rect 9965 18037 9999 18071
rect 10333 18037 10367 18071
rect 14335 18037 14369 18071
rect 15025 18037 15059 18071
rect 15117 18037 15151 18071
rect 15485 18037 15519 18071
rect 16037 18037 16071 18071
rect 9551 17833 9585 17867
rect 5457 17765 5491 17799
rect 2083 17697 2117 17731
rect 2237 17697 2271 17731
rect 4537 17697 4571 17731
rect 7757 17697 7791 17731
rect 9965 17697 9999 17731
rect 12909 17697 12943 17731
rect 15025 17697 15059 17731
rect 8125 17629 8159 17663
rect 13369 17629 13403 17663
rect 15301 17629 15335 17663
rect 16773 17629 16807 17663
rect 17233 17629 17267 17663
rect 6745 17561 6779 17595
rect 2053 17493 2087 17527
rect 3249 17493 3283 17527
rect 11253 17493 11287 17527
rect 17877 17493 17911 17527
rect 1961 17289 1995 17323
rect 2605 17289 2639 17323
rect 12357 17289 12391 17323
rect 1731 17221 1765 17255
rect 857 17153 891 17187
rect 1869 17153 1903 17187
rect 2513 17153 2547 17187
rect 3617 17153 3651 17187
rect 6377 17153 6411 17187
rect 11253 17153 11287 17187
rect 12081 17153 12115 17187
rect 12265 17153 12299 17187
rect 13001 17153 13035 17187
rect 17509 17153 17543 17187
rect 765 17085 799 17119
rect 1593 17085 1627 17119
rect 2053 17085 2087 17119
rect 2329 17085 2363 17119
rect 2973 17085 3007 17119
rect 3157 17085 3191 17119
rect 4261 17085 4295 17119
rect 4445 17085 4479 17119
rect 4813 17085 4847 17119
rect 5273 17085 5307 17119
rect 6009 17085 6043 17119
rect 6745 17085 6779 17119
rect 11345 17085 11379 17119
rect 12357 17085 12391 17119
rect 12633 17085 12667 17119
rect 12787 17085 12821 17119
rect 13553 17085 13587 17119
rect 13737 17085 13771 17119
rect 14197 17085 14231 17119
rect 17785 17085 17819 17119
rect 2697 17017 2731 17051
rect 5825 17017 5859 17051
rect 9045 17017 9079 17051
rect 10609 17017 10643 17051
rect 14841 17017 14875 17051
rect 1133 16949 1167 16983
rect 2421 16949 2455 16983
rect 3065 16949 3099 16983
rect 4721 16949 4755 16983
rect 5365 16949 5399 16983
rect 5457 16949 5491 16983
rect 8171 16949 8205 16983
rect 11713 16949 11747 16983
rect 16037 16949 16071 16983
rect 2789 16745 2823 16779
rect 7711 16745 7745 16779
rect 12633 16745 12667 16779
rect 13369 16745 13403 16779
rect 15117 16745 15151 16779
rect 15485 16745 15519 16779
rect 18245 16745 18279 16779
rect 5273 16677 5307 16711
rect 9965 16677 9999 16711
rect 13001 16677 13035 16711
rect 15853 16677 15887 16711
rect 9505 16609 9539 16643
rect 12357 16609 12391 16643
rect 12909 16609 12943 16643
rect 13093 16609 13127 16643
rect 13645 16609 13679 16643
rect 14289 16609 14323 16643
rect 15761 16609 15795 16643
rect 17969 16609 18003 16643
rect 18429 16609 18463 16643
rect 4261 16541 4295 16575
rect 4537 16541 4571 16575
rect 9137 16541 9171 16575
rect 12633 16541 12667 16575
rect 13369 16541 13403 16575
rect 14841 16541 14875 16575
rect 15025 16541 15059 16575
rect 11253 16473 11287 16507
rect 6745 16405 6779 16439
rect 12449 16405 12483 16439
rect 13553 16405 13587 16439
rect 14197 16405 14231 16439
rect 5825 16201 5859 16235
rect 7205 16201 7239 16235
rect 9413 16201 9447 16235
rect 10057 16201 10091 16235
rect 12449 16201 12483 16235
rect 13829 16201 13863 16235
rect 2697 16133 2731 16167
rect 1777 16065 1811 16099
rect 4445 16065 4479 16099
rect 6653 16065 6687 16099
rect 7481 16065 7515 16099
rect 8769 16065 8803 16099
rect 15945 16065 15979 16099
rect 2605 15997 2639 16031
rect 2789 15997 2823 16031
rect 4701 15997 4735 16031
rect 6837 15997 6871 16031
rect 7573 15997 7607 16031
rect 10057 15997 10091 16031
rect 16313 15997 16347 16031
rect 1869 15929 1903 15963
rect 11161 15929 11195 15963
rect 15301 15929 15335 15963
rect 1961 15861 1995 15895
rect 2329 15861 2363 15895
rect 6745 15861 6779 15895
rect 17739 15861 17773 15895
rect 1501 15657 1535 15691
rect 1961 15657 1995 15691
rect 5733 15657 5767 15691
rect 8309 15657 8343 15691
rect 11621 15657 11655 15691
rect 13093 15657 13127 15691
rect 14013 15657 14047 15691
rect 17141 15657 17175 15691
rect 7021 15589 7055 15623
rect 9597 15589 9631 15623
rect 949 15521 983 15555
rect 1593 15521 1627 15555
rect 9965 15521 9999 15555
rect 10057 15521 10091 15555
rect 10333 15521 10367 15555
rect 10517 15521 10551 15555
rect 12689 15521 12723 15555
rect 12797 15527 12831 15561
rect 12905 15521 12939 15555
rect 16497 15521 16531 15555
rect 18429 15521 18463 15555
rect 1409 15453 1443 15487
rect 11713 15453 11747 15487
rect 11897 15453 11931 15487
rect 13829 15453 13863 15487
rect 13921 15453 13955 15487
rect 17785 15453 17819 15487
rect 10333 15385 10367 15419
rect 18245 15385 18279 15419
rect 857 15317 891 15351
rect 11253 15317 11287 15351
rect 14381 15317 14415 15351
rect 15209 15317 15243 15351
rect 3525 15113 3559 15147
rect 9505 15113 9539 15147
rect 10149 15113 10183 15147
rect 11161 15113 11195 15147
rect 17923 15113 17957 15147
rect 4997 15045 5031 15079
rect 13737 15045 13771 15079
rect 1777 14977 1811 15011
rect 6377 14977 6411 15011
rect 8125 14977 8159 15011
rect 8953 14977 8987 15011
rect 11621 14977 11655 15011
rect 11713 14977 11747 15011
rect 14289 14977 14323 15011
rect 15393 14977 15427 15011
rect 16129 14977 16163 15011
rect 3985 14909 4019 14943
rect 4169 14909 4203 14943
rect 4813 14909 4847 14943
rect 5917 14909 5951 14943
rect 10240 14909 10274 14943
rect 10333 14909 10367 14943
rect 11529 14909 11563 14943
rect 12265 14909 12299 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 13185 14909 13219 14943
rect 14105 14909 14139 14943
rect 15117 14909 15151 14943
rect 15209 14909 15243 14943
rect 15301 14909 15335 14943
rect 16497 14909 16531 14943
rect 2053 14841 2087 14875
rect 6653 14841 6687 14875
rect 4169 14773 4203 14807
rect 5365 14773 5399 14807
rect 9045 14773 9079 14807
rect 9137 14773 9171 14807
rect 12633 14773 12667 14807
rect 13093 14773 13127 14807
rect 14197 14773 14231 14807
rect 15577 14773 15611 14807
rect 18429 14773 18463 14807
rect 3341 14569 3375 14603
rect 7021 14569 7055 14603
rect 8585 14569 8619 14603
rect 9137 14569 9171 14603
rect 1133 14501 1167 14535
rect 3525 14501 3559 14535
rect 5549 14501 5583 14535
rect 12633 14501 12667 14535
rect 1225 14433 1259 14467
rect 3617 14433 3651 14467
rect 5273 14433 5307 14467
rect 8217 14433 8251 14467
rect 9229 14433 9263 14467
rect 11345 14433 11379 14467
rect 12357 14433 12391 14467
rect 13093 14433 13127 14467
rect 13185 14433 13219 14467
rect 14289 14433 14323 14467
rect 16773 14433 16807 14467
rect 18061 14433 18095 14467
rect 18245 14433 18279 14467
rect 1041 14365 1075 14399
rect 3157 14365 3191 14399
rect 3709 14365 3743 14399
rect 8309 14365 8343 14399
rect 9045 14365 9079 14399
rect 13369 14365 13403 14399
rect 14013 14365 14047 14399
rect 16497 14365 16531 14399
rect 17141 14365 17175 14399
rect 17693 14365 17727 14399
rect 9597 14297 9631 14331
rect 1593 14229 1627 14263
rect 10057 14229 10091 14263
rect 11345 14229 11379 14263
rect 13277 14229 13311 14263
rect 15025 14229 15059 14263
rect 18153 14229 18187 14263
rect 3525 14025 3559 14059
rect 7113 14025 7147 14059
rect 9321 14025 9355 14059
rect 16484 14025 16518 14059
rect 17969 14025 18003 14059
rect 2145 13889 2179 13923
rect 4169 13889 4203 13923
rect 7665 13889 7699 13923
rect 11161 13889 11195 13923
rect 11529 13889 11563 13923
rect 13001 13889 13035 13923
rect 14841 13889 14875 13923
rect 15025 13889 15059 13923
rect 15209 13889 15243 13923
rect 15301 13889 15335 13923
rect 16221 13889 16255 13923
rect 1777 13821 1811 13855
rect 4537 13821 4571 13855
rect 5963 13821 5997 13855
rect 8769 13821 8803 13855
rect 8861 13821 8895 13855
rect 14473 13821 14507 13855
rect 15117 13753 15151 13787
rect 15393 13685 15427 13719
rect 1133 13481 1167 13515
rect 1593 13481 1627 13515
rect 3617 13481 3651 13515
rect 8309 13481 8343 13515
rect 10057 13481 10091 13515
rect 10885 13481 10919 13515
rect 13553 13481 13587 13515
rect 16497 13481 16531 13515
rect 1501 13413 1535 13447
rect 9597 13413 9631 13447
rect 12817 13413 12851 13447
rect 13369 13413 13403 13447
rect 15025 13413 15059 13447
rect 17509 13413 17543 13447
rect 3341 13345 3375 13379
rect 5273 13345 5307 13379
rect 5540 13345 5574 13379
rect 9965 13345 9999 13379
rect 10241 13345 10275 13379
rect 10977 13345 11011 13379
rect 11161 13345 11195 13379
rect 11805 13345 11839 13379
rect 12725 13345 12759 13379
rect 13645 13345 13679 13379
rect 17601 13345 17635 13379
rect 1777 13277 1811 13311
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 12909 13277 12943 13311
rect 11897 13209 11931 13243
rect 13369 13209 13403 13243
rect 6653 13141 6687 13175
rect 10425 13141 10459 13175
rect 12357 13141 12391 13175
rect 9689 12937 9723 12971
rect 13829 12937 13863 12971
rect 10701 12869 10735 12903
rect 16313 12869 16347 12903
rect 4077 12801 4111 12835
rect 7849 12801 7883 12835
rect 10057 12801 10091 12835
rect 10241 12801 10275 12835
rect 12909 12801 12943 12835
rect 13185 12801 13219 12835
rect 15577 12801 15611 12835
rect 17601 12801 17635 12835
rect 1685 12733 1719 12767
rect 2053 12733 2087 12767
rect 7757 12733 7791 12767
rect 9229 12733 9263 12767
rect 9321 12733 9355 12767
rect 9505 12733 9539 12767
rect 15945 12733 15979 12767
rect 16313 12733 16347 12767
rect 16405 12733 16439 12767
rect 16773 12733 16807 12767
rect 17417 12733 17451 12767
rect 4344 12665 4378 12699
rect 5733 12665 5767 12699
rect 15301 12665 15335 12699
rect 17233 12665 17267 12699
rect 3479 12597 3513 12631
rect 5457 12597 5491 12631
rect 8125 12597 8159 12631
rect 10333 12597 10367 12631
rect 11437 12597 11471 12631
rect 17233 12393 17267 12427
rect 1777 12325 1811 12359
rect 6101 12325 6135 12359
rect 6469 12325 6503 12359
rect 6653 12325 6687 12359
rect 16129 12325 16163 12359
rect 765 12257 799 12291
rect 2145 12257 2179 12291
rect 5733 12257 5767 12291
rect 5826 12257 5860 12291
rect 6377 12257 6411 12291
rect 9321 12257 9355 12291
rect 10425 12257 10459 12291
rect 11069 12257 11103 12291
rect 13093 12257 13127 12291
rect 13829 12257 13863 12291
rect 14105 12257 14139 12291
rect 15945 12257 15979 12291
rect 17141 12257 17175 12291
rect 17325 12257 17359 12291
rect 857 12189 891 12223
rect 9045 12189 9079 12223
rect 10793 12189 10827 12223
rect 10977 12189 11011 12223
rect 12725 12189 12759 12223
rect 13369 12189 13403 12223
rect 16221 12189 16255 12223
rect 7573 12121 7607 12155
rect 1041 12053 1075 12087
rect 6377 12053 6411 12087
rect 10149 12053 10183 12087
rect 11437 12053 11471 12087
rect 14841 12053 14875 12087
rect 10793 11849 10827 11883
rect 15301 11849 15335 11883
rect 17923 11849 17957 11883
rect 5641 11781 5675 11815
rect 2237 11713 2271 11747
rect 9045 11713 9079 11747
rect 10149 11713 10183 11747
rect 16497 11713 16531 11747
rect 1961 11645 1995 11679
rect 5273 11645 5307 11679
rect 5427 11645 5461 11679
rect 9229 11645 9263 11679
rect 10425 11645 10459 11679
rect 11161 11645 11195 11679
rect 13553 11645 13587 11679
rect 16129 11645 16163 11679
rect 8125 11577 8159 11611
rect 13829 11577 13863 11611
rect 1593 11509 1627 11543
rect 2053 11509 2087 11543
rect 6837 11509 6871 11543
rect 9137 11509 9171 11543
rect 9597 11509 9631 11543
rect 10333 11509 10367 11543
rect 11345 11509 11379 11543
rect 1593 11305 1627 11339
rect 2053 11305 2087 11339
rect 8217 11305 8251 11339
rect 8861 11305 8895 11339
rect 9229 11305 9263 11339
rect 11759 11305 11793 11339
rect 14749 11305 14783 11339
rect 16037 11305 16071 11339
rect 17141 11305 17175 11339
rect 18245 11305 18279 11339
rect 1685 11237 1719 11271
rect 9965 11169 9999 11203
rect 10333 11169 10367 11203
rect 15025 11169 15059 11203
rect 15577 11169 15611 11203
rect 15761 11169 15795 11203
rect 16405 11169 16439 11203
rect 17969 11169 18003 11203
rect 18429 11169 18463 11203
rect 1501 11101 1535 11135
rect 4261 11101 4295 11135
rect 4537 11101 4571 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 8677 11101 8711 11135
rect 8769 11101 8803 11135
rect 14749 11101 14783 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 2789 11033 2823 11067
rect 14933 11033 14967 11067
rect 15761 11033 15795 11067
rect 6929 10965 6963 10999
rect 17509 10965 17543 10999
rect 1869 10761 1903 10795
rect 10609 10761 10643 10795
rect 11437 10761 11471 10795
rect 16313 10761 16347 10795
rect 7573 10693 7607 10727
rect 3341 10625 3375 10659
rect 7021 10625 7055 10659
rect 8217 10625 8251 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 13553 10625 13587 10659
rect 3617 10557 3651 10591
rect 3985 10557 4019 10591
rect 7113 10557 7147 10591
rect 7941 10557 7975 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 16313 10557 16347 10591
rect 17417 10557 17451 10591
rect 17510 10557 17544 10591
rect 4252 10489 4286 10523
rect 8125 10489 8159 10523
rect 15301 10489 15335 10523
rect 5365 10421 5399 10455
rect 7205 10421 7239 10455
rect 17141 10421 17175 10455
rect 17785 10421 17819 10455
rect 18429 10421 18463 10455
rect 2053 10217 2087 10251
rect 2421 10217 2455 10251
rect 3249 10217 3283 10251
rect 5733 10217 5767 10251
rect 9413 10217 9447 10251
rect 4537 10149 4571 10183
rect 581 10081 615 10115
rect 1041 10081 1075 10115
rect 5181 10081 5215 10115
rect 5457 10081 5491 10115
rect 5549 10081 5583 10115
rect 6193 10081 6227 10115
rect 7205 10081 7239 10115
rect 9597 10081 9631 10115
rect 13828 10081 13862 10115
rect 13921 10081 13955 10115
rect 17325 10081 17359 10115
rect 18275 10081 18309 10115
rect 18429 10081 18463 10115
rect 1869 10013 1903 10047
rect 1961 10013 1995 10047
rect 6009 10013 6043 10047
rect 14749 10013 14783 10047
rect 15117 10013 15151 10047
rect 17601 10013 17635 10047
rect 7021 9945 7055 9979
rect 13553 9945 13587 9979
rect 18061 9945 18095 9979
rect 765 9877 799 9911
rect 5273 9877 5307 9911
rect 16543 9877 16577 9911
rect 17325 9673 17359 9707
rect 857 9605 891 9639
rect 2421 9605 2455 9639
rect 13921 9605 13955 9639
rect 15301 9605 15335 9639
rect 765 9537 799 9571
rect 1869 9537 1903 9571
rect 2789 9537 2823 9571
rect 6929 9537 6963 9571
rect 10793 9537 10827 9571
rect 12909 9537 12943 9571
rect 14013 9537 14047 9571
rect 1041 9469 1075 9503
rect 2697 9469 2731 9503
rect 2881 9469 2915 9503
rect 4261 9469 4295 9503
rect 4445 9469 4479 9503
rect 4905 9469 4939 9503
rect 5089 9469 5123 9503
rect 6561 9469 6595 9503
rect 13737 9469 13771 9503
rect 15301 9469 15335 9503
rect 15577 9469 15611 9503
rect 15945 9469 15979 9503
rect 17785 9469 17819 9503
rect 17877 9469 17911 9503
rect 2053 9401 2087 9435
rect 10517 9401 10551 9435
rect 12633 9401 12667 9435
rect 16212 9401 16246 9435
rect 17601 9401 17635 9435
rect 1225 9333 1259 9367
rect 1961 9333 1995 9367
rect 4629 9333 4663 9367
rect 4997 9333 5031 9367
rect 8355 9333 8389 9367
rect 9045 9333 9079 9367
rect 11161 9333 11195 9367
rect 13553 9333 13587 9367
rect 14381 9333 14415 9367
rect 15485 9333 15519 9367
rect 17693 9333 17727 9367
rect 18337 9333 18371 9367
rect 2973 9129 3007 9163
rect 4445 9129 4479 9163
rect 5641 9129 5675 9163
rect 6009 9129 6043 9163
rect 8033 9129 8067 9163
rect 12817 9129 12851 9163
rect 17325 9129 17359 9163
rect 3249 9061 3283 9095
rect 14105 9061 14139 9095
rect 16497 9061 16531 9095
rect 1869 8993 1903 9027
rect 2053 8993 2087 9027
rect 2973 8993 3007 9027
rect 4629 8993 4663 9027
rect 4721 8993 4755 9027
rect 5917 8993 5951 9027
rect 6101 8993 6135 9027
rect 6837 8993 6871 9027
rect 7573 8993 7607 9027
rect 8033 8993 8067 9027
rect 8585 8993 8619 9027
rect 8861 8993 8895 9027
rect 11713 8993 11747 9027
rect 12817 8993 12851 9027
rect 12909 8993 12943 9027
rect 17233 8993 17267 9027
rect 17877 8993 17911 9027
rect 4445 8925 4479 8959
rect 6561 8925 6595 8959
rect 9965 8925 9999 8959
rect 11437 8925 11471 8959
rect 13093 8925 13127 8959
rect 13829 8925 13863 8959
rect 18153 8925 18187 8959
rect 1777 8857 1811 8891
rect 3065 8857 3099 8891
rect 7711 8857 7745 8891
rect 13461 8857 13495 8891
rect 7849 8789 7883 8823
rect 15209 8789 15243 8823
rect 2329 8585 2363 8619
rect 7849 8585 7883 8619
rect 8309 8585 8343 8619
rect 13553 8585 13587 8619
rect 15301 8585 15335 8619
rect 17785 8585 17819 8619
rect 18429 8585 18463 8619
rect 1777 8449 1811 8483
rect 1869 8449 1903 8483
rect 2973 8449 3007 8483
rect 3341 8449 3375 8483
rect 8953 8449 8987 8483
rect 10793 8449 10827 8483
rect 13921 8449 13955 8483
rect 15209 8449 15243 8483
rect 16405 8449 16439 8483
rect 949 8381 983 8415
rect 3157 8381 3191 8415
rect 3433 8381 3467 8415
rect 5641 8381 5675 8415
rect 7481 8381 7515 8415
rect 7665 8381 7699 8415
rect 8125 8381 8159 8415
rect 8309 8381 8343 8415
rect 10425 8381 10459 8415
rect 11621 8381 11655 8415
rect 14473 8381 14507 8415
rect 14749 8381 14783 8415
rect 14933 8381 14967 8415
rect 15393 8381 15427 8415
rect 15485 8381 15519 8415
rect 16672 8381 16706 8415
rect 1961 8313 1995 8347
rect 5273 8313 5307 8347
rect 11345 8313 11379 8347
rect 857 8245 891 8279
rect 16037 8245 16071 8279
rect 1225 8041 1259 8075
rect 7665 8041 7699 8075
rect 8769 8041 8803 8075
rect 10195 8041 10229 8075
rect 14749 8041 14783 8075
rect 857 7973 891 8007
rect 17969 7973 18003 8007
rect 1041 7905 1075 7939
rect 1317 7905 1351 7939
rect 5181 7905 5215 7939
rect 11989 7905 12023 7939
rect 12725 7905 12759 7939
rect 16497 7905 16531 7939
rect 17325 7905 17359 7939
rect 17417 7905 17451 7939
rect 17693 7905 17727 7939
rect 18245 7905 18279 7939
rect 5549 7837 5583 7871
rect 6975 7837 7009 7871
rect 11621 7837 11655 7871
rect 12449 7837 12483 7871
rect 16221 7837 16255 7871
rect 17141 7837 17175 7871
rect 17969 7837 18003 7871
rect 12633 7769 12667 7803
rect 14381 7769 14415 7803
rect 12541 7701 12575 7735
rect 17601 7701 17635 7735
rect 18153 7701 18187 7735
rect 5089 7497 5123 7531
rect 5457 7497 5491 7531
rect 5825 7497 5859 7531
rect 7573 7497 7607 7531
rect 8953 7497 8987 7531
rect 13810 7497 13844 7531
rect 17785 7497 17819 7531
rect 18429 7497 18463 7531
rect 9321 7429 9355 7463
rect 11437 7429 11471 7463
rect 1869 7361 1903 7395
rect 5549 7361 5583 7395
rect 9045 7361 9079 7395
rect 13553 7361 13587 7395
rect 16129 7361 16163 7395
rect 5273 7293 5307 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 9505 7293 9539 7327
rect 9597 7293 9631 7327
rect 11253 7293 11287 7327
rect 17969 7293 18003 7327
rect 2145 7225 2179 7259
rect 4077 7225 4111 7259
rect 4813 7225 4847 7259
rect 9321 7225 9355 7259
rect 15577 7225 15611 7259
rect 16396 7225 16430 7259
rect 3617 7157 3651 7191
rect 17509 7157 17543 7191
rect 1501 6953 1535 6987
rect 17969 6953 18003 6987
rect 18337 6953 18371 6987
rect 2881 6817 2915 6851
rect 7021 6817 7055 6851
rect 11529 6817 11563 6851
rect 12909 6817 12943 6851
rect 13369 6817 13403 6851
rect 17785 6817 17819 6851
rect 18245 6817 18279 6851
rect 18429 6817 18463 6851
rect 1225 6749 1259 6783
rect 1409 6749 1443 6783
rect 3157 6749 3191 6783
rect 7757 6749 7791 6783
rect 8125 6749 8159 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 16313 6749 16347 6783
rect 17601 6749 17635 6783
rect 1869 6681 1903 6715
rect 4629 6681 4663 6715
rect 11345 6681 11379 6715
rect 16681 6681 16715 6715
rect 17233 6681 17267 6715
rect 5733 6613 5767 6647
rect 9505 6613 9539 6647
rect 15393 6613 15427 6647
rect 15945 6613 15979 6647
rect 1685 6409 1719 6443
rect 3985 6409 4019 6443
rect 11161 6409 11195 6443
rect 12651 6409 12685 6443
rect 18337 6409 18371 6443
rect 5917 6341 5951 6375
rect 9229 6341 9263 6375
rect 14749 6341 14783 6375
rect 2053 6273 2087 6307
rect 4445 6273 4479 6307
rect 4537 6273 4571 6307
rect 6377 6273 6411 6307
rect 12909 6273 12943 6307
rect 15301 6273 15335 6307
rect 16129 6273 16163 6307
rect 16497 6273 16531 6307
rect 1961 6205 1995 6239
rect 2421 6205 2455 6239
rect 5181 6205 5215 6239
rect 5641 6205 5675 6239
rect 5825 6205 5859 6239
rect 6005 6205 6039 6239
rect 14013 6205 14047 6239
rect 14289 6205 14323 6239
rect 14473 6205 14507 6239
rect 14841 6205 14875 6239
rect 14933 6205 14967 6239
rect 4353 6137 4387 6171
rect 6653 6137 6687 6171
rect 9045 6137 9079 6171
rect 8125 6069 8159 6103
rect 9689 6069 9723 6103
rect 17923 6069 17957 6103
rect 10885 5865 10919 5899
rect 18245 5865 18279 5899
rect 2237 5797 2271 5831
rect 7849 5797 7883 5831
rect 2053 5729 2087 5763
rect 2329 5729 2363 5763
rect 3341 5729 3375 5763
rect 3893 5729 3927 5763
rect 5549 5729 5583 5763
rect 10977 5729 11011 5763
rect 11161 5729 11195 5763
rect 11529 5729 11563 5763
rect 11621 5729 11655 5763
rect 11805 5729 11839 5763
rect 16773 5729 16807 5763
rect 17969 5729 18003 5763
rect 18429 5729 18463 5763
rect 3525 5661 3559 5695
rect 3801 5661 3835 5695
rect 4721 5661 4755 5695
rect 5181 5661 5215 5695
rect 7573 5661 7607 5695
rect 9597 5661 9631 5695
rect 11713 5661 11747 5695
rect 11989 5661 12023 5695
rect 13829 5661 13863 5695
rect 14197 5661 14231 5695
rect 16405 5661 16439 5695
rect 2973 5593 3007 5627
rect 10701 5593 10735 5627
rect 12449 5593 12483 5627
rect 2053 5525 2087 5559
rect 6929 5525 6963 5559
rect 10057 5525 10091 5559
rect 15025 5525 15059 5559
rect 1685 5321 1719 5355
rect 3157 5321 3191 5355
rect 5365 5321 5399 5355
rect 7849 5321 7883 5355
rect 8125 5321 8159 5355
rect 11161 5321 11195 5355
rect 14013 5321 14047 5355
rect 1777 5253 1811 5287
rect 4077 5253 4111 5287
rect 9045 5253 9079 5287
rect 1869 5185 1903 5219
rect 11805 5185 11839 5219
rect 1593 5117 1627 5151
rect 3065 5117 3099 5151
rect 3985 5117 4019 5151
rect 4261 5117 4295 5151
rect 4445 5117 4479 5151
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 8769 5117 8803 5151
rect 8953 5117 8987 5151
rect 9229 5117 9263 5151
rect 9597 5117 9631 5151
rect 9781 5117 9815 5151
rect 10517 5117 10551 5151
rect 15301 5117 15335 5151
rect 6377 5049 6411 5083
rect 10241 5049 10275 5083
rect 4353 4981 4387 5015
rect 4721 4981 4755 5015
rect 7297 4981 7331 5015
rect 11529 4981 11563 5015
rect 11621 4981 11655 5015
rect 12265 4981 12299 5015
rect 857 4777 891 4811
rect 1777 4777 1811 4811
rect 4537 4777 4571 4811
rect 5273 4777 5307 4811
rect 7021 4777 7055 4811
rect 8401 4777 8435 4811
rect 10977 4777 11011 4811
rect 12909 4777 12943 4811
rect 4353 4709 4387 4743
rect 7757 4709 7791 4743
rect 8769 4709 8803 4743
rect 10149 4709 10183 4743
rect 17141 4709 17175 4743
rect 949 4641 983 4675
rect 1501 4641 1535 4675
rect 1593 4641 1627 4675
rect 4261 4641 4295 4675
rect 4721 4641 4755 4675
rect 4813 4641 4847 4675
rect 6653 4641 6687 4675
rect 6807 4641 6841 4675
rect 8125 4641 8159 4675
rect 8677 4641 8711 4675
rect 8861 4641 8895 4675
rect 10425 4641 10459 4675
rect 11345 4641 11379 4675
rect 12633 4641 12667 4675
rect 12817 4641 12851 4675
rect 13461 4641 13495 4675
rect 13553 4641 13587 4675
rect 13737 4641 13771 4675
rect 16773 4641 16807 4675
rect 17749 4641 17783 4675
rect 17877 4641 17911 4675
rect 17969 4641 18003 4675
rect 1777 4573 1811 4607
rect 7849 4573 7883 4607
rect 8217 4573 8251 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 16497 4573 16531 4607
rect 13645 4505 13679 4539
rect 13093 4437 13127 4471
rect 13921 4437 13955 4471
rect 15025 4437 15059 4471
rect 18153 4437 18187 4471
rect 2605 4233 2639 4267
rect 5825 4233 5859 4267
rect 7573 4233 7607 4267
rect 8769 4233 8803 4267
rect 9781 4233 9815 4267
rect 11897 4233 11931 4267
rect 12265 4233 12299 4267
rect 15313 4233 15347 4267
rect 2237 4097 2271 4131
rect 6009 4097 6043 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 9321 4097 9355 4131
rect 13829 4097 13863 4131
rect 15577 4097 15611 4131
rect 16773 4097 16807 4131
rect 17325 4097 17359 4131
rect 2789 4029 2823 4063
rect 2881 4007 2915 4041
rect 3009 4029 3043 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 6745 4029 6779 4063
rect 7665 4029 7699 4063
rect 7941 4029 7975 4063
rect 8125 4029 8159 4063
rect 9781 4029 9815 4063
rect 9965 4029 9999 4063
rect 17693 4029 17727 4063
rect 17785 4029 17819 4063
rect 6009 3961 6043 3995
rect 7021 3961 7055 3995
rect 7113 3961 7147 3995
rect 7389 3961 7423 3995
rect 9229 3961 9263 3995
rect 10241 3961 10275 3995
rect 1593 3893 1627 3927
rect 1961 3893 1995 3927
rect 2053 3893 2087 3927
rect 6469 3893 6503 3927
rect 9137 3893 9171 3927
rect 13185 3893 13219 3927
rect 16221 3893 16255 3927
rect 16589 3893 16623 3927
rect 16681 3893 16715 3927
rect 17969 3893 18003 3927
rect 2789 3689 2823 3723
rect 3893 3689 3927 3723
rect 4629 3689 4663 3723
rect 5181 3689 5215 3723
rect 11253 3689 11287 3723
rect 12357 3689 12391 3723
rect 13553 3689 13587 3723
rect 17141 3689 17175 3723
rect 18153 3689 18187 3723
rect 11621 3621 11655 3655
rect 12725 3621 12759 3655
rect 17509 3621 17543 3655
rect 2973 3553 3007 3587
rect 3065 3553 3099 3587
rect 3157 3553 3191 3587
rect 3525 3553 3559 3587
rect 3663 3553 3697 3587
rect 4169 3553 4203 3587
rect 4721 3553 4755 3587
rect 5457 3553 5491 3587
rect 5641 3553 5675 3587
rect 11713 3553 11747 3587
rect 13921 3553 13955 3587
rect 14013 3553 14047 3587
rect 14749 3553 14783 3587
rect 17601 3553 17635 3587
rect 18153 3553 18187 3587
rect 18337 3553 18371 3587
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 11897 3485 11931 3519
rect 12817 3485 12851 3519
rect 13001 3485 13035 3519
rect 14197 3485 14231 3519
rect 15025 3485 15059 3519
rect 17693 3485 17727 3519
rect 4353 3417 4387 3451
rect 4261 3349 4295 3383
rect 16497 3349 16531 3383
rect 949 3145 983 3179
rect 2329 3145 2363 3179
rect 4077 3145 4111 3179
rect 5273 3145 5307 3179
rect 9413 3145 9447 3179
rect 12449 3145 12483 3179
rect 13185 3145 13219 3179
rect 16681 3145 16715 3179
rect 17785 3145 17819 3179
rect 18337 3145 18371 3179
rect 16957 3077 16991 3111
rect 1777 3009 1811 3043
rect 5917 3009 5951 3043
rect 9965 3009 9999 3043
rect 16129 3009 16163 3043
rect 1041 2941 1075 2975
rect 1869 2941 1903 2975
rect 3985 2941 4019 2975
rect 4169 2941 4203 2975
rect 5733 2941 5767 2975
rect 6377 2941 6411 2975
rect 9873 2941 9907 2975
rect 10425 2941 10459 2975
rect 12081 2941 12115 2975
rect 13001 2941 13035 2975
rect 13185 2941 13219 2975
rect 13737 2941 13771 2975
rect 13829 2941 13863 2975
rect 14105 2941 14139 2975
rect 17509 2941 17543 2975
rect 17969 2941 18003 2975
rect 1961 2805 1995 2839
rect 5641 2805 5675 2839
rect 9781 2805 9815 2839
rect 13645 2805 13679 2839
rect 14473 2805 14507 2839
rect 16221 2805 16255 2839
rect 16313 2805 16347 2839
rect 1685 2601 1719 2635
rect 5273 2601 5307 2635
rect 6469 2601 6503 2635
rect 6837 2601 6871 2635
rect 7757 2601 7791 2635
rect 8217 2601 8251 2635
rect 9321 2601 9355 2635
rect 14105 2601 14139 2635
rect 15669 2601 15703 2635
rect 17233 2601 17267 2635
rect 2145 2533 2179 2567
rect 6929 2533 6963 2567
rect 8125 2533 8159 2567
rect 10793 2533 10827 2567
rect 13645 2533 13679 2567
rect 14933 2533 14967 2567
rect 15301 2533 15335 2567
rect 2053 2465 2087 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 9321 2465 9355 2499
rect 9597 2465 9631 2499
rect 10241 2465 10275 2499
rect 10517 2465 10551 2499
rect 13737 2465 13771 2499
rect 17233 2465 17267 2499
rect 17509 2465 17543 2499
rect 17877 2465 17911 2499
rect 2329 2397 2363 2431
rect 7021 2397 7055 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 9965 2397 9999 2431
rect 13553 2397 13587 2431
rect 15117 2397 15151 2431
rect 15209 2397 15243 2431
rect 17325 2397 17359 2431
rect 18337 2397 18371 2431
rect 10149 2329 10183 2363
rect 10609 2329 10643 2363
rect 17969 2329 18003 2363
rect 10057 2261 10091 2295
rect 10517 2261 10551 2295
rect 14933 2261 14967 2295
rect 1915 2057 1949 2091
rect 2881 2057 2915 2091
rect 5273 2057 5307 2091
rect 6377 2057 6411 2091
rect 6929 2057 6963 2091
rect 9229 2057 9263 2091
rect 13737 2057 13771 2091
rect 15255 2057 15289 2091
rect 16129 2057 16163 2091
rect 10241 1989 10275 2023
rect 12173 1989 12207 2023
rect 13001 1989 13035 2023
rect 14197 1989 14231 2023
rect 15117 1989 15151 2023
rect 3525 1921 3559 1955
rect 5825 1921 5859 1955
rect 7481 1921 7515 1955
rect 10517 1921 10551 1955
rect 11897 1921 11931 1955
rect 13553 1921 13587 1955
rect 16773 1921 16807 1955
rect 17693 1921 17727 1955
rect 2018 1853 2052 1887
rect 3985 1853 4019 1887
rect 4353 1853 4387 1887
rect 4813 1853 4847 1887
rect 7389 1853 7423 1887
rect 9045 1853 9079 1887
rect 10609 1853 10643 1887
rect 11805 1853 11839 1887
rect 12817 1853 12851 1887
rect 13093 1853 13127 1887
rect 13829 1853 13863 1887
rect 14933 1853 14967 1887
rect 15393 1853 15427 1887
rect 16589 1853 16623 1887
rect 17969 1853 18003 1887
rect 3341 1785 3375 1819
rect 5733 1785 5767 1819
rect 3249 1717 3283 1751
rect 4537 1717 4571 1751
rect 5641 1717 5675 1751
rect 7297 1717 7331 1751
rect 13093 1717 13127 1751
rect 13553 1717 13587 1751
rect 15025 1717 15059 1751
rect 16497 1717 16531 1751
rect 18429 1717 18463 1751
rect 3157 1513 3191 1547
rect 5917 1513 5951 1547
rect 8033 1513 8067 1547
rect 8493 1513 8527 1547
rect 13461 1513 13495 1547
rect 15485 1513 15519 1547
rect 15945 1513 15979 1547
rect 16773 1513 16807 1547
rect 3801 1445 3835 1479
rect 3432 1377 3466 1411
rect 3525 1377 3559 1411
rect 3985 1377 4019 1411
rect 4077 1377 4111 1411
rect 4353 1377 4387 1411
rect 4629 1377 4663 1411
rect 5549 1377 5583 1411
rect 8401 1377 8435 1411
rect 10179 1377 10213 1411
rect 10333 1377 10367 1411
rect 13093 1377 13127 1411
rect 13247 1377 13281 1411
rect 15024 1377 15058 1411
rect 15117 1377 15151 1411
rect 16773 1377 16807 1411
rect 17509 1377 17543 1411
rect 3801 1309 3835 1343
rect 5457 1309 5491 1343
rect 8677 1309 8711 1343
rect 9965 1309 9999 1343
rect 14749 1309 14783 1343
rect 16497 1309 16531 1343
rect 17601 1309 17635 1343
rect 4353 1241 4387 1275
rect 4445 1241 4479 1275
rect 16681 1241 16715 1275
rect 17141 1241 17175 1275
<< metal1 >>
rect 184 18522 18860 18544
rect 184 18470 1556 18522
rect 1608 18470 1620 18522
rect 1672 18470 1684 18522
rect 1736 18470 1748 18522
rect 1800 18470 1812 18522
rect 1864 18470 4656 18522
rect 4708 18470 4720 18522
rect 4772 18470 4784 18522
rect 4836 18470 4848 18522
rect 4900 18470 4912 18522
rect 4964 18470 7756 18522
rect 7808 18470 7820 18522
rect 7872 18470 7884 18522
rect 7936 18470 7948 18522
rect 8000 18470 8012 18522
rect 8064 18470 10856 18522
rect 10908 18470 10920 18522
rect 10972 18470 10984 18522
rect 11036 18470 11048 18522
rect 11100 18470 11112 18522
rect 11164 18470 13956 18522
rect 14008 18470 14020 18522
rect 14072 18470 14084 18522
rect 14136 18470 14148 18522
rect 14200 18470 14212 18522
rect 14264 18470 17056 18522
rect 17108 18470 17120 18522
rect 17172 18470 17184 18522
rect 17236 18470 17248 18522
rect 17300 18470 17312 18522
rect 17364 18470 18860 18522
rect 184 18448 18860 18470
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4246 18408 4252 18420
rect 3651 18380 4252 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 4338 18368 4344 18420
rect 4396 18408 4402 18420
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 4396 18380 4629 18408
rect 4396 18368 4402 18380
rect 4617 18377 4629 18380
rect 4663 18377 4675 18411
rect 18414 18408 18420 18420
rect 18375 18380 18420 18408
rect 4617 18371 4675 18377
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 5994 18340 6000 18352
rect 4264 18312 6000 18340
rect 4264 18281 4292 18312
rect 5994 18300 6000 18312
rect 6052 18340 6058 18352
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 6052 18312 17785 18340
rect 6052 18300 6058 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 6687 18244 7205 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 7193 18241 7205 18244
rect 7239 18272 7251 18275
rect 8662 18272 8668 18284
rect 7239 18244 8668 18272
rect 7239 18241 7251 18244
rect 7193 18235 7251 18241
rect 1394 18164 1400 18216
rect 1452 18204 1458 18216
rect 1581 18207 1639 18213
rect 1581 18204 1593 18207
rect 1452 18176 1593 18204
rect 1452 18164 1458 18176
rect 1581 18173 1593 18176
rect 1627 18204 1639 18207
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1627 18176 2053 18204
rect 1627 18173 1639 18176
rect 1581 18167 1639 18173
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 5261 18207 5319 18213
rect 5261 18173 5273 18207
rect 5307 18204 5319 18207
rect 5997 18207 6055 18213
rect 5997 18204 6009 18207
rect 5307 18176 6009 18204
rect 5307 18173 5319 18176
rect 5261 18167 5319 18173
rect 5997 18173 6009 18176
rect 6043 18204 6055 18207
rect 6656 18204 6684 18235
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 10502 18272 10508 18284
rect 10463 18244 10508 18272
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 14642 18232 14648 18284
rect 14700 18272 14706 18284
rect 14829 18275 14887 18281
rect 14829 18272 14841 18275
rect 14700 18244 14841 18272
rect 14700 18232 14706 18244
rect 14829 18241 14841 18244
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 6043 18176 6684 18204
rect 6825 18207 6883 18213
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 8202 18204 8208 18216
rect 6871 18176 8064 18204
rect 8163 18176 8208 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 5442 18136 5448 18148
rect 4632 18108 5448 18136
rect 4632 18077 4660 18108
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 5718 18136 5724 18148
rect 5679 18108 5724 18136
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 7834 18136 7840 18148
rect 7795 18108 7840 18136
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 8036 18136 8064 18176
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 8444 18176 9321 18204
rect 8444 18164 8450 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 9732 18176 11253 18204
rect 9732 18164 9738 18176
rect 11241 18173 11253 18176
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 12894 18204 12900 18216
rect 11747 18176 12900 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 14220 18207 14278 18213
rect 14220 18204 14232 18207
rect 13504 18176 14232 18204
rect 13504 18164 13510 18176
rect 14220 18173 14232 18176
rect 14266 18173 14278 18207
rect 14220 18167 14278 18173
rect 16114 18164 16120 18216
rect 16172 18204 16178 18216
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 16172 18176 16221 18204
rect 16172 18164 16178 18176
rect 16209 18173 16221 18176
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 18414 18204 18420 18216
rect 18003 18176 18420 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 8110 18136 8116 18148
rect 8036 18108 8116 18136
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 10413 18139 10471 18145
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 13814 18136 13820 18148
rect 10459 18108 13820 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 13814 18096 13820 18108
rect 13872 18136 13878 18148
rect 14918 18136 14924 18148
rect 13872 18108 14924 18136
rect 13872 18096 13878 18108
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 15028 18108 16068 18136
rect 15028 18080 15056 18108
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 4617 18071 4675 18077
rect 4617 18068 4629 18071
rect 1811 18040 4629 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 4617 18037 4629 18040
rect 4663 18037 4675 18071
rect 4617 18031 4675 18037
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4982 18068 4988 18080
rect 4847 18040 4988 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8757 18071 8815 18077
rect 8757 18068 8769 18071
rect 8352 18040 8769 18068
rect 8352 18028 8358 18040
rect 8757 18037 8769 18040
rect 8803 18037 8815 18071
rect 9950 18068 9956 18080
rect 9911 18040 9956 18068
rect 8757 18031 8815 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 14323 18071 14381 18077
rect 14323 18037 14335 18071
rect 14369 18068 14381 18071
rect 14826 18068 14832 18080
rect 14369 18040 14832 18068
rect 14369 18037 14381 18040
rect 14323 18031 14381 18037
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15194 18068 15200 18080
rect 15151 18040 15200 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 16040 18077 16068 18108
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15436 18040 15485 18068
rect 15436 18028 15442 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 15473 18031 15531 18037
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 184 17978 18920 18000
rect 184 17926 3106 17978
rect 3158 17926 3170 17978
rect 3222 17926 3234 17978
rect 3286 17926 3298 17978
rect 3350 17926 3362 17978
rect 3414 17926 6206 17978
rect 6258 17926 6270 17978
rect 6322 17926 6334 17978
rect 6386 17926 6398 17978
rect 6450 17926 6462 17978
rect 6514 17926 9306 17978
rect 9358 17926 9370 17978
rect 9422 17926 9434 17978
rect 9486 17926 9498 17978
rect 9550 17926 9562 17978
rect 9614 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 12534 17978
rect 12586 17926 12598 17978
rect 12650 17926 12662 17978
rect 12714 17926 15506 17978
rect 15558 17926 15570 17978
rect 15622 17926 15634 17978
rect 15686 17926 15698 17978
rect 15750 17926 15762 17978
rect 15814 17926 18606 17978
rect 18658 17926 18670 17978
rect 18722 17926 18734 17978
rect 18786 17926 18798 17978
rect 18850 17926 18862 17978
rect 18914 17926 18920 17978
rect 184 17904 18920 17926
rect 9539 17867 9597 17873
rect 9539 17833 9551 17867
rect 9585 17864 9597 17867
rect 9674 17864 9680 17876
rect 9585 17836 9680 17864
rect 9585 17833 9597 17836
rect 9539 17827 9597 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 4246 17756 4252 17808
rect 4304 17796 4310 17808
rect 5445 17799 5503 17805
rect 5445 17796 5457 17799
rect 4304 17768 5457 17796
rect 4304 17756 4310 17768
rect 5445 17765 5457 17768
rect 5491 17765 5503 17799
rect 5445 17759 5503 17765
rect 8662 17756 8668 17808
rect 8720 17756 8726 17808
rect 16850 17796 16856 17808
rect 16514 17768 16856 17796
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 1946 17688 1952 17740
rect 2004 17728 2010 17740
rect 2071 17731 2129 17737
rect 2071 17728 2083 17731
rect 2004 17700 2083 17728
rect 2004 17688 2010 17700
rect 2071 17697 2083 17700
rect 2117 17697 2129 17731
rect 2071 17691 2129 17697
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2406 17728 2412 17740
rect 2271 17700 2412 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17728 4583 17731
rect 5166 17728 5172 17740
rect 4571 17700 5172 17728
rect 4571 17697 4583 17700
rect 4525 17691 4583 17697
rect 5166 17688 5172 17700
rect 5224 17728 5230 17740
rect 7745 17731 7803 17737
rect 5224 17700 6776 17728
rect 5224 17688 5230 17700
rect 4338 17552 4344 17604
rect 4396 17592 4402 17604
rect 5350 17592 5356 17604
rect 4396 17564 5356 17592
rect 4396 17552 4402 17564
rect 5350 17552 5356 17564
rect 5408 17552 5414 17604
rect 6748 17601 6776 17700
rect 7745 17697 7757 17731
rect 7791 17728 7803 17731
rect 7834 17728 7840 17740
rect 7791 17700 7840 17728
rect 7791 17697 7803 17700
rect 7745 17691 7803 17697
rect 7834 17688 7840 17700
rect 7892 17688 7898 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9232 17700 9965 17728
rect 9232 17672 9260 17700
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 12894 17728 12900 17740
rect 12855 17700 12900 17728
rect 9953 17691 10011 17697
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 15013 17731 15071 17737
rect 15013 17728 15025 17731
rect 14976 17700 15025 17728
rect 14976 17688 14982 17700
rect 15013 17697 15025 17700
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8294 17660 8300 17672
rect 8159 17632 8300 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 9214 17620 9220 17672
rect 9272 17620 9278 17672
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12860 17632 13369 17660
rect 12860 17620 12866 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 16666 17660 16672 17672
rect 15335 17632 16672 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 16807 17632 17233 17660
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 17221 17629 17233 17632
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 6733 17595 6791 17601
rect 6733 17561 6745 17595
rect 6779 17561 6791 17595
rect 6733 17555 6791 17561
rect 2041 17527 2099 17533
rect 2041 17493 2053 17527
rect 2087 17524 2099 17527
rect 2866 17524 2872 17536
rect 2087 17496 2872 17524
rect 2087 17493 2099 17496
rect 2041 17487 2099 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3237 17527 3295 17533
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 5258 17524 5264 17536
rect 3283 17496 5264 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 9732 17496 11253 17524
rect 9732 17484 9738 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11241 17487 11299 17493
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 17552 17496 17877 17524
rect 17552 17484 17558 17496
rect 17865 17493 17877 17496
rect 17911 17493 17923 17527
rect 17865 17487 17923 17493
rect 184 17434 18860 17456
rect 184 17382 1556 17434
rect 1608 17382 1620 17434
rect 1672 17382 1684 17434
rect 1736 17382 1748 17434
rect 1800 17382 1812 17434
rect 1864 17382 4656 17434
rect 4708 17382 4720 17434
rect 4772 17382 4784 17434
rect 4836 17382 4848 17434
rect 4900 17382 4912 17434
rect 4964 17382 7756 17434
rect 7808 17382 7820 17434
rect 7872 17382 7884 17434
rect 7936 17382 7948 17434
rect 8000 17382 8012 17434
rect 8064 17382 10856 17434
rect 10908 17382 10920 17434
rect 10972 17382 10984 17434
rect 11036 17382 11048 17434
rect 11100 17382 11112 17434
rect 11164 17382 13956 17434
rect 14008 17382 14020 17434
rect 14072 17382 14084 17434
rect 14136 17382 14148 17434
rect 14200 17382 14212 17434
rect 14264 17382 17056 17434
rect 17108 17382 17120 17434
rect 17172 17382 17184 17434
rect 17236 17382 17248 17434
rect 17300 17382 17312 17434
rect 17364 17382 18860 17434
rect 184 17360 18860 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 2148 17292 2605 17320
rect 1719 17255 1777 17261
rect 1719 17252 1731 17255
rect 768 17224 1731 17252
rect 768 17125 796 17224
rect 1719 17221 1731 17224
rect 1765 17252 1777 17255
rect 2148 17252 2176 17292
rect 2593 17289 2605 17292
rect 2639 17320 2651 17323
rect 2682 17320 2688 17332
rect 2639 17292 2688 17320
rect 2639 17289 2651 17292
rect 2593 17283 2651 17289
rect 2682 17280 2688 17292
rect 2740 17320 2746 17332
rect 2740 17292 3188 17320
rect 2740 17280 2746 17292
rect 1765 17224 2176 17252
rect 1765 17221 1777 17224
rect 1719 17215 1777 17221
rect 845 17187 903 17193
rect 845 17153 857 17187
rect 891 17184 903 17187
rect 1857 17187 1915 17193
rect 1857 17184 1869 17187
rect 891 17156 1869 17184
rect 891 17153 903 17156
rect 845 17147 903 17153
rect 1857 17153 1869 17156
rect 1903 17184 1915 17187
rect 1946 17184 1952 17196
rect 1903 17156 1952 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 1946 17144 1952 17156
rect 2004 17184 2010 17196
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 2004 17156 2513 17184
rect 2004 17144 2010 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 753 17119 811 17125
rect 753 17085 765 17119
rect 799 17085 811 17119
rect 753 17079 811 17085
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 2087 17088 2329 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 2317 17085 2329 17088
rect 2363 17116 2375 17119
rect 2958 17116 2964 17128
rect 2363 17088 2964 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 1596 17048 1624 17079
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3160 17125 3188 17292
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 5718 17320 5724 17332
rect 4488 17292 5724 17320
rect 4488 17280 4494 17292
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 12345 17323 12403 17329
rect 12345 17289 12357 17323
rect 12391 17320 12403 17323
rect 12391 17292 12664 17320
rect 12391 17289 12403 17292
rect 12345 17283 12403 17289
rect 12526 17252 12532 17264
rect 5184 17224 6316 17252
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 5184 17184 5212 17224
rect 3651 17156 5212 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4430 17116 4436 17128
rect 4391 17088 4436 17116
rect 4249 17079 4307 17085
rect 2685 17051 2743 17057
rect 2685 17048 2697 17051
rect 1596 17020 2697 17048
rect 2608 16992 2636 17020
rect 2685 17017 2697 17020
rect 2731 17017 2743 17051
rect 4264 17048 4292 17079
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 4847 17088 5212 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5074 17048 5080 17060
rect 4264 17020 5080 17048
rect 2685 17011 2743 17017
rect 5074 17008 5080 17020
rect 5132 17008 5138 17060
rect 5184 17048 5212 17088
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5994 17116 6000 17128
rect 5316 17088 5361 17116
rect 5955 17088 6000 17116
rect 5316 17076 5322 17088
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 6288 17116 6316 17224
rect 12084 17224 12532 17252
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 7466 17184 7472 17196
rect 6411 17156 7472 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 12084 17193 12112 17224
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 11241 17187 11299 17193
rect 11241 17153 11253 17187
rect 11287 17153 11299 17187
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11241 17147 11299 17153
rect 11348 17156 12081 17184
rect 6733 17119 6791 17125
rect 6733 17116 6745 17119
rect 6288 17088 6745 17116
rect 6733 17085 6745 17088
rect 6779 17085 6791 17119
rect 6733 17079 6791 17085
rect 5813 17051 5871 17057
rect 5813 17048 5825 17051
rect 5184 17020 5825 17048
rect 5813 17017 5825 17020
rect 5859 17017 5871 17051
rect 8018 17048 8024 17060
rect 7774 17020 8024 17048
rect 5813 17011 5871 17017
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 9030 17048 9036 17060
rect 8991 17020 9036 17048
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 10594 17048 10600 17060
rect 10555 17020 10600 17048
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 11256 17048 11284 17147
rect 11348 17125 11376 17156
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12253 17187 12311 17193
rect 12253 17184 12265 17187
rect 12216 17156 12265 17184
rect 12216 17144 12222 17156
rect 12253 17153 12265 17156
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12406 17156 12572 17184
rect 12406 17128 12434 17156
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 12342 17116 12348 17128
rect 12303 17088 12348 17116
rect 11333 17079 11391 17085
rect 12342 17076 12348 17088
rect 12400 17088 12434 17128
rect 12400 17076 12406 17088
rect 12158 17048 12164 17060
rect 11256 17020 12164 17048
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 12544 17048 12572 17156
rect 12636 17125 12664 17292
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17184 13047 17187
rect 14274 17184 14280 17196
rect 13035 17156 14280 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 17494 17184 17500 17196
rect 17455 17156 17500 17184
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 12802 17125 12808 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12775 17119 12808 17125
rect 12775 17085 12787 17119
rect 12775 17079 12808 17085
rect 12802 17076 12808 17079
rect 12860 17076 12866 17128
rect 13446 17076 13452 17128
rect 13504 17116 13510 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 13504 17088 13553 17116
rect 13504 17076 13510 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13688 17088 13737 17116
rect 13688 17076 13694 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17085 14243 17119
rect 14185 17079 14243 17085
rect 14200 17048 14228 17079
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 17828 17088 17873 17116
rect 17828 17076 17834 17088
rect 12544 17020 14228 17048
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 14792 17020 14841 17048
rect 14792 17008 14798 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 14829 17011 14887 17017
rect 16482 17008 16488 17060
rect 16540 17008 16546 17060
rect 1118 16980 1124 16992
rect 1079 16952 1124 16980
rect 1118 16940 1124 16952
rect 1176 16940 1182 16992
rect 2406 16980 2412 16992
rect 2367 16952 2412 16980
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 2590 16940 2596 16992
rect 2648 16940 2654 16992
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 2832 16952 3065 16980
rect 2832 16940 2838 16952
rect 3053 16949 3065 16952
rect 3099 16949 3111 16983
rect 3053 16943 3111 16949
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 4709 16983 4767 16989
rect 4709 16980 4721 16983
rect 4580 16952 4721 16980
rect 4580 16940 4586 16952
rect 4709 16949 4721 16952
rect 4755 16949 4767 16983
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 4709 16943 4767 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 8159 16983 8217 16989
rect 5500 16952 5545 16980
rect 5500 16940 5506 16952
rect 8159 16949 8171 16983
rect 8205 16980 8217 16983
rect 8754 16980 8760 16992
rect 8205 16952 8760 16980
rect 8205 16949 8217 16952
rect 8159 16943 8217 16949
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 13078 16980 13084 16992
rect 12584 16952 13084 16980
rect 12584 16940 12590 16952
rect 13078 16940 13084 16952
rect 13136 16980 13142 16992
rect 13630 16980 13636 16992
rect 13136 16952 13636 16980
rect 13136 16940 13142 16952
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 16025 16983 16083 16989
rect 16025 16980 16037 16983
rect 14516 16952 16037 16980
rect 14516 16940 14522 16952
rect 16025 16949 16037 16952
rect 16071 16949 16083 16983
rect 16025 16943 16083 16949
rect 184 16890 18920 16912
rect 184 16838 3106 16890
rect 3158 16838 3170 16890
rect 3222 16838 3234 16890
rect 3286 16838 3298 16890
rect 3350 16838 3362 16890
rect 3414 16838 6206 16890
rect 6258 16838 6270 16890
rect 6322 16838 6334 16890
rect 6386 16838 6398 16890
rect 6450 16838 6462 16890
rect 6514 16838 9306 16890
rect 9358 16838 9370 16890
rect 9422 16838 9434 16890
rect 9486 16838 9498 16890
rect 9550 16838 9562 16890
rect 9614 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 12534 16890
rect 12586 16838 12598 16890
rect 12650 16838 12662 16890
rect 12714 16838 15506 16890
rect 15558 16838 15570 16890
rect 15622 16838 15634 16890
rect 15686 16838 15698 16890
rect 15750 16838 15762 16890
rect 15814 16838 18606 16890
rect 18658 16838 18670 16890
rect 18722 16838 18734 16890
rect 18786 16838 18798 16890
rect 18850 16838 18862 16890
rect 18914 16838 18920 16890
rect 184 16816 18920 16838
rect 2777 16779 2835 16785
rect 2777 16745 2789 16779
rect 2823 16776 2835 16779
rect 2958 16776 2964 16788
rect 2823 16748 2964 16776
rect 2823 16745 2835 16748
rect 2777 16739 2835 16745
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 4430 16736 4436 16788
rect 4488 16736 4494 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5718 16776 5724 16788
rect 5132 16748 5724 16776
rect 5132 16736 5138 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 7699 16779 7757 16785
rect 7699 16745 7711 16779
rect 7745 16776 7757 16779
rect 8386 16776 8392 16788
rect 7745 16748 8392 16776
rect 7745 16745 7757 16748
rect 7699 16739 7757 16745
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 12621 16779 12679 16785
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12802 16776 12808 16788
rect 12667 16748 12808 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13357 16779 13415 16785
rect 13357 16745 13369 16779
rect 13403 16776 13415 16779
rect 13403 16748 14596 16776
rect 13403 16745 13415 16748
rect 13357 16739 13415 16745
rect 3786 16668 3792 16720
rect 3844 16708 3850 16720
rect 4448 16708 4476 16736
rect 3844 16680 4476 16708
rect 3844 16668 3850 16680
rect 5166 16668 5172 16720
rect 5224 16708 5230 16720
rect 5261 16711 5319 16717
rect 5261 16708 5273 16711
rect 5224 16680 5273 16708
rect 5224 16668 5230 16680
rect 5261 16677 5273 16680
rect 5307 16677 5319 16711
rect 5261 16671 5319 16677
rect 8110 16668 8116 16720
rect 8168 16668 8174 16720
rect 9950 16708 9956 16720
rect 9911 16680 9956 16708
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12989 16711 13047 16717
rect 12989 16708 13001 16711
rect 12124 16680 13001 16708
rect 12124 16668 12130 16680
rect 12989 16677 13001 16680
rect 13035 16677 13047 16711
rect 12989 16671 13047 16677
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 10042 16640 10048 16652
rect 9539 16612 10048 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 12250 16600 12256 16652
rect 12308 16600 12314 16652
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12894 16640 12900 16652
rect 12391 16612 12756 16640
rect 12855 16612 12900 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 2866 16532 2872 16584
rect 2924 16572 2930 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 2924 16544 4261 16572
rect 2924 16532 2930 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16541 4583 16575
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 4525 16535 4583 16541
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 4540 16436 4568 16535
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 12268 16572 12296 16600
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 12268 16544 12633 16572
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12728 16572 12756 16612
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 13078 16640 13084 16652
rect 13004 16612 13084 16640
rect 13004 16572 13032 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 14277 16643 14335 16649
rect 13679 16612 14228 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 13354 16572 13360 16584
rect 12728 16544 13032 16572
rect 13315 16544 13360 16572
rect 12621 16535 12679 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 9916 16476 11253 16504
rect 9916 16464 9922 16476
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 14200 16504 14228 16612
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14458 16640 14464 16652
rect 14323 16612 14464 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 14568 16640 14596 16748
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15105 16779 15163 16785
rect 15105 16776 15117 16779
rect 14884 16748 15117 16776
rect 14884 16736 14890 16748
rect 15105 16745 15117 16748
rect 15151 16745 15163 16779
rect 15105 16739 15163 16745
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 15252 16748 15485 16776
rect 15252 16736 15258 16748
rect 15473 16745 15485 16748
rect 15519 16745 15531 16779
rect 15473 16739 15531 16745
rect 16666 16736 16672 16788
rect 16724 16776 16730 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 16724 16748 18245 16776
rect 16724 16736 16730 16748
rect 18233 16745 18245 16748
rect 18279 16745 18291 16779
rect 18233 16739 18291 16745
rect 15841 16711 15899 16717
rect 15841 16708 15853 16711
rect 15304 16680 15853 16708
rect 15194 16640 15200 16652
rect 14568 16612 15200 16640
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 14829 16575 14887 16581
rect 14829 16572 14841 16575
rect 14792 16544 14841 16572
rect 14792 16532 14798 16544
rect 14829 16541 14841 16544
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15013 16575 15071 16581
rect 15013 16572 15025 16575
rect 14976 16544 15025 16572
rect 14976 16532 14982 16544
rect 15013 16541 15025 16544
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 15304 16504 15332 16680
rect 15841 16677 15853 16680
rect 15887 16677 15899 16711
rect 15841 16671 15899 16677
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15436 16612 15761 16640
rect 15436 16600 15442 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16640 18015 16643
rect 18414 16640 18420 16652
rect 18003 16612 18420 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 14200 16476 15332 16504
rect 11241 16467 11299 16473
rect 4488 16408 4568 16436
rect 6733 16439 6791 16445
rect 4488 16396 4494 16408
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 6822 16436 6828 16448
rect 6779 16408 6828 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 12437 16439 12495 16445
rect 12437 16436 12449 16439
rect 12216 16408 12449 16436
rect 12216 16396 12222 16408
rect 12437 16405 12449 16408
rect 12483 16436 12495 16439
rect 12802 16436 12808 16448
rect 12483 16408 12808 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 12802 16396 12808 16408
rect 12860 16436 12866 16448
rect 13446 16436 13452 16448
rect 12860 16408 13452 16436
rect 12860 16396 12866 16408
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 14185 16439 14243 16445
rect 13596 16408 13641 16436
rect 13596 16396 13602 16408
rect 14185 16405 14197 16439
rect 14231 16436 14243 16439
rect 14366 16436 14372 16448
rect 14231 16408 14372 16436
rect 14231 16405 14243 16408
rect 14185 16399 14243 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 184 16346 18860 16368
rect 184 16294 1556 16346
rect 1608 16294 1620 16346
rect 1672 16294 1684 16346
rect 1736 16294 1748 16346
rect 1800 16294 1812 16346
rect 1864 16294 4656 16346
rect 4708 16294 4720 16346
rect 4772 16294 4784 16346
rect 4836 16294 4848 16346
rect 4900 16294 4912 16346
rect 4964 16294 7756 16346
rect 7808 16294 7820 16346
rect 7872 16294 7884 16346
rect 7936 16294 7948 16346
rect 8000 16294 8012 16346
rect 8064 16294 10856 16346
rect 10908 16294 10920 16346
rect 10972 16294 10984 16346
rect 11036 16294 11048 16346
rect 11100 16294 11112 16346
rect 11164 16294 13956 16346
rect 14008 16294 14020 16346
rect 14072 16294 14084 16346
rect 14136 16294 14148 16346
rect 14200 16294 14212 16346
rect 14264 16294 17056 16346
rect 17108 16294 17120 16346
rect 17172 16294 17184 16346
rect 17236 16294 17248 16346
rect 17300 16294 17312 16346
rect 17364 16294 18860 16346
rect 184 16272 18860 16294
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5776 16204 5825 16232
rect 5776 16192 5782 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 5813 16195 5871 16201
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 9030 16232 9036 16244
rect 7239 16204 9036 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9401 16235 9459 16241
rect 9401 16232 9413 16235
rect 9180 16204 9413 16232
rect 9180 16192 9186 16204
rect 9401 16201 9413 16204
rect 9447 16201 9459 16235
rect 10042 16232 10048 16244
rect 10003 16204 10048 16232
rect 9401 16195 9459 16201
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 10376 16204 12449 16232
rect 10376 16192 10382 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 12437 16195 12495 16201
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 1394 16124 1400 16176
rect 1452 16164 1458 16176
rect 2685 16167 2743 16173
rect 2685 16164 2697 16167
rect 1452 16136 2697 16164
rect 1452 16124 1458 16136
rect 2685 16133 2697 16136
rect 2731 16133 2743 16167
rect 2685 16127 2743 16133
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2130 16096 2136 16108
rect 1811 16068 2136 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 2130 16056 2136 16068
rect 2188 16096 2194 16108
rect 2498 16096 2504 16108
rect 2188 16068 2504 16096
rect 2188 16056 2194 16068
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 4430 16096 4436 16108
rect 4391 16068 4436 16096
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16096 6699 16099
rect 7282 16096 7288 16108
rect 6687 16068 7288 16096
rect 6687 16065 6699 16068
rect 6641 16059 6699 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7466 16096 7472 16108
rect 7427 16068 7472 16096
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 8754 16096 8760 16108
rect 8715 16068 8760 16096
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 13832 16096 13860 16192
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 13832 16068 15945 16096
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 934 15988 940 16040
rect 992 16028 998 16040
rect 1946 16028 1952 16040
rect 992 16000 1952 16028
rect 992 15988 998 16000
rect 1946 15988 1952 16000
rect 2004 16028 2010 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2004 16000 2605 16028
rect 2004 15988 2010 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 2832 16000 2877 16028
rect 2832 15988 2838 16000
rect 4522 15988 4528 16040
rect 4580 16028 4586 16040
rect 4689 16031 4747 16037
rect 4689 16028 4701 16031
rect 4580 16000 4701 16028
rect 4580 15988 4586 16000
rect 4689 15997 4701 16000
rect 4735 15997 4747 16031
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 4689 15991 4747 15997
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 7248 16000 7573 16028
rect 7248 15988 7254 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 15997 10103 16031
rect 16298 16028 16304 16040
rect 16259 16000 16304 16028
rect 10045 15991 10103 15997
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15960 1915 15963
rect 2038 15960 2044 15972
rect 1903 15932 2044 15960
rect 1903 15929 1915 15932
rect 1857 15923 1915 15929
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 10060 15960 10088 15991
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 8260 15932 10088 15960
rect 11149 15963 11207 15969
rect 8260 15920 8266 15932
rect 11149 15929 11161 15963
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2314 15892 2320 15904
rect 2004 15864 2049 15892
rect 2275 15864 2320 15892
rect 2004 15852 2010 15864
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 6733 15895 6791 15901
rect 6733 15861 6745 15895
rect 6779 15892 6791 15895
rect 7006 15892 7012 15904
rect 6779 15864 7012 15892
rect 6779 15861 6791 15864
rect 6733 15855 6791 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10594 15892 10600 15904
rect 9916 15864 10600 15892
rect 9916 15852 9922 15864
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 11164 15892 11192 15923
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 15289 15963 15347 15969
rect 15289 15960 15301 15963
rect 15068 15932 15301 15960
rect 15068 15920 15074 15932
rect 15289 15929 15301 15932
rect 15335 15929 15347 15963
rect 15289 15923 15347 15929
rect 16850 15920 16856 15972
rect 16908 15920 16914 15972
rect 10652 15864 11192 15892
rect 10652 15852 10658 15864
rect 17678 15852 17684 15904
rect 17736 15901 17742 15904
rect 17736 15895 17785 15901
rect 17736 15861 17739 15895
rect 17773 15861 17785 15895
rect 17736 15855 17785 15861
rect 17736 15852 17742 15855
rect 184 15802 18920 15824
rect 184 15750 3106 15802
rect 3158 15750 3170 15802
rect 3222 15750 3234 15802
rect 3286 15750 3298 15802
rect 3350 15750 3362 15802
rect 3414 15750 6206 15802
rect 6258 15750 6270 15802
rect 6322 15750 6334 15802
rect 6386 15750 6398 15802
rect 6450 15750 6462 15802
rect 6514 15750 9306 15802
rect 9358 15750 9370 15802
rect 9422 15750 9434 15802
rect 9486 15750 9498 15802
rect 9550 15750 9562 15802
rect 9614 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 12534 15802
rect 12586 15750 12598 15802
rect 12650 15750 12662 15802
rect 12714 15750 15506 15802
rect 15558 15750 15570 15802
rect 15622 15750 15634 15802
rect 15686 15750 15698 15802
rect 15750 15750 15762 15802
rect 15814 15750 18606 15802
rect 18658 15750 18670 15802
rect 18722 15750 18734 15802
rect 18786 15750 18798 15802
rect 18850 15750 18862 15802
rect 18914 15750 18920 15802
rect 184 15728 18920 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 1176 15660 1501 15688
rect 1176 15648 1182 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1489 15651 1547 15657
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 5721 15691 5779 15697
rect 5721 15657 5733 15691
rect 5767 15688 5779 15691
rect 7190 15688 7196 15700
rect 5767 15660 7196 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 8260 15660 8309 15688
rect 8260 15648 8266 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 11609 15691 11667 15697
rect 11609 15657 11621 15691
rect 11655 15688 11667 15691
rect 11698 15688 11704 15700
rect 11655 15660 11704 15688
rect 11655 15657 11667 15660
rect 11609 15651 11667 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12802 15688 12808 15700
rect 12790 15648 12808 15688
rect 12860 15648 12866 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13354 15688 13360 15700
rect 13127 15660 13360 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 14001 15691 14059 15697
rect 14001 15657 14013 15691
rect 14047 15688 14059 15691
rect 14274 15688 14280 15700
rect 14047 15660 14280 15688
rect 14047 15657 14059 15660
rect 14001 15651 14059 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 16298 15648 16304 15700
rect 16356 15688 16362 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 16356 15660 17141 15688
rect 16356 15648 16362 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 7009 15623 7067 15629
rect 7009 15589 7021 15623
rect 7055 15620 7067 15623
rect 9585 15623 9643 15629
rect 9585 15620 9597 15623
rect 7055 15592 9597 15620
rect 7055 15589 7067 15592
rect 7009 15583 7067 15589
rect 9585 15589 9597 15592
rect 9631 15620 9643 15623
rect 9674 15620 9680 15632
rect 9631 15592 9680 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 12790 15567 12818 15648
rect 934 15552 940 15564
rect 895 15524 940 15552
rect 934 15512 940 15524
rect 992 15512 998 15564
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 2866 15552 2872 15564
rect 1627 15524 2872 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 9968 15484 9996 15515
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10318 15552 10324 15564
rect 10100 15524 10145 15552
rect 10279 15524 10324 15552
rect 10100 15512 10106 15524
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 12066 15552 12072 15564
rect 10551 15524 12072 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12785 15561 12843 15567
rect 12894 15561 12900 15564
rect 12677 15555 12735 15561
rect 12677 15552 12689 15555
rect 12216 15524 12689 15552
rect 12216 15512 12222 15524
rect 12677 15521 12689 15524
rect 12723 15521 12735 15555
rect 12785 15527 12797 15561
rect 12831 15527 12843 15561
rect 12785 15521 12843 15527
rect 12677 15515 12735 15521
rect 12893 15515 12900 15561
rect 12952 15552 12958 15564
rect 14734 15552 14740 15564
rect 12952 15524 12993 15552
rect 13832 15524 14740 15552
rect 12894 15512 12900 15515
rect 12952 15512 12958 15524
rect 11330 15484 11336 15496
rect 9968 15456 11336 15484
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 13832 15493 13860 15524
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 16298 15512 16304 15564
rect 16356 15552 16362 15564
rect 16485 15555 16543 15561
rect 16485 15552 16497 15555
rect 16356 15524 16497 15552
rect 16356 15512 16362 15524
rect 16485 15521 16497 15524
rect 16531 15521 16543 15555
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 16485 15515 16543 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15484 11943 15487
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 11931 15456 13829 15484
rect 11931 15453 11943 15456
rect 11885 15447 11943 15453
rect 13817 15453 13829 15456
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 14274 15484 14280 15496
rect 13955 15456 14280 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 10321 15419 10379 15425
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 11514 15416 11520 15428
rect 10367 15388 11520 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 11514 15376 11520 15388
rect 11572 15376 11578 15428
rect 11606 15376 11612 15428
rect 11664 15416 11670 15428
rect 11716 15416 11744 15447
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 17678 15484 17684 15496
rect 16500 15456 17684 15484
rect 16500 15416 16528 15456
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 17773 15487 17831 15493
rect 17773 15453 17785 15487
rect 17819 15484 17831 15487
rect 17862 15484 17868 15496
rect 17819 15456 17868 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 11664 15388 16528 15416
rect 11664 15376 11670 15388
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 18233 15419 18291 15425
rect 18233 15416 18245 15419
rect 16632 15388 18245 15416
rect 16632 15376 16638 15388
rect 18233 15385 18245 15388
rect 18279 15385 18291 15419
rect 18233 15379 18291 15385
rect 845 15351 903 15357
rect 845 15317 857 15351
rect 891 15348 903 15351
rect 1302 15348 1308 15360
rect 891 15320 1308 15348
rect 891 15317 903 15320
rect 845 15311 903 15317
rect 1302 15308 1308 15320
rect 1360 15308 1366 15360
rect 11238 15348 11244 15360
rect 11199 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 14366 15348 14372 15360
rect 14327 15320 14372 15348
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 15197 15351 15255 15357
rect 15197 15348 15209 15351
rect 15068 15320 15209 15348
rect 15068 15308 15074 15320
rect 15197 15317 15209 15320
rect 15243 15317 15255 15351
rect 15197 15311 15255 15317
rect 184 15258 18860 15280
rect 184 15206 1556 15258
rect 1608 15206 1620 15258
rect 1672 15206 1684 15258
rect 1736 15206 1748 15258
rect 1800 15206 1812 15258
rect 1864 15206 4656 15258
rect 4708 15206 4720 15258
rect 4772 15206 4784 15258
rect 4836 15206 4848 15258
rect 4900 15206 4912 15258
rect 4964 15206 7756 15258
rect 7808 15206 7820 15258
rect 7872 15206 7884 15258
rect 7936 15206 7948 15258
rect 8000 15206 8012 15258
rect 8064 15206 10856 15258
rect 10908 15206 10920 15258
rect 10972 15206 10984 15258
rect 11036 15206 11048 15258
rect 11100 15206 11112 15258
rect 11164 15206 13956 15258
rect 14008 15206 14020 15258
rect 14072 15206 14084 15258
rect 14136 15206 14148 15258
rect 14200 15206 14212 15258
rect 14264 15206 17056 15258
rect 17108 15206 17120 15258
rect 17172 15206 17184 15258
rect 17236 15206 17248 15258
rect 17300 15206 17312 15258
rect 17364 15206 18860 15258
rect 184 15184 18860 15206
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2682 15144 2688 15156
rect 2096 15116 2688 15144
rect 2096 15104 2102 15116
rect 2682 15104 2688 15116
rect 2740 15144 2746 15156
rect 3513 15147 3571 15153
rect 3513 15144 3525 15147
rect 2740 15116 3525 15144
rect 2740 15104 2746 15116
rect 3513 15113 3525 15116
rect 3559 15113 3571 15147
rect 3513 15107 3571 15113
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 9272 15116 9505 15144
rect 9272 15104 9278 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9493 15107 9551 15113
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10100 15116 10149 15144
rect 10100 15104 10106 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 11149 15147 11207 15153
rect 11149 15113 11161 15147
rect 11195 15144 11207 15147
rect 11330 15144 11336 15156
rect 11195 15116 11336 15144
rect 11195 15113 11207 15116
rect 11149 15107 11207 15113
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 16942 15144 16948 15156
rect 16540 15116 16948 15144
rect 16540 15104 16546 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17862 15104 17868 15156
rect 17920 15153 17926 15156
rect 17920 15147 17969 15153
rect 17920 15113 17923 15147
rect 17957 15113 17969 15147
rect 17920 15107 17969 15113
rect 17920 15104 17926 15107
rect 4985 15079 5043 15085
rect 4985 15045 4997 15079
rect 5031 15076 5043 15079
rect 5031 15048 6500 15076
rect 5031 15045 5043 15048
rect 4985 15039 5043 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2038 15008 2044 15020
rect 1811 14980 2044 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 4430 14968 4436 15020
rect 4488 15008 4494 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 4488 14980 6377 15008
rect 4488 14968 4494 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6472 15008 6500 15048
rect 10318 15036 10324 15088
rect 10376 15076 10382 15088
rect 10376 15048 11744 15076
rect 10376 15036 10382 15048
rect 8113 15011 8171 15017
rect 6472 14980 7880 15008
rect 6365 14971 6423 14977
rect 3970 14940 3976 14952
rect 3931 14912 3976 14940
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4154 14940 4160 14952
rect 4115 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 4982 14940 4988 14952
rect 4847 14912 4988 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5776 14912 5917 14940
rect 5776 14900 5782 14912
rect 5905 14909 5917 14912
rect 5951 14909 5963 14943
rect 5905 14903 5963 14909
rect 2041 14875 2099 14881
rect 2041 14841 2053 14875
rect 2087 14872 2099 14875
rect 2314 14872 2320 14884
rect 2087 14844 2320 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2314 14832 2320 14844
rect 2372 14832 2378 14884
rect 3786 14872 3792 14884
rect 3266 14844 3792 14872
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 6914 14872 6920 14884
rect 6687 14844 6920 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7852 14872 7880 14980
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8159 14980 8953 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8941 14977 8953 14980
rect 8987 15008 8999 15011
rect 10502 15008 10508 15020
rect 8987 14980 10508 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 11606 15008 11612 15020
rect 11567 14980 11612 15008
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 11716 15017 11744 15048
rect 12250 15036 12256 15088
rect 12308 15076 12314 15088
rect 13725 15079 13783 15085
rect 12308 15048 12388 15076
rect 12308 15036 12314 15048
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 12360 15008 12388 15048
rect 13725 15045 13737 15079
rect 13771 15045 13783 15079
rect 13725 15039 13783 15045
rect 12360 14980 13124 15008
rect 10228 14943 10286 14949
rect 10228 14909 10240 14943
rect 10274 14909 10286 14943
rect 10228 14903 10286 14909
rect 8110 14872 8116 14884
rect 7852 14858 8116 14872
rect 7866 14844 8116 14858
rect 8110 14832 8116 14844
rect 8168 14832 8174 14884
rect 10243 14872 10271 14903
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10376 14912 10421 14940
rect 10376 14900 10382 14912
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11296 14912 11529 14940
rect 11296 14900 11302 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11716 14940 11744 14971
rect 12158 14940 12164 14952
rect 11716 14912 12164 14940
rect 11517 14903 11575 14909
rect 12158 14900 12164 14912
rect 12216 14940 12222 14952
rect 12360 14949 12388 14980
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 12216 14912 12265 14940
rect 12216 14900 12222 14912
rect 12253 14909 12265 14912
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 12894 14940 12900 14952
rect 12483 14912 12900 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 11790 14872 11796 14884
rect 10243 14844 11796 14872
rect 11790 14832 11796 14844
rect 11848 14872 11854 14884
rect 12452 14872 12480 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 11848 14844 12480 14872
rect 13096 14872 13124 14980
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13740 14940 13768 15039
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14056 14980 14289 15008
rect 14056 14968 14062 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 14976 14980 15393 15008
rect 14976 14968 14982 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16758 15008 16764 15020
rect 16163 14980 16764 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 13219 14912 13768 14940
rect 14093 14943 14151 14949
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14366 14940 14372 14952
rect 14139 14912 14372 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15102 14940 15108 14952
rect 15063 14912 15108 14940
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15838 14940 15844 14952
rect 15335 14912 15844 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 13096 14844 14596 14872
rect 11848 14832 11854 14844
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4522 14804 4528 14816
rect 4203 14776 4528 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 5353 14807 5411 14813
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5534 14804 5540 14816
rect 5399 14776 5540 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 9030 14804 9036 14816
rect 8991 14776 9036 14804
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 9180 14776 9225 14804
rect 9180 14764 9186 14776
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 10318 14804 10324 14816
rect 9824 14776 10324 14804
rect 9824 14764 9830 14776
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 12621 14807 12679 14813
rect 12621 14773 12633 14807
rect 12667 14804 12679 14807
rect 12894 14804 12900 14816
rect 12667 14776 12900 14804
rect 12667 14773 12679 14776
rect 12621 14767 12679 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13078 14804 13084 14816
rect 13039 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 14182 14804 14188 14816
rect 14143 14776 14188 14804
rect 14182 14764 14188 14776
rect 14240 14804 14246 14816
rect 14458 14804 14464 14816
rect 14240 14776 14464 14804
rect 14240 14764 14246 14776
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14568 14804 14596 14844
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 15212 14872 15240 14903
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16485 14943 16543 14949
rect 16485 14909 16497 14943
rect 16531 14940 16543 14943
rect 16574 14940 16580 14952
rect 16531 14912 16580 14940
rect 16531 14909 16543 14912
rect 16485 14903 16543 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 14792 14844 15240 14872
rect 14792 14832 14798 14844
rect 16850 14832 16856 14884
rect 16908 14832 16914 14884
rect 15378 14804 15384 14816
rect 14568 14776 15384 14804
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 18046 14804 18052 14816
rect 15611 14776 18052 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18414 14804 18420 14816
rect 18327 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14804 18478 14816
rect 19058 14804 19064 14816
rect 18472 14776 19064 14804
rect 18472 14764 18478 14776
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 184 14714 18920 14736
rect 184 14662 3106 14714
rect 3158 14662 3170 14714
rect 3222 14662 3234 14714
rect 3286 14662 3298 14714
rect 3350 14662 3362 14714
rect 3414 14662 6206 14714
rect 6258 14662 6270 14714
rect 6322 14662 6334 14714
rect 6386 14662 6398 14714
rect 6450 14662 6462 14714
rect 6514 14662 9306 14714
rect 9358 14662 9370 14714
rect 9422 14662 9434 14714
rect 9486 14662 9498 14714
rect 9550 14662 9562 14714
rect 9614 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 12534 14714
rect 12586 14662 12598 14714
rect 12650 14662 12662 14714
rect 12714 14662 15506 14714
rect 15558 14662 15570 14714
rect 15622 14662 15634 14714
rect 15686 14662 15698 14714
rect 15750 14662 15762 14714
rect 15814 14662 18606 14714
rect 18658 14662 18670 14714
rect 18722 14662 18734 14714
rect 18786 14662 18798 14714
rect 18850 14662 18862 14714
rect 18914 14662 18920 14714
rect 184 14640 18920 14662
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 4154 14600 4160 14612
rect 3375 14572 4160 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 7006 14600 7012 14612
rect 6967 14572 7012 14600
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14600 8631 14603
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8619 14572 9137 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 16942 14600 16948 14612
rect 9125 14563 9183 14569
rect 12360 14572 16948 14600
rect 934 14492 940 14544
rect 992 14532 998 14544
rect 1121 14535 1179 14541
rect 1121 14532 1133 14535
rect 992 14504 1133 14532
rect 992 14492 998 14504
rect 1121 14501 1133 14504
rect 1167 14532 1179 14535
rect 1167 14504 2360 14532
rect 1167 14501 1179 14504
rect 1121 14495 1179 14501
rect 1210 14464 1216 14476
rect 1171 14436 1216 14464
rect 1210 14424 1216 14436
rect 1268 14424 1274 14476
rect 2332 14464 2360 14504
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 3513 14535 3571 14541
rect 3513 14532 3525 14535
rect 2832 14504 3525 14532
rect 2832 14492 2838 14504
rect 3513 14501 3525 14504
rect 3559 14501 3571 14535
rect 5534 14532 5540 14544
rect 5495 14504 5540 14532
rect 3513 14495 3571 14501
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5810 14492 5816 14544
rect 5868 14532 5874 14544
rect 5868 14504 6026 14532
rect 5868 14492 5874 14504
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 12360 14532 12388 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 12618 14532 12624 14544
rect 8168 14504 12388 14532
rect 12531 14504 12624 14532
rect 8168 14492 8174 14504
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 2332 14436 3617 14464
rect 3528 14408 3556 14436
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 5261 14467 5319 14473
rect 5261 14464 5273 14467
rect 4488 14436 5273 14464
rect 4488 14424 4494 14436
rect 5261 14433 5273 14436
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14464 8263 14467
rect 9217 14467 9275 14473
rect 8251 14436 9168 14464
rect 8251 14433 8263 14436
rect 8205 14427 8263 14433
rect 1029 14399 1087 14405
rect 1029 14365 1041 14399
rect 1075 14396 1087 14399
rect 2130 14396 2136 14408
rect 1075 14368 2136 14396
rect 1075 14365 1087 14368
rect 1029 14359 1087 14365
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 2958 14396 2964 14408
rect 2188 14368 2964 14396
rect 2188 14356 2194 14368
rect 2958 14356 2964 14368
rect 3016 14396 3022 14408
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 3016 14368 3157 14396
rect 3016 14356 3022 14368
rect 3145 14365 3157 14368
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3510 14356 3516 14408
rect 3568 14356 3574 14408
rect 3697 14399 3755 14405
rect 3697 14365 3709 14399
rect 3743 14365 3755 14399
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 3697 14359 3755 14365
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 3712 14328 3740 14359
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 9140 14396 9168 14436
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 10042 14464 10048 14476
rect 9263 14436 10048 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 12360 14473 12388 14504
rect 12618 14492 12624 14504
rect 12676 14532 12682 14544
rect 12676 14504 14136 14532
rect 12676 14492 12682 14504
rect 11333 14467 11391 14473
rect 11333 14464 11345 14467
rect 11296 14436 11345 14464
rect 11296 14424 11302 14436
rect 11333 14433 11345 14436
rect 11379 14433 11391 14467
rect 11333 14427 11391 14433
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14433 12403 14467
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 12345 14427 12403 14433
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13538 14464 13544 14476
rect 13219 14436 13544 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 9140 14368 10272 14396
rect 9033 14359 9091 14365
rect 3660 14300 3740 14328
rect 3660 14288 3666 14300
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 2130 14260 2136 14272
rect 1627 14232 2136 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 9048 14260 9076 14359
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 10134 14328 10140 14340
rect 9631 14300 10140 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10244 14328 10272 14368
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 12952 14368 13369 14396
rect 12952 14356 12958 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13998 14396 14004 14408
rect 13504 14368 14004 14396
rect 13504 14356 13510 14368
rect 13998 14356 14004 14368
rect 14056 14356 14062 14408
rect 14108 14396 14136 14504
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 16850 14532 16856 14544
rect 16080 14504 16856 14532
rect 16080 14492 16086 14504
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14458 14464 14464 14476
rect 14323 14436 14464 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 17770 14464 17776 14476
rect 16816 14436 17776 14464
rect 16816 14424 16822 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18046 14464 18052 14476
rect 18007 14436 18052 14464
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 18233 14467 18291 14473
rect 18233 14433 18245 14467
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 16022 14396 16028 14408
rect 14108 14368 16028 14396
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14396 16543 14399
rect 17129 14399 17187 14405
rect 17129 14396 17141 14399
rect 16531 14368 17141 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 17129 14365 17141 14368
rect 17175 14365 17187 14399
rect 17129 14359 17187 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 17954 14396 17960 14408
rect 17727 14368 17960 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 13722 14328 13728 14340
rect 10244 14300 13728 14328
rect 9766 14260 9772 14272
rect 9048 14232 9772 14260
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 10045 14263 10103 14269
rect 10045 14229 10057 14263
rect 10091 14260 10103 14263
rect 10244 14260 10272 14300
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 14016 14328 14044 14356
rect 15378 14328 15384 14340
rect 14016 14300 15384 14328
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 18248 14328 18276 14427
rect 16908 14300 18276 14328
rect 16908 14288 16914 14300
rect 11330 14260 11336 14272
rect 10091 14232 10272 14260
rect 11291 14232 11336 14260
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14260 13323 14263
rect 13814 14260 13820 14272
rect 13311 14232 13820 14260
rect 13311 14229 13323 14232
rect 13265 14223 13323 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 15013 14263 15071 14269
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 16114 14260 16120 14272
rect 15059 14232 16120 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 16114 14220 16120 14232
rect 16172 14260 16178 14272
rect 17678 14260 17684 14272
rect 16172 14232 17684 14260
rect 16172 14220 16178 14232
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 18138 14260 18144 14272
rect 18099 14232 18144 14260
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 184 14170 18860 14192
rect 184 14118 1556 14170
rect 1608 14118 1620 14170
rect 1672 14118 1684 14170
rect 1736 14118 1748 14170
rect 1800 14118 1812 14170
rect 1864 14118 4656 14170
rect 4708 14118 4720 14170
rect 4772 14118 4784 14170
rect 4836 14118 4848 14170
rect 4900 14118 4912 14170
rect 4964 14118 7756 14170
rect 7808 14118 7820 14170
rect 7872 14118 7884 14170
rect 7936 14118 7948 14170
rect 8000 14118 8012 14170
rect 8064 14118 10856 14170
rect 10908 14118 10920 14170
rect 10972 14118 10984 14170
rect 11036 14118 11048 14170
rect 11100 14118 11112 14170
rect 11164 14118 13956 14170
rect 14008 14118 14020 14170
rect 14072 14118 14084 14170
rect 14136 14118 14148 14170
rect 14200 14118 14212 14170
rect 14264 14118 17056 14170
rect 17108 14118 17120 14170
rect 17172 14118 17184 14170
rect 17236 14118 17248 14170
rect 17300 14118 17312 14170
rect 17364 14118 18860 14170
rect 184 14096 18860 14118
rect 3510 14056 3516 14068
rect 3471 14028 3516 14056
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3660 14028 5304 14056
rect 3660 14016 3666 14028
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4430 13920 4436 13932
rect 4203 13892 4436 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 2038 13852 2044 13864
rect 1811 13824 2044 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 4522 13852 4528 13864
rect 4483 13824 4528 13852
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 5276 13852 5304 14028
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 6972 14028 7113 14056
rect 6972 14016 6978 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 8352 14028 9321 14056
rect 8352 14016 8358 14028
rect 9309 14025 9321 14028
rect 9355 14056 9367 14059
rect 12894 14056 12900 14068
rect 9355 14028 12900 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 15838 14056 15844 14068
rect 15120 14028 15844 14056
rect 13630 13948 13636 14000
rect 13688 13988 13694 14000
rect 15120 13988 15148 14028
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16472 14059 16530 14065
rect 16472 14025 16484 14059
rect 16518 14056 16530 14059
rect 17954 14056 17960 14068
rect 16518 14028 17816 14056
rect 17915 14028 17960 14056
rect 16518 14025 16530 14028
rect 16472 14019 16530 14025
rect 13688 13960 15148 13988
rect 17788 13988 17816 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18230 13988 18236 14000
rect 17788 13960 18236 13988
rect 13688 13948 13694 13960
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 7650 13920 7656 13932
rect 7340 13892 7656 13920
rect 7340 13880 7346 13892
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11330 13920 11336 13932
rect 11195 13892 11336 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 11514 13920 11520 13932
rect 11475 13892 11520 13920
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 12986 13920 12992 13932
rect 12947 13892 12992 13920
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 15028 13929 15056 13960
rect 18230 13948 18236 13960
rect 18288 13948 18294 14000
rect 14829 13923 14887 13929
rect 14829 13920 14841 13923
rect 14792 13892 14841 13920
rect 14792 13880 14798 13892
rect 14829 13889 14841 13892
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15197 13923 15255 13929
rect 15197 13920 15209 13923
rect 15160 13892 15209 13920
rect 15160 13880 15166 13892
rect 15197 13889 15209 13892
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15378 13920 15384 13932
rect 15335 13892 15384 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 5951 13855 6009 13861
rect 5951 13852 5963 13855
rect 5276 13824 5963 13852
rect 5951 13821 5963 13824
rect 5997 13852 6009 13855
rect 7098 13852 7104 13864
rect 5997 13824 7104 13852
rect 5997 13821 6009 13824
rect 5951 13815 6009 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13852 8907 13855
rect 10042 13852 10048 13864
rect 8895 13824 10048 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 14424 13824 14473 13852
rect 14424 13812 14430 13824
rect 14461 13821 14473 13824
rect 14507 13821 14519 13855
rect 14461 13815 14519 13821
rect 14918 13812 14924 13864
rect 14976 13852 14982 13864
rect 14976 13824 15148 13852
rect 14976 13812 14982 13824
rect 3786 13784 3792 13796
rect 3174 13756 3792 13784
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 5810 13784 5816 13796
rect 5566 13756 5816 13784
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 12618 13784 12624 13796
rect 12558 13756 12624 13784
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 15120 13793 15148 13824
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13753 15163 13787
rect 15212 13784 15240 13883
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 16209 13923 16267 13929
rect 16209 13889 16221 13923
rect 16255 13920 16267 13923
rect 16574 13920 16580 13932
rect 16255 13892 16580 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 15396 13824 16252 13852
rect 15396 13784 15424 13824
rect 15212 13756 15424 13784
rect 16224 13784 16252 13824
rect 16758 13784 16764 13796
rect 16224 13756 16764 13784
rect 15105 13747 15163 13753
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 16942 13744 16948 13796
rect 17000 13744 17006 13796
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12636 13716 12664 13744
rect 12216 13688 12664 13716
rect 15381 13719 15439 13725
rect 12216 13676 12222 13688
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 16850 13716 16856 13728
rect 15427 13688 16856 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 184 13626 18920 13648
rect 184 13574 3106 13626
rect 3158 13574 3170 13626
rect 3222 13574 3234 13626
rect 3286 13574 3298 13626
rect 3350 13574 3362 13626
rect 3414 13574 6206 13626
rect 6258 13574 6270 13626
rect 6322 13574 6334 13626
rect 6386 13574 6398 13626
rect 6450 13574 6462 13626
rect 6514 13574 9306 13626
rect 9358 13574 9370 13626
rect 9422 13574 9434 13626
rect 9486 13574 9498 13626
rect 9550 13574 9562 13626
rect 9614 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 12534 13626
rect 12586 13574 12598 13626
rect 12650 13574 12662 13626
rect 12714 13574 15506 13626
rect 15558 13574 15570 13626
rect 15622 13574 15634 13626
rect 15686 13574 15698 13626
rect 15750 13574 15762 13626
rect 15814 13574 18606 13626
rect 18658 13574 18670 13626
rect 18722 13574 18734 13626
rect 18786 13574 18798 13626
rect 18850 13574 18862 13626
rect 18914 13574 18920 13626
rect 184 13552 18920 13574
rect 1121 13515 1179 13521
rect 1121 13481 1133 13515
rect 1167 13512 1179 13515
rect 1210 13512 1216 13524
rect 1167 13484 1216 13512
rect 1167 13481 1179 13484
rect 1121 13475 1179 13481
rect 1210 13472 1216 13484
rect 1268 13472 1274 13524
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1360 13484 1593 13512
rect 1360 13472 1366 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 3970 13512 3976 13524
rect 3651 13484 3976 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 9122 13512 9128 13524
rect 8343 13484 9128 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 10042 13512 10048 13524
rect 10003 13484 10048 13512
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10152 13484 10885 13512
rect 1489 13447 1547 13453
rect 1489 13413 1501 13447
rect 1535 13444 1547 13447
rect 5350 13444 5356 13456
rect 1535 13416 5356 13444
rect 1535 13413 1547 13416
rect 1489 13407 1547 13413
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 9585 13447 9643 13453
rect 9585 13413 9597 13447
rect 9631 13444 9643 13447
rect 9858 13444 9864 13456
rect 9631 13416 9864 13444
rect 9631 13413 9643 13416
rect 9585 13407 9643 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 2958 13336 2964 13388
rect 3016 13376 3022 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 3016 13348 3341 13376
rect 3016 13336 3022 13348
rect 3329 13345 3341 13348
rect 3375 13376 3387 13379
rect 3375 13348 4384 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1452 13280 1777 13308
rect 1452 13268 1458 13280
rect 1765 13277 1777 13280
rect 1811 13308 1823 13311
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 1811 13280 3433 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3602 13308 3608 13320
rect 3563 13280 3608 13308
rect 3421 13271 3479 13277
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 4356 13308 4384 13348
rect 4430 13336 4436 13388
rect 4488 13376 4494 13388
rect 5258 13376 5264 13388
rect 4488 13348 5264 13376
rect 4488 13336 4494 13348
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5528 13379 5586 13385
rect 5528 13376 5540 13379
rect 5368 13348 5540 13376
rect 5368 13308 5396 13348
rect 5528 13345 5540 13348
rect 5574 13376 5586 13379
rect 7282 13376 7288 13388
rect 5574 13348 7288 13376
rect 5574 13345 5586 13348
rect 5528 13339 5586 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10152 13376 10180 13484
rect 10873 13481 10885 13484
rect 10919 13512 10931 13515
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 10919 13484 13553 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 13541 13481 13553 13484
rect 13587 13512 13599 13515
rect 13630 13512 13636 13524
rect 13587 13484 13636 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 16482 13512 16488 13524
rect 16443 13484 16488 13512
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 12066 13404 12072 13456
rect 12124 13444 12130 13456
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 12124 13416 12817 13444
rect 12124 13404 12130 13416
rect 12805 13413 12817 13416
rect 12851 13444 12863 13447
rect 13357 13447 13415 13453
rect 13357 13444 13369 13447
rect 12851 13416 13369 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 13357 13413 13369 13416
rect 13403 13444 13415 13447
rect 13446 13444 13452 13456
rect 13403 13416 13452 13444
rect 13403 13413 13415 13416
rect 13357 13407 13415 13413
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 15010 13444 15016 13456
rect 14971 13416 15016 13444
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 17497 13447 17555 13453
rect 17497 13444 17509 13447
rect 16816 13416 17509 13444
rect 16816 13404 16822 13416
rect 17497 13413 17509 13416
rect 17543 13413 17555 13447
rect 17497 13407 17555 13413
rect 9999 13348 10180 13376
rect 10229 13379 10287 13385
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11514 13376 11520 13388
rect 11195 13348 11520 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 4356 13280 5396 13308
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 10244 13308 10272 13339
rect 9732 13280 10272 13308
rect 10980 13308 11008 13339
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 11790 13376 11796 13388
rect 11751 13348 11796 13376
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 13262 13376 13268 13388
rect 12759 13348 13268 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 14550 13376 14556 13388
rect 13679 13348 14556 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 14550 13336 14556 13348
rect 14608 13376 14614 13388
rect 14918 13376 14924 13388
rect 14608 13348 14924 13376
rect 14608 13336 14614 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 17586 13376 17592 13388
rect 17547 13348 17592 13376
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 11422 13308 11428 13320
rect 10980 13280 11428 13308
rect 9732 13268 9738 13280
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 11885 13243 11943 13249
rect 11885 13209 11897 13243
rect 11931 13240 11943 13243
rect 12912 13240 12940 13271
rect 11931 13212 12940 13240
rect 13357 13243 13415 13249
rect 11931 13209 11943 13212
rect 11885 13203 11943 13209
rect 13357 13209 13369 13243
rect 13403 13240 13415 13243
rect 13538 13240 13544 13252
rect 13403 13212 13544 13240
rect 13403 13209 13415 13212
rect 13357 13203 13415 13209
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 6638 13172 6644 13184
rect 6599 13144 6644 13172
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 10778 13172 10784 13184
rect 10560 13144 10784 13172
rect 10560 13132 10566 13144
rect 10778 13132 10784 13144
rect 10836 13172 10842 13184
rect 12345 13175 12403 13181
rect 12345 13172 12357 13175
rect 10836 13144 12357 13172
rect 10836 13132 10842 13144
rect 12345 13141 12357 13144
rect 12391 13141 12403 13175
rect 12345 13135 12403 13141
rect 184 13082 18860 13104
rect 184 13030 1556 13082
rect 1608 13030 1620 13082
rect 1672 13030 1684 13082
rect 1736 13030 1748 13082
rect 1800 13030 1812 13082
rect 1864 13030 4656 13082
rect 4708 13030 4720 13082
rect 4772 13030 4784 13082
rect 4836 13030 4848 13082
rect 4900 13030 4912 13082
rect 4964 13030 7756 13082
rect 7808 13030 7820 13082
rect 7872 13030 7884 13082
rect 7936 13030 7948 13082
rect 8000 13030 8012 13082
rect 8064 13030 10856 13082
rect 10908 13030 10920 13082
rect 10972 13030 10984 13082
rect 11036 13030 11048 13082
rect 11100 13030 11112 13082
rect 11164 13030 13956 13082
rect 14008 13030 14020 13082
rect 14072 13030 14084 13082
rect 14136 13030 14148 13082
rect 14200 13030 14212 13082
rect 14264 13030 17056 13082
rect 17108 13030 17120 13082
rect 17172 13030 17184 13082
rect 17236 13030 17248 13082
rect 17300 13030 17312 13082
rect 17364 13030 18860 13082
rect 184 13008 18860 13030
rect 4430 12968 4436 12980
rect 4080 12940 4436 12968
rect 4080 12841 4108 12940
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 12860 12940 13829 12968
rect 12860 12928 12866 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 10502 12900 10508 12912
rect 10060 12872 10508 12900
rect 10060 12844 10088 12872
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 10689 12903 10747 12909
rect 10689 12869 10701 12903
rect 10735 12869 10747 12903
rect 16298 12900 16304 12912
rect 16259 12872 16304 12900
rect 10689 12863 10747 12869
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12832 4123 12835
rect 7837 12835 7895 12841
rect 4111 12804 4200 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 4172 12776 4200 12804
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8754 12832 8760 12844
rect 7883 12804 8760 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 10042 12832 10048 12844
rect 9955 12804 10048 12832
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 10192 12804 10241 12832
rect 10192 12792 10198 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10704 12832 10732 12863
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 10704 12804 12909 12832
rect 10229 12795 10287 12801
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 13170 12832 13176 12844
rect 13083 12804 13176 12832
rect 12897 12795 12955 12801
rect 13170 12792 13176 12804
rect 13228 12832 13234 12844
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 13228 12804 15577 12832
rect 13228 12792 13234 12804
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 17586 12832 17592 12844
rect 15565 12795 15623 12801
rect 15764 12804 16436 12832
rect 17547 12804 17592 12832
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 1946 12724 1952 12776
rect 2004 12764 2010 12776
rect 2041 12767 2099 12773
rect 2041 12764 2053 12767
rect 2004 12736 2053 12764
rect 2004 12724 2010 12736
rect 2041 12733 2053 12736
rect 2087 12733 2099 12767
rect 2041 12727 2099 12733
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 9214 12764 9220 12776
rect 7791 12736 9220 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 11422 12764 11428 12776
rect 9539 12736 11428 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3786 12696 3792 12708
rect 3108 12668 3792 12696
rect 3108 12656 3114 12668
rect 3786 12656 3792 12668
rect 3844 12656 3850 12708
rect 4332 12699 4390 12705
rect 4332 12665 4344 12699
rect 4378 12696 4390 12699
rect 5626 12696 5632 12708
rect 4378 12668 5632 12696
rect 4378 12665 4390 12668
rect 4332 12659 4390 12665
rect 5626 12656 5632 12668
rect 5684 12696 5690 12708
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 5684 12668 5733 12696
rect 5684 12656 5690 12668
rect 5721 12665 5733 12668
rect 5767 12665 5779 12699
rect 5721 12659 5779 12665
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 9324 12696 9352 12727
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 8812 12668 9352 12696
rect 8812 12656 8818 12668
rect 1486 12588 1492 12640
rect 1544 12628 1550 12640
rect 2130 12628 2136 12640
rect 1544 12600 2136 12628
rect 1544 12588 1550 12600
rect 2130 12588 2136 12600
rect 2188 12628 2194 12640
rect 3467 12631 3525 12637
rect 3467 12628 3479 12631
rect 2188 12600 3479 12628
rect 2188 12588 2194 12600
rect 3467 12597 3479 12600
rect 3513 12597 3525 12631
rect 5442 12628 5448 12640
rect 5403 12600 5448 12628
rect 3467 12591 3525 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8846 12628 8852 12640
rect 8159 12600 8852 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9324 12628 9352 12668
rect 12158 12656 12164 12708
rect 12216 12656 12222 12708
rect 14858 12668 14964 12696
rect 14936 12640 14964 12668
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 15252 12668 15301 12696
rect 15252 12656 15258 12668
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9324 12600 10333 12628
rect 10321 12597 10333 12600
rect 10367 12628 10379 12631
rect 11425 12631 11483 12637
rect 11425 12628 11437 12631
rect 10367 12600 11437 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 11425 12597 11437 12600
rect 11471 12597 11483 12631
rect 11425 12591 11483 12597
rect 14918 12588 14924 12640
rect 14976 12588 14982 12640
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 15764 12628 15792 12804
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 16114 12764 16120 12776
rect 15979 12736 16120 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16408 12773 16436 12804
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12733 16451 12767
rect 16758 12764 16764 12776
rect 16719 12736 16764 12764
rect 16393 12727 16451 12733
rect 16316 12696 16344 12727
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 17184 12736 17417 12764
rect 17184 12724 17190 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17221 12699 17279 12705
rect 17221 12696 17233 12699
rect 16316 12668 17233 12696
rect 17221 12665 17233 12668
rect 17267 12665 17279 12699
rect 17221 12659 17279 12665
rect 15068 12600 15792 12628
rect 15068 12588 15074 12600
rect 184 12538 18920 12560
rect 184 12486 3106 12538
rect 3158 12486 3170 12538
rect 3222 12486 3234 12538
rect 3286 12486 3298 12538
rect 3350 12486 3362 12538
rect 3414 12486 6206 12538
rect 6258 12486 6270 12538
rect 6322 12486 6334 12538
rect 6386 12486 6398 12538
rect 6450 12486 6462 12538
rect 6514 12486 9306 12538
rect 9358 12486 9370 12538
rect 9422 12486 9434 12538
rect 9486 12486 9498 12538
rect 9550 12486 9562 12538
rect 9614 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 12534 12538
rect 12586 12486 12598 12538
rect 12650 12486 12662 12538
rect 12714 12486 15506 12538
rect 15558 12486 15570 12538
rect 15622 12486 15634 12538
rect 15686 12486 15698 12538
rect 15750 12486 15762 12538
rect 15814 12486 18606 12538
rect 18658 12486 18670 12538
rect 18722 12486 18734 12538
rect 18786 12486 18798 12538
rect 18850 12486 18862 12538
rect 18914 12486 18920 12538
rect 184 12464 18920 12486
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5316 12396 9352 12424
rect 5316 12384 5322 12396
rect 1670 12316 1676 12368
rect 1728 12356 1734 12368
rect 1765 12359 1823 12365
rect 1765 12356 1777 12359
rect 1728 12328 1777 12356
rect 1728 12316 1734 12328
rect 1765 12325 1777 12328
rect 1811 12325 1823 12359
rect 1765 12319 1823 12325
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 6089 12359 6147 12365
rect 5408 12328 5856 12356
rect 5408 12316 5414 12328
rect 5828 12300 5856 12328
rect 6089 12325 6101 12359
rect 6135 12356 6147 12359
rect 6457 12359 6515 12365
rect 6457 12356 6469 12359
rect 6135 12328 6469 12356
rect 6135 12325 6147 12328
rect 6089 12319 6147 12325
rect 6457 12325 6469 12328
rect 6503 12325 6515 12359
rect 6638 12356 6644 12368
rect 6599 12328 6644 12356
rect 6457 12319 6515 12325
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 8570 12316 8576 12368
rect 8628 12316 8634 12368
rect 753 12291 811 12297
rect 753 12257 765 12291
rect 799 12288 811 12291
rect 1486 12288 1492 12300
rect 799 12260 1492 12288
rect 799 12257 811 12260
rect 753 12251 811 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2133 12291 2191 12297
rect 2133 12288 2145 12291
rect 2096 12260 2145 12288
rect 2096 12248 2102 12260
rect 2133 12257 2145 12260
rect 2179 12288 2191 12291
rect 4154 12288 4160 12300
rect 2179 12260 4160 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5500 12260 5733 12288
rect 5500 12248 5506 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 6362 12288 6368 12300
rect 5868 12260 5961 12288
rect 6323 12260 6368 12288
rect 5868 12248 5874 12260
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 9324 12297 9352 12396
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 15194 12424 15200 12436
rect 14424 12396 15200 12424
rect 14424 12384 14430 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 16816 12396 17233 12424
rect 16816 12384 16822 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 17221 12387 17279 12393
rect 11238 12356 11244 12368
rect 10428 12328 11244 12356
rect 10428 12297 10456 12328
rect 11238 12316 11244 12328
rect 11296 12356 11302 12368
rect 13170 12356 13176 12368
rect 11296 12328 13176 12356
rect 11296 12316 11302 12328
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13538 12316 13544 12368
rect 13596 12316 13602 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14826 12356 14832 12368
rect 13780 12328 14832 12356
rect 13780 12316 13786 12328
rect 9309 12291 9367 12297
rect 9309 12257 9321 12291
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12257 10471 12291
rect 10413 12251 10471 12257
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 11057 12291 11115 12297
rect 10744 12260 11008 12288
rect 10744 12248 10750 12260
rect 845 12223 903 12229
rect 845 12189 857 12223
rect 891 12220 903 12223
rect 1394 12220 1400 12232
rect 891 12192 1400 12220
rect 891 12189 903 12192
rect 845 12183 903 12189
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 8570 12220 8576 12232
rect 6886 12192 8576 12220
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 6886 12152 6914 12192
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12220 9091 12223
rect 10778 12220 10784 12232
rect 9079 12192 10640 12220
rect 10739 12192 10784 12220
rect 9079 12189 9091 12192
rect 9033 12183 9091 12189
rect 5776 12124 6914 12152
rect 7561 12155 7619 12161
rect 5776 12112 5782 12124
rect 7561 12121 7573 12155
rect 7607 12152 7619 12155
rect 7650 12152 7656 12164
rect 7607 12124 7656 12152
rect 7607 12121 7619 12124
rect 7561 12115 7619 12121
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 10612 12152 10640 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10980 12229 11008 12260
rect 11057 12257 11069 12291
rect 11103 12288 11115 12291
rect 11422 12288 11428 12300
rect 11103 12260 11428 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13556 12288 13584 12316
rect 13832 12297 13860 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 16114 12356 16120 12368
rect 16075 12328 16120 12356
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 13127 12260 13584 12288
rect 13817 12291 13875 12297
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12288 14151 12291
rect 14274 12288 14280 12300
rect 14139 12260 14280 12288
rect 14139 12257 14151 12260
rect 14093 12251 14151 12257
rect 14274 12248 14280 12260
rect 14332 12288 14338 12300
rect 15010 12288 15016 12300
rect 14332 12260 15016 12288
rect 14332 12248 14338 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 11848 12192 12725 12220
rect 11848 12180 11854 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 14734 12220 14740 12232
rect 13403 12192 14740 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 14734 12180 14740 12192
rect 14792 12220 14798 12232
rect 15948 12220 15976 12251
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 17126 12288 17132 12300
rect 16632 12260 17132 12288
rect 16632 12248 16638 12260
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17402 12288 17408 12300
rect 17359 12260 17408 12288
rect 17359 12257 17371 12260
rect 17313 12251 17371 12257
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 14792 12192 15976 12220
rect 14792 12180 14798 12192
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 16080 12192 16221 12220
rect 16080 12180 16086 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 12802 12152 12808 12164
rect 10612 12124 12808 12152
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 1026 12084 1032 12096
rect 987 12056 1032 12084
rect 1026 12044 1032 12056
rect 1084 12044 1090 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 6365 12087 6423 12093
rect 6365 12084 6377 12087
rect 5592 12056 6377 12084
rect 5592 12044 5598 12056
rect 6365 12053 6377 12056
rect 6411 12053 6423 12087
rect 6365 12047 6423 12053
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10137 12087 10195 12093
rect 10137 12084 10149 12087
rect 10008 12056 10149 12084
rect 10008 12044 10014 12056
rect 10137 12053 10149 12056
rect 10183 12053 10195 12087
rect 10137 12047 10195 12053
rect 11425 12087 11483 12093
rect 11425 12053 11437 12087
rect 11471 12084 11483 12087
rect 12894 12084 12900 12096
rect 11471 12056 12900 12084
rect 11471 12053 11483 12056
rect 11425 12047 11483 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 14826 12084 14832 12096
rect 14787 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 184 11994 18860 12016
rect 184 11942 1556 11994
rect 1608 11942 1620 11994
rect 1672 11942 1684 11994
rect 1736 11942 1748 11994
rect 1800 11942 1812 11994
rect 1864 11942 4656 11994
rect 4708 11942 4720 11994
rect 4772 11942 4784 11994
rect 4836 11942 4848 11994
rect 4900 11942 4912 11994
rect 4964 11942 7756 11994
rect 7808 11942 7820 11994
rect 7872 11942 7884 11994
rect 7936 11942 7948 11994
rect 8000 11942 8012 11994
rect 8064 11942 10856 11994
rect 10908 11942 10920 11994
rect 10972 11942 10984 11994
rect 11036 11942 11048 11994
rect 11100 11942 11112 11994
rect 11164 11942 13956 11994
rect 14008 11942 14020 11994
rect 14072 11942 14084 11994
rect 14136 11942 14148 11994
rect 14200 11942 14212 11994
rect 14264 11942 17056 11994
rect 17108 11942 17120 11994
rect 17172 11942 17184 11994
rect 17236 11942 17248 11994
rect 17300 11942 17312 11994
rect 17364 11942 18860 11994
rect 184 11920 18860 11942
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 10744 11852 10793 11880
rect 10744 11840 10750 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 10781 11843 10839 11849
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15378 11880 15384 11892
rect 15335 11852 15384 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 17402 11840 17408 11892
rect 17460 11880 17466 11892
rect 17911 11883 17969 11889
rect 17911 11880 17923 11883
rect 17460 11852 17923 11880
rect 17460 11840 17466 11852
rect 17911 11849 17923 11852
rect 17957 11849 17969 11883
rect 17911 11843 17969 11849
rect 5629 11815 5687 11821
rect 5629 11781 5641 11815
rect 5675 11812 5687 11815
rect 6362 11812 6368 11824
rect 5675 11784 6368 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 6362 11772 6368 11784
rect 6420 11772 6426 11824
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 9824 11784 10180 11812
rect 9824 11772 9830 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2406 11744 2412 11756
rect 2271 11716 2412 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11744 9091 11747
rect 10042 11744 10048 11756
rect 9079 11716 10048 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10152 11753 10180 11784
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11713 10195 11747
rect 11514 11744 11520 11756
rect 10137 11707 10195 11713
rect 10244 11716 11520 11744
rect 1026 11636 1032 11688
rect 1084 11676 1090 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1084 11648 1961 11676
rect 1084 11636 1090 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 5258 11676 5264 11688
rect 5219 11648 5264 11676
rect 1949 11639 2007 11645
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5442 11685 5448 11688
rect 5415 11679 5448 11685
rect 5415 11645 5427 11679
rect 5415 11639 5448 11645
rect 5442 11636 5448 11639
rect 5500 11636 5506 11688
rect 9214 11676 9220 11688
rect 9127 11648 9220 11676
rect 9214 11636 9220 11648
rect 9272 11676 9278 11688
rect 10244 11676 10272 11716
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 15286 11744 15292 11756
rect 12406 11716 15292 11744
rect 10410 11676 10416 11688
rect 9272 11648 10272 11676
rect 10371 11648 10416 11676
rect 9272 11636 9278 11648
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11330 11676 11336 11688
rect 11195 11648 11336 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 8113 11611 8171 11617
rect 8113 11577 8125 11611
rect 8159 11608 8171 11611
rect 8202 11608 8208 11620
rect 8159 11580 8208 11608
rect 8159 11577 8171 11580
rect 8113 11571 8171 11577
rect 8202 11568 8208 11580
rect 8260 11608 8266 11620
rect 12406 11608 12434 11716
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 18138 11744 18144 11756
rect 16531 11716 18144 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 13228 11648 13553 11676
rect 13228 11636 13234 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 13541 11639 13599 11645
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 13814 11608 13820 11620
rect 8260 11580 12434 11608
rect 13775 11580 13820 11608
rect 8260 11568 8266 11580
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 15102 11608 15108 11620
rect 15015 11580 15108 11608
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 16776 11580 16882 11608
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2038 11540 2044 11552
rect 1999 11512 2044 11540
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7006 11540 7012 11552
rect 6871 11512 7012 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 9122 11540 9128 11552
rect 9083 11512 9128 11540
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 10226 11540 10232 11552
rect 9631 11512 10232 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10321 11543 10379 11549
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10686 11540 10692 11552
rect 10367 11512 10692 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11296 11512 11345 11540
rect 11296 11500 11302 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11333 11503 11391 11509
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 15120 11540 15148 11568
rect 16776 11540 16804 11580
rect 14240 11512 16804 11540
rect 14240 11500 14246 11512
rect 184 11450 18920 11472
rect 184 11398 3106 11450
rect 3158 11398 3170 11450
rect 3222 11398 3234 11450
rect 3286 11398 3298 11450
rect 3350 11398 3362 11450
rect 3414 11398 6206 11450
rect 6258 11398 6270 11450
rect 6322 11398 6334 11450
rect 6386 11398 6398 11450
rect 6450 11398 6462 11450
rect 6514 11398 9306 11450
rect 9358 11398 9370 11450
rect 9422 11398 9434 11450
rect 9486 11398 9498 11450
rect 9550 11398 9562 11450
rect 9614 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 12534 11450
rect 12586 11398 12598 11450
rect 12650 11398 12662 11450
rect 12714 11398 15506 11450
rect 15558 11398 15570 11450
rect 15622 11398 15634 11450
rect 15686 11398 15698 11450
rect 15750 11398 15762 11450
rect 15814 11398 18606 11450
rect 18658 11398 18670 11450
rect 18722 11398 18734 11450
rect 18786 11398 18798 11450
rect 18850 11398 18862 11450
rect 18914 11398 18920 11450
rect 184 11376 18920 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2041 11339 2099 11345
rect 2041 11336 2053 11339
rect 2004 11308 2053 11336
rect 2004 11296 2010 11308
rect 2041 11305 2053 11308
rect 2087 11305 2099 11339
rect 8202 11336 8208 11348
rect 8163 11308 8208 11336
rect 2041 11299 2099 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 9180 11308 9229 11336
rect 9180 11296 9186 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 9324 11308 10640 11336
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11268 1731 11271
rect 2130 11268 2136 11280
rect 1719 11240 2136 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 1964 11212 1992 11240
rect 2130 11228 2136 11240
rect 2188 11228 2194 11280
rect 2958 11228 2964 11280
rect 3016 11268 3022 11280
rect 3016 11240 3082 11268
rect 3016 11228 3022 11240
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 5776 11240 5934 11268
rect 5776 11228 5782 11240
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 9324 11268 9352 11308
rect 8628 11240 9352 11268
rect 10612 11268 10640 11308
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 11747 11339 11805 11345
rect 11747 11336 11759 11339
rect 11572 11308 11759 11336
rect 11572 11296 11578 11308
rect 11747 11305 11759 11308
rect 11793 11305 11805 11339
rect 11747 11299 11805 11305
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 13872 11308 14749 11336
rect 13872 11296 13878 11308
rect 14737 11305 14749 11308
rect 14783 11336 14795 11339
rect 14918 11336 14924 11348
rect 14783 11308 14924 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16022 11336 16028 11348
rect 15983 11308 16028 11336
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16448 11308 17141 11336
rect 16448 11296 16454 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 18230 11336 18236 11348
rect 18191 11308 18236 11336
rect 17129 11299 17187 11305
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 10612 11240 10718 11268
rect 8628 11228 8634 11240
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 16408 11268 16436 11296
rect 15252 11240 16436 11268
rect 15252 11228 15258 11240
rect 1946 11160 1952 11212
rect 2004 11160 2010 11212
rect 9766 11200 9772 11212
rect 8680 11172 9772 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 2222 11132 2228 11144
rect 1535 11104 2228 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5442 11132 5448 11144
rect 5215 11104 5304 11132
rect 5403 11104 5448 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2777 11067 2835 11073
rect 2777 11064 2789 11067
rect 2188 11036 2789 11064
rect 2188 11024 2194 11036
rect 2777 11033 2789 11036
rect 2823 11033 2835 11067
rect 2777 11027 2835 11033
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 4154 10996 4160 11008
rect 3660 10968 4160 10996
rect 3660 10956 3666 10968
rect 4154 10956 4160 10968
rect 4212 10996 4218 11008
rect 4540 10996 4568 11095
rect 4212 10968 4568 10996
rect 5276 10996 5304 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 8680 11141 8708 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10284 11172 10333 11200
rect 10284 11160 10290 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 15010 11200 15016 11212
rect 14971 11172 15016 11200
rect 10321 11163 10379 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15580 11209 15608 11240
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 16942 11200 16948 11212
rect 16439 11172 16948 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 10594 11132 10600 11144
rect 8803 11104 10600 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 14734 11132 14740 11144
rect 14695 11104 14740 11132
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 15764 11132 15792 11163
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11200 18015 11203
rect 18414 11200 18420 11212
rect 18003 11172 18420 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 16482 11132 16488 11144
rect 14884 11104 15792 11132
rect 16443 11104 16488 11132
rect 14884 11092 14890 11104
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 14918 11064 14924 11076
rect 14879 11036 14924 11064
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 15749 11067 15807 11073
rect 15749 11033 15761 11067
rect 15795 11064 15807 11067
rect 16592 11064 16620 11095
rect 15795 11036 16620 11064
rect 15795 11033 15807 11036
rect 15749 11027 15807 11033
rect 6546 10996 6552 11008
rect 5276 10968 6552 10996
rect 4212 10956 4218 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 17494 10996 17500 11008
rect 6972 10968 7017 10996
rect 17455 10968 17500 10996
rect 6972 10956 6978 10968
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 184 10906 18860 10928
rect 184 10854 1556 10906
rect 1608 10854 1620 10906
rect 1672 10854 1684 10906
rect 1736 10854 1748 10906
rect 1800 10854 1812 10906
rect 1864 10854 4656 10906
rect 4708 10854 4720 10906
rect 4772 10854 4784 10906
rect 4836 10854 4848 10906
rect 4900 10854 4912 10906
rect 4964 10854 7756 10906
rect 7808 10854 7820 10906
rect 7872 10854 7884 10906
rect 7936 10854 7948 10906
rect 8000 10854 8012 10906
rect 8064 10854 10856 10906
rect 10908 10854 10920 10906
rect 10972 10854 10984 10906
rect 11036 10854 11048 10906
rect 11100 10854 11112 10906
rect 11164 10854 13956 10906
rect 14008 10854 14020 10906
rect 14072 10854 14084 10906
rect 14136 10854 14148 10906
rect 14200 10854 14212 10906
rect 14264 10854 17056 10906
rect 17108 10854 17120 10906
rect 17172 10854 17184 10906
rect 17236 10854 17248 10906
rect 17300 10854 17312 10906
rect 17364 10854 18860 10906
rect 184 10832 18860 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1857 10795 1915 10801
rect 1857 10792 1869 10795
rect 1452 10764 1869 10792
rect 1452 10752 1458 10764
rect 1857 10761 1869 10764
rect 1903 10761 1915 10795
rect 10594 10792 10600 10804
rect 10555 10764 10600 10792
rect 1857 10755 1915 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 16172 10764 16313 10792
rect 16172 10752 16178 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 7607 10696 8248 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2924 10628 3341 10656
rect 2924 10616 2930 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7190 10656 7196 10668
rect 7055 10628 7196 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 8220 10665 8248 10696
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 8205 10619 8263 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10656 13234 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13228 10628 13553 10656
rect 13228 10616 13234 10628
rect 13541 10625 13553 10628
rect 13587 10656 13599 10659
rect 16482 10656 16488 10668
rect 13587 10628 16488 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 3602 10588 3608 10600
rect 3563 10560 3608 10588
rect 3602 10548 3608 10560
rect 3660 10588 3666 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3660 10560 3985 10588
rect 3660 10548 3666 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 3973 10551 4031 10557
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 6604 10560 7113 10588
rect 6604 10548 6610 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7340 10560 7941 10588
rect 7340 10548 7346 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 10686 10588 10692 10600
rect 10643 10560 10692 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 11422 10588 11428 10600
rect 10827 10560 11428 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 16316 10597 16344 10628
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10557 16359 10591
rect 17402 10588 17408 10600
rect 17363 10560 17408 10588
rect 16301 10551 16359 10557
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 17494 10548 17500 10600
rect 17552 10588 17558 10600
rect 17552 10560 17645 10588
rect 17552 10548 17558 10560
rect 4240 10523 4298 10529
rect 2898 10492 3004 10520
rect 2976 10464 3004 10492
rect 4240 10489 4252 10523
rect 4286 10520 4298 10523
rect 5902 10520 5908 10532
rect 4286 10492 5908 10520
rect 4286 10489 4298 10492
rect 4240 10483 4298 10489
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 8110 10520 8116 10532
rect 8071 10492 8116 10520
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 12158 10480 12164 10532
rect 12216 10480 12222 10532
rect 15286 10520 15292 10532
rect 15247 10492 15292 10520
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 17512 10520 17540 10548
rect 17144 10492 17540 10520
rect 17144 10464 17172 10492
rect 2958 10412 2964 10464
rect 3016 10412 3022 10464
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 5040 10424 5365 10452
rect 5040 10412 5046 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 7156 10424 7205 10452
rect 7156 10412 7162 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 7193 10415 7251 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 184 10362 18920 10384
rect 184 10310 3106 10362
rect 3158 10310 3170 10362
rect 3222 10310 3234 10362
rect 3286 10310 3298 10362
rect 3350 10310 3362 10362
rect 3414 10310 6206 10362
rect 6258 10310 6270 10362
rect 6322 10310 6334 10362
rect 6386 10310 6398 10362
rect 6450 10310 6462 10362
rect 6514 10310 9306 10362
rect 9358 10310 9370 10362
rect 9422 10310 9434 10362
rect 9486 10310 9498 10362
rect 9550 10310 9562 10362
rect 9614 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 12534 10362
rect 12586 10310 12598 10362
rect 12650 10310 12662 10362
rect 12714 10310 15506 10362
rect 15558 10310 15570 10362
rect 15622 10310 15634 10362
rect 15686 10310 15698 10362
rect 15750 10310 15762 10362
rect 15814 10310 18606 10362
rect 18658 10310 18670 10362
rect 18722 10310 18734 10362
rect 18786 10310 18798 10362
rect 18850 10310 18862 10362
rect 18914 10310 18920 10362
rect 184 10288 18920 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2130 10248 2136 10260
rect 2087 10220 2136 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3602 10248 3608 10260
rect 3283 10220 3608 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 2424 10180 2452 10211
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5500 10220 5733 10248
rect 5500 10208 5506 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 9088 10220 9413 10248
rect 9088 10208 9094 10220
rect 9401 10217 9413 10220
rect 9447 10248 9459 10251
rect 10778 10248 10784 10260
rect 9447 10220 10784 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 15068 10220 17356 10248
rect 15068 10208 15074 10220
rect 4246 10180 4252 10192
rect 2424 10152 4252 10180
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 4525 10183 4583 10189
rect 4525 10149 4537 10183
rect 4571 10180 4583 10183
rect 7006 10180 7012 10192
rect 4571 10152 7012 10180
rect 4571 10149 4583 10152
rect 4525 10143 4583 10149
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 16022 10140 16028 10192
rect 16080 10140 16086 10192
rect 17328 10180 17356 10220
rect 17862 10180 17868 10192
rect 17328 10152 17868 10180
rect 569 10115 627 10121
rect 569 10081 581 10115
rect 615 10112 627 10115
rect 934 10112 940 10124
rect 615 10084 940 10112
rect 615 10081 627 10084
rect 569 10075 627 10081
rect 934 10072 940 10084
rect 992 10112 998 10124
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 992 10084 1041 10112
rect 992 10072 998 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 2464 10084 5181 10112
rect 2464 10072 2470 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5169 10075 5227 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2314 10044 2320 10056
rect 1995 10016 2320 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 1872 9976 1900 10007
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 5184 10044 5212 10075
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 6181 10115 6239 10121
rect 5592 10084 5637 10112
rect 5592 10072 5598 10084
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6914 10112 6920 10124
rect 6227 10084 6920 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 9585 10115 9643 10121
rect 7239 10084 9444 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5184 10016 6009 10044
rect 5997 10013 6009 10016
rect 6043 10044 6055 10047
rect 7650 10044 7656 10056
rect 6043 10016 7656 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 9416 10044 9444 10084
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 11238 10112 11244 10124
rect 9631 10084 11244 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 14458 10112 14464 10124
rect 13955 10084 14464 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 17328 10121 17356 10152
rect 17862 10140 17868 10152
rect 17920 10140 17926 10192
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 18263 10115 18321 10121
rect 18263 10112 18275 10115
rect 17460 10084 18275 10112
rect 17460 10072 17466 10084
rect 18263 10081 18275 10084
rect 18309 10081 18321 10115
rect 18263 10075 18321 10081
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18472 10084 18565 10112
rect 18472 10072 18478 10084
rect 9858 10044 9864 10056
rect 9416 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 13228 10016 14749 10044
rect 13228 10004 13234 10016
rect 14737 10013 14749 10016
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10044 15163 10047
rect 15378 10044 15384 10056
rect 15151 10016 15384 10044
rect 15151 10013 15163 10016
rect 15105 10007 15163 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 17126 10004 17132 10056
rect 17184 10044 17190 10056
rect 17589 10047 17647 10053
rect 17589 10044 17601 10047
rect 17184 10016 17601 10044
rect 17184 10004 17190 10016
rect 17589 10013 17601 10016
rect 17635 10044 17647 10047
rect 17954 10044 17960 10056
rect 17635 10016 17960 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17954 10004 17960 10016
rect 18012 10044 18018 10056
rect 18432 10044 18460 10072
rect 18012 10016 18460 10044
rect 18012 10004 18018 10016
rect 2222 9976 2228 9988
rect 1872 9948 2228 9976
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 7282 9976 7288 9988
rect 7055 9948 7288 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 13262 9936 13268 9988
rect 13320 9976 13326 9988
rect 13538 9976 13544 9988
rect 13320 9948 13544 9976
rect 13320 9936 13326 9948
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 17862 9936 17868 9988
rect 17920 9976 17926 9988
rect 18049 9979 18107 9985
rect 18049 9976 18061 9979
rect 17920 9948 18061 9976
rect 17920 9936 17926 9948
rect 18049 9945 18061 9948
rect 18095 9945 18107 9979
rect 18049 9939 18107 9945
rect 753 9911 811 9917
rect 753 9877 765 9911
rect 799 9908 811 9911
rect 4338 9908 4344 9920
rect 799 9880 4344 9908
rect 799 9877 811 9880
rect 753 9871 811 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4430 9868 4436 9920
rect 4488 9908 4494 9920
rect 5261 9911 5319 9917
rect 5261 9908 5273 9911
rect 4488 9880 5273 9908
rect 4488 9868 4494 9880
rect 5261 9877 5273 9880
rect 5307 9877 5319 9911
rect 5261 9871 5319 9877
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 15838 9908 15844 9920
rect 15620 9880 15844 9908
rect 15620 9868 15626 9880
rect 15838 9868 15844 9880
rect 15896 9908 15902 9920
rect 16574 9917 16580 9920
rect 16531 9911 16580 9917
rect 16531 9908 16543 9911
rect 15896 9880 16543 9908
rect 15896 9868 15902 9880
rect 16531 9877 16543 9880
rect 16577 9877 16580 9911
rect 16531 9871 16580 9877
rect 16574 9868 16580 9871
rect 16632 9868 16638 9920
rect 184 9818 18860 9840
rect 184 9766 1556 9818
rect 1608 9766 1620 9818
rect 1672 9766 1684 9818
rect 1736 9766 1748 9818
rect 1800 9766 1812 9818
rect 1864 9766 4656 9818
rect 4708 9766 4720 9818
rect 4772 9766 4784 9818
rect 4836 9766 4848 9818
rect 4900 9766 4912 9818
rect 4964 9766 7756 9818
rect 7808 9766 7820 9818
rect 7872 9766 7884 9818
rect 7936 9766 7948 9818
rect 8000 9766 8012 9818
rect 8064 9766 10856 9818
rect 10908 9766 10920 9818
rect 10972 9766 10984 9818
rect 11036 9766 11048 9818
rect 11100 9766 11112 9818
rect 11164 9766 13956 9818
rect 14008 9766 14020 9818
rect 14072 9766 14084 9818
rect 14136 9766 14148 9818
rect 14200 9766 14212 9818
rect 14264 9766 17056 9818
rect 17108 9766 17120 9818
rect 17172 9766 17184 9818
rect 17236 9766 17248 9818
rect 17300 9766 17312 9818
rect 17364 9766 18860 9818
rect 184 9744 18860 9766
rect 10686 9664 10692 9716
rect 10744 9664 10750 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 17313 9707 17371 9713
rect 14516 9676 15148 9704
rect 14516 9664 14522 9676
rect 845 9639 903 9645
rect 845 9605 857 9639
rect 891 9636 903 9639
rect 1394 9636 1400 9648
rect 891 9608 1400 9636
rect 891 9605 903 9608
rect 845 9599 903 9605
rect 1394 9596 1400 9608
rect 1452 9596 1458 9648
rect 2222 9636 2228 9648
rect 1872 9608 2228 9636
rect 753 9571 811 9577
rect 753 9537 765 9571
rect 799 9568 811 9571
rect 1762 9568 1768 9580
rect 799 9540 1768 9568
rect 799 9537 811 9540
rect 753 9531 811 9537
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 1872 9577 1900 9608
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2866 9636 2872 9648
rect 2455 9608 2872 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 10704 9636 10732 9664
rect 11606 9636 11612 9648
rect 10704 9608 11612 9636
rect 11606 9596 11612 9608
rect 11664 9596 11670 9648
rect 13909 9639 13967 9645
rect 13909 9605 13921 9639
rect 13955 9636 13967 9639
rect 14734 9636 14740 9648
rect 13955 9608 14740 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2096 9540 2789 9568
rect 2096 9528 2102 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 8938 9568 8944 9580
rect 6963 9540 8944 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 11940 9540 12909 9568
rect 11940 9528 11946 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 15010 9568 15016 9580
rect 14047 9540 15016 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 15120 9568 15148 9676
rect 17313 9673 17325 9707
rect 17359 9704 17371 9707
rect 17402 9704 17408 9716
rect 17359 9676 17408 9704
rect 17359 9673 17371 9676
rect 17313 9667 17371 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 15252 9608 15301 9636
rect 15252 9596 15258 9608
rect 15289 9605 15301 9608
rect 15335 9605 15347 9639
rect 15289 9599 15347 9605
rect 15120 9540 16068 9568
rect 1029 9503 1087 9509
rect 1029 9469 1041 9503
rect 1075 9500 1087 9503
rect 2130 9500 2136 9512
rect 1075 9472 2136 9500
rect 1075 9469 1087 9472
rect 1029 9463 1087 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4479 9472 4905 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4893 9469 4905 9472
rect 4939 9500 4951 9503
rect 4982 9500 4988 9512
rect 4939 9472 4988 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 1394 9392 1400 9444
rect 1452 9432 1458 9444
rect 2041 9435 2099 9441
rect 2041 9432 2053 9435
rect 1452 9404 2053 9432
rect 1452 9392 1458 9404
rect 2041 9401 2053 9404
rect 2087 9401 2099 9435
rect 2041 9395 2099 9401
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 4264 9432 4292 9463
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5092 9432 5120 9463
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6546 9500 6552 9512
rect 5776 9472 6552 9500
rect 5776 9460 5782 9472
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14366 9500 14372 9512
rect 13771 9472 14372 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 15212 9500 15240 9540
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 15212 9472 15301 9500
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15562 9500 15568 9512
rect 15523 9472 15568 9500
rect 15289 9463 15347 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16040 9500 16068 9540
rect 17310 9500 17316 9512
rect 16040 9472 17316 9500
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17770 9500 17776 9512
rect 17731 9472 17776 9500
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 17920 9472 17965 9500
rect 17920 9460 17926 9472
rect 6638 9432 6644 9444
rect 2832 9404 6644 9432
rect 2832 9392 2838 9404
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 8662 9432 8668 9444
rect 7958 9404 8668 9432
rect 8662 9392 8668 9404
rect 8720 9432 8726 9444
rect 10505 9435 10563 9441
rect 8720 9404 9338 9432
rect 8720 9392 8726 9404
rect 10505 9401 10517 9435
rect 10551 9401 10563 9435
rect 10505 9395 10563 9401
rect 1026 9324 1032 9376
rect 1084 9364 1090 9376
rect 1213 9367 1271 9373
rect 1213 9364 1225 9367
rect 1084 9336 1225 9364
rect 1084 9324 1090 9336
rect 1213 9333 1225 9336
rect 1259 9333 1271 9367
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1213 9327 1271 9333
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 8386 9373 8392 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4764 9336 4997 9364
rect 4764 9324 4770 9336
rect 4985 9333 4997 9336
rect 5031 9333 5043 9367
rect 4985 9327 5043 9333
rect 8343 9367 8392 9373
rect 8343 9333 8355 9367
rect 8389 9333 8392 9367
rect 8343 9327 8392 9333
rect 8386 9324 8392 9327
rect 8444 9324 8450 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10520 9364 10548 9395
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 16206 9441 16212 9444
rect 12621 9435 12679 9441
rect 10836 9404 11454 9432
rect 10836 9392 10842 9404
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 12667 9404 16160 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10520 9336 11161 9364
rect 11149 9333 11161 9336
rect 11195 9333 11207 9367
rect 11149 9327 11207 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 11664 9336 13553 9364
rect 11664 9324 11670 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 14366 9364 14372 9376
rect 14327 9336 14372 9364
rect 13541 9327 13599 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 15068 9336 15485 9364
rect 15068 9324 15074 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 16132 9364 16160 9404
rect 16200 9395 16212 9441
rect 16264 9432 16270 9444
rect 17586 9432 17592 9444
rect 16264 9404 16300 9432
rect 17547 9404 17592 9432
rect 16206 9392 16212 9395
rect 16264 9392 16270 9404
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 16850 9364 16856 9376
rect 16132 9336 16856 9364
rect 15473 9327 15531 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 17460 9336 17693 9364
rect 17460 9324 17466 9336
rect 17681 9333 17693 9336
rect 17727 9333 17739 9367
rect 17681 9327 17739 9333
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18012 9336 18337 9364
rect 18012 9324 18018 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 184 9274 18920 9296
rect 184 9222 3106 9274
rect 3158 9222 3170 9274
rect 3222 9222 3234 9274
rect 3286 9222 3298 9274
rect 3350 9222 3362 9274
rect 3414 9222 6206 9274
rect 6258 9222 6270 9274
rect 6322 9222 6334 9274
rect 6386 9222 6398 9274
rect 6450 9222 6462 9274
rect 6514 9222 9306 9274
rect 9358 9222 9370 9274
rect 9422 9222 9434 9274
rect 9486 9222 9498 9274
rect 9550 9222 9562 9274
rect 9614 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 12534 9274
rect 12586 9222 12598 9274
rect 12650 9222 12662 9274
rect 12714 9222 15506 9274
rect 15558 9222 15570 9274
rect 15622 9222 15634 9274
rect 15686 9222 15698 9274
rect 15750 9222 15762 9274
rect 15814 9222 18606 9274
rect 18658 9222 18670 9274
rect 18722 9222 18734 9274
rect 18786 9222 18798 9274
rect 18850 9222 18862 9274
rect 18914 9222 18920 9274
rect 184 9200 18920 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2924 9132 2973 9160
rect 2924 9120 2930 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 5442 9160 5448 9172
rect 4479 9132 5448 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5626 9160 5632 9172
rect 5587 9132 5632 9160
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 5997 9163 6055 9169
rect 5997 9129 6009 9163
rect 6043 9160 6055 9163
rect 7190 9160 7196 9172
rect 6043 9132 7196 9160
rect 6043 9129 6055 9132
rect 5997 9123 6055 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 11330 9160 11336 9172
rect 8067 9132 11336 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 11480 9132 12817 9160
rect 11480 9120 11486 9132
rect 12805 9129 12817 9132
rect 12851 9129 12863 9163
rect 17310 9160 17316 9172
rect 17271 9132 17316 9160
rect 12805 9123 12863 9129
rect 17310 9120 17316 9132
rect 17368 9160 17374 9172
rect 17494 9160 17500 9172
rect 17368 9132 17500 9160
rect 17368 9120 17374 9132
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 2130 9092 2136 9104
rect 1872 9064 2136 9092
rect 1872 9033 1900 9064
rect 2130 9052 2136 9064
rect 2188 9052 2194 9104
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 3237 9095 3295 9101
rect 3237 9092 3249 9095
rect 2832 9064 3249 9092
rect 2832 9052 2838 9064
rect 3237 9061 3249 9064
rect 3283 9061 3295 9095
rect 5644 9092 5672 9120
rect 9030 9092 9036 9104
rect 5644 9064 6132 9092
rect 3237 9055 3295 9061
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 8993 1915 9027
rect 2038 9024 2044 9036
rect 1999 8996 2044 9024
rect 1857 8987 1915 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 4154 9024 4160 9036
rect 3007 8996 4160 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5902 9024 5908 9036
rect 4764 8996 4809 9024
rect 5863 8996 5908 9024
rect 4764 8984 4770 8996
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6104 9033 6132 9064
rect 6840 9064 9036 9092
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6840 9033 6868 9064
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 10778 9052 10784 9104
rect 10836 9052 10842 9104
rect 12986 9092 12992 9104
rect 12820 9064 12992 9092
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6696 8996 6837 9024
rect 6696 8984 6702 8996
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8110 9024 8116 9036
rect 8067 8996 8116 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5920 8956 5948 8984
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 5920 8928 6561 8956
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 7576 8956 7604 8987
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 9024 8631 9027
rect 8662 9024 8668 9036
rect 8619 8996 8668 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 8662 8984 8668 8996
rect 8720 9024 8726 9036
rect 8849 9027 8907 9033
rect 8849 9024 8861 9027
rect 8720 8996 8861 9024
rect 8720 8984 8726 8996
rect 8849 8993 8861 8996
rect 8895 8993 8907 9027
rect 8849 8987 8907 8993
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 11882 9024 11888 9036
rect 11747 8996 11888 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12820 9033 12848 9064
rect 12986 9052 12992 9064
rect 13044 9092 13050 9104
rect 14093 9095 14151 9101
rect 14093 9092 14105 9095
rect 13044 9064 14105 9092
rect 13044 9052 13050 9064
rect 14093 9061 14105 9064
rect 14139 9061 14151 9095
rect 14093 9055 14151 9061
rect 16485 9095 16543 9101
rect 16485 9061 16497 9095
rect 16531 9092 16543 9095
rect 18506 9092 18512 9104
rect 16531 9064 18512 9092
rect 16531 9061 16543 9064
rect 16485 9055 16543 9061
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 9024 12955 9027
rect 12943 8996 13860 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 8294 8956 8300 8968
rect 7576 8928 8300 8956
rect 6549 8919 6607 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9916 8928 9965 8956
rect 9916 8916 9922 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 13832 8965 13860 8996
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 14700 8996 17233 9024
rect 14700 8984 14706 8996
rect 17221 8993 17233 8996
rect 17267 8993 17279 9027
rect 17221 8987 17279 8993
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17736 8996 17877 9024
rect 17736 8984 17742 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11388 8928 11437 8956
rect 11388 8916 11394 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8956 13875 8959
rect 14826 8956 14832 8968
rect 13863 8928 14832 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 2038 8888 2044 8900
rect 1811 8860 2044 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 2038 8848 2044 8860
rect 2096 8848 2102 8900
rect 3053 8891 3111 8897
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3418 8888 3424 8900
rect 3099 8860 3424 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3418 8848 3424 8860
rect 3476 8888 3482 8900
rect 5810 8888 5816 8900
rect 3476 8860 5816 8888
rect 3476 8848 3482 8860
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 7699 8891 7757 8897
rect 7699 8888 7711 8891
rect 6052 8860 7711 8888
rect 6052 8848 6058 8860
rect 7699 8857 7711 8860
rect 7745 8857 7757 8891
rect 13096 8888 13124 8919
rect 14826 8916 14832 8928
rect 14884 8956 14890 8968
rect 16206 8956 16212 8968
rect 14884 8928 16212 8956
rect 14884 8916 14890 8928
rect 16206 8916 16212 8928
rect 16264 8956 16270 8968
rect 17954 8956 17960 8968
rect 16264 8928 17960 8956
rect 16264 8916 16270 8928
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 13449 8891 13507 8897
rect 13449 8888 13461 8891
rect 13096 8860 13461 8888
rect 7699 8851 7757 8857
rect 13449 8857 13461 8860
rect 13495 8888 13507 8891
rect 14366 8888 14372 8900
rect 13495 8860 14372 8888
rect 13495 8857 13507 8860
rect 13449 8851 13507 8857
rect 14366 8848 14372 8860
rect 14424 8888 14430 8900
rect 15562 8888 15568 8900
rect 14424 8860 15568 8888
rect 14424 8848 14430 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 8110 8820 8116 8832
rect 7883 8792 8116 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15286 8820 15292 8832
rect 15243 8792 15292 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 18156 8820 18184 8919
rect 18414 8820 18420 8832
rect 16632 8792 18420 8820
rect 16632 8780 16638 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 184 8730 18860 8752
rect 184 8678 1556 8730
rect 1608 8678 1620 8730
rect 1672 8678 1684 8730
rect 1736 8678 1748 8730
rect 1800 8678 1812 8730
rect 1864 8678 4656 8730
rect 4708 8678 4720 8730
rect 4772 8678 4784 8730
rect 4836 8678 4848 8730
rect 4900 8678 4912 8730
rect 4964 8678 7756 8730
rect 7808 8678 7820 8730
rect 7872 8678 7884 8730
rect 7936 8678 7948 8730
rect 8000 8678 8012 8730
rect 8064 8678 10856 8730
rect 10908 8678 10920 8730
rect 10972 8678 10984 8730
rect 11036 8678 11048 8730
rect 11100 8678 11112 8730
rect 11164 8678 13956 8730
rect 14008 8678 14020 8730
rect 14072 8678 14084 8730
rect 14136 8678 14148 8730
rect 14200 8678 14212 8730
rect 14264 8678 17056 8730
rect 17108 8678 17120 8730
rect 17172 8678 17184 8730
rect 17236 8678 17248 8730
rect 17300 8678 17312 8730
rect 17364 8678 18860 8730
rect 184 8656 18860 8678
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8294 8616 8300 8628
rect 8255 8588 8300 8616
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13044 8588 13553 8616
rect 13044 8576 13050 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 5868 8520 8984 8548
rect 5868 8508 5874 8520
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2682 8480 2688 8492
rect 1903 8452 2688 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 937 8415 995 8421
rect 937 8381 949 8415
rect 983 8412 995 8415
rect 1394 8412 1400 8424
rect 983 8384 1400 8412
rect 983 8381 995 8384
rect 937 8375 995 8381
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1780 8412 1808 8443
rect 2682 8440 2688 8452
rect 2740 8480 2746 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2740 8452 2973 8480
rect 2740 8440 2746 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 4154 8480 4160 8492
rect 3375 8452 4160 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 5166 8480 5172 8492
rect 4212 8452 5172 8480
rect 4212 8440 4218 8452
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 8956 8489 8984 8520
rect 8941 8483 8999 8489
rect 7484 8452 8156 8480
rect 2406 8412 2412 8424
rect 1780 8384 2412 8412
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3418 8412 3424 8424
rect 3379 8384 3424 8412
rect 3145 8375 3203 8381
rect 1118 8304 1124 8356
rect 1176 8344 1182 8356
rect 1949 8347 2007 8353
rect 1949 8344 1961 8347
rect 1176 8316 1961 8344
rect 1176 8304 1182 8316
rect 1949 8313 1961 8316
rect 1995 8313 2007 8347
rect 3160 8344 3188 8375
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 5718 8412 5724 8424
rect 5675 8384 5724 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7484 8421 7512 8452
rect 8128 8421 8156 8452
rect 8941 8449 8953 8483
rect 8987 8480 8999 8483
rect 10502 8480 10508 8492
rect 8987 8452 10508 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11882 8480 11888 8492
rect 10827 8452 11888 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 6972 8384 7481 8412
rect 6972 8372 6978 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 8294 8412 8300 8424
rect 8255 8384 8300 8412
rect 8113 8375 8171 8381
rect 3786 8344 3792 8356
rect 3160 8316 3792 8344
rect 1949 8307 2007 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 5258 8344 5264 8356
rect 5219 8316 5264 8344
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 7668 8344 7696 8375
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 10410 8412 10416 8424
rect 10371 8384 10416 8412
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8412 11667 8415
rect 12250 8412 12256 8424
rect 11655 8384 12256 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 12250 8372 12256 8384
rect 12308 8412 12314 8424
rect 13556 8412 13584 8579
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17644 8588 17785 8616
rect 17644 8576 17650 8588
rect 17773 8585 17785 8588
rect 17819 8585 17831 8619
rect 17773 8579 17831 8585
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 18506 8616 18512 8628
rect 18463 8588 18512 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13872 8452 13921 8480
rect 13872 8440 13878 8452
rect 13909 8449 13921 8452
rect 13955 8480 13967 8483
rect 14550 8480 14556 8492
rect 13955 8452 14556 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 15194 8480 15200 8492
rect 15155 8452 15200 8480
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 15988 8452 16405 8480
rect 15988 8440 15994 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 16393 8443 16451 8449
rect 14458 8412 14464 8424
rect 12308 8384 12388 8412
rect 13556 8384 14464 8412
rect 12308 8372 12314 8384
rect 8312 8344 8340 8372
rect 7668 8316 8340 8344
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 8720 8316 9430 8344
rect 8720 8304 8726 8316
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 10928 8316 11345 8344
rect 10928 8304 10934 8316
rect 11333 8313 11345 8316
rect 11379 8344 11391 8347
rect 12158 8344 12164 8356
rect 11379 8316 12164 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 12360 8344 12388 8384
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8412 14795 8415
rect 14826 8412 14832 8424
rect 14783 8384 14832 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 14936 8344 14964 8375
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15068 8384 15393 8412
rect 15068 8372 15074 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15838 8412 15844 8424
rect 15519 8384 15844 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16408 8412 16436 8443
rect 16482 8412 16488 8424
rect 16408 8384 16488 8412
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 16666 8421 16672 8424
rect 16660 8412 16672 8421
rect 16627 8384 16672 8412
rect 16660 8375 16672 8384
rect 16666 8372 16672 8375
rect 16724 8372 16730 8424
rect 15562 8344 15568 8356
rect 12360 8316 13768 8344
rect 14936 8316 15568 8344
rect 845 8279 903 8285
rect 845 8245 857 8279
rect 891 8276 903 8279
rect 1210 8276 1216 8288
rect 891 8248 1216 8276
rect 891 8245 903 8248
rect 845 8239 903 8245
rect 1210 8236 1216 8248
rect 1268 8236 1274 8288
rect 13740 8276 13768 8316
rect 15562 8304 15568 8316
rect 15620 8344 15626 8356
rect 15620 8316 16068 8344
rect 15620 8304 15626 8316
rect 14274 8276 14280 8288
rect 13740 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 16040 8285 16068 8316
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 16390 8276 16396 8288
rect 16071 8248 16396 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 184 8186 18920 8208
rect 184 8134 3106 8186
rect 3158 8134 3170 8186
rect 3222 8134 3234 8186
rect 3286 8134 3298 8186
rect 3350 8134 3362 8186
rect 3414 8134 6206 8186
rect 6258 8134 6270 8186
rect 6322 8134 6334 8186
rect 6386 8134 6398 8186
rect 6450 8134 6462 8186
rect 6514 8134 9306 8186
rect 9358 8134 9370 8186
rect 9422 8134 9434 8186
rect 9486 8134 9498 8186
rect 9550 8134 9562 8186
rect 9614 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 12534 8186
rect 12586 8134 12598 8186
rect 12650 8134 12662 8186
rect 12714 8134 15506 8186
rect 15558 8134 15570 8186
rect 15622 8134 15634 8186
rect 15686 8134 15698 8186
rect 15750 8134 15762 8186
rect 15814 8134 18606 8186
rect 18658 8134 18670 8186
rect 18722 8134 18734 8186
rect 18786 8134 18798 8186
rect 18850 8134 18862 8186
rect 18914 8134 18920 8186
rect 184 8112 18920 8134
rect 1210 8072 1216 8084
rect 1171 8044 1216 8072
rect 1210 8032 1216 8044
rect 1268 8032 1274 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7616 8044 7665 8072
rect 7616 8032 7622 8044
rect 7653 8041 7665 8044
rect 7699 8072 7711 8075
rect 8662 8072 8668 8084
rect 7699 8044 8668 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 8662 8032 8668 8044
rect 8720 8072 8726 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8720 8044 8769 8072
rect 8720 8032 8726 8044
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 10183 8075 10241 8081
rect 10183 8041 10195 8075
rect 10229 8072 10241 8075
rect 10410 8072 10416 8084
rect 10229 8044 10416 8072
rect 10229 8041 10241 8044
rect 10183 8035 10241 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 14737 8075 14795 8081
rect 14737 8072 14749 8075
rect 14700 8044 14749 8072
rect 14700 8032 14706 8044
rect 14737 8041 14749 8044
rect 14783 8041 14795 8075
rect 18322 8072 18328 8084
rect 14737 8035 14795 8041
rect 14936 8044 18328 8072
rect 845 8007 903 8013
rect 845 7973 857 8007
rect 891 8004 903 8007
rect 1118 8004 1124 8016
rect 891 7976 1124 8004
rect 891 7973 903 7976
rect 845 7967 903 7973
rect 1118 7964 1124 7976
rect 1176 7964 1182 8016
rect 6546 7964 6552 8016
rect 6604 7964 6610 8016
rect 10870 7964 10876 8016
rect 10928 7964 10934 8016
rect 14936 8004 14964 8044
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 15930 8004 15936 8016
rect 12406 7976 14964 8004
rect 15778 7976 15936 8004
rect 1026 7936 1032 7948
rect 987 7908 1032 7936
rect 1026 7896 1032 7908
rect 1084 7896 1090 7948
rect 1305 7939 1363 7945
rect 1305 7905 1317 7939
rect 1351 7936 1363 7939
rect 2038 7936 2044 7948
rect 1351 7908 2044 7936
rect 1351 7905 1363 7908
rect 1305 7899 1363 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5258 7936 5264 7948
rect 5215 7908 5264 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11940 7908 11989 7936
rect 11940 7896 11946 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 12406 7936 12434 7976
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 17957 8007 18015 8013
rect 17957 8004 17969 8007
rect 17420 7976 17969 8004
rect 11977 7899 12035 7905
rect 12360 7908 12434 7936
rect 12713 7939 12771 7945
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5040 7840 5549 7868
rect 5040 7828 5046 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 6914 7828 6920 7880
rect 6972 7877 6978 7880
rect 6972 7871 7021 7877
rect 6972 7837 6975 7871
rect 7009 7837 7021 7871
rect 6972 7831 7021 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 12360 7868 12388 7908
rect 12713 7905 12725 7939
rect 12759 7936 12771 7939
rect 12986 7936 12992 7948
rect 12759 7908 12992 7936
rect 12759 7905 12771 7908
rect 12713 7899 12771 7905
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 17310 7936 17316 7948
rect 16540 7908 16585 7936
rect 17271 7908 17316 7936
rect 16540 7896 16546 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 17420 7945 17448 7976
rect 17957 7973 17969 7976
rect 18003 7973 18015 8007
rect 17957 7967 18015 7973
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17552 7908 17693 7936
rect 17552 7896 17558 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 18230 7936 18236 7948
rect 18191 7908 18236 7936
rect 17681 7899 17739 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 11655 7840 12388 7868
rect 12437 7871 12495 7877
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12802 7868 12808 7880
rect 12483 7840 12808 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 6972 7828 6978 7831
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 16255 7840 17141 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17129 7831 17187 7837
rect 17604 7840 17969 7868
rect 12621 7803 12679 7809
rect 12621 7769 12633 7803
rect 12667 7800 12679 7803
rect 13538 7800 13544 7812
rect 12667 7772 13544 7800
rect 12667 7769 12679 7772
rect 12621 7763 12679 7769
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 14369 7803 14427 7809
rect 14369 7769 14381 7803
rect 14415 7800 14427 7803
rect 14826 7800 14832 7812
rect 14415 7772 14832 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 14826 7760 14832 7772
rect 14884 7760 14890 7812
rect 12526 7732 12532 7744
rect 12487 7704 12532 7732
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 17604 7741 17632 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 14608 7704 17601 7732
rect 14608 7692 14614 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 18196 7704 18241 7732
rect 18196 7692 18202 7704
rect 184 7642 18860 7664
rect 184 7590 1556 7642
rect 1608 7590 1620 7642
rect 1672 7590 1684 7642
rect 1736 7590 1748 7642
rect 1800 7590 1812 7642
rect 1864 7590 4656 7642
rect 4708 7590 4720 7642
rect 4772 7590 4784 7642
rect 4836 7590 4848 7642
rect 4900 7590 4912 7642
rect 4964 7590 7756 7642
rect 7808 7590 7820 7642
rect 7872 7590 7884 7642
rect 7936 7590 7948 7642
rect 8000 7590 8012 7642
rect 8064 7590 10856 7642
rect 10908 7590 10920 7642
rect 10972 7590 10984 7642
rect 11036 7590 11048 7642
rect 11100 7590 11112 7642
rect 11164 7590 13956 7642
rect 14008 7590 14020 7642
rect 14072 7590 14084 7642
rect 14136 7590 14148 7642
rect 14200 7590 14212 7642
rect 14264 7590 17056 7642
rect 17108 7590 17120 7642
rect 17172 7590 17184 7642
rect 17236 7590 17248 7642
rect 17300 7590 17312 7642
rect 17364 7590 18860 7642
rect 184 7568 18860 7590
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 5074 7528 5080 7540
rect 4488 7500 5080 7528
rect 4488 7488 4494 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 5408 7500 5457 7528
rect 5408 7488 5414 7500
rect 5445 7497 5457 7500
rect 5491 7528 5503 7531
rect 5626 7528 5632 7540
rect 5491 7500 5632 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 5626 7488 5632 7500
rect 5684 7528 5690 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5684 7500 5825 7528
rect 5684 7488 5690 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 7558 7528 7564 7540
rect 7519 7500 7564 7528
rect 5813 7491 5871 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 8938 7528 8944 7540
rect 8899 7500 8944 7528
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 13798 7531 13856 7537
rect 13798 7528 13810 7531
rect 12584 7500 13810 7528
rect 12584 7488 12590 7500
rect 13798 7497 13810 7500
rect 13844 7497 13856 7531
rect 16482 7528 16488 7540
rect 13798 7491 13856 7497
rect 16132 7500 16488 7528
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7429 9367 7463
rect 11422 7460 11428 7472
rect 11335 7432 11428 7460
rect 9309 7423 9367 7429
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2866 7392 2872 7404
rect 1903 7364 2872 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5902 7392 5908 7404
rect 5583 7364 5908 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9324 7392 9352 7423
rect 11422 7420 11428 7432
rect 11480 7460 11486 7472
rect 11882 7460 11888 7472
rect 11480 7432 11888 7460
rect 11480 7420 11486 7432
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 16132 7404 16160 7500
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 16908 7500 17785 7528
rect 16908 7488 16914 7500
rect 17773 7497 17785 7500
rect 17819 7497 17831 7531
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 17773 7491 17831 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 9079 7364 9352 7392
rect 13541 7395 13599 7401
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 16114 7392 16120 7404
rect 13587 7364 16120 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 5258 7324 5264 7336
rect 5219 7296 5264 7324
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8352 7296 8769 7324
rect 8352 7284 8358 7296
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 2130 7256 2136 7268
rect 2091 7228 2136 7256
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3358 7228 4077 7256
rect 4065 7225 4077 7228
rect 4111 7256 4123 7259
rect 4154 7256 4160 7268
rect 4111 7228 4160 7256
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 4154 7216 4160 7228
rect 4212 7256 4218 7268
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4212 7228 4813 7256
rect 4212 7216 4218 7228
rect 4801 7225 4813 7228
rect 4847 7256 4859 7259
rect 5902 7256 5908 7268
rect 4847 7228 5908 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5902 7216 5908 7228
rect 5960 7256 5966 7268
rect 6546 7256 6552 7268
rect 5960 7228 6552 7256
rect 5960 7216 5966 7228
rect 6546 7216 6552 7228
rect 6604 7256 6610 7268
rect 7558 7256 7564 7268
rect 6604 7228 7564 7256
rect 6604 7216 6610 7228
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 8772 7256 8800 7287
rect 8846 7284 8852 7336
rect 8904 7324 8910 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 8904 7296 9505 7324
rect 8904 7284 8910 7296
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7293 9643 7327
rect 11238 7324 11244 7336
rect 11199 7296 11244 7324
rect 9585 7287 9643 7293
rect 8772 7228 9168 7256
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 9140 7188 9168 7228
rect 9214 7216 9220 7268
rect 9272 7256 9278 7268
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 9272 7228 9321 7256
rect 9272 7216 9278 7228
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 9309 7219 9367 7225
rect 9600 7188 9628 7287
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 14274 7216 14280 7268
rect 14332 7216 14338 7268
rect 16390 7265 16396 7268
rect 15565 7259 15623 7265
rect 15565 7225 15577 7259
rect 15611 7225 15623 7259
rect 16384 7256 16396 7265
rect 16351 7228 16396 7256
rect 15565 7219 15623 7225
rect 16384 7219 16396 7228
rect 9140 7160 9628 7188
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 15580 7188 15608 7219
rect 16390 7216 16396 7219
rect 16448 7216 16454 7268
rect 17494 7188 17500 7200
rect 14608 7160 15608 7188
rect 17455 7160 17500 7188
rect 14608 7148 14614 7160
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 184 7098 18920 7120
rect 184 7046 3106 7098
rect 3158 7046 3170 7098
rect 3222 7046 3234 7098
rect 3286 7046 3298 7098
rect 3350 7046 3362 7098
rect 3414 7046 6206 7098
rect 6258 7046 6270 7098
rect 6322 7046 6334 7098
rect 6386 7046 6398 7098
rect 6450 7046 6462 7098
rect 6514 7046 9306 7098
rect 9358 7046 9370 7098
rect 9422 7046 9434 7098
rect 9486 7046 9498 7098
rect 9550 7046 9562 7098
rect 9614 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 12534 7098
rect 12586 7046 12598 7098
rect 12650 7046 12662 7098
rect 12714 7046 15506 7098
rect 15558 7046 15570 7098
rect 15622 7046 15634 7098
rect 15686 7046 15698 7098
rect 15750 7046 15762 7098
rect 15814 7046 18606 7098
rect 18658 7046 18670 7098
rect 18722 7046 18734 7098
rect 18786 7046 18798 7098
rect 18850 7046 18862 7098
rect 18914 7046 18920 7098
rect 184 7024 18920 7046
rect 1210 6944 1216 6996
rect 1268 6984 1274 6996
rect 1489 6987 1547 6993
rect 1489 6984 1501 6987
rect 1268 6956 1501 6984
rect 1268 6944 1274 6956
rect 1489 6953 1501 6956
rect 1535 6953 1547 6987
rect 1489 6947 1547 6953
rect 17957 6987 18015 6993
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18138 6984 18144 6996
rect 18003 6956 18144 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18325 6987 18383 6993
rect 18325 6984 18337 6987
rect 18288 6956 18337 6984
rect 18288 6944 18294 6956
rect 18325 6953 18337 6956
rect 18371 6953 18383 6987
rect 18325 6947 18383 6953
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 8662 6876 8668 6928
rect 8720 6876 8726 6928
rect 2406 6848 2412 6860
rect 1228 6820 2412 6848
rect 1228 6789 1256 6820
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 7006 6848 7012 6860
rect 6967 6820 7012 6848
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 8202 6848 8208 6860
rect 7708 6820 8208 6848
rect 7708 6808 7714 6820
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 11514 6848 11520 6860
rect 11475 6820 11520 6848
rect 11514 6808 11520 6820
rect 11572 6808 11578 6860
rect 12894 6848 12900 6860
rect 12855 6820 12900 6848
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 16758 6848 16764 6860
rect 13403 6820 16764 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 17552 6820 17785 6848
rect 17552 6808 17558 6820
rect 17773 6817 17785 6820
rect 17819 6848 17831 6851
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 17819 6820 18245 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 18233 6817 18245 6820
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6817 18475 6851
rect 18417 6811 18475 6817
rect 1213 6783 1271 6789
rect 1213 6749 1225 6783
rect 1259 6749 1271 6783
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1213 6743 1271 6749
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2832 6752 3157 6780
rect 2832 6740 2838 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8386 6780 8392 6792
rect 8159 6752 8392 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 1946 6712 1952 6724
rect 1903 6684 1952 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 4212 6684 4629 6712
rect 4212 6672 4218 6684
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 6822 6712 6828 6724
rect 4617 6675 4675 6681
rect 5736 6684 6828 6712
rect 5736 6656 5764 6684
rect 6822 6672 6828 6684
rect 6880 6712 6886 6724
rect 7760 6712 7788 6743
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 11238 6780 11244 6792
rect 11199 6752 11244 6780
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6780 11483 6783
rect 11606 6780 11612 6792
rect 11471 6752 11612 6780
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 11606 6740 11612 6752
rect 11664 6780 11670 6792
rect 13814 6780 13820 6792
rect 11664 6752 13820 6780
rect 11664 6740 11670 6752
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 14516 6752 16313 6780
rect 14516 6740 14522 6752
rect 16301 6749 16313 6752
rect 16347 6780 16359 6783
rect 16574 6780 16580 6792
rect 16347 6752 16580 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 18432 6780 18460 6811
rect 17635 6752 18460 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 6880 6684 7788 6712
rect 11333 6715 11391 6721
rect 6880 6672 6886 6684
rect 11333 6681 11345 6715
rect 11379 6712 11391 6715
rect 12802 6712 12808 6724
rect 11379 6684 12808 6712
rect 11379 6681 11391 6684
rect 11333 6675 11391 6681
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 15746 6712 15752 6724
rect 15120 6684 15752 6712
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 5718 6644 5724 6656
rect 2924 6616 5724 6644
rect 2924 6604 2930 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6638 6644 6644 6656
rect 5868 6616 6644 6644
rect 5868 6604 5874 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9493 6647 9551 6653
rect 9493 6644 9505 6647
rect 8996 6616 9505 6644
rect 8996 6604 9002 6616
rect 9493 6613 9505 6616
rect 9539 6613 9551 6647
rect 9493 6607 9551 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 15120 6644 15148 6684
rect 15746 6672 15752 6684
rect 15804 6672 15810 6724
rect 16390 6712 16396 6724
rect 16040 6684 16396 6712
rect 15378 6644 15384 6656
rect 12216 6616 15148 6644
rect 15339 6616 15384 6644
rect 12216 6604 12222 6616
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 15933 6647 15991 6653
rect 15933 6644 15945 6647
rect 15896 6616 15945 6644
rect 15896 6604 15902 6616
rect 15933 6613 15945 6616
rect 15979 6644 15991 6647
rect 16040 6644 16068 6684
rect 16390 6672 16396 6684
rect 16448 6712 16454 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16448 6684 16681 6712
rect 16448 6672 16454 6684
rect 16669 6681 16681 6684
rect 16715 6712 16727 6715
rect 17221 6715 17279 6721
rect 17221 6712 17233 6715
rect 16715 6684 17233 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 17221 6681 17233 6684
rect 17267 6712 17279 6715
rect 17604 6712 17632 6743
rect 17267 6684 17632 6712
rect 17267 6681 17279 6684
rect 17221 6675 17279 6681
rect 15979 6616 16068 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 184 6554 18860 6576
rect 184 6502 1556 6554
rect 1608 6502 1620 6554
rect 1672 6502 1684 6554
rect 1736 6502 1748 6554
rect 1800 6502 1812 6554
rect 1864 6502 4656 6554
rect 4708 6502 4720 6554
rect 4772 6502 4784 6554
rect 4836 6502 4848 6554
rect 4900 6502 4912 6554
rect 4964 6502 7756 6554
rect 7808 6502 7820 6554
rect 7872 6502 7884 6554
rect 7936 6502 7948 6554
rect 8000 6502 8012 6554
rect 8064 6502 10856 6554
rect 10908 6502 10920 6554
rect 10972 6502 10984 6554
rect 11036 6502 11048 6554
rect 11100 6502 11112 6554
rect 11164 6502 13956 6554
rect 14008 6502 14020 6554
rect 14072 6502 14084 6554
rect 14136 6502 14148 6554
rect 14200 6502 14212 6554
rect 14264 6502 17056 6554
rect 17108 6502 17120 6554
rect 17172 6502 17184 6554
rect 17236 6502 17248 6554
rect 17300 6502 17312 6554
rect 17364 6502 18860 6554
rect 184 6480 18860 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1673 6443 1731 6449
rect 1673 6440 1685 6443
rect 1452 6412 1685 6440
rect 1452 6400 1458 6412
rect 1673 6409 1685 6412
rect 1719 6409 1731 6443
rect 1673 6403 1731 6409
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 2280 6412 3985 6440
rect 2280 6400 2286 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 5626 6440 5632 6452
rect 3973 6403 4031 6409
rect 4540 6412 5632 6440
rect 4540 6372 4568 6412
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11330 6440 11336 6452
rect 11195 6412 11336 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 12639 6443 12697 6449
rect 12639 6409 12651 6443
rect 12685 6440 12697 6443
rect 17586 6440 17592 6452
rect 12685 6412 17592 6440
rect 12685 6409 12697 6412
rect 12639 6403 12697 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18012 6412 18337 6440
rect 18012 6400 18018 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 4448 6344 4568 6372
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2222 6304 2228 6316
rect 2087 6276 2228 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 4448 6313 4476 6344
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5810 6372 5816 6384
rect 5592 6344 5816 6372
rect 5592 6332 5598 6344
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 5905 6375 5963 6381
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 5994 6372 6000 6384
rect 5951 6344 6000 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 8754 6372 8760 6384
rect 7668 6344 8760 6372
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4580 6276 4625 6304
rect 4580 6264 4586 6276
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 6365 6307 6423 6313
rect 5316 6276 6040 6304
rect 5316 6264 5322 6276
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2409 6239 2467 6245
rect 2409 6236 2421 6239
rect 1995 6208 2421 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2409 6205 2421 6208
rect 2455 6236 2467 6239
rect 3878 6236 3884 6248
rect 2455 6208 3884 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 3878 6196 3884 6208
rect 3936 6236 3942 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 3936 6208 5181 6236
rect 3936 6196 3942 6208
rect 5169 6205 5181 6208
rect 5215 6236 5227 6239
rect 5350 6236 5356 6248
rect 5215 6208 5356 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5350 6196 5356 6208
rect 5408 6236 5414 6248
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5408 6208 5641 6236
rect 5408 6196 5414 6208
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 5629 6199 5687 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6012 6245 6040 6276
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 5993 6239 6051 6245
rect 5993 6205 6005 6239
rect 6039 6205 6051 6239
rect 5993 6199 6051 6205
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 4387 6140 5672 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 5534 6100 5540 6112
rect 3844 6072 5540 6100
rect 3844 6060 3850 6072
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5644 6100 5672 6140
rect 5718 6128 5724 6180
rect 5776 6168 5782 6180
rect 6380 6168 6408 6267
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 7668 6304 7696 6344
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 9214 6372 9220 6384
rect 9175 6344 9220 6372
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 15010 6372 15016 6384
rect 14783 6344 15016 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 6696 6276 7696 6304
rect 6696 6264 6702 6276
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 9232 6304 9260 6332
rect 8536 6276 9260 6304
rect 8536 6264 8542 6276
rect 11422 6264 11428 6316
rect 11480 6304 11486 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 11480 6276 12909 6304
rect 11480 6264 11486 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 14424 6276 15301 6304
rect 14424 6264 14430 6276
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13228 6208 14013 6236
rect 13228 6196 13234 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14458 6236 14464 6248
rect 14419 6208 14464 6236
rect 14277 6199 14335 6205
rect 6638 6168 6644 6180
rect 5776 6140 6408 6168
rect 6599 6140 6644 6168
rect 5776 6128 5782 6140
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 8018 6168 8024 6180
rect 7866 6140 8024 6168
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 8260 6140 9045 6168
rect 8260 6128 8266 6140
rect 9033 6137 9045 6140
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 12158 6128 12164 6180
rect 12216 6128 12222 6180
rect 14292 6168 14320 6199
rect 14458 6196 14464 6208
rect 14516 6236 14522 6248
rect 14642 6236 14648 6248
rect 14516 6208 14648 6236
rect 14516 6196 14522 6208
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 14826 6236 14832 6248
rect 14739 6208 14832 6236
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 14936 6245 14964 6276
rect 15289 6273 15301 6276
rect 15335 6304 15347 6307
rect 15838 6304 15844 6316
rect 15335 6276 15844 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 18046 6304 18052 6316
rect 16531 6276 18052 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 14550 6168 14556 6180
rect 14292 6140 14556 6168
rect 14550 6128 14556 6140
rect 14608 6128 14614 6180
rect 14844 6168 14872 6196
rect 15378 6168 15384 6180
rect 14844 6140 15384 6168
rect 15378 6128 15384 6140
rect 15436 6128 15442 6180
rect 16776 6140 16882 6168
rect 7006 6100 7012 6112
rect 5644 6072 7012 6100
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 7616 6072 8125 6100
rect 7616 6060 7622 6072
rect 8113 6069 8125 6072
rect 8159 6069 8171 6103
rect 8113 6063 8171 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9272 6072 9689 6100
rect 9272 6060 9278 6072
rect 9677 6069 9689 6072
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16776 6100 16804 6140
rect 15988 6072 16804 6100
rect 15988 6060 15994 6072
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17911 6103 17969 6109
rect 17911 6100 17923 6103
rect 17000 6072 17923 6100
rect 17000 6060 17006 6072
rect 17911 6069 17923 6072
rect 17957 6069 17969 6103
rect 17911 6063 17969 6069
rect 184 6010 18920 6032
rect 184 5958 3106 6010
rect 3158 5958 3170 6010
rect 3222 5958 3234 6010
rect 3286 5958 3298 6010
rect 3350 5958 3362 6010
rect 3414 5958 6206 6010
rect 6258 5958 6270 6010
rect 6322 5958 6334 6010
rect 6386 5958 6398 6010
rect 6450 5958 6462 6010
rect 6514 5958 9306 6010
rect 9358 5958 9370 6010
rect 9422 5958 9434 6010
rect 9486 5958 9498 6010
rect 9550 5958 9562 6010
rect 9614 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 12534 6010
rect 12586 5958 12598 6010
rect 12650 5958 12662 6010
rect 12714 5958 15506 6010
rect 15558 5958 15570 6010
rect 15622 5958 15634 6010
rect 15686 5958 15698 6010
rect 15750 5958 15762 6010
rect 15814 5958 18606 6010
rect 18658 5958 18670 6010
rect 18722 5958 18734 6010
rect 18786 5958 18798 6010
rect 18850 5958 18862 6010
rect 18914 5958 18920 6010
rect 184 5936 18920 5958
rect 2038 5856 2044 5908
rect 2096 5856 2102 5908
rect 8018 5896 8024 5908
rect 5828 5868 8024 5896
rect 2056 5828 2084 5856
rect 2225 5831 2283 5837
rect 2225 5828 2237 5831
rect 2056 5800 2237 5828
rect 2225 5797 2237 5800
rect 2271 5828 2283 5831
rect 4430 5828 4436 5840
rect 2271 5800 4436 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 2004 5732 2053 5760
rect 2004 5720 2010 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 3234 5760 3240 5772
rect 2363 5732 3240 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3344 5769 3372 5800
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 5828 5828 5856 5868
rect 8018 5856 8024 5868
rect 8076 5896 8082 5908
rect 10873 5899 10931 5905
rect 8076 5868 9168 5896
rect 8076 5856 8082 5868
rect 5902 5828 5908 5840
rect 5828 5800 5908 5828
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7432 5800 7849 5828
rect 7432 5788 7438 5800
rect 7837 5797 7849 5800
rect 7883 5797 7895 5831
rect 9140 5828 9168 5868
rect 10873 5865 10885 5899
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 9214 5828 9220 5840
rect 9062 5800 9220 5828
rect 7837 5791 7895 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 10888 5828 10916 5859
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 18233 5899 18291 5905
rect 16172 5868 16804 5896
rect 16172 5856 16178 5868
rect 10888 5800 11560 5828
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5729 3387 5763
rect 3878 5760 3884 5772
rect 3839 5732 3884 5760
rect 3329 5723 3387 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 4396 5732 5549 5760
rect 4396 5720 4402 5732
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11422 5760 11428 5772
rect 11195 5732 11428 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 2280 5664 3525 5692
rect 2280 5652 2286 5664
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2740 5596 2973 5624
rect 2740 5584 2746 5596
rect 2961 5593 2973 5596
rect 3007 5593 3019 5627
rect 2961 5587 3019 5593
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 3160 5556 3188 5664
rect 3513 5661 3525 5664
rect 3559 5661 3571 5695
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3513 5655 3571 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 3896 5692 3924 5720
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 3896 5664 4721 5692
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 5166 5692 5172 5704
rect 5127 5664 5172 5692
rect 4709 5655 4767 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 6880 5664 7573 5692
rect 6880 5652 6886 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 9582 5692 9588 5704
rect 9543 5664 9588 5692
rect 7561 5655 7619 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 10980 5692 11008 5723
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 11532 5769 11560 5800
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 12216 5800 12834 5828
rect 12216 5788 12222 5800
rect 15930 5788 15936 5840
rect 15988 5788 15994 5840
rect 16776 5772 16804 5868
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18322 5896 18328 5908
rect 18279 5868 18328 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 11664 5732 11709 5760
rect 11664 5720 11670 5732
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 16758 5760 16764 5772
rect 11848 5732 11893 5760
rect 16671 5732 16764 5760
rect 11848 5720 11854 5732
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18414 5760 18420 5772
rect 18003 5732 18420 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18414 5720 18420 5732
rect 18472 5720 18478 5772
rect 11624 5692 11652 5720
rect 10980 5664 11652 5692
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 12023 5664 13829 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13817 5655 13875 5661
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5692 14243 5695
rect 14274 5692 14280 5704
rect 14231 5664 14280 5692
rect 14231 5661 14243 5664
rect 14185 5655 14243 5661
rect 3234 5584 3240 5636
rect 3292 5624 3298 5636
rect 5074 5624 5080 5636
rect 3292 5596 5080 5624
rect 3292 5584 3298 5596
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 10689 5627 10747 5633
rect 10689 5593 10701 5627
rect 10735 5624 10747 5627
rect 11238 5624 11244 5636
rect 10735 5596 11244 5624
rect 10735 5593 10747 5596
rect 10689 5587 10747 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11716 5624 11744 5655
rect 14274 5652 14280 5664
rect 14332 5692 14338 5704
rect 16114 5692 16120 5704
rect 14332 5664 16120 5692
rect 14332 5652 14338 5664
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 16264 5664 16405 5692
rect 16264 5652 16270 5664
rect 16393 5661 16405 5664
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 12250 5624 12256 5636
rect 11716 5596 12256 5624
rect 12250 5584 12256 5596
rect 12308 5624 12314 5636
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 12308 5596 12449 5624
rect 12308 5584 12314 5596
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 4246 5556 4252 5568
rect 3160 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5556 4310 5568
rect 5350 5556 5356 5568
rect 4304 5528 5356 5556
rect 4304 5516 4310 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7098 5556 7104 5568
rect 6963 5528 7104 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 10226 5556 10232 5568
rect 10091 5528 10232 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 14826 5516 14832 5568
rect 14884 5556 14890 5568
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14884 5528 15025 5556
rect 14884 5516 14890 5528
rect 15013 5525 15025 5528
rect 15059 5525 15071 5559
rect 15013 5519 15071 5525
rect 184 5466 18860 5488
rect 184 5414 1556 5466
rect 1608 5414 1620 5466
rect 1672 5414 1684 5466
rect 1736 5414 1748 5466
rect 1800 5414 1812 5466
rect 1864 5414 4656 5466
rect 4708 5414 4720 5466
rect 4772 5414 4784 5466
rect 4836 5414 4848 5466
rect 4900 5414 4912 5466
rect 4964 5414 7756 5466
rect 7808 5414 7820 5466
rect 7872 5414 7884 5466
rect 7936 5414 7948 5466
rect 8000 5414 8012 5466
rect 8064 5414 10856 5466
rect 10908 5414 10920 5466
rect 10972 5414 10984 5466
rect 11036 5414 11048 5466
rect 11100 5414 11112 5466
rect 11164 5414 13956 5466
rect 14008 5414 14020 5466
rect 14072 5414 14084 5466
rect 14136 5414 14148 5466
rect 14200 5414 14212 5466
rect 14264 5414 17056 5466
rect 17108 5414 17120 5466
rect 17172 5414 17184 5466
rect 17236 5414 17248 5466
rect 17300 5414 17312 5466
rect 17364 5414 18860 5466
rect 184 5392 18860 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 1673 5355 1731 5361
rect 1673 5352 1685 5355
rect 1636 5324 1685 5352
rect 1636 5312 1642 5324
rect 1673 5321 1685 5324
rect 1719 5352 1731 5355
rect 2038 5352 2044 5364
rect 1719 5324 2044 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 4522 5352 4528 5364
rect 3191 5324 4528 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 5224 5324 5365 5352
rect 5224 5312 5230 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8110 5352 8116 5364
rect 7883 5324 8116 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 11238 5352 11244 5364
rect 11195 5324 11244 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14274 5352 14280 5364
rect 14047 5324 14280 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2130 5284 2136 5296
rect 1811 5256 2136 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2130 5244 2136 5256
rect 2188 5244 2194 5296
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 4065 5287 4123 5293
rect 4065 5284 4077 5287
rect 3936 5256 4077 5284
rect 3936 5244 3942 5256
rect 4065 5253 4077 5256
rect 4111 5253 4123 5287
rect 4065 5247 4123 5253
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8904 5256 9045 5284
rect 8904 5244 8910 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2774 5216 2780 5228
rect 1903 5188 2780 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 7282 5216 7288 5228
rect 5316 5188 7288 5216
rect 5316 5176 5322 5188
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 11790 5216 11796 5228
rect 7340 5188 9076 5216
rect 11751 5188 11796 5216
rect 7340 5176 7346 5188
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 900 5120 1593 5148
rect 900 5108 906 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 3053 5151 3111 5157
rect 3053 5148 3065 5151
rect 2740 5120 3065 5148
rect 2740 5108 2746 5120
rect 3053 5117 3065 5120
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3936 5120 3985 5148
rect 3936 5108 3942 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 4246 5148 4252 5160
rect 4207 5120 4252 5148
rect 3973 5111 4031 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4430 5148 4436 5160
rect 4391 5120 4436 5148
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5718 5148 5724 5160
rect 5675 5120 5724 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 6914 5148 6920 5160
rect 6871 5120 6920 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 8202 5148 8208 5160
rect 7423 5120 8208 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8754 5148 8760 5160
rect 8352 5120 8760 5148
rect 8352 5108 8358 5120
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8904 5120 8953 5148
rect 8904 5108 8910 5120
rect 8941 5117 8953 5120
rect 8987 5117 8999 5151
rect 9048 5148 9076 5188
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 9214 5148 9220 5160
rect 9048 5120 9220 5148
rect 8941 5111 8999 5117
rect 9214 5108 9220 5120
rect 9272 5148 9278 5160
rect 9582 5148 9588 5160
rect 9272 5120 9365 5148
rect 9543 5120 9588 5148
rect 9272 5108 9278 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 15286 5148 15292 5160
rect 15247 5120 15292 5148
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 4798 5040 4804 5092
rect 4856 5080 4862 5092
rect 5442 5080 5448 5092
rect 4856 5052 5448 5080
rect 4856 5040 4862 5052
rect 5442 5040 5448 5052
rect 5500 5080 5506 5092
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 5500 5052 6377 5080
rect 5500 5040 5506 5052
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 9030 5040 9036 5092
rect 9088 5080 9094 5092
rect 9600 5080 9628 5108
rect 10226 5080 10232 5092
rect 9088 5052 9628 5080
rect 10187 5052 10232 5080
rect 9088 5040 9094 5052
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4522 5012 4528 5024
rect 4387 4984 4528 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6880 4984 7297 5012
rect 6880 4972 6886 4984
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 7285 4975 7343 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11655 4984 12265 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 12253 4981 12265 4984
rect 12299 5012 12311 5015
rect 12894 5012 12900 5024
rect 12299 4984 12900 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 184 4922 18920 4944
rect 184 4870 3106 4922
rect 3158 4870 3170 4922
rect 3222 4870 3234 4922
rect 3286 4870 3298 4922
rect 3350 4870 3362 4922
rect 3414 4870 6206 4922
rect 6258 4870 6270 4922
rect 6322 4870 6334 4922
rect 6386 4870 6398 4922
rect 6450 4870 6462 4922
rect 6514 4870 9306 4922
rect 9358 4870 9370 4922
rect 9422 4870 9434 4922
rect 9486 4870 9498 4922
rect 9550 4870 9562 4922
rect 9614 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 12534 4922
rect 12586 4870 12598 4922
rect 12650 4870 12662 4922
rect 12714 4870 15506 4922
rect 15558 4870 15570 4922
rect 15622 4870 15634 4922
rect 15686 4870 15698 4922
rect 15750 4870 15762 4922
rect 15814 4870 18606 4922
rect 18658 4870 18670 4922
rect 18722 4870 18734 4922
rect 18786 4870 18798 4922
rect 18850 4870 18862 4922
rect 18914 4870 18920 4922
rect 184 4848 18920 4870
rect 842 4808 848 4820
rect 803 4780 848 4808
rect 842 4768 848 4780
rect 900 4768 906 4820
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 2866 4808 2872 4820
rect 1811 4780 2872 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4982 4808 4988 4820
rect 4571 4780 4988 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4808 5414 4820
rect 5810 4808 5816 4820
rect 5408 4780 5816 4808
rect 5408 4768 5414 4780
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 7006 4768 7012 4780
rect 7064 4808 7070 4820
rect 7190 4808 7196 4820
rect 7064 4780 7196 4808
rect 7064 4768 7070 4780
rect 7190 4768 7196 4780
rect 7248 4808 7254 4820
rect 8386 4808 8392 4820
rect 7248 4780 7788 4808
rect 8347 4780 8392 4808
rect 7248 4768 7254 4780
rect 4341 4743 4399 4749
rect 4341 4709 4353 4743
rect 4387 4740 4399 4743
rect 5166 4740 5172 4752
rect 4387 4712 5172 4740
rect 4387 4709 4399 4712
rect 4341 4703 4399 4709
rect 5166 4700 5172 4712
rect 5224 4700 5230 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 7760 4749 7788 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11330 4808 11336 4820
rect 11011 4780 11336 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4777 12955 4811
rect 17402 4808 17408 4820
rect 12897 4771 12955 4777
rect 14660 4780 17408 4808
rect 7745 4743 7803 4749
rect 6052 4712 6868 4740
rect 6052 4700 6058 4712
rect 934 4672 940 4684
rect 895 4644 940 4672
rect 934 4632 940 4644
rect 992 4632 998 4684
rect 1026 4632 1032 4684
rect 1084 4672 1090 4684
rect 1489 4675 1547 4681
rect 1489 4672 1501 4675
rect 1084 4644 1501 4672
rect 1084 4632 1090 4644
rect 1489 4641 1501 4644
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 4246 4672 4252 4684
rect 1636 4644 1681 4672
rect 4207 4644 4252 4672
rect 1636 4632 1642 4644
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 4706 4672 4712 4684
rect 4667 4644 4712 4672
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 6840 4681 6868 4712
rect 7745 4709 7757 4743
rect 7791 4709 7803 4743
rect 8757 4743 8815 4749
rect 8757 4740 8769 4743
rect 7745 4703 7803 4709
rect 8220 4712 8769 4740
rect 6641 4675 6699 4681
rect 4856 4644 4901 4672
rect 4856 4632 4862 4644
rect 6641 4641 6653 4675
rect 6687 4641 6699 4675
rect 6795 4675 6868 4681
rect 6795 4672 6807 4675
rect 6735 4644 6807 4672
rect 6641 4635 6699 4641
rect 6795 4641 6807 4644
rect 6841 4672 6868 4675
rect 7466 4672 7472 4684
rect 6841 4644 7472 4672
rect 6841 4641 6853 4644
rect 6795 4635 6853 4641
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2590 4604 2596 4616
rect 1811 4576 2596 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 6656 4604 6684 4635
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 8113 4675 8171 4681
rect 7576 4644 7972 4672
rect 7576 4604 7604 4644
rect 6656 4576 6868 4604
rect 6840 4548 6868 4576
rect 6932 4576 7604 4604
rect 7837 4607 7895 4613
rect 6822 4496 6828 4548
rect 6880 4496 6886 4548
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 6932 4468 6960 4576
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7944 4604 7972 4644
rect 8113 4641 8125 4675
rect 8159 4673 8171 4675
rect 8220 4673 8248 4712
rect 8757 4709 8769 4712
rect 8803 4709 8815 4743
rect 8757 4703 8815 4709
rect 9214 4700 9220 4752
rect 9272 4740 9278 4752
rect 10137 4743 10195 4749
rect 10137 4740 10149 4743
rect 9272 4712 10149 4740
rect 9272 4700 9278 4712
rect 10137 4709 10149 4712
rect 10183 4709 10195 4743
rect 10137 4703 10195 4709
rect 8159 4645 8248 4673
rect 8665 4675 8723 4681
rect 8159 4641 8171 4645
rect 8113 4635 8171 4641
rect 8665 4641 8677 4675
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 8849 4675 8907 4681
rect 8849 4641 8861 4675
rect 8895 4672 8907 4675
rect 8938 4672 8944 4684
rect 8895 4644 8944 4672
rect 8895 4641 8907 4644
rect 8849 4635 8907 4641
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 7944 4576 8217 4604
rect 7837 4567 7895 4573
rect 8205 4573 8217 4576
rect 8251 4604 8263 4607
rect 8478 4604 8484 4616
rect 8251 4576 8484 4604
rect 8251 4573 8263 4576
rect 8205 4567 8263 4573
rect 7852 4536 7880 4567
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8680 4604 8708 4635
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 10008 4644 10425 4672
rect 10008 4632 10014 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 10413 4635 10471 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11790 4672 11796 4684
rect 11624 4644 11796 4672
rect 11422 4604 11428 4616
rect 8680 4576 8892 4604
rect 11383 4576 11428 4604
rect 8754 4536 8760 4548
rect 7852 4508 8760 4536
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 5776 4440 6960 4468
rect 5776 4428 5782 4440
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8864 4468 8892 4576
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11624 4613 11652 4644
rect 11790 4632 11796 4644
rect 11848 4672 11854 4684
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 11848 4644 12633 4672
rect 11848 4632 11854 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4641 12863 4675
rect 12912 4672 12940 4771
rect 13814 4740 13820 4752
rect 13556 4712 13820 4740
rect 13556 4681 13584 4712
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 12912 4644 13461 4672
rect 12805 4635 12863 4641
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4641 13599 4675
rect 13541 4635 13599 4641
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4672 13783 4675
rect 14274 4672 14280 4684
rect 13771 4644 14280 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 12636 4536 12664 4635
rect 12820 4604 12848 4635
rect 13556 4604 13584 4635
rect 12820 4576 13584 4604
rect 12636 4508 13216 4536
rect 13078 4468 13084 4480
rect 7524 4440 8892 4468
rect 13039 4440 13084 4468
rect 7524 4428 7530 4440
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13188 4468 13216 4508
rect 13630 4496 13636 4548
rect 13688 4536 13694 4548
rect 13688 4508 13733 4536
rect 13688 4496 13694 4508
rect 13832 4468 13860 4644
rect 14274 4632 14280 4644
rect 14332 4672 14338 4684
rect 14660 4672 14688 4780
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 15930 4700 15936 4752
rect 15988 4700 15994 4752
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 17129 4743 17187 4749
rect 17129 4740 17141 4743
rect 16632 4712 17141 4740
rect 16632 4700 16638 4712
rect 17129 4709 17141 4712
rect 17175 4709 17187 4743
rect 17129 4703 17187 4709
rect 14332 4644 14688 4672
rect 14332 4632 14338 4644
rect 16758 4632 16764 4684
rect 16816 4672 16822 4684
rect 16816 4644 16861 4672
rect 16816 4632 16822 4644
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17737 4675 17795 4681
rect 17737 4672 17749 4675
rect 17000 4644 17749 4672
rect 17000 4632 17006 4644
rect 17737 4641 17749 4644
rect 17783 4641 17795 4675
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17737 4635 17795 4641
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 17957 4675 18015 4681
rect 17957 4641 17969 4675
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 17972 4604 18000 4635
rect 16531 4576 16712 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 16684 4480 16712 4576
rect 17788 4576 18000 4604
rect 17788 4548 17816 4576
rect 17770 4496 17776 4548
rect 17828 4496 17834 4548
rect 13188 4440 13860 4468
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14918 4468 14924 4480
rect 13955 4440 14924 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15010 4428 15016 4480
rect 15068 4468 15074 4480
rect 15068 4440 15113 4468
rect 15068 4428 15074 4440
rect 16666 4428 16672 4480
rect 16724 4428 16730 4480
rect 18138 4468 18144 4480
rect 18099 4440 18144 4468
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 184 4378 18860 4400
rect 184 4326 1556 4378
rect 1608 4326 1620 4378
rect 1672 4326 1684 4378
rect 1736 4326 1748 4378
rect 1800 4326 1812 4378
rect 1864 4326 4656 4378
rect 4708 4326 4720 4378
rect 4772 4326 4784 4378
rect 4836 4326 4848 4378
rect 4900 4326 4912 4378
rect 4964 4326 7756 4378
rect 7808 4326 7820 4378
rect 7872 4326 7884 4378
rect 7936 4326 7948 4378
rect 8000 4326 8012 4378
rect 8064 4326 10856 4378
rect 10908 4326 10920 4378
rect 10972 4326 10984 4378
rect 11036 4326 11048 4378
rect 11100 4326 11112 4378
rect 11164 4326 13956 4378
rect 14008 4326 14020 4378
rect 14072 4326 14084 4378
rect 14136 4326 14148 4378
rect 14200 4326 14212 4378
rect 14264 4326 17056 4378
rect 17108 4326 17120 4378
rect 17172 4326 17184 4378
rect 17236 4326 17248 4378
rect 17300 4326 17312 4378
rect 17364 4326 18860 4378
rect 184 4304 18860 4326
rect 2590 4264 2596 4276
rect 2551 4236 2596 4264
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 5813 4267 5871 4273
rect 5813 4264 5825 4267
rect 5132 4236 5825 4264
rect 5132 4224 5138 4236
rect 5813 4233 5825 4236
rect 5859 4233 5871 4267
rect 5813 4227 5871 4233
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7248 4236 7573 4264
rect 7248 4224 7254 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 8754 4264 8760 4276
rect 8715 4236 8760 4264
rect 7561 4227 7619 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9766 4264 9772 4276
rect 8996 4236 9628 4264
rect 9727 4236 9772 4264
rect 8996 4224 9002 4236
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 4154 4196 4160 4208
rect 2924 4168 4160 4196
rect 2924 4156 2930 4168
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 6880 4168 9352 4196
rect 6880 4156 6886 4168
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2225 4131 2283 4137
rect 2225 4128 2237 4131
rect 2004 4100 2237 4128
rect 2004 4088 2010 4100
rect 2225 4097 2237 4100
rect 2271 4128 2283 4131
rect 2314 4128 2320 4140
rect 2271 4100 2320 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2314 4088 2320 4100
rect 2372 4128 2378 4140
rect 5994 4128 6000 4140
rect 2372 4100 3004 4128
rect 5955 4100 6000 4128
rect 2372 4088 2378 4100
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 2976 4069 3004 4100
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 9324 4137 9352 4168
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6564 4100 7389 4128
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2740 4032 2789 4060
rect 2740 4020 2746 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2976 4063 3055 4069
rect 2777 4023 2835 4029
rect 2869 4041 2927 4047
rect 2869 4007 2881 4041
rect 2915 4007 2927 4041
rect 2976 4032 3009 4063
rect 2997 4029 3009 4032
rect 3043 4060 3055 4063
rect 3510 4060 3516 4072
rect 3043 4032 3516 4060
rect 3043 4029 3055 4032
rect 2997 4023 3055 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 5718 4060 5724 4072
rect 5679 4032 5724 4060
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 2869 4001 2927 4007
rect 2884 3936 2912 4001
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6564 3992 6592 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7377 4091 7435 4097
rect 7484 4100 8033 4128
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4060 6791 4063
rect 7484 4060 7512 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9600 4128 9628 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11480 4236 11897 4264
rect 11480 4224 11486 4236
rect 11885 4233 11897 4236
rect 11931 4264 11943 4267
rect 12253 4267 12311 4273
rect 12253 4264 12265 4267
rect 11931 4236 12265 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12253 4233 12265 4236
rect 12299 4264 12311 4267
rect 14642 4264 14648 4276
rect 12299 4236 14648 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 15301 4267 15359 4273
rect 15301 4264 15313 4267
rect 14976 4236 15313 4264
rect 14976 4224 14982 4236
rect 15301 4233 15313 4236
rect 15347 4233 15359 4267
rect 15301 4227 15359 4233
rect 16758 4224 16764 4276
rect 16816 4224 16822 4276
rect 16776 4196 16804 4224
rect 16546 4168 16804 4196
rect 9674 4128 9680 4140
rect 9587 4100 9680 4128
rect 9309 4091 9367 4097
rect 9674 4088 9680 4100
rect 9732 4128 9738 4140
rect 9732 4100 9996 4128
rect 9732 4088 9738 4100
rect 6779 4032 7512 4060
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 6043 3964 6592 3992
rect 6656 3992 6684 4023
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7929 4063 7987 4069
rect 7708 4032 7753 4060
rect 7708 4020 7714 4032
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7929 4023 7987 4029
rect 8036 4032 8125 4060
rect 6822 3992 6828 4004
rect 6656 3964 6828 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 7006 3992 7012 4004
rect 6967 3964 7012 3992
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 7101 3995 7159 4001
rect 7101 3961 7113 3995
rect 7147 3992 7159 3995
rect 7190 3992 7196 4004
rect 7147 3964 7196 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 7374 3992 7380 4004
rect 7335 3964 7380 3992
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 7944 3992 7972 4023
rect 7524 3964 7972 3992
rect 7524 3952 7530 3964
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 992 3896 1593 3924
rect 992 3884 998 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1946 3924 1952 3936
rect 1907 3896 1952 3924
rect 1581 3887 1639 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2096 3896 2141 3924
rect 2096 3884 2102 3896
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6638 3924 6644 3936
rect 6503 3896 6644 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8036 3924 8064 4032
rect 8113 4029 8125 4032
rect 8159 4060 8171 4063
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 8159 4032 9781 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 9769 4029 9781 4032
rect 9815 4060 9827 4063
rect 9858 4060 9864 4072
rect 9815 4032 9864 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 9968 4069 9996 4100
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13688 4100 13829 4128
rect 13688 4088 13694 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15565 4131 15623 4137
rect 15565 4128 15577 4131
rect 14976 4100 15577 4128
rect 14976 4088 14982 4100
rect 15565 4097 15577 4100
rect 15611 4128 15623 4131
rect 16546 4128 16574 4168
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 15611 4100 16574 4128
rect 16684 4100 16773 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16684 4060 16712 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 16942 4088 16948 4140
rect 17000 4128 17006 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17000 4100 17325 4128
rect 17000 4088 17006 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17862 4128 17868 4140
rect 17313 4091 17371 4097
rect 17696 4100 17868 4128
rect 17696 4069 17724 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 16632 4032 16712 4060
rect 16776 4032 17693 4060
rect 16632 4020 16638 4032
rect 8938 3952 8944 4004
rect 8996 3992 9002 4004
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 8996 3964 9229 3992
rect 8996 3952 9002 3964
rect 9217 3961 9229 3964
rect 9263 3992 9275 3995
rect 10226 3992 10232 4004
rect 9263 3964 10232 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 15930 3992 15936 4004
rect 14858 3964 15936 3992
rect 15930 3952 15936 3964
rect 15988 3952 15994 4004
rect 16776 3936 16804 4032
rect 17681 4029 17693 4032
rect 17727 4029 17739 4063
rect 17681 4023 17739 4029
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 17828 4032 17873 4060
rect 17828 4020 17834 4032
rect 9122 3924 9128 3936
rect 7616 3896 8064 3924
rect 9083 3896 9128 3924
rect 7616 3884 7622 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12952 3896 13185 3924
rect 12952 3884 12958 3896
rect 13173 3893 13185 3896
rect 13219 3924 13231 3927
rect 15378 3924 15384 3936
rect 13219 3896 15384 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 16206 3924 16212 3936
rect 16167 3896 16212 3924
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 16574 3924 16580 3936
rect 16535 3896 16580 3924
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16669 3927 16727 3933
rect 16669 3893 16681 3927
rect 16715 3924 16727 3927
rect 16758 3924 16764 3936
rect 16715 3896 16764 3924
rect 16715 3893 16727 3896
rect 16669 3887 16727 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 17957 3927 18015 3933
rect 17957 3893 17969 3927
rect 18003 3924 18015 3927
rect 18322 3924 18328 3936
rect 18003 3896 18328 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 184 3834 18920 3856
rect 184 3782 3106 3834
rect 3158 3782 3170 3834
rect 3222 3782 3234 3834
rect 3286 3782 3298 3834
rect 3350 3782 3362 3834
rect 3414 3782 6206 3834
rect 6258 3782 6270 3834
rect 6322 3782 6334 3834
rect 6386 3782 6398 3834
rect 6450 3782 6462 3834
rect 6514 3782 9306 3834
rect 9358 3782 9370 3834
rect 9422 3782 9434 3834
rect 9486 3782 9498 3834
rect 9550 3782 9562 3834
rect 9614 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 12534 3834
rect 12586 3782 12598 3834
rect 12650 3782 12662 3834
rect 12714 3782 15506 3834
rect 15558 3782 15570 3834
rect 15622 3782 15634 3834
rect 15686 3782 15698 3834
rect 15750 3782 15762 3834
rect 15814 3782 18606 3834
rect 18658 3782 18670 3834
rect 18722 3782 18734 3834
rect 18786 3782 18798 3834
rect 18850 3782 18862 3834
rect 18914 3782 18920 3834
rect 184 3760 18920 3782
rect 2774 3720 2780 3732
rect 2735 3692 2780 3720
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3602 3680 3608 3732
rect 3660 3680 3666 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4246 3720 4252 3732
rect 3927 3692 4252 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4246 3680 4252 3692
rect 4304 3720 4310 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4304 3692 4629 3720
rect 4304 3680 4310 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 4617 3683 4675 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 11330 3720 11336 3732
rect 11287 3692 11336 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 11572 3692 12357 3720
rect 11572 3680 11578 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12986 3720 12992 3732
rect 12345 3683 12403 3689
rect 12636 3692 12992 3720
rect 3620 3652 3648 3680
rect 11609 3655 11667 3661
rect 3068 3624 4660 3652
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 2958 3584 2964 3596
rect 2740 3556 2964 3584
rect 2740 3544 2746 3556
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3068 3593 3096 3624
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3584 3203 3587
rect 3510 3584 3516 3596
rect 3191 3556 3516 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 3436 3380 3464 3556
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 3694 3593 3700 3596
rect 3651 3587 3700 3593
rect 3651 3553 3663 3587
rect 3697 3553 3700 3587
rect 3651 3547 3700 3553
rect 3682 3546 3700 3547
rect 3694 3544 3700 3546
rect 3752 3544 3758 3596
rect 4154 3584 4160 3596
rect 4115 3556 4160 3584
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 4632 3516 4660 3624
rect 11609 3621 11621 3655
rect 11655 3652 11667 3655
rect 12526 3652 12532 3664
rect 11655 3624 12532 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 12526 3612 12532 3624
rect 12584 3652 12590 3664
rect 12636 3652 12664 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 13136 3692 13553 3720
rect 13136 3680 13142 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 13541 3683 13599 3689
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16632 3692 17141 3720
rect 16632 3680 16638 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18104 3692 18153 3720
rect 18104 3680 18110 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 12584 3624 12664 3652
rect 12713 3655 12771 3661
rect 12584 3612 12590 3624
rect 12713 3621 12725 3655
rect 12759 3652 12771 3655
rect 12802 3652 12808 3664
rect 12759 3624 12808 3652
rect 12759 3621 12771 3624
rect 12713 3615 12771 3621
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 14918 3652 14924 3664
rect 14752 3624 14924 3652
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 5258 3584 5264 3596
rect 4755 3556 5264 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5626 3584 5632 3596
rect 5587 3556 5632 3584
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11480 3556 11713 3584
rect 11480 3544 11486 3556
rect 11701 3553 11713 3556
rect 11747 3553 11759 3587
rect 11701 3547 11759 3553
rect 11900 3556 13032 3584
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4632 3488 5365 3516
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 11900 3525 11928 3556
rect 11885 3519 11943 3525
rect 5592 3488 5637 3516
rect 5592 3476 5598 3488
rect 11885 3485 11897 3519
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3516 12863 3519
rect 12894 3516 12900 3528
rect 12851 3488 12900 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13004 3525 13032 3556
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13872 3556 13921 3584
rect 13872 3544 13878 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14001 3587 14059 3593
rect 14001 3553 14013 3587
rect 14047 3584 14059 3587
rect 14366 3584 14372 3596
rect 14047 3556 14372 3584
rect 14047 3553 14059 3556
rect 14001 3547 14059 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 14752 3593 14780 3624
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 16022 3612 16028 3664
rect 16080 3612 16086 3664
rect 17497 3655 17555 3661
rect 17497 3621 17509 3655
rect 17543 3652 17555 3655
rect 17678 3652 17684 3664
rect 17543 3624 17684 3652
rect 17543 3621 17555 3624
rect 17497 3615 17555 3621
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 17862 3584 17868 3596
rect 17635 3556 17868 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13538 3516 13544 3528
rect 13035 3488 13544 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3516 14243 3519
rect 14274 3516 14280 3528
rect 14231 3488 14280 3516
rect 14231 3485 14243 3488
rect 14185 3479 14243 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14752 3488 15025 3516
rect 14752 3460 14780 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 17604 3516 17632 3547
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 15436 3488 17632 3516
rect 17681 3519 17739 3525
rect 15436 3476 15442 3488
rect 17681 3485 17693 3519
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 4338 3448 4344 3460
rect 4299 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 14734 3408 14740 3460
rect 14792 3408 14798 3460
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 17696 3448 17724 3479
rect 16908 3420 17724 3448
rect 16908 3408 16914 3420
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 3436 3352 4261 3380
rect 4249 3349 4261 3352
rect 4295 3380 4307 3383
rect 5718 3380 5724 3392
rect 4295 3352 5724 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 16482 3380 16488 3392
rect 16443 3352 16488 3380
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 184 3290 18860 3312
rect 184 3238 1556 3290
rect 1608 3238 1620 3290
rect 1672 3238 1684 3290
rect 1736 3238 1748 3290
rect 1800 3238 1812 3290
rect 1864 3238 4656 3290
rect 4708 3238 4720 3290
rect 4772 3238 4784 3290
rect 4836 3238 4848 3290
rect 4900 3238 4912 3290
rect 4964 3238 7756 3290
rect 7808 3238 7820 3290
rect 7872 3238 7884 3290
rect 7936 3238 7948 3290
rect 8000 3238 8012 3290
rect 8064 3238 10856 3290
rect 10908 3238 10920 3290
rect 10972 3238 10984 3290
rect 11036 3238 11048 3290
rect 11100 3238 11112 3290
rect 11164 3238 13956 3290
rect 14008 3238 14020 3290
rect 14072 3238 14084 3290
rect 14136 3238 14148 3290
rect 14200 3238 14212 3290
rect 14264 3238 17056 3290
rect 17108 3238 17120 3290
rect 17172 3238 17184 3290
rect 17236 3238 17248 3290
rect 17300 3238 17312 3290
rect 17364 3238 18860 3290
rect 184 3216 18860 3238
rect 937 3179 995 3185
rect 937 3145 949 3179
rect 983 3176 995 3179
rect 1026 3176 1032 3188
rect 983 3148 1032 3176
rect 983 3145 995 3148
rect 937 3139 995 3145
rect 1026 3136 1032 3148
rect 1084 3136 1090 3188
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2317 3179 2375 3185
rect 2317 3176 2329 3179
rect 2004 3148 2329 3176
rect 2004 3136 2010 3148
rect 2317 3145 2329 3148
rect 2363 3145 2375 3179
rect 2317 3139 2375 3145
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4154 3176 4160 3188
rect 4111 3148 4160 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9180 3148 9413 3176
rect 9180 3136 9186 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12526 3176 12532 3188
rect 12483 3148 12532 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 16666 3176 16672 3188
rect 16627 3148 16672 3176
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17644 3148 17785 3176
rect 17644 3136 17650 3148
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 17920 3148 18337 3176
rect 17920 3136 17926 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 18325 3139 18383 3145
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 8938 3108 8944 3120
rect 6420 3080 8944 3108
rect 6420 3068 6426 3080
rect 8938 3068 8944 3080
rect 8996 3108 9002 3120
rect 12544 3108 12572 3136
rect 13722 3108 13728 3120
rect 8996 3080 9168 3108
rect 12544 3080 13728 3108
rect 8996 3068 9002 3080
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3040 1823 3043
rect 2774 3040 2780 3052
rect 1811 3012 2780 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5684 3012 5917 3040
rect 5684 3000 5690 3012
rect 5905 3009 5917 3012
rect 5951 3040 5963 3043
rect 6822 3040 6828 3052
rect 5951 3012 6828 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 1026 2972 1032 2984
rect 987 2944 1032 2972
rect 1026 2932 1032 2944
rect 1084 2932 1090 2984
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2038 2972 2044 2984
rect 1903 2944 2044 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2958 2932 2964 2984
rect 3016 2972 3022 2984
rect 3694 2972 3700 2984
rect 3016 2944 3700 2972
rect 3016 2932 3022 2944
rect 3694 2932 3700 2944
rect 3752 2972 3758 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3752 2944 3985 2972
rect 3752 2932 3758 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 5350 2972 5356 2984
rect 4203 2944 5356 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 5810 2972 5816 2984
rect 5767 2944 5816 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 5810 2932 5816 2944
rect 5868 2972 5874 2984
rect 6362 2972 6368 2984
rect 5868 2944 6368 2972
rect 5868 2932 5874 2944
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 9140 2972 9168 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 16574 3108 16580 3120
rect 16132 3080 16580 3108
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9272 3012 9965 3040
rect 9272 3000 9278 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 13630 3040 13636 3052
rect 9953 3003 10011 3009
rect 13188 3012 13636 3040
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9140 2944 9873 2972
rect 9861 2941 9873 2944
rect 9907 2972 9919 2975
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 9907 2944 10425 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 10413 2935 10471 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 13188 2981 13216 3012
rect 13630 3000 13636 3012
rect 13688 3040 13694 3052
rect 16132 3049 16160 3080
rect 16574 3068 16580 3080
rect 16632 3108 16638 3120
rect 16945 3111 17003 3117
rect 16945 3108 16957 3111
rect 16632 3080 16957 3108
rect 16632 3068 16638 3080
rect 16945 3077 16957 3080
rect 16991 3108 17003 3111
rect 17494 3108 17500 3120
rect 16991 3080 17500 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 16117 3043 16175 3049
rect 13688 3012 13860 3040
rect 13688 3000 13694 3012
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13173 2975 13231 2981
rect 13035 2944 13124 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13096 2904 13124 2944
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13173 2935 13231 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 13832 2981 13860 3012
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17543 2944 17969 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 17957 2941 17969 2944
rect 18003 2972 18015 2975
rect 19058 2972 19064 2984
rect 18003 2944 19064 2972
rect 18003 2941 18015 2944
rect 17957 2935 18015 2941
rect 14108 2904 14136 2935
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 13096 2876 14136 2904
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 5626 2836 5632 2848
rect 2004 2808 2049 2836
rect 5587 2808 5632 2836
rect 2004 2796 2010 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12986 2836 12992 2848
rect 12492 2808 12992 2836
rect 12492 2796 12498 2808
rect 12986 2796 12992 2808
rect 13044 2836 13050 2848
rect 13096 2836 13124 2876
rect 13044 2808 13124 2836
rect 13044 2796 13050 2808
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 13633 2839 13691 2845
rect 13633 2836 13645 2839
rect 13596 2808 13645 2836
rect 13596 2796 13602 2808
rect 13633 2805 13645 2808
rect 13679 2805 13691 2839
rect 13633 2799 13691 2805
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14366 2836 14372 2848
rect 13964 2808 14372 2836
rect 13964 2796 13970 2808
rect 14366 2796 14372 2808
rect 14424 2836 14430 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14424 2808 14473 2836
rect 14424 2796 14430 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16206 2836 16212 2848
rect 15252 2808 16212 2836
rect 15252 2796 15258 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 16356 2808 16401 2836
rect 16356 2796 16362 2808
rect 184 2746 18920 2768
rect 184 2694 3106 2746
rect 3158 2694 3170 2746
rect 3222 2694 3234 2746
rect 3286 2694 3298 2746
rect 3350 2694 3362 2746
rect 3414 2694 6206 2746
rect 6258 2694 6270 2746
rect 6322 2694 6334 2746
rect 6386 2694 6398 2746
rect 6450 2694 6462 2746
rect 6514 2694 9306 2746
rect 9358 2694 9370 2746
rect 9422 2694 9434 2746
rect 9486 2694 9498 2746
rect 9550 2694 9562 2746
rect 9614 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 12534 2746
rect 12586 2694 12598 2746
rect 12650 2694 12662 2746
rect 12714 2694 15506 2746
rect 15558 2694 15570 2746
rect 15622 2694 15634 2746
rect 15686 2694 15698 2746
rect 15750 2694 15762 2746
rect 15814 2694 18606 2746
rect 18658 2694 18670 2746
rect 18722 2694 18734 2746
rect 18786 2694 18798 2746
rect 18850 2694 18862 2746
rect 18914 2694 18920 2746
rect 184 2672 18920 2694
rect 1026 2592 1032 2644
rect 1084 2632 1090 2644
rect 1673 2635 1731 2641
rect 1673 2632 1685 2635
rect 1084 2604 1685 2632
rect 1084 2592 1090 2604
rect 1673 2601 1685 2604
rect 1719 2601 1731 2635
rect 1673 2595 1731 2601
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5534 2632 5540 2644
rect 5307 2604 5540 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 6052 2604 6469 2632
rect 6052 2592 6058 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 6871 2604 7757 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 7745 2595 7803 2601
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 8076 2604 8217 2632
rect 8076 2592 8082 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 9309 2635 9367 2641
rect 9309 2632 9321 2635
rect 9272 2604 9321 2632
rect 9272 2592 9278 2604
rect 9309 2601 9321 2604
rect 9355 2601 9367 2635
rect 9309 2595 9367 2601
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 13872 2604 14105 2632
rect 13872 2592 13878 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 15378 2632 15384 2644
rect 15291 2604 15384 2632
rect 14093 2595 14151 2601
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 3326 2564 3332 2576
rect 2179 2536 3332 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 3326 2524 3332 2536
rect 3384 2564 3390 2576
rect 3878 2564 3884 2576
rect 3384 2536 3884 2564
rect 3384 2524 3390 2536
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 6917 2567 6975 2573
rect 6917 2533 6929 2567
rect 6963 2564 6975 2567
rect 7282 2564 7288 2576
rect 6963 2536 7288 2564
rect 6963 2533 6975 2536
rect 6917 2527 6975 2533
rect 7282 2524 7288 2536
rect 7340 2564 7346 2576
rect 7340 2536 7604 2564
rect 7340 2524 7346 2536
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 2866 2496 2872 2508
rect 2087 2468 2872 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 4120 2468 5181 2496
rect 4120 2456 4126 2468
rect 5169 2465 5181 2468
rect 5215 2465 5227 2499
rect 5169 2459 5227 2465
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 7098 2496 7104 2508
rect 5408 2468 7104 2496
rect 5408 2456 5414 2468
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7576 2496 7604 2536
rect 7650 2524 7656 2576
rect 7708 2564 7714 2576
rect 8113 2567 8171 2573
rect 8113 2564 8125 2567
rect 7708 2536 8125 2564
rect 7708 2524 7714 2536
rect 8113 2533 8125 2536
rect 8159 2533 8171 2567
rect 8662 2564 8668 2576
rect 8113 2527 8171 2533
rect 8404 2536 8668 2564
rect 8018 2496 8024 2508
rect 7576 2468 8024 2496
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 2314 2428 2320 2440
rect 2275 2400 2320 2428
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 5776 2400 7021 2428
rect 5776 2388 5782 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 8128 2360 8156 2527
rect 8404 2437 8432 2536
rect 8662 2524 8668 2536
rect 8720 2564 8726 2576
rect 9232 2564 9260 2592
rect 9858 2564 9864 2576
rect 8720 2536 9260 2564
rect 9324 2536 9864 2564
rect 8720 2524 8726 2536
rect 9324 2505 9352 2536
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 10594 2564 10600 2576
rect 10244 2536 10600 2564
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9674 2496 9680 2508
rect 9631 2468 9680 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9674 2456 9680 2468
rect 9732 2496 9738 2508
rect 10244 2505 10272 2536
rect 10594 2524 10600 2536
rect 10652 2564 10658 2576
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 10652 2536 10793 2564
rect 10652 2524 10658 2536
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 13906 2564 13912 2576
rect 13679 2536 13912 2564
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 15304 2573 15332 2604
rect 15378 2592 15384 2604
rect 15436 2632 15442 2644
rect 15657 2635 15715 2641
rect 15657 2632 15669 2635
rect 15436 2604 15669 2632
rect 15436 2592 15442 2604
rect 15657 2601 15669 2604
rect 15703 2632 15715 2635
rect 16574 2632 16580 2644
rect 15703 2604 16580 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 17770 2632 17776 2644
rect 17267 2604 17776 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14884 2536 14933 2564
rect 14884 2524 14890 2536
rect 14921 2533 14933 2536
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2533 15347 2567
rect 16758 2564 16764 2576
rect 15289 2527 15347 2533
rect 16546 2536 16764 2564
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9732 2468 10241 2496
rect 9732 2456 9738 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2465 10563 2499
rect 13722 2496 13728 2508
rect 13683 2468 13728 2496
rect 10505 2459 10563 2465
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9140 2360 9168 2391
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9916 2400 9965 2428
rect 9916 2388 9922 2400
rect 9953 2397 9965 2400
rect 9999 2428 10011 2431
rect 10520 2428 10548 2459
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 14936 2496 14964 2527
rect 16546 2496 16574 2536
rect 16758 2524 16764 2536
rect 16816 2564 16822 2576
rect 16816 2536 17908 2564
rect 16816 2524 16822 2536
rect 17880 2508 17908 2536
rect 14936 2468 16574 2496
rect 17221 2499 17279 2505
rect 17221 2465 17233 2499
rect 17267 2496 17279 2499
rect 17402 2496 17408 2508
rect 17267 2468 17408 2496
rect 17267 2465 17279 2468
rect 17221 2459 17279 2465
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 17494 2456 17500 2508
rect 17552 2496 17558 2508
rect 17862 2496 17868 2508
rect 17552 2468 17597 2496
rect 17823 2468 17868 2496
rect 17552 2456 17558 2468
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 13538 2428 13544 2440
rect 9999 2400 10548 2428
rect 13499 2400 13544 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 13538 2388 13544 2400
rect 13596 2388 13602 2440
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 15068 2400 15117 2428
rect 15068 2388 15074 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 16482 2428 16488 2440
rect 15252 2400 16488 2428
rect 15252 2388 15258 2400
rect 16482 2388 16488 2400
rect 16540 2428 16546 2440
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 16540 2400 17325 2428
rect 16540 2388 16546 2400
rect 17313 2397 17325 2400
rect 17359 2397 17371 2431
rect 17512 2428 17540 2456
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17512 2400 18337 2428
rect 17313 2391 17371 2397
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 9214 2360 9220 2372
rect 8128 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 9876 2332 10149 2360
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9876 2292 9904 2332
rect 10137 2329 10149 2332
rect 10183 2360 10195 2363
rect 10597 2363 10655 2369
rect 10597 2360 10609 2363
rect 10183 2332 10609 2360
rect 10183 2329 10195 2332
rect 10137 2323 10195 2329
rect 10597 2329 10609 2332
rect 10643 2329 10655 2363
rect 10597 2323 10655 2329
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17678 2360 17684 2372
rect 16816 2332 17684 2360
rect 16816 2320 16822 2332
rect 17678 2320 17684 2332
rect 17736 2360 17742 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17736 2332 17969 2360
rect 17736 2320 17742 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 17957 2323 18015 2329
rect 10042 2292 10048 2304
rect 9088 2264 9904 2292
rect 10003 2264 10048 2292
rect 9088 2252 9094 2264
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 14918 2292 14924 2304
rect 14879 2264 14924 2292
rect 10505 2255 10563 2261
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 184 2202 18860 2224
rect 184 2150 1556 2202
rect 1608 2150 1620 2202
rect 1672 2150 1684 2202
rect 1736 2150 1748 2202
rect 1800 2150 1812 2202
rect 1864 2150 4656 2202
rect 4708 2150 4720 2202
rect 4772 2150 4784 2202
rect 4836 2150 4848 2202
rect 4900 2150 4912 2202
rect 4964 2150 7756 2202
rect 7808 2150 7820 2202
rect 7872 2150 7884 2202
rect 7936 2150 7948 2202
rect 8000 2150 8012 2202
rect 8064 2150 10856 2202
rect 10908 2150 10920 2202
rect 10972 2150 10984 2202
rect 11036 2150 11048 2202
rect 11100 2150 11112 2202
rect 11164 2150 13956 2202
rect 14008 2150 14020 2202
rect 14072 2150 14084 2202
rect 14136 2150 14148 2202
rect 14200 2150 14212 2202
rect 14264 2150 17056 2202
rect 17108 2150 17120 2202
rect 17172 2150 17184 2202
rect 17236 2150 17248 2202
rect 17300 2150 17312 2202
rect 17364 2150 18860 2202
rect 184 2128 18860 2150
rect 1946 2097 1952 2100
rect 1903 2091 1952 2097
rect 1903 2057 1915 2091
rect 1949 2057 1952 2091
rect 1903 2051 1952 2057
rect 1946 2048 1952 2051
rect 2004 2048 2010 2100
rect 2866 2088 2872 2100
rect 2827 2060 2872 2088
rect 2866 2048 2872 2060
rect 2924 2048 2930 2100
rect 5261 2091 5319 2097
rect 5261 2057 5273 2091
rect 5307 2088 5319 2091
rect 5626 2088 5632 2100
rect 5307 2060 5632 2088
rect 5307 2057 5319 2060
rect 5261 2051 5319 2057
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 6365 2091 6423 2097
rect 6365 2088 6377 2091
rect 5868 2060 6377 2088
rect 5868 2048 5874 2060
rect 6365 2057 6377 2060
rect 6411 2057 6423 2091
rect 6365 2051 6423 2057
rect 6917 2091 6975 2097
rect 6917 2057 6929 2091
rect 6963 2088 6975 2091
rect 7006 2088 7012 2100
rect 6963 2060 7012 2088
rect 6963 2057 6975 2060
rect 6917 2051 6975 2057
rect 7006 2048 7012 2060
rect 7064 2048 7070 2100
rect 9214 2088 9220 2100
rect 9175 2060 9220 2088
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 13725 2091 13783 2097
rect 13725 2088 13737 2091
rect 13004 2060 13737 2088
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 10229 2023 10287 2029
rect 10229 2020 10241 2023
rect 9824 1992 10241 2020
rect 9824 1980 9830 1992
rect 10229 1989 10241 1992
rect 10275 1989 10287 2023
rect 10229 1983 10287 1989
rect 12161 2023 12219 2029
rect 12161 1989 12173 2023
rect 12207 2020 12219 2023
rect 12802 2020 12808 2032
rect 12207 1992 12808 2020
rect 12207 1989 12219 1992
rect 12161 1983 12219 1989
rect 12802 1980 12808 1992
rect 12860 1980 12866 2032
rect 13004 2029 13032 2060
rect 13725 2057 13737 2060
rect 13771 2088 13783 2091
rect 14550 2088 14556 2100
rect 13771 2060 14556 2088
rect 13771 2057 13783 2060
rect 13725 2051 13783 2057
rect 14550 2048 14556 2060
rect 14608 2048 14614 2100
rect 15010 2048 15016 2100
rect 15068 2088 15074 2100
rect 15243 2091 15301 2097
rect 15243 2088 15255 2091
rect 15068 2060 15255 2088
rect 15068 2048 15074 2060
rect 15243 2057 15255 2060
rect 15289 2057 15301 2091
rect 15243 2051 15301 2057
rect 16117 2091 16175 2097
rect 16117 2057 16129 2091
rect 16163 2088 16175 2091
rect 16298 2088 16304 2100
rect 16163 2060 16304 2088
rect 16163 2057 16175 2060
rect 16117 2051 16175 2057
rect 16298 2048 16304 2060
rect 16356 2048 16362 2100
rect 12989 2023 13047 2029
rect 12989 1989 13001 2023
rect 13035 1989 13047 2023
rect 12989 1983 13047 1989
rect 2774 1912 2780 1964
rect 2832 1952 2838 1964
rect 3513 1955 3571 1961
rect 3513 1952 3525 1955
rect 2832 1924 3525 1952
rect 2832 1912 2838 1924
rect 3513 1921 3525 1924
rect 3559 1952 3571 1955
rect 4522 1952 4528 1964
rect 3559 1924 4528 1952
rect 3559 1921 3571 1924
rect 3513 1915 3571 1921
rect 4522 1912 4528 1924
rect 4580 1952 4586 1964
rect 5813 1955 5871 1961
rect 5813 1952 5825 1955
rect 4580 1924 5825 1952
rect 4580 1912 4586 1924
rect 5813 1921 5825 1924
rect 5859 1921 5871 1955
rect 5813 1915 5871 1921
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 7469 1955 7527 1961
rect 7469 1952 7481 1955
rect 6972 1924 7481 1952
rect 6972 1912 6978 1924
rect 7469 1921 7481 1924
rect 7515 1921 7527 1955
rect 7469 1915 7527 1921
rect 10505 1955 10563 1961
rect 10505 1921 10517 1955
rect 10551 1921 10563 1955
rect 10505 1915 10563 1921
rect 11885 1955 11943 1961
rect 11885 1921 11897 1955
rect 11931 1952 11943 1955
rect 12066 1952 12072 1964
rect 11931 1924 12072 1952
rect 11931 1921 11943 1924
rect 11885 1915 11943 1921
rect 2006 1887 2064 1893
rect 2006 1853 2018 1887
rect 2052 1884 2064 1887
rect 3602 1884 3608 1896
rect 2052 1856 3608 1884
rect 2052 1853 2064 1856
rect 2006 1847 2064 1853
rect 3602 1844 3608 1856
rect 3660 1884 3666 1896
rect 3970 1884 3976 1896
rect 3660 1856 3976 1884
rect 3660 1844 3666 1856
rect 3970 1844 3976 1856
rect 4028 1844 4034 1896
rect 4062 1844 4068 1896
rect 4120 1884 4126 1896
rect 4338 1884 4344 1896
rect 4120 1856 4344 1884
rect 4120 1844 4126 1856
rect 4338 1844 4344 1856
rect 4396 1844 4402 1896
rect 4801 1887 4859 1893
rect 4801 1853 4813 1887
rect 4847 1884 4859 1887
rect 5350 1884 5356 1896
rect 4847 1856 5356 1884
rect 4847 1853 4859 1856
rect 4801 1847 4859 1853
rect 5350 1844 5356 1856
rect 5408 1844 5414 1896
rect 7377 1887 7435 1893
rect 7377 1853 7389 1887
rect 7423 1884 7435 1887
rect 8294 1884 8300 1896
rect 7423 1856 8300 1884
rect 7423 1853 7435 1856
rect 7377 1847 7435 1853
rect 8294 1844 8300 1856
rect 8352 1844 8358 1896
rect 9030 1884 9036 1896
rect 8991 1856 9036 1884
rect 9030 1844 9036 1856
rect 9088 1884 9094 1896
rect 10520 1884 10548 1915
rect 12066 1912 12072 1924
rect 12124 1952 12130 1964
rect 13004 1952 13032 1983
rect 13814 1980 13820 2032
rect 13872 2020 13878 2032
rect 14185 2023 14243 2029
rect 14185 2020 14197 2023
rect 13872 1992 14197 2020
rect 13872 1980 13878 1992
rect 14185 1989 14197 1992
rect 14231 1989 14243 2023
rect 14185 1983 14243 1989
rect 12124 1924 13032 1952
rect 13541 1955 13599 1961
rect 12124 1912 12130 1924
rect 13541 1921 13553 1955
rect 13587 1952 13599 1955
rect 13630 1952 13636 1964
rect 13587 1924 13636 1952
rect 13587 1921 13599 1924
rect 13541 1915 13599 1921
rect 9088 1856 10548 1884
rect 9088 1844 9094 1856
rect 10594 1844 10600 1896
rect 10652 1884 10658 1896
rect 11793 1887 11851 1893
rect 10652 1856 10697 1884
rect 10652 1844 10658 1856
rect 11793 1853 11805 1887
rect 11839 1884 11851 1887
rect 12805 1887 12863 1893
rect 12805 1884 12817 1887
rect 11839 1856 12817 1884
rect 11839 1853 11851 1856
rect 11793 1847 11851 1853
rect 12805 1853 12817 1856
rect 12851 1884 12863 1887
rect 12986 1884 12992 1896
rect 12851 1856 12992 1884
rect 12851 1853 12863 1856
rect 12805 1847 12863 1853
rect 12986 1844 12992 1856
rect 13044 1844 13050 1896
rect 13081 1887 13139 1893
rect 13081 1853 13093 1887
rect 13127 1884 13139 1887
rect 13556 1884 13584 1915
rect 13630 1912 13636 1924
rect 13688 1912 13694 1964
rect 13127 1856 13584 1884
rect 13817 1887 13875 1893
rect 13127 1853 13139 1856
rect 13081 1847 13139 1853
rect 13817 1853 13829 1887
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 3326 1816 3332 1828
rect 3287 1788 3332 1816
rect 3326 1776 3332 1788
rect 3384 1776 3390 1828
rect 5721 1819 5779 1825
rect 5721 1785 5733 1819
rect 5767 1816 5779 1819
rect 5810 1816 5816 1828
rect 5767 1788 5816 1816
rect 5767 1785 5779 1788
rect 5721 1779 5779 1785
rect 5810 1776 5816 1788
rect 5868 1776 5874 1828
rect 13004 1816 13032 1844
rect 13832 1816 13860 1847
rect 13004 1788 13860 1816
rect 14200 1816 14228 1983
rect 14826 1980 14832 2032
rect 14884 2020 14890 2032
rect 15105 2023 15163 2029
rect 15105 2020 15117 2023
rect 14884 1992 15117 2020
rect 14884 1980 14890 1992
rect 15105 1989 15117 1992
rect 15151 1989 15163 2023
rect 15105 1983 15163 1989
rect 15194 1952 15200 1964
rect 14936 1924 15200 1952
rect 14936 1893 14964 1924
rect 15194 1912 15200 1924
rect 15252 1912 15258 1964
rect 16761 1955 16819 1961
rect 16761 1921 16773 1955
rect 16807 1952 16819 1955
rect 16850 1952 16856 1964
rect 16807 1924 16856 1952
rect 16807 1921 16819 1924
rect 16761 1915 16819 1921
rect 16850 1912 16856 1924
rect 16908 1912 16914 1964
rect 16942 1912 16948 1964
rect 17000 1952 17006 1964
rect 17681 1955 17739 1961
rect 17681 1952 17693 1955
rect 17000 1924 17693 1952
rect 17000 1912 17006 1924
rect 17681 1921 17693 1924
rect 17727 1921 17739 1955
rect 17681 1915 17739 1921
rect 14921 1887 14979 1893
rect 14921 1853 14933 1887
rect 14967 1853 14979 1887
rect 14921 1847 14979 1853
rect 15378 1844 15384 1896
rect 15436 1884 15442 1896
rect 15930 1884 15936 1896
rect 15436 1856 15481 1884
rect 15580 1856 15936 1884
rect 15436 1844 15442 1856
rect 15580 1816 15608 1856
rect 15930 1844 15936 1856
rect 15988 1884 15994 1896
rect 16577 1887 16635 1893
rect 16577 1884 16589 1887
rect 15988 1856 16589 1884
rect 15988 1844 15994 1856
rect 16577 1853 16589 1856
rect 16623 1853 16635 1887
rect 16577 1847 16635 1853
rect 17957 1887 18015 1893
rect 17957 1853 17969 1887
rect 18003 1884 18015 1887
rect 18003 1856 18460 1884
rect 18003 1853 18015 1856
rect 17957 1847 18015 1853
rect 14200 1788 15608 1816
rect 16206 1776 16212 1828
rect 16264 1816 16270 1828
rect 17402 1816 17408 1828
rect 16264 1788 17408 1816
rect 16264 1776 16270 1788
rect 17402 1776 17408 1788
rect 17460 1776 17466 1828
rect 18432 1760 18460 1856
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 3237 1751 3295 1757
rect 3237 1748 3249 1751
rect 3016 1720 3249 1748
rect 3016 1708 3022 1720
rect 3237 1717 3249 1720
rect 3283 1717 3295 1751
rect 4522 1748 4528 1760
rect 4483 1720 4528 1748
rect 3237 1711 3295 1717
rect 4522 1708 4528 1720
rect 4580 1708 4586 1760
rect 5626 1748 5632 1760
rect 5587 1720 5632 1748
rect 5626 1708 5632 1720
rect 5684 1708 5690 1760
rect 7282 1748 7288 1760
rect 7243 1720 7288 1748
rect 7282 1708 7288 1720
rect 7340 1708 7346 1760
rect 13078 1748 13084 1760
rect 13039 1720 13084 1748
rect 13078 1708 13084 1720
rect 13136 1708 13142 1760
rect 13538 1748 13544 1760
rect 13499 1720 13544 1748
rect 13538 1708 13544 1720
rect 13596 1708 13602 1760
rect 15010 1748 15016 1760
rect 14971 1720 15016 1748
rect 15010 1708 15016 1720
rect 15068 1708 15074 1760
rect 16482 1748 16488 1760
rect 16443 1720 16488 1748
rect 16482 1708 16488 1720
rect 16540 1708 16546 1760
rect 18414 1748 18420 1760
rect 18375 1720 18420 1748
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 184 1658 18920 1680
rect 184 1606 3106 1658
rect 3158 1606 3170 1658
rect 3222 1606 3234 1658
rect 3286 1606 3298 1658
rect 3350 1606 3362 1658
rect 3414 1606 6206 1658
rect 6258 1606 6270 1658
rect 6322 1606 6334 1658
rect 6386 1606 6398 1658
rect 6450 1606 6462 1658
rect 6514 1606 9306 1658
rect 9358 1606 9370 1658
rect 9422 1606 9434 1658
rect 9486 1606 9498 1658
rect 9550 1606 9562 1658
rect 9614 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 12534 1658
rect 12586 1606 12598 1658
rect 12650 1606 12662 1658
rect 12714 1606 15506 1658
rect 15558 1606 15570 1658
rect 15622 1606 15634 1658
rect 15686 1606 15698 1658
rect 15750 1606 15762 1658
rect 15814 1606 18606 1658
rect 18658 1606 18670 1658
rect 18722 1606 18734 1658
rect 18786 1606 18798 1658
rect 18850 1606 18862 1658
rect 18914 1606 18920 1658
rect 184 1584 18920 1606
rect 2958 1504 2964 1556
rect 3016 1544 3022 1556
rect 3145 1547 3203 1553
rect 3145 1544 3157 1547
rect 3016 1516 3157 1544
rect 3016 1504 3022 1516
rect 3145 1513 3157 1516
rect 3191 1513 3203 1547
rect 3145 1507 3203 1513
rect 5626 1504 5632 1556
rect 5684 1544 5690 1556
rect 5905 1547 5963 1553
rect 5905 1544 5917 1547
rect 5684 1516 5917 1544
rect 5684 1504 5690 1516
rect 5905 1513 5917 1516
rect 5951 1513 5963 1547
rect 5905 1507 5963 1513
rect 7282 1504 7288 1556
rect 7340 1544 7346 1556
rect 8021 1547 8079 1553
rect 8021 1544 8033 1547
rect 7340 1516 8033 1544
rect 7340 1504 7346 1516
rect 8021 1513 8033 1516
rect 8067 1513 8079 1547
rect 8021 1507 8079 1513
rect 8294 1504 8300 1556
rect 8352 1544 8358 1556
rect 8481 1547 8539 1553
rect 8481 1544 8493 1547
rect 8352 1516 8493 1544
rect 8352 1504 8358 1516
rect 8481 1513 8493 1516
rect 8527 1513 8539 1547
rect 8481 1507 8539 1513
rect 13449 1547 13507 1553
rect 13449 1513 13461 1547
rect 13495 1544 13507 1547
rect 13722 1544 13728 1556
rect 13495 1516 13728 1544
rect 13495 1513 13507 1516
rect 13449 1507 13507 1513
rect 13722 1504 13728 1516
rect 13780 1504 13786 1556
rect 15378 1504 15384 1556
rect 15436 1544 15442 1556
rect 15473 1547 15531 1553
rect 15473 1544 15485 1547
rect 15436 1516 15485 1544
rect 15436 1504 15442 1516
rect 15473 1513 15485 1516
rect 15519 1513 15531 1547
rect 15930 1544 15936 1556
rect 15891 1516 15936 1544
rect 15473 1507 15531 1513
rect 15930 1504 15936 1516
rect 15988 1504 15994 1556
rect 16761 1547 16819 1553
rect 16761 1513 16773 1547
rect 16807 1544 16819 1547
rect 16850 1544 16856 1556
rect 16807 1516 16856 1544
rect 16807 1513 16819 1516
rect 16761 1507 16819 1513
rect 16850 1504 16856 1516
rect 16908 1504 16914 1556
rect 3789 1479 3847 1485
rect 3789 1476 3801 1479
rect 3436 1448 3801 1476
rect 3436 1417 3464 1448
rect 3789 1445 3801 1448
rect 3835 1445 3847 1479
rect 3789 1439 3847 1445
rect 4080 1448 4660 1476
rect 3420 1411 3478 1417
rect 3420 1377 3432 1411
rect 3466 1377 3478 1411
rect 3420 1371 3478 1377
rect 3513 1411 3571 1417
rect 3513 1377 3525 1411
rect 3559 1377 3571 1411
rect 3970 1408 3976 1420
rect 3931 1380 3976 1408
rect 3513 1371 3571 1377
rect 3528 1272 3556 1371
rect 3970 1368 3976 1380
rect 4028 1368 4034 1420
rect 4080 1417 4108 1448
rect 4065 1411 4123 1417
rect 4065 1377 4077 1411
rect 4111 1377 4123 1411
rect 4338 1408 4344 1420
rect 4299 1380 4344 1408
rect 4065 1371 4123 1377
rect 4338 1368 4344 1380
rect 4396 1368 4402 1420
rect 4632 1417 4660 1448
rect 14918 1436 14924 1488
rect 14976 1476 14982 1488
rect 14976 1448 15148 1476
rect 14976 1436 14982 1448
rect 4617 1411 4675 1417
rect 4617 1377 4629 1411
rect 4663 1408 4675 1411
rect 5350 1408 5356 1420
rect 4663 1380 5356 1408
rect 4663 1377 4675 1380
rect 4617 1371 4675 1377
rect 5350 1368 5356 1380
rect 5408 1408 5414 1420
rect 5537 1411 5595 1417
rect 5537 1408 5549 1411
rect 5408 1380 5549 1408
rect 5408 1368 5414 1380
rect 5537 1377 5549 1380
rect 5583 1377 5595 1411
rect 5537 1371 5595 1377
rect 8389 1411 8447 1417
rect 8389 1377 8401 1411
rect 8435 1408 8447 1411
rect 8435 1380 9352 1408
rect 8435 1377 8447 1380
rect 8389 1371 8447 1377
rect 3789 1343 3847 1349
rect 3789 1309 3801 1343
rect 3835 1340 3847 1343
rect 4356 1340 4384 1368
rect 3835 1312 4384 1340
rect 5445 1343 5503 1349
rect 3835 1309 3847 1312
rect 3789 1303 3847 1309
rect 5445 1309 5457 1343
rect 5491 1309 5503 1343
rect 8662 1340 8668 1352
rect 8623 1312 8668 1340
rect 5445 1303 5503 1309
rect 4341 1275 4399 1281
rect 4341 1272 4353 1275
rect 3528 1244 4353 1272
rect 4341 1241 4353 1244
rect 4387 1241 4399 1275
rect 4341 1235 4399 1241
rect 4433 1275 4491 1281
rect 4433 1241 4445 1275
rect 4479 1272 4491 1275
rect 5460 1272 5488 1303
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 9324 1340 9352 1380
rect 10042 1368 10048 1420
rect 10100 1408 10106 1420
rect 10167 1411 10225 1417
rect 10167 1408 10179 1411
rect 10100 1380 10179 1408
rect 10100 1368 10106 1380
rect 10167 1377 10179 1380
rect 10213 1377 10225 1411
rect 10167 1371 10225 1377
rect 10318 1368 10324 1420
rect 10376 1408 10382 1420
rect 13078 1408 13084 1420
rect 10376 1380 10421 1408
rect 13039 1380 13084 1408
rect 10376 1368 10382 1380
rect 13078 1368 13084 1380
rect 13136 1368 13142 1420
rect 13235 1411 13293 1417
rect 13235 1377 13247 1411
rect 13281 1408 13293 1411
rect 13538 1408 13544 1420
rect 13281 1380 13544 1408
rect 13281 1377 13293 1380
rect 13235 1371 13293 1377
rect 13538 1368 13544 1380
rect 13596 1368 13602 1420
rect 15010 1408 15016 1420
rect 14971 1380 15016 1408
rect 15010 1368 15016 1380
rect 15068 1368 15074 1420
rect 15120 1417 15148 1448
rect 16482 1436 16488 1488
rect 16540 1476 16546 1488
rect 16540 1436 16574 1476
rect 15105 1411 15163 1417
rect 15105 1377 15117 1411
rect 15151 1377 15163 1411
rect 15105 1371 15163 1377
rect 16390 1368 16396 1420
rect 16448 1368 16454 1420
rect 16546 1408 16574 1436
rect 16546 1380 16620 1408
rect 9953 1343 10011 1349
rect 9953 1340 9965 1343
rect 9324 1312 9965 1340
rect 9953 1309 9965 1312
rect 9999 1309 10011 1343
rect 14734 1340 14740 1352
rect 14695 1312 14740 1340
rect 9953 1303 10011 1309
rect 14734 1300 14740 1312
rect 14792 1300 14798 1352
rect 16408 1340 16436 1368
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 16408 1312 16497 1340
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16592 1340 16620 1380
rect 16758 1368 16764 1420
rect 16816 1408 16822 1420
rect 16816 1380 16861 1408
rect 16816 1368 16822 1380
rect 17402 1368 17408 1420
rect 17460 1408 17466 1420
rect 17497 1411 17555 1417
rect 17497 1408 17509 1411
rect 17460 1380 17509 1408
rect 17460 1368 17466 1380
rect 17497 1377 17509 1380
rect 17543 1377 17555 1411
rect 17497 1371 17555 1377
rect 17589 1343 17647 1349
rect 16592 1312 17172 1340
rect 16485 1303 16543 1309
rect 17144 1281 17172 1312
rect 17589 1309 17601 1343
rect 17635 1340 17647 1343
rect 17862 1340 17868 1352
rect 17635 1312 17868 1340
rect 17635 1309 17647 1312
rect 17589 1303 17647 1309
rect 17862 1300 17868 1312
rect 17920 1300 17926 1352
rect 4479 1244 5488 1272
rect 16669 1275 16727 1281
rect 4479 1241 4491 1244
rect 4433 1235 4491 1241
rect 16669 1241 16681 1275
rect 16715 1241 16727 1275
rect 16669 1235 16727 1241
rect 17129 1275 17187 1281
rect 17129 1241 17141 1275
rect 17175 1241 17187 1275
rect 17129 1235 17187 1241
rect 3970 1164 3976 1216
rect 4028 1204 4034 1216
rect 4448 1204 4476 1235
rect 4028 1176 4476 1204
rect 16684 1204 16712 1235
rect 17402 1204 17408 1216
rect 16684 1176 17408 1204
rect 4028 1164 4034 1176
rect 17402 1164 17408 1176
rect 17460 1164 17466 1216
rect 184 1114 18860 1136
rect 184 1062 1556 1114
rect 1608 1062 1620 1114
rect 1672 1062 1684 1114
rect 1736 1062 1748 1114
rect 1800 1062 1812 1114
rect 1864 1062 4656 1114
rect 4708 1062 4720 1114
rect 4772 1062 4784 1114
rect 4836 1062 4848 1114
rect 4900 1062 4912 1114
rect 4964 1062 7756 1114
rect 7808 1062 7820 1114
rect 7872 1062 7884 1114
rect 7936 1062 7948 1114
rect 8000 1062 8012 1114
rect 8064 1062 10856 1114
rect 10908 1062 10920 1114
rect 10972 1062 10984 1114
rect 11036 1062 11048 1114
rect 11100 1062 11112 1114
rect 11164 1062 13956 1114
rect 14008 1062 14020 1114
rect 14072 1062 14084 1114
rect 14136 1062 14148 1114
rect 14200 1062 14212 1114
rect 14264 1062 17056 1114
rect 17108 1062 17120 1114
rect 17172 1062 17184 1114
rect 17236 1062 17248 1114
rect 17300 1062 17312 1114
rect 17364 1062 18860 1114
rect 184 1040 18860 1062
rect 184 570 18920 592
rect 184 518 3106 570
rect 3158 518 3170 570
rect 3222 518 3234 570
rect 3286 518 3298 570
rect 3350 518 3362 570
rect 3414 518 6206 570
rect 6258 518 6270 570
rect 6322 518 6334 570
rect 6386 518 6398 570
rect 6450 518 6462 570
rect 6514 518 9306 570
rect 9358 518 9370 570
rect 9422 518 9434 570
rect 9486 518 9498 570
rect 9550 518 9562 570
rect 9614 518 12406 570
rect 12458 518 12470 570
rect 12522 518 12534 570
rect 12586 518 12598 570
rect 12650 518 12662 570
rect 12714 518 15506 570
rect 15558 518 15570 570
rect 15622 518 15634 570
rect 15686 518 15698 570
rect 15750 518 15762 570
rect 15814 518 18606 570
rect 18658 518 18670 570
rect 18722 518 18734 570
rect 18786 518 18798 570
rect 18850 518 18862 570
rect 18914 518 18920 570
rect 184 496 18920 518
<< via1 >>
rect 1556 18470 1608 18522
rect 1620 18470 1672 18522
rect 1684 18470 1736 18522
rect 1748 18470 1800 18522
rect 1812 18470 1864 18522
rect 4656 18470 4708 18522
rect 4720 18470 4772 18522
rect 4784 18470 4836 18522
rect 4848 18470 4900 18522
rect 4912 18470 4964 18522
rect 7756 18470 7808 18522
rect 7820 18470 7872 18522
rect 7884 18470 7936 18522
rect 7948 18470 8000 18522
rect 8012 18470 8064 18522
rect 10856 18470 10908 18522
rect 10920 18470 10972 18522
rect 10984 18470 11036 18522
rect 11048 18470 11100 18522
rect 11112 18470 11164 18522
rect 13956 18470 14008 18522
rect 14020 18470 14072 18522
rect 14084 18470 14136 18522
rect 14148 18470 14200 18522
rect 14212 18470 14264 18522
rect 17056 18470 17108 18522
rect 17120 18470 17172 18522
rect 17184 18470 17236 18522
rect 17248 18470 17300 18522
rect 17312 18470 17364 18522
rect 4252 18368 4304 18420
rect 4344 18368 4396 18420
rect 18420 18411 18472 18420
rect 18420 18377 18429 18411
rect 18429 18377 18463 18411
rect 18463 18377 18472 18411
rect 18420 18368 18472 18377
rect 6000 18300 6052 18352
rect 1400 18164 1452 18216
rect 8668 18232 8720 18284
rect 10508 18275 10560 18284
rect 10508 18241 10517 18275
rect 10517 18241 10551 18275
rect 10551 18241 10560 18275
rect 10508 18232 10560 18241
rect 14648 18232 14700 18284
rect 8208 18207 8260 18216
rect 5448 18096 5500 18148
rect 5724 18139 5776 18148
rect 5724 18105 5733 18139
rect 5733 18105 5767 18139
rect 5767 18105 5776 18139
rect 5724 18096 5776 18105
rect 7840 18139 7892 18148
rect 7840 18105 7849 18139
rect 7849 18105 7883 18139
rect 7883 18105 7892 18139
rect 7840 18096 7892 18105
rect 8208 18173 8217 18207
rect 8217 18173 8251 18207
rect 8251 18173 8260 18207
rect 8208 18164 8260 18173
rect 8392 18164 8444 18216
rect 9680 18164 9732 18216
rect 12900 18164 12952 18216
rect 13452 18164 13504 18216
rect 16120 18164 16172 18216
rect 18420 18164 18472 18216
rect 8116 18096 8168 18148
rect 13820 18096 13872 18148
rect 14924 18096 14976 18148
rect 4988 18028 5040 18080
rect 8300 18028 8352 18080
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 14832 18028 14884 18080
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 15200 18028 15252 18080
rect 15384 18028 15436 18080
rect 3106 17926 3158 17978
rect 3170 17926 3222 17978
rect 3234 17926 3286 17978
rect 3298 17926 3350 17978
rect 3362 17926 3414 17978
rect 6206 17926 6258 17978
rect 6270 17926 6322 17978
rect 6334 17926 6386 17978
rect 6398 17926 6450 17978
rect 6462 17926 6514 17978
rect 9306 17926 9358 17978
rect 9370 17926 9422 17978
rect 9434 17926 9486 17978
rect 9498 17926 9550 17978
rect 9562 17926 9614 17978
rect 12406 17926 12458 17978
rect 12470 17926 12522 17978
rect 12534 17926 12586 17978
rect 12598 17926 12650 17978
rect 12662 17926 12714 17978
rect 15506 17926 15558 17978
rect 15570 17926 15622 17978
rect 15634 17926 15686 17978
rect 15698 17926 15750 17978
rect 15762 17926 15814 17978
rect 18606 17926 18658 17978
rect 18670 17926 18722 17978
rect 18734 17926 18786 17978
rect 18798 17926 18850 17978
rect 18862 17926 18914 17978
rect 9680 17824 9732 17876
rect 4252 17756 4304 17808
rect 8668 17756 8720 17808
rect 16856 17756 16908 17808
rect 1952 17688 2004 17740
rect 2412 17688 2464 17740
rect 5172 17688 5224 17740
rect 4344 17552 4396 17604
rect 5356 17552 5408 17604
rect 7840 17688 7892 17740
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 14924 17688 14976 17740
rect 8300 17620 8352 17672
rect 9220 17620 9272 17672
rect 12808 17620 12860 17672
rect 16672 17620 16724 17672
rect 2872 17484 2924 17536
rect 5264 17484 5316 17536
rect 9680 17484 9732 17536
rect 17500 17484 17552 17536
rect 1556 17382 1608 17434
rect 1620 17382 1672 17434
rect 1684 17382 1736 17434
rect 1748 17382 1800 17434
rect 1812 17382 1864 17434
rect 4656 17382 4708 17434
rect 4720 17382 4772 17434
rect 4784 17382 4836 17434
rect 4848 17382 4900 17434
rect 4912 17382 4964 17434
rect 7756 17382 7808 17434
rect 7820 17382 7872 17434
rect 7884 17382 7936 17434
rect 7948 17382 8000 17434
rect 8012 17382 8064 17434
rect 10856 17382 10908 17434
rect 10920 17382 10972 17434
rect 10984 17382 11036 17434
rect 11048 17382 11100 17434
rect 11112 17382 11164 17434
rect 13956 17382 14008 17434
rect 14020 17382 14072 17434
rect 14084 17382 14136 17434
rect 14148 17382 14200 17434
rect 14212 17382 14264 17434
rect 17056 17382 17108 17434
rect 17120 17382 17172 17434
rect 17184 17382 17236 17434
rect 17248 17382 17300 17434
rect 17312 17382 17364 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2688 17280 2740 17332
rect 1952 17144 2004 17196
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 4436 17280 4488 17332
rect 5724 17280 5776 17332
rect 4436 17119 4488 17128
rect 4436 17085 4445 17119
rect 4445 17085 4479 17119
rect 4479 17085 4488 17119
rect 4436 17076 4488 17085
rect 5080 17008 5132 17060
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 6000 17119 6052 17128
rect 5264 17076 5316 17085
rect 6000 17085 6009 17119
rect 6009 17085 6043 17119
rect 6043 17085 6052 17119
rect 6000 17076 6052 17085
rect 7472 17144 7524 17196
rect 12532 17212 12584 17264
rect 8024 17008 8076 17060
rect 9036 17051 9088 17060
rect 9036 17017 9045 17051
rect 9045 17017 9079 17051
rect 9079 17017 9088 17051
rect 9036 17008 9088 17017
rect 10600 17051 10652 17060
rect 10600 17017 10609 17051
rect 10609 17017 10643 17051
rect 10643 17017 10652 17051
rect 10600 17008 10652 17017
rect 12164 17144 12216 17196
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 12164 17008 12216 17060
rect 14280 17144 14332 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 12808 17119 12860 17128
rect 12808 17085 12821 17119
rect 12821 17085 12860 17119
rect 12808 17076 12860 17085
rect 13452 17076 13504 17128
rect 13636 17076 13688 17128
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 14740 17008 14792 17060
rect 16488 17008 16540 17060
rect 1124 16983 1176 16992
rect 1124 16949 1133 16983
rect 1133 16949 1167 16983
rect 1167 16949 1176 16983
rect 1124 16940 1176 16949
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 2596 16940 2648 16992
rect 2780 16940 2832 16992
rect 4528 16940 4580 16992
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 8760 16940 8812 16992
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 12532 16940 12584 16992
rect 13084 16940 13136 16992
rect 13636 16940 13688 16992
rect 14464 16940 14516 16992
rect 3106 16838 3158 16890
rect 3170 16838 3222 16890
rect 3234 16838 3286 16890
rect 3298 16838 3350 16890
rect 3362 16838 3414 16890
rect 6206 16838 6258 16890
rect 6270 16838 6322 16890
rect 6334 16838 6386 16890
rect 6398 16838 6450 16890
rect 6462 16838 6514 16890
rect 9306 16838 9358 16890
rect 9370 16838 9422 16890
rect 9434 16838 9486 16890
rect 9498 16838 9550 16890
rect 9562 16838 9614 16890
rect 12406 16838 12458 16890
rect 12470 16838 12522 16890
rect 12534 16838 12586 16890
rect 12598 16838 12650 16890
rect 12662 16838 12714 16890
rect 15506 16838 15558 16890
rect 15570 16838 15622 16890
rect 15634 16838 15686 16890
rect 15698 16838 15750 16890
rect 15762 16838 15814 16890
rect 18606 16838 18658 16890
rect 18670 16838 18722 16890
rect 18734 16838 18786 16890
rect 18798 16838 18850 16890
rect 18862 16838 18914 16890
rect 2964 16736 3016 16788
rect 4436 16736 4488 16788
rect 5080 16736 5132 16788
rect 5724 16736 5776 16788
rect 8392 16736 8444 16788
rect 12808 16736 12860 16788
rect 3792 16668 3844 16720
rect 5172 16668 5224 16720
rect 8116 16668 8168 16720
rect 9956 16711 10008 16720
rect 9956 16677 9965 16711
rect 9965 16677 9999 16711
rect 9999 16677 10008 16711
rect 9956 16668 10008 16677
rect 12072 16668 12124 16720
rect 10048 16600 10100 16652
rect 12256 16600 12308 16652
rect 12900 16643 12952 16652
rect 2872 16532 2924 16584
rect 9128 16575 9180 16584
rect 4436 16396 4488 16448
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 12900 16609 12909 16643
rect 12909 16609 12943 16643
rect 12943 16609 12952 16643
rect 12900 16600 12952 16609
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 9864 16464 9916 16516
rect 14464 16600 14516 16652
rect 14832 16736 14884 16788
rect 15200 16736 15252 16788
rect 16672 16736 16724 16788
rect 15200 16600 15252 16652
rect 14740 16532 14792 16584
rect 14924 16532 14976 16584
rect 15384 16600 15436 16652
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 6828 16396 6880 16448
rect 12164 16396 12216 16448
rect 12808 16396 12860 16448
rect 13452 16396 13504 16448
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 14372 16396 14424 16448
rect 1556 16294 1608 16346
rect 1620 16294 1672 16346
rect 1684 16294 1736 16346
rect 1748 16294 1800 16346
rect 1812 16294 1864 16346
rect 4656 16294 4708 16346
rect 4720 16294 4772 16346
rect 4784 16294 4836 16346
rect 4848 16294 4900 16346
rect 4912 16294 4964 16346
rect 7756 16294 7808 16346
rect 7820 16294 7872 16346
rect 7884 16294 7936 16346
rect 7948 16294 8000 16346
rect 8012 16294 8064 16346
rect 10856 16294 10908 16346
rect 10920 16294 10972 16346
rect 10984 16294 11036 16346
rect 11048 16294 11100 16346
rect 11112 16294 11164 16346
rect 13956 16294 14008 16346
rect 14020 16294 14072 16346
rect 14084 16294 14136 16346
rect 14148 16294 14200 16346
rect 14212 16294 14264 16346
rect 17056 16294 17108 16346
rect 17120 16294 17172 16346
rect 17184 16294 17236 16346
rect 17248 16294 17300 16346
rect 17312 16294 17364 16346
rect 5724 16192 5776 16244
rect 9036 16192 9088 16244
rect 9128 16192 9180 16244
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 10324 16192 10376 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 1400 16124 1452 16176
rect 2136 16056 2188 16108
rect 2504 16056 2556 16108
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 7288 16056 7340 16108
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 940 15988 992 16040
rect 1952 15988 2004 16040
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 4528 15988 4580 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7196 15988 7248 16040
rect 16304 16031 16356 16040
rect 2044 15920 2096 15972
rect 8208 15920 8260 15972
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 2320 15895 2372 15904
rect 1952 15852 2004 15861
rect 2320 15861 2329 15895
rect 2329 15861 2363 15895
rect 2363 15861 2372 15895
rect 2320 15852 2372 15861
rect 7012 15852 7064 15904
rect 9864 15852 9916 15904
rect 10600 15852 10652 15904
rect 15016 15920 15068 15972
rect 16856 15920 16908 15972
rect 17684 15852 17736 15904
rect 3106 15750 3158 15802
rect 3170 15750 3222 15802
rect 3234 15750 3286 15802
rect 3298 15750 3350 15802
rect 3362 15750 3414 15802
rect 6206 15750 6258 15802
rect 6270 15750 6322 15802
rect 6334 15750 6386 15802
rect 6398 15750 6450 15802
rect 6462 15750 6514 15802
rect 9306 15750 9358 15802
rect 9370 15750 9422 15802
rect 9434 15750 9486 15802
rect 9498 15750 9550 15802
rect 9562 15750 9614 15802
rect 12406 15750 12458 15802
rect 12470 15750 12522 15802
rect 12534 15750 12586 15802
rect 12598 15750 12650 15802
rect 12662 15750 12714 15802
rect 15506 15750 15558 15802
rect 15570 15750 15622 15802
rect 15634 15750 15686 15802
rect 15698 15750 15750 15802
rect 15762 15750 15814 15802
rect 18606 15750 18658 15802
rect 18670 15750 18722 15802
rect 18734 15750 18786 15802
rect 18798 15750 18850 15802
rect 18862 15750 18914 15802
rect 1124 15648 1176 15700
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 7196 15648 7248 15700
rect 8208 15648 8260 15700
rect 11704 15648 11756 15700
rect 12808 15648 12860 15700
rect 13360 15648 13412 15700
rect 14280 15648 14332 15700
rect 16304 15648 16356 15700
rect 9680 15580 9732 15632
rect 940 15555 992 15564
rect 940 15521 949 15555
rect 949 15521 983 15555
rect 983 15521 992 15555
rect 940 15512 992 15521
rect 2872 15512 2924 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10324 15555 10376 15564
rect 10048 15512 10100 15521
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 12072 15512 12124 15564
rect 12164 15512 12216 15564
rect 12900 15555 12952 15564
rect 12900 15521 12905 15555
rect 12905 15521 12939 15555
rect 12939 15521 12952 15555
rect 12900 15512 12952 15521
rect 11336 15444 11388 15496
rect 14740 15512 14792 15564
rect 16304 15512 16356 15564
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 11520 15376 11572 15428
rect 11612 15376 11664 15428
rect 14280 15444 14332 15496
rect 17684 15444 17736 15496
rect 17868 15444 17920 15496
rect 16580 15376 16632 15428
rect 1308 15308 1360 15360
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 15016 15308 15068 15360
rect 1556 15206 1608 15258
rect 1620 15206 1672 15258
rect 1684 15206 1736 15258
rect 1748 15206 1800 15258
rect 1812 15206 1864 15258
rect 4656 15206 4708 15258
rect 4720 15206 4772 15258
rect 4784 15206 4836 15258
rect 4848 15206 4900 15258
rect 4912 15206 4964 15258
rect 7756 15206 7808 15258
rect 7820 15206 7872 15258
rect 7884 15206 7936 15258
rect 7948 15206 8000 15258
rect 8012 15206 8064 15258
rect 10856 15206 10908 15258
rect 10920 15206 10972 15258
rect 10984 15206 11036 15258
rect 11048 15206 11100 15258
rect 11112 15206 11164 15258
rect 13956 15206 14008 15258
rect 14020 15206 14072 15258
rect 14084 15206 14136 15258
rect 14148 15206 14200 15258
rect 14212 15206 14264 15258
rect 17056 15206 17108 15258
rect 17120 15206 17172 15258
rect 17184 15206 17236 15258
rect 17248 15206 17300 15258
rect 17312 15206 17364 15258
rect 2044 15104 2096 15156
rect 2688 15104 2740 15156
rect 9220 15104 9272 15156
rect 10048 15104 10100 15156
rect 11336 15104 11388 15156
rect 16488 15104 16540 15156
rect 16948 15104 17000 15156
rect 17868 15104 17920 15156
rect 2044 14968 2096 15020
rect 4436 14968 4488 15020
rect 10324 15036 10376 15088
rect 3976 14943 4028 14952
rect 3976 14909 3985 14943
rect 3985 14909 4019 14943
rect 4019 14909 4028 14943
rect 3976 14900 4028 14909
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 4988 14900 5040 14952
rect 5724 14900 5776 14952
rect 2320 14832 2372 14884
rect 3792 14832 3844 14884
rect 6920 14832 6972 14884
rect 10508 14968 10560 15020
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 12256 15036 12308 15088
rect 8116 14832 8168 14884
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 10324 14900 10376 14909
rect 11244 14900 11296 14952
rect 12164 14900 12216 14952
rect 11796 14832 11848 14884
rect 12900 14900 12952 14952
rect 14004 14968 14056 15020
rect 14924 14968 14976 15020
rect 16764 14968 16816 15020
rect 14372 14900 14424 14952
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 4528 14764 4580 14816
rect 5540 14764 5592 14816
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 9772 14764 9824 14816
rect 10324 14764 10376 14816
rect 12900 14764 12952 14816
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14464 14764 14516 14816
rect 14740 14832 14792 14884
rect 15844 14900 15896 14952
rect 16580 14900 16632 14952
rect 16856 14832 16908 14884
rect 15384 14764 15436 14816
rect 18052 14764 18104 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 19064 14764 19116 14816
rect 3106 14662 3158 14714
rect 3170 14662 3222 14714
rect 3234 14662 3286 14714
rect 3298 14662 3350 14714
rect 3362 14662 3414 14714
rect 6206 14662 6258 14714
rect 6270 14662 6322 14714
rect 6334 14662 6386 14714
rect 6398 14662 6450 14714
rect 6462 14662 6514 14714
rect 9306 14662 9358 14714
rect 9370 14662 9422 14714
rect 9434 14662 9486 14714
rect 9498 14662 9550 14714
rect 9562 14662 9614 14714
rect 12406 14662 12458 14714
rect 12470 14662 12522 14714
rect 12534 14662 12586 14714
rect 12598 14662 12650 14714
rect 12662 14662 12714 14714
rect 15506 14662 15558 14714
rect 15570 14662 15622 14714
rect 15634 14662 15686 14714
rect 15698 14662 15750 14714
rect 15762 14662 15814 14714
rect 18606 14662 18658 14714
rect 18670 14662 18722 14714
rect 18734 14662 18786 14714
rect 18798 14662 18850 14714
rect 18862 14662 18914 14714
rect 4160 14560 4212 14612
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 940 14492 992 14544
rect 1216 14467 1268 14476
rect 1216 14433 1225 14467
rect 1225 14433 1259 14467
rect 1259 14433 1268 14467
rect 1216 14424 1268 14433
rect 2780 14492 2832 14544
rect 5540 14535 5592 14544
rect 5540 14501 5549 14535
rect 5549 14501 5583 14535
rect 5583 14501 5592 14535
rect 5540 14492 5592 14501
rect 5816 14492 5868 14544
rect 8116 14492 8168 14544
rect 16948 14560 17000 14612
rect 12624 14535 12676 14544
rect 4436 14424 4488 14476
rect 2136 14356 2188 14408
rect 2964 14356 3016 14408
rect 3516 14356 3568 14408
rect 8300 14399 8352 14408
rect 3608 14288 3660 14340
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 10048 14424 10100 14476
rect 11244 14424 11296 14476
rect 12624 14501 12633 14535
rect 12633 14501 12667 14535
rect 12667 14501 12676 14535
rect 12624 14492 12676 14501
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13544 14424 13596 14476
rect 2136 14220 2188 14272
rect 10140 14288 10192 14340
rect 12900 14356 12952 14408
rect 13452 14356 13504 14408
rect 14004 14399 14056 14408
rect 14004 14365 14013 14399
rect 14013 14365 14047 14399
rect 14047 14365 14056 14399
rect 14004 14356 14056 14365
rect 16028 14492 16080 14544
rect 16856 14492 16908 14544
rect 14464 14424 14516 14476
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 17776 14424 17828 14476
rect 18052 14467 18104 14476
rect 18052 14433 18061 14467
rect 18061 14433 18095 14467
rect 18095 14433 18104 14467
rect 18052 14424 18104 14433
rect 16028 14356 16080 14408
rect 17960 14356 18012 14408
rect 9772 14220 9824 14272
rect 13728 14288 13780 14340
rect 15384 14288 15436 14340
rect 16856 14288 16908 14340
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 13820 14220 13872 14272
rect 16120 14220 16172 14272
rect 17684 14220 17736 14272
rect 18144 14263 18196 14272
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 1556 14118 1608 14170
rect 1620 14118 1672 14170
rect 1684 14118 1736 14170
rect 1748 14118 1800 14170
rect 1812 14118 1864 14170
rect 4656 14118 4708 14170
rect 4720 14118 4772 14170
rect 4784 14118 4836 14170
rect 4848 14118 4900 14170
rect 4912 14118 4964 14170
rect 7756 14118 7808 14170
rect 7820 14118 7872 14170
rect 7884 14118 7936 14170
rect 7948 14118 8000 14170
rect 8012 14118 8064 14170
rect 10856 14118 10908 14170
rect 10920 14118 10972 14170
rect 10984 14118 11036 14170
rect 11048 14118 11100 14170
rect 11112 14118 11164 14170
rect 13956 14118 14008 14170
rect 14020 14118 14072 14170
rect 14084 14118 14136 14170
rect 14148 14118 14200 14170
rect 14212 14118 14264 14170
rect 17056 14118 17108 14170
rect 17120 14118 17172 14170
rect 17184 14118 17236 14170
rect 17248 14118 17300 14170
rect 17312 14118 17364 14170
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 3608 14016 3660 14068
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 4436 13880 4488 13932
rect 2044 13812 2096 13864
rect 4528 13855 4580 13864
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 6920 14016 6972 14068
rect 8300 14016 8352 14068
rect 12900 14016 12952 14068
rect 13636 13948 13688 14000
rect 15844 14016 15896 14068
rect 17960 14059 18012 14068
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 7288 13880 7340 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 11336 13880 11388 13932
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14740 13880 14792 13932
rect 18236 13948 18288 14000
rect 15108 13880 15160 13932
rect 7104 13812 7156 13864
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 10048 13812 10100 13864
rect 14372 13812 14424 13864
rect 14924 13812 14976 13864
rect 3792 13744 3844 13796
rect 5816 13744 5868 13796
rect 12624 13744 12676 13796
rect 15384 13880 15436 13932
rect 16580 13880 16632 13932
rect 16764 13744 16816 13796
rect 16948 13744 17000 13796
rect 12164 13676 12216 13728
rect 16856 13676 16908 13728
rect 3106 13574 3158 13626
rect 3170 13574 3222 13626
rect 3234 13574 3286 13626
rect 3298 13574 3350 13626
rect 3362 13574 3414 13626
rect 6206 13574 6258 13626
rect 6270 13574 6322 13626
rect 6334 13574 6386 13626
rect 6398 13574 6450 13626
rect 6462 13574 6514 13626
rect 9306 13574 9358 13626
rect 9370 13574 9422 13626
rect 9434 13574 9486 13626
rect 9498 13574 9550 13626
rect 9562 13574 9614 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 12534 13574 12586 13626
rect 12598 13574 12650 13626
rect 12662 13574 12714 13626
rect 15506 13574 15558 13626
rect 15570 13574 15622 13626
rect 15634 13574 15686 13626
rect 15698 13574 15750 13626
rect 15762 13574 15814 13626
rect 18606 13574 18658 13626
rect 18670 13574 18722 13626
rect 18734 13574 18786 13626
rect 18798 13574 18850 13626
rect 18862 13574 18914 13626
rect 1216 13472 1268 13524
rect 1308 13472 1360 13524
rect 3976 13472 4028 13524
rect 9128 13472 9180 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 5356 13404 5408 13456
rect 9864 13404 9916 13456
rect 2964 13336 3016 13388
rect 1400 13268 1452 13320
rect 3608 13311 3660 13320
rect 3608 13277 3617 13311
rect 3617 13277 3651 13311
rect 3651 13277 3660 13311
rect 3608 13268 3660 13277
rect 4436 13336 4488 13388
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 7288 13336 7340 13388
rect 13636 13472 13688 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 12072 13404 12124 13456
rect 13452 13404 13504 13456
rect 15016 13447 15068 13456
rect 15016 13413 15025 13447
rect 15025 13413 15059 13447
rect 15059 13413 15068 13447
rect 15016 13404 15068 13413
rect 16764 13404 16816 13456
rect 9680 13268 9732 13320
rect 11520 13336 11572 13388
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 13268 13336 13320 13388
rect 14556 13336 14608 13388
rect 14924 13336 14976 13388
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 11428 13268 11480 13320
rect 13544 13200 13596 13252
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 10508 13132 10560 13184
rect 10784 13132 10836 13184
rect 1556 13030 1608 13082
rect 1620 13030 1672 13082
rect 1684 13030 1736 13082
rect 1748 13030 1800 13082
rect 1812 13030 1864 13082
rect 4656 13030 4708 13082
rect 4720 13030 4772 13082
rect 4784 13030 4836 13082
rect 4848 13030 4900 13082
rect 4912 13030 4964 13082
rect 7756 13030 7808 13082
rect 7820 13030 7872 13082
rect 7884 13030 7936 13082
rect 7948 13030 8000 13082
rect 8012 13030 8064 13082
rect 10856 13030 10908 13082
rect 10920 13030 10972 13082
rect 10984 13030 11036 13082
rect 11048 13030 11100 13082
rect 11112 13030 11164 13082
rect 13956 13030 14008 13082
rect 14020 13030 14072 13082
rect 14084 13030 14136 13082
rect 14148 13030 14200 13082
rect 14212 13030 14264 13082
rect 17056 13030 17108 13082
rect 17120 13030 17172 13082
rect 17184 13030 17236 13082
rect 17248 13030 17300 13082
rect 17312 13030 17364 13082
rect 4436 12928 4488 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 12808 12928 12860 12980
rect 10508 12860 10560 12912
rect 16304 12903 16356 12912
rect 8760 12792 8812 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10140 12792 10192 12844
rect 16304 12869 16313 12903
rect 16313 12869 16347 12903
rect 16347 12869 16356 12903
rect 16304 12860 16356 12869
rect 13176 12835 13228 12844
rect 13176 12801 13185 12835
rect 13185 12801 13219 12835
rect 13219 12801 13228 12835
rect 13176 12792 13228 12801
rect 17592 12835 17644 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 1952 12724 2004 12776
rect 4160 12724 4212 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 3056 12656 3108 12708
rect 3792 12656 3844 12708
rect 5632 12656 5684 12708
rect 8760 12656 8812 12708
rect 11428 12724 11480 12776
rect 1492 12588 1544 12640
rect 2136 12588 2188 12640
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 8852 12588 8904 12640
rect 12164 12656 12216 12708
rect 15200 12656 15252 12708
rect 14924 12588 14976 12640
rect 15016 12588 15068 12640
rect 16120 12724 16172 12776
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 17132 12724 17184 12776
rect 3106 12486 3158 12538
rect 3170 12486 3222 12538
rect 3234 12486 3286 12538
rect 3298 12486 3350 12538
rect 3362 12486 3414 12538
rect 6206 12486 6258 12538
rect 6270 12486 6322 12538
rect 6334 12486 6386 12538
rect 6398 12486 6450 12538
rect 6462 12486 6514 12538
rect 9306 12486 9358 12538
rect 9370 12486 9422 12538
rect 9434 12486 9486 12538
rect 9498 12486 9550 12538
rect 9562 12486 9614 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 12534 12486 12586 12538
rect 12598 12486 12650 12538
rect 12662 12486 12714 12538
rect 15506 12486 15558 12538
rect 15570 12486 15622 12538
rect 15634 12486 15686 12538
rect 15698 12486 15750 12538
rect 15762 12486 15814 12538
rect 18606 12486 18658 12538
rect 18670 12486 18722 12538
rect 18734 12486 18786 12538
rect 18798 12486 18850 12538
rect 18862 12486 18914 12538
rect 5264 12384 5316 12436
rect 1676 12316 1728 12368
rect 5356 12316 5408 12368
rect 6644 12359 6696 12368
rect 6644 12325 6653 12359
rect 6653 12325 6687 12359
rect 6687 12325 6696 12359
rect 6644 12316 6696 12325
rect 8576 12316 8628 12368
rect 1492 12248 1544 12300
rect 2044 12248 2096 12300
rect 4160 12248 4212 12300
rect 5448 12248 5500 12300
rect 5816 12291 5868 12300
rect 5816 12257 5826 12291
rect 5826 12257 5860 12291
rect 5860 12257 5868 12291
rect 6368 12291 6420 12300
rect 5816 12248 5868 12257
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 14372 12384 14424 12436
rect 15200 12384 15252 12436
rect 16764 12384 16816 12436
rect 11244 12316 11296 12368
rect 13176 12316 13228 12368
rect 13544 12316 13596 12368
rect 13728 12316 13780 12368
rect 10692 12248 10744 12300
rect 1400 12180 1452 12232
rect 5724 12112 5776 12164
rect 8576 12180 8628 12232
rect 10784 12223 10836 12232
rect 7656 12112 7708 12164
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11428 12248 11480 12300
rect 14832 12316 14884 12368
rect 16120 12359 16172 12368
rect 16120 12325 16129 12359
rect 16129 12325 16163 12359
rect 16163 12325 16172 12359
rect 16120 12316 16172 12325
rect 14280 12248 14332 12300
rect 15016 12248 15068 12300
rect 11796 12180 11848 12232
rect 14740 12180 14792 12232
rect 16580 12248 16632 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17408 12248 17460 12300
rect 16028 12180 16080 12232
rect 12808 12112 12860 12164
rect 1032 12087 1084 12096
rect 1032 12053 1041 12087
rect 1041 12053 1075 12087
rect 1075 12053 1084 12087
rect 1032 12044 1084 12053
rect 5540 12044 5592 12096
rect 9956 12044 10008 12096
rect 12900 12044 12952 12096
rect 14832 12087 14884 12096
rect 14832 12053 14841 12087
rect 14841 12053 14875 12087
rect 14875 12053 14884 12087
rect 14832 12044 14884 12053
rect 1556 11942 1608 11994
rect 1620 11942 1672 11994
rect 1684 11942 1736 11994
rect 1748 11942 1800 11994
rect 1812 11942 1864 11994
rect 4656 11942 4708 11994
rect 4720 11942 4772 11994
rect 4784 11942 4836 11994
rect 4848 11942 4900 11994
rect 4912 11942 4964 11994
rect 7756 11942 7808 11994
rect 7820 11942 7872 11994
rect 7884 11942 7936 11994
rect 7948 11942 8000 11994
rect 8012 11942 8064 11994
rect 10856 11942 10908 11994
rect 10920 11942 10972 11994
rect 10984 11942 11036 11994
rect 11048 11942 11100 11994
rect 11112 11942 11164 11994
rect 13956 11942 14008 11994
rect 14020 11942 14072 11994
rect 14084 11942 14136 11994
rect 14148 11942 14200 11994
rect 14212 11942 14264 11994
rect 17056 11942 17108 11994
rect 17120 11942 17172 11994
rect 17184 11942 17236 11994
rect 17248 11942 17300 11994
rect 17312 11942 17364 11994
rect 10692 11840 10744 11892
rect 15384 11840 15436 11892
rect 17408 11840 17460 11892
rect 6368 11772 6420 11824
rect 9772 11772 9824 11824
rect 2412 11704 2464 11756
rect 10048 11704 10100 11756
rect 1032 11636 1084 11688
rect 5264 11679 5316 11688
rect 5264 11645 5273 11679
rect 5273 11645 5307 11679
rect 5307 11645 5316 11679
rect 5264 11636 5316 11645
rect 5448 11679 5500 11688
rect 5448 11645 5461 11679
rect 5461 11645 5500 11679
rect 5448 11636 5500 11645
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 11520 11704 11572 11756
rect 10416 11679 10468 11688
rect 9220 11636 9272 11645
rect 10416 11645 10425 11679
rect 10425 11645 10459 11679
rect 10459 11645 10468 11679
rect 10416 11636 10468 11645
rect 11336 11636 11388 11688
rect 8208 11568 8260 11620
rect 15292 11704 15344 11756
rect 18144 11704 18196 11756
rect 13176 11636 13228 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 13820 11611 13872 11620
rect 13820 11577 13829 11611
rect 13829 11577 13863 11611
rect 13863 11577 13872 11611
rect 13820 11568 13872 11577
rect 15108 11568 15160 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 7012 11500 7064 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10232 11500 10284 11552
rect 10692 11500 10744 11552
rect 11244 11500 11296 11552
rect 14188 11500 14240 11552
rect 3106 11398 3158 11450
rect 3170 11398 3222 11450
rect 3234 11398 3286 11450
rect 3298 11398 3350 11450
rect 3362 11398 3414 11450
rect 6206 11398 6258 11450
rect 6270 11398 6322 11450
rect 6334 11398 6386 11450
rect 6398 11398 6450 11450
rect 6462 11398 6514 11450
rect 9306 11398 9358 11450
rect 9370 11398 9422 11450
rect 9434 11398 9486 11450
rect 9498 11398 9550 11450
rect 9562 11398 9614 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 12534 11398 12586 11450
rect 12598 11398 12650 11450
rect 12662 11398 12714 11450
rect 15506 11398 15558 11450
rect 15570 11398 15622 11450
rect 15634 11398 15686 11450
rect 15698 11398 15750 11450
rect 15762 11398 15814 11450
rect 18606 11398 18658 11450
rect 18670 11398 18722 11450
rect 18734 11398 18786 11450
rect 18798 11398 18850 11450
rect 18862 11398 18914 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 1952 11296 2004 11348
rect 8208 11339 8260 11348
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 9128 11296 9180 11348
rect 2136 11228 2188 11280
rect 2964 11228 3016 11280
rect 5724 11228 5776 11280
rect 8576 11228 8628 11280
rect 11520 11296 11572 11348
rect 13820 11296 13872 11348
rect 14924 11296 14976 11348
rect 16028 11339 16080 11348
rect 16028 11305 16037 11339
rect 16037 11305 16071 11339
rect 16071 11305 16080 11339
rect 16028 11296 16080 11305
rect 16396 11296 16448 11348
rect 18236 11339 18288 11348
rect 18236 11305 18245 11339
rect 18245 11305 18279 11339
rect 18279 11305 18288 11339
rect 18236 11296 18288 11305
rect 15200 11228 15252 11280
rect 1952 11160 2004 11212
rect 2228 11092 2280 11144
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 5448 11135 5500 11144
rect 2136 11024 2188 11076
rect 3608 10956 3660 11008
rect 4160 10956 4212 11008
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 9772 11160 9824 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10232 11160 10284 11212
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 10600 11092 10652 11144
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 14832 11092 14884 11144
rect 16948 11160 17000 11212
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 6552 10956 6604 11008
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 17500 10999 17552 11008
rect 6920 10956 6972 10965
rect 17500 10965 17509 10999
rect 17509 10965 17543 10999
rect 17543 10965 17552 10999
rect 17500 10956 17552 10965
rect 1556 10854 1608 10906
rect 1620 10854 1672 10906
rect 1684 10854 1736 10906
rect 1748 10854 1800 10906
rect 1812 10854 1864 10906
rect 4656 10854 4708 10906
rect 4720 10854 4772 10906
rect 4784 10854 4836 10906
rect 4848 10854 4900 10906
rect 4912 10854 4964 10906
rect 7756 10854 7808 10906
rect 7820 10854 7872 10906
rect 7884 10854 7936 10906
rect 7948 10854 8000 10906
rect 8012 10854 8064 10906
rect 10856 10854 10908 10906
rect 10920 10854 10972 10906
rect 10984 10854 11036 10906
rect 11048 10854 11100 10906
rect 11112 10854 11164 10906
rect 13956 10854 14008 10906
rect 14020 10854 14072 10906
rect 14084 10854 14136 10906
rect 14148 10854 14200 10906
rect 14212 10854 14264 10906
rect 17056 10854 17108 10906
rect 17120 10854 17172 10906
rect 17184 10854 17236 10906
rect 17248 10854 17300 10906
rect 17312 10854 17364 10906
rect 1400 10752 1452 10804
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 16120 10752 16172 10804
rect 2872 10616 2924 10668
rect 7196 10616 7248 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 6552 10548 6604 10600
rect 7288 10548 7340 10600
rect 10692 10548 10744 10600
rect 11428 10548 11480 10600
rect 16488 10616 16540 10668
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 17500 10591 17552 10600
rect 17500 10557 17510 10591
rect 17510 10557 17544 10591
rect 17544 10557 17552 10591
rect 17500 10548 17552 10557
rect 5908 10480 5960 10532
rect 8116 10523 8168 10532
rect 8116 10489 8125 10523
rect 8125 10489 8159 10523
rect 8159 10489 8168 10523
rect 8116 10480 8168 10489
rect 12164 10480 12216 10532
rect 15292 10523 15344 10532
rect 15292 10489 15301 10523
rect 15301 10489 15335 10523
rect 15335 10489 15344 10523
rect 15292 10480 15344 10489
rect 2964 10412 3016 10464
rect 4988 10412 5040 10464
rect 7104 10412 7156 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 3106 10310 3158 10362
rect 3170 10310 3222 10362
rect 3234 10310 3286 10362
rect 3298 10310 3350 10362
rect 3362 10310 3414 10362
rect 6206 10310 6258 10362
rect 6270 10310 6322 10362
rect 6334 10310 6386 10362
rect 6398 10310 6450 10362
rect 6462 10310 6514 10362
rect 9306 10310 9358 10362
rect 9370 10310 9422 10362
rect 9434 10310 9486 10362
rect 9498 10310 9550 10362
rect 9562 10310 9614 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 12534 10310 12586 10362
rect 12598 10310 12650 10362
rect 12662 10310 12714 10362
rect 15506 10310 15558 10362
rect 15570 10310 15622 10362
rect 15634 10310 15686 10362
rect 15698 10310 15750 10362
rect 15762 10310 15814 10362
rect 18606 10310 18658 10362
rect 18670 10310 18722 10362
rect 18734 10310 18786 10362
rect 18798 10310 18850 10362
rect 18862 10310 18914 10362
rect 2136 10208 2188 10260
rect 3608 10208 3660 10260
rect 5448 10208 5500 10260
rect 9036 10208 9088 10260
rect 10784 10208 10836 10260
rect 15016 10208 15068 10260
rect 4252 10140 4304 10192
rect 7012 10140 7064 10192
rect 16028 10140 16080 10192
rect 940 10072 992 10124
rect 2412 10072 2464 10124
rect 5448 10115 5500 10124
rect 2320 10004 2372 10056
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6920 10072 6972 10124
rect 7656 10004 7708 10056
rect 11244 10072 11296 10124
rect 13820 10115 13872 10124
rect 13820 10081 13828 10115
rect 13828 10081 13862 10115
rect 13862 10081 13872 10115
rect 13820 10072 13872 10081
rect 14464 10072 14516 10124
rect 17868 10140 17920 10192
rect 17408 10072 17460 10124
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 9864 10004 9916 10056
rect 13176 10004 13228 10056
rect 15384 10004 15436 10056
rect 17132 10004 17184 10056
rect 17960 10004 18012 10056
rect 2228 9936 2280 9988
rect 7288 9936 7340 9988
rect 13268 9936 13320 9988
rect 13544 9979 13596 9988
rect 13544 9945 13553 9979
rect 13553 9945 13587 9979
rect 13587 9945 13596 9979
rect 13544 9936 13596 9945
rect 17868 9936 17920 9988
rect 4344 9868 4396 9920
rect 4436 9868 4488 9920
rect 15568 9868 15620 9920
rect 15844 9868 15896 9920
rect 16580 9868 16632 9920
rect 1556 9766 1608 9818
rect 1620 9766 1672 9818
rect 1684 9766 1736 9818
rect 1748 9766 1800 9818
rect 1812 9766 1864 9818
rect 4656 9766 4708 9818
rect 4720 9766 4772 9818
rect 4784 9766 4836 9818
rect 4848 9766 4900 9818
rect 4912 9766 4964 9818
rect 7756 9766 7808 9818
rect 7820 9766 7872 9818
rect 7884 9766 7936 9818
rect 7948 9766 8000 9818
rect 8012 9766 8064 9818
rect 10856 9766 10908 9818
rect 10920 9766 10972 9818
rect 10984 9766 11036 9818
rect 11048 9766 11100 9818
rect 11112 9766 11164 9818
rect 13956 9766 14008 9818
rect 14020 9766 14072 9818
rect 14084 9766 14136 9818
rect 14148 9766 14200 9818
rect 14212 9766 14264 9818
rect 17056 9766 17108 9818
rect 17120 9766 17172 9818
rect 17184 9766 17236 9818
rect 17248 9766 17300 9818
rect 17312 9766 17364 9818
rect 10692 9664 10744 9716
rect 14464 9664 14516 9716
rect 1400 9596 1452 9648
rect 1768 9528 1820 9580
rect 2228 9596 2280 9648
rect 2872 9596 2924 9648
rect 11612 9596 11664 9648
rect 14740 9596 14792 9648
rect 2044 9528 2096 9580
rect 8944 9528 8996 9580
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 11888 9528 11940 9580
rect 15016 9528 15068 9580
rect 17408 9664 17460 9716
rect 15200 9596 15252 9648
rect 2136 9460 2188 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 1400 9392 1452 9444
rect 2780 9392 2832 9444
rect 4988 9460 5040 9512
rect 5724 9460 5776 9512
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 14372 9460 14424 9512
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 17316 9460 17368 9512
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 6644 9392 6696 9444
rect 8668 9392 8720 9444
rect 1032 9324 1084 9376
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 4712 9324 4764 9376
rect 8392 9324 8444 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 10784 9392 10836 9444
rect 11612 9324 11664 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 15016 9324 15068 9376
rect 16212 9435 16264 9444
rect 16212 9401 16246 9435
rect 16246 9401 16264 9435
rect 17592 9435 17644 9444
rect 16212 9392 16264 9401
rect 17592 9401 17601 9435
rect 17601 9401 17635 9435
rect 17635 9401 17644 9435
rect 17592 9392 17644 9401
rect 16856 9324 16908 9376
rect 17408 9324 17460 9376
rect 17960 9324 18012 9376
rect 3106 9222 3158 9274
rect 3170 9222 3222 9274
rect 3234 9222 3286 9274
rect 3298 9222 3350 9274
rect 3362 9222 3414 9274
rect 6206 9222 6258 9274
rect 6270 9222 6322 9274
rect 6334 9222 6386 9274
rect 6398 9222 6450 9274
rect 6462 9222 6514 9274
rect 9306 9222 9358 9274
rect 9370 9222 9422 9274
rect 9434 9222 9486 9274
rect 9498 9222 9550 9274
rect 9562 9222 9614 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 12534 9222 12586 9274
rect 12598 9222 12650 9274
rect 12662 9222 12714 9274
rect 15506 9222 15558 9274
rect 15570 9222 15622 9274
rect 15634 9222 15686 9274
rect 15698 9222 15750 9274
rect 15762 9222 15814 9274
rect 18606 9222 18658 9274
rect 18670 9222 18722 9274
rect 18734 9222 18786 9274
rect 18798 9222 18850 9274
rect 18862 9222 18914 9274
rect 2872 9120 2924 9172
rect 5448 9120 5500 9172
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 7196 9120 7248 9172
rect 11336 9120 11388 9172
rect 11428 9120 11480 9172
rect 17316 9163 17368 9172
rect 17316 9129 17325 9163
rect 17325 9129 17359 9163
rect 17359 9129 17368 9163
rect 17316 9120 17368 9129
rect 17500 9120 17552 9172
rect 2136 9052 2188 9104
rect 2780 9052 2832 9104
rect 2044 9027 2096 9036
rect 2044 8993 2053 9027
rect 2053 8993 2087 9027
rect 2087 8993 2096 9027
rect 2044 8984 2096 8993
rect 4160 8984 4212 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 5908 9027 5960 9036
rect 4712 8984 4764 8993
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6644 8984 6696 9036
rect 9036 9052 9088 9104
rect 10784 9052 10836 9104
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 8116 8984 8168 9036
rect 8668 8984 8720 9036
rect 11888 8984 11940 9036
rect 12992 9052 13044 9104
rect 18512 9052 18564 9104
rect 8300 8916 8352 8968
rect 9864 8916 9916 8968
rect 11336 8916 11388 8968
rect 14648 8984 14700 9036
rect 17684 8984 17736 9036
rect 2044 8848 2096 8900
rect 3424 8848 3476 8900
rect 5816 8848 5868 8900
rect 6000 8848 6052 8900
rect 14832 8916 14884 8968
rect 16212 8916 16264 8968
rect 17960 8916 18012 8968
rect 14372 8848 14424 8900
rect 15568 8848 15620 8900
rect 8116 8780 8168 8832
rect 15292 8780 15344 8832
rect 16580 8780 16632 8832
rect 18420 8780 18472 8832
rect 1556 8678 1608 8730
rect 1620 8678 1672 8730
rect 1684 8678 1736 8730
rect 1748 8678 1800 8730
rect 1812 8678 1864 8730
rect 4656 8678 4708 8730
rect 4720 8678 4772 8730
rect 4784 8678 4836 8730
rect 4848 8678 4900 8730
rect 4912 8678 4964 8730
rect 7756 8678 7808 8730
rect 7820 8678 7872 8730
rect 7884 8678 7936 8730
rect 7948 8678 8000 8730
rect 8012 8678 8064 8730
rect 10856 8678 10908 8730
rect 10920 8678 10972 8730
rect 10984 8678 11036 8730
rect 11048 8678 11100 8730
rect 11112 8678 11164 8730
rect 13956 8678 14008 8730
rect 14020 8678 14072 8730
rect 14084 8678 14136 8730
rect 14148 8678 14200 8730
rect 14212 8678 14264 8730
rect 17056 8678 17108 8730
rect 17120 8678 17172 8730
rect 17184 8678 17236 8730
rect 17248 8678 17300 8730
rect 17312 8678 17364 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 8116 8576 8168 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 12992 8576 13044 8628
rect 5816 8508 5868 8560
rect 1400 8372 1452 8424
rect 2688 8440 2740 8492
rect 4160 8440 4212 8492
rect 5172 8440 5224 8492
rect 2412 8372 2464 8424
rect 3424 8415 3476 8424
rect 1124 8304 1176 8356
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 5724 8372 5776 8424
rect 6920 8372 6972 8424
rect 10508 8440 10560 8492
rect 11888 8440 11940 8492
rect 8300 8415 8352 8424
rect 3792 8304 3844 8356
rect 5264 8347 5316 8356
rect 5264 8313 5273 8347
rect 5273 8313 5307 8347
rect 5307 8313 5316 8347
rect 5264 8304 5316 8313
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 12256 8372 12308 8424
rect 15384 8576 15436 8628
rect 17592 8576 17644 8628
rect 18512 8576 18564 8628
rect 13820 8440 13872 8492
rect 14556 8440 14608 8492
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15936 8440 15988 8492
rect 14464 8415 14516 8424
rect 8668 8304 8720 8356
rect 10876 8304 10928 8356
rect 12164 8304 12216 8356
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14832 8372 14884 8424
rect 15016 8372 15068 8424
rect 15844 8372 15896 8424
rect 16488 8372 16540 8424
rect 16672 8415 16724 8424
rect 16672 8381 16706 8415
rect 16706 8381 16724 8415
rect 16672 8372 16724 8381
rect 1216 8236 1268 8288
rect 15568 8304 15620 8356
rect 14280 8236 14332 8288
rect 16396 8236 16448 8288
rect 3106 8134 3158 8186
rect 3170 8134 3222 8186
rect 3234 8134 3286 8186
rect 3298 8134 3350 8186
rect 3362 8134 3414 8186
rect 6206 8134 6258 8186
rect 6270 8134 6322 8186
rect 6334 8134 6386 8186
rect 6398 8134 6450 8186
rect 6462 8134 6514 8186
rect 9306 8134 9358 8186
rect 9370 8134 9422 8186
rect 9434 8134 9486 8186
rect 9498 8134 9550 8186
rect 9562 8134 9614 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 12534 8134 12586 8186
rect 12598 8134 12650 8186
rect 12662 8134 12714 8186
rect 15506 8134 15558 8186
rect 15570 8134 15622 8186
rect 15634 8134 15686 8186
rect 15698 8134 15750 8186
rect 15762 8134 15814 8186
rect 18606 8134 18658 8186
rect 18670 8134 18722 8186
rect 18734 8134 18786 8186
rect 18798 8134 18850 8186
rect 18862 8134 18914 8186
rect 1216 8075 1268 8084
rect 1216 8041 1225 8075
rect 1225 8041 1259 8075
rect 1259 8041 1268 8075
rect 1216 8032 1268 8041
rect 7564 8032 7616 8084
rect 8668 8032 8720 8084
rect 10416 8032 10468 8084
rect 14648 8032 14700 8084
rect 1124 7964 1176 8016
rect 6552 7964 6604 8016
rect 10876 7964 10928 8016
rect 18328 8032 18380 8084
rect 1032 7939 1084 7948
rect 1032 7905 1041 7939
rect 1041 7905 1075 7939
rect 1075 7905 1084 7939
rect 1032 7896 1084 7905
rect 2044 7896 2096 7948
rect 5264 7896 5316 7948
rect 11888 7896 11940 7948
rect 15936 7964 15988 8016
rect 4988 7828 5040 7880
rect 6920 7828 6972 7880
rect 12992 7896 13044 7948
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 17316 7939 17368 7948
rect 16488 7896 16540 7905
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 17500 7896 17552 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 12808 7828 12860 7880
rect 13544 7760 13596 7812
rect 14832 7760 14884 7812
rect 12532 7735 12584 7744
rect 12532 7701 12541 7735
rect 12541 7701 12575 7735
rect 12575 7701 12584 7735
rect 12532 7692 12584 7701
rect 14556 7692 14608 7744
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 1556 7590 1608 7642
rect 1620 7590 1672 7642
rect 1684 7590 1736 7642
rect 1748 7590 1800 7642
rect 1812 7590 1864 7642
rect 4656 7590 4708 7642
rect 4720 7590 4772 7642
rect 4784 7590 4836 7642
rect 4848 7590 4900 7642
rect 4912 7590 4964 7642
rect 7756 7590 7808 7642
rect 7820 7590 7872 7642
rect 7884 7590 7936 7642
rect 7948 7590 8000 7642
rect 8012 7590 8064 7642
rect 10856 7590 10908 7642
rect 10920 7590 10972 7642
rect 10984 7590 11036 7642
rect 11048 7590 11100 7642
rect 11112 7590 11164 7642
rect 13956 7590 14008 7642
rect 14020 7590 14072 7642
rect 14084 7590 14136 7642
rect 14148 7590 14200 7642
rect 14212 7590 14264 7642
rect 17056 7590 17108 7642
rect 17120 7590 17172 7642
rect 17184 7590 17236 7642
rect 17248 7590 17300 7642
rect 17312 7590 17364 7642
rect 4436 7488 4488 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5356 7488 5408 7540
rect 5632 7488 5684 7540
rect 7564 7531 7616 7540
rect 7564 7497 7573 7531
rect 7573 7497 7607 7531
rect 7607 7497 7616 7531
rect 7564 7488 7616 7497
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 12532 7488 12584 7540
rect 11428 7463 11480 7472
rect 2872 7352 2924 7404
rect 5908 7352 5960 7404
rect 11428 7429 11437 7463
rect 11437 7429 11471 7463
rect 11471 7429 11480 7463
rect 11428 7420 11480 7429
rect 11888 7420 11940 7472
rect 16488 7488 16540 7540
rect 16856 7488 16908 7540
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 8300 7284 8352 7336
rect 2136 7259 2188 7268
rect 2136 7225 2145 7259
rect 2145 7225 2179 7259
rect 2179 7225 2188 7259
rect 2136 7216 2188 7225
rect 4160 7216 4212 7268
rect 5908 7216 5960 7268
rect 6552 7216 6604 7268
rect 7564 7216 7616 7268
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 11244 7327 11296 7336
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 9220 7216 9272 7268
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 14280 7216 14332 7268
rect 16396 7259 16448 7268
rect 16396 7225 16430 7259
rect 16430 7225 16448 7259
rect 14556 7148 14608 7200
rect 16396 7216 16448 7225
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 3106 7046 3158 7098
rect 3170 7046 3222 7098
rect 3234 7046 3286 7098
rect 3298 7046 3350 7098
rect 3362 7046 3414 7098
rect 6206 7046 6258 7098
rect 6270 7046 6322 7098
rect 6334 7046 6386 7098
rect 6398 7046 6450 7098
rect 6462 7046 6514 7098
rect 9306 7046 9358 7098
rect 9370 7046 9422 7098
rect 9434 7046 9486 7098
rect 9498 7046 9550 7098
rect 9562 7046 9614 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 12534 7046 12586 7098
rect 12598 7046 12650 7098
rect 12662 7046 12714 7098
rect 15506 7046 15558 7098
rect 15570 7046 15622 7098
rect 15634 7046 15686 7098
rect 15698 7046 15750 7098
rect 15762 7046 15814 7098
rect 18606 7046 18658 7098
rect 18670 7046 18722 7098
rect 18734 7046 18786 7098
rect 18798 7046 18850 7098
rect 18862 7046 18914 7098
rect 1216 6944 1268 6996
rect 18144 6944 18196 6996
rect 18236 6944 18288 6996
rect 4160 6876 4212 6928
rect 8668 6876 8720 6928
rect 2412 6808 2464 6860
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7656 6808 7708 6860
rect 8208 6808 8260 6860
rect 11520 6851 11572 6860
rect 11520 6817 11529 6851
rect 11529 6817 11563 6851
rect 11563 6817 11572 6851
rect 11520 6808 11572 6817
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 16764 6808 16816 6860
rect 17500 6808 17552 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2780 6740 2832 6792
rect 1952 6672 2004 6724
rect 4160 6672 4212 6724
rect 6828 6672 6880 6724
rect 8392 6740 8444 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11612 6740 11664 6792
rect 13820 6740 13872 6792
rect 14464 6740 14516 6792
rect 16580 6740 16632 6792
rect 12808 6672 12860 6724
rect 2872 6604 2924 6656
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 5816 6604 5868 6656
rect 6644 6604 6696 6656
rect 8944 6604 8996 6656
rect 12164 6604 12216 6656
rect 15752 6672 15804 6724
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 15844 6604 15896 6656
rect 16396 6672 16448 6724
rect 1556 6502 1608 6554
rect 1620 6502 1672 6554
rect 1684 6502 1736 6554
rect 1748 6502 1800 6554
rect 1812 6502 1864 6554
rect 4656 6502 4708 6554
rect 4720 6502 4772 6554
rect 4784 6502 4836 6554
rect 4848 6502 4900 6554
rect 4912 6502 4964 6554
rect 7756 6502 7808 6554
rect 7820 6502 7872 6554
rect 7884 6502 7936 6554
rect 7948 6502 8000 6554
rect 8012 6502 8064 6554
rect 10856 6502 10908 6554
rect 10920 6502 10972 6554
rect 10984 6502 11036 6554
rect 11048 6502 11100 6554
rect 11112 6502 11164 6554
rect 13956 6502 14008 6554
rect 14020 6502 14072 6554
rect 14084 6502 14136 6554
rect 14148 6502 14200 6554
rect 14212 6502 14264 6554
rect 17056 6502 17108 6554
rect 17120 6502 17172 6554
rect 17184 6502 17236 6554
rect 17248 6502 17300 6554
rect 17312 6502 17364 6554
rect 1400 6400 1452 6452
rect 2228 6400 2280 6452
rect 5632 6400 5684 6452
rect 11336 6400 11388 6452
rect 17592 6400 17644 6452
rect 17960 6400 18012 6452
rect 2228 6264 2280 6316
rect 5540 6332 5592 6384
rect 5816 6332 5868 6384
rect 6000 6332 6052 6384
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5264 6264 5316 6316
rect 3884 6196 3936 6248
rect 5356 6196 5408 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 3792 6060 3844 6112
rect 5540 6060 5592 6112
rect 5724 6128 5776 6180
rect 6644 6264 6696 6316
rect 8760 6332 8812 6384
rect 9220 6375 9272 6384
rect 9220 6341 9229 6375
rect 9229 6341 9263 6375
rect 9263 6341 9272 6375
rect 9220 6332 9272 6341
rect 15016 6332 15068 6384
rect 8484 6264 8536 6316
rect 11428 6264 11480 6316
rect 14372 6264 14424 6316
rect 13176 6196 13228 6248
rect 14464 6239 14516 6248
rect 6644 6171 6696 6180
rect 6644 6137 6653 6171
rect 6653 6137 6687 6171
rect 6687 6137 6696 6171
rect 6644 6128 6696 6137
rect 8024 6128 8076 6180
rect 8208 6128 8260 6180
rect 12164 6128 12216 6180
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 14648 6196 14700 6248
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 15844 6264 15896 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 18052 6264 18104 6316
rect 14556 6128 14608 6180
rect 15384 6128 15436 6180
rect 7012 6060 7064 6112
rect 7564 6060 7616 6112
rect 9220 6060 9272 6112
rect 15936 6060 15988 6112
rect 16948 6060 17000 6112
rect 3106 5958 3158 6010
rect 3170 5958 3222 6010
rect 3234 5958 3286 6010
rect 3298 5958 3350 6010
rect 3362 5958 3414 6010
rect 6206 5958 6258 6010
rect 6270 5958 6322 6010
rect 6334 5958 6386 6010
rect 6398 5958 6450 6010
rect 6462 5958 6514 6010
rect 9306 5958 9358 6010
rect 9370 5958 9422 6010
rect 9434 5958 9486 6010
rect 9498 5958 9550 6010
rect 9562 5958 9614 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 12534 5958 12586 6010
rect 12598 5958 12650 6010
rect 12662 5958 12714 6010
rect 15506 5958 15558 6010
rect 15570 5958 15622 6010
rect 15634 5958 15686 6010
rect 15698 5958 15750 6010
rect 15762 5958 15814 6010
rect 18606 5958 18658 6010
rect 18670 5958 18722 6010
rect 18734 5958 18786 6010
rect 18798 5958 18850 6010
rect 18862 5958 18914 6010
rect 2044 5856 2096 5908
rect 1952 5720 2004 5772
rect 3240 5720 3292 5772
rect 4436 5788 4488 5840
rect 8024 5856 8076 5908
rect 5908 5788 5960 5840
rect 7380 5788 7432 5840
rect 9220 5788 9272 5840
rect 16120 5856 16172 5908
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 4344 5720 4396 5772
rect 2228 5652 2280 5704
rect 2688 5584 2740 5636
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 6828 5652 6880 5704
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 11428 5720 11480 5772
rect 12164 5788 12216 5840
rect 15936 5788 15988 5840
rect 18328 5856 18380 5908
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 16764 5763 16816 5772
rect 11796 5720 11848 5729
rect 16764 5729 16773 5763
rect 16773 5729 16807 5763
rect 16807 5729 16816 5763
rect 16764 5720 16816 5729
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 3240 5584 3292 5636
rect 5080 5584 5132 5636
rect 11244 5584 11296 5636
rect 14280 5652 14332 5704
rect 16120 5652 16172 5704
rect 16212 5652 16264 5704
rect 12256 5584 12308 5636
rect 4252 5516 4304 5568
rect 5356 5516 5408 5568
rect 7104 5516 7156 5568
rect 10232 5516 10284 5568
rect 14832 5516 14884 5568
rect 1556 5414 1608 5466
rect 1620 5414 1672 5466
rect 1684 5414 1736 5466
rect 1748 5414 1800 5466
rect 1812 5414 1864 5466
rect 4656 5414 4708 5466
rect 4720 5414 4772 5466
rect 4784 5414 4836 5466
rect 4848 5414 4900 5466
rect 4912 5414 4964 5466
rect 7756 5414 7808 5466
rect 7820 5414 7872 5466
rect 7884 5414 7936 5466
rect 7948 5414 8000 5466
rect 8012 5414 8064 5466
rect 10856 5414 10908 5466
rect 10920 5414 10972 5466
rect 10984 5414 11036 5466
rect 11048 5414 11100 5466
rect 11112 5414 11164 5466
rect 13956 5414 14008 5466
rect 14020 5414 14072 5466
rect 14084 5414 14136 5466
rect 14148 5414 14200 5466
rect 14212 5414 14264 5466
rect 17056 5414 17108 5466
rect 17120 5414 17172 5466
rect 17184 5414 17236 5466
rect 17248 5414 17300 5466
rect 17312 5414 17364 5466
rect 1584 5312 1636 5364
rect 2044 5312 2096 5364
rect 4528 5312 4580 5364
rect 5172 5312 5224 5364
rect 8116 5355 8168 5364
rect 8116 5321 8125 5355
rect 8125 5321 8159 5355
rect 8159 5321 8168 5355
rect 8116 5312 8168 5321
rect 11244 5312 11296 5364
rect 14280 5312 14332 5364
rect 2136 5244 2188 5296
rect 3884 5244 3936 5296
rect 8852 5244 8904 5296
rect 2780 5176 2832 5228
rect 5264 5176 5316 5228
rect 7288 5176 7340 5228
rect 11796 5219 11848 5228
rect 848 5108 900 5160
rect 2688 5108 2740 5160
rect 3884 5108 3936 5160
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 4436 5151 4488 5160
rect 4436 5117 4445 5151
rect 4445 5117 4479 5151
rect 4479 5117 4488 5151
rect 4436 5108 4488 5117
rect 5724 5108 5776 5160
rect 6920 5108 6972 5160
rect 8208 5108 8260 5160
rect 8300 5108 8352 5160
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 8852 5108 8904 5160
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9588 5151 9640 5160
rect 9220 5108 9272 5117
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 4804 5040 4856 5092
rect 5448 5040 5500 5092
rect 9036 5040 9088 5092
rect 10232 5083 10284 5092
rect 10232 5049 10241 5083
rect 10241 5049 10275 5083
rect 10275 5049 10284 5083
rect 10232 5040 10284 5049
rect 4528 4972 4580 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 6828 4972 6880 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 12900 4972 12952 5024
rect 3106 4870 3158 4922
rect 3170 4870 3222 4922
rect 3234 4870 3286 4922
rect 3298 4870 3350 4922
rect 3362 4870 3414 4922
rect 6206 4870 6258 4922
rect 6270 4870 6322 4922
rect 6334 4870 6386 4922
rect 6398 4870 6450 4922
rect 6462 4870 6514 4922
rect 9306 4870 9358 4922
rect 9370 4870 9422 4922
rect 9434 4870 9486 4922
rect 9498 4870 9550 4922
rect 9562 4870 9614 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 12534 4870 12586 4922
rect 12598 4870 12650 4922
rect 12662 4870 12714 4922
rect 15506 4870 15558 4922
rect 15570 4870 15622 4922
rect 15634 4870 15686 4922
rect 15698 4870 15750 4922
rect 15762 4870 15814 4922
rect 18606 4870 18658 4922
rect 18670 4870 18722 4922
rect 18734 4870 18786 4922
rect 18798 4870 18850 4922
rect 18862 4870 18914 4922
rect 848 4811 900 4820
rect 848 4777 857 4811
rect 857 4777 891 4811
rect 891 4777 900 4811
rect 848 4768 900 4777
rect 2872 4768 2924 4820
rect 4988 4768 5040 4820
rect 5356 4768 5408 4820
rect 5816 4768 5868 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7196 4768 7248 4820
rect 8392 4811 8444 4820
rect 5172 4700 5224 4752
rect 6000 4700 6052 4752
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 11336 4768 11388 4820
rect 940 4675 992 4684
rect 940 4641 949 4675
rect 949 4641 983 4675
rect 983 4641 992 4675
rect 940 4632 992 4641
rect 1032 4632 1084 4684
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 4252 4675 4304 4684
rect 1584 4632 1636 4641
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 4712 4675 4764 4684
rect 4712 4641 4721 4675
rect 4721 4641 4755 4675
rect 4755 4641 4764 4675
rect 4712 4632 4764 4641
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 2596 4564 2648 4616
rect 7472 4632 7524 4684
rect 6828 4496 6880 4548
rect 5724 4428 5776 4480
rect 9220 4700 9272 4752
rect 8484 4564 8536 4616
rect 8944 4632 8996 4684
rect 9956 4632 10008 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 11428 4607 11480 4616
rect 8760 4496 8812 4548
rect 7472 4428 7524 4480
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11796 4632 11848 4684
rect 13820 4700 13872 4752
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 13636 4539 13688 4548
rect 13636 4505 13645 4539
rect 13645 4505 13679 4539
rect 13679 4505 13688 4539
rect 13636 4496 13688 4505
rect 14280 4632 14332 4684
rect 17408 4768 17460 4820
rect 15936 4700 15988 4752
rect 16580 4700 16632 4752
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 16948 4632 17000 4684
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 17776 4496 17828 4548
rect 14924 4428 14976 4480
rect 15016 4471 15068 4480
rect 15016 4437 15025 4471
rect 15025 4437 15059 4471
rect 15059 4437 15068 4471
rect 15016 4428 15068 4437
rect 16672 4428 16724 4480
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 1556 4326 1608 4378
rect 1620 4326 1672 4378
rect 1684 4326 1736 4378
rect 1748 4326 1800 4378
rect 1812 4326 1864 4378
rect 4656 4326 4708 4378
rect 4720 4326 4772 4378
rect 4784 4326 4836 4378
rect 4848 4326 4900 4378
rect 4912 4326 4964 4378
rect 7756 4326 7808 4378
rect 7820 4326 7872 4378
rect 7884 4326 7936 4378
rect 7948 4326 8000 4378
rect 8012 4326 8064 4378
rect 10856 4326 10908 4378
rect 10920 4326 10972 4378
rect 10984 4326 11036 4378
rect 11048 4326 11100 4378
rect 11112 4326 11164 4378
rect 13956 4326 14008 4378
rect 14020 4326 14072 4378
rect 14084 4326 14136 4378
rect 14148 4326 14200 4378
rect 14212 4326 14264 4378
rect 17056 4326 17108 4378
rect 17120 4326 17172 4378
rect 17184 4326 17236 4378
rect 17248 4326 17300 4378
rect 17312 4326 17364 4378
rect 2596 4267 2648 4276
rect 2596 4233 2605 4267
rect 2605 4233 2639 4267
rect 2639 4233 2648 4267
rect 2596 4224 2648 4233
rect 5080 4224 5132 4276
rect 7196 4224 7248 4276
rect 8760 4267 8812 4276
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 8944 4224 8996 4276
rect 9772 4267 9824 4276
rect 2872 4156 2924 4208
rect 4160 4156 4212 4208
rect 6828 4156 6880 4208
rect 1952 4088 2004 4140
rect 2320 4088 2372 4140
rect 6000 4131 6052 4140
rect 2688 4020 2740 4072
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 3516 4020 3568 4072
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 11428 4224 11480 4276
rect 14648 4224 14700 4276
rect 14924 4224 14976 4276
rect 16764 4224 16816 4276
rect 9680 4088 9732 4140
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 6828 3952 6880 4004
rect 7012 3995 7064 4004
rect 7012 3961 7021 3995
rect 7021 3961 7055 3995
rect 7055 3961 7064 3995
rect 7012 3952 7064 3961
rect 7196 3952 7248 4004
rect 7380 3995 7432 4004
rect 7380 3961 7389 3995
rect 7389 3961 7423 3995
rect 7423 3961 7432 3995
rect 7380 3952 7432 3961
rect 7472 3952 7524 4004
rect 940 3884 992 3936
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 2872 3884 2924 3936
rect 6644 3884 6696 3936
rect 7564 3884 7616 3936
rect 9864 4020 9916 4072
rect 13636 4088 13688 4140
rect 14924 4088 14976 4140
rect 16580 4020 16632 4072
rect 16948 4088 17000 4140
rect 17868 4088 17920 4140
rect 8944 3952 8996 4004
rect 10232 3995 10284 4004
rect 10232 3961 10241 3995
rect 10241 3961 10275 3995
rect 10275 3961 10284 3995
rect 10232 3952 10284 3961
rect 15936 3952 15988 4004
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 12900 3884 12952 3936
rect 15384 3884 15436 3936
rect 16212 3927 16264 3936
rect 16212 3893 16221 3927
rect 16221 3893 16255 3927
rect 16255 3893 16264 3927
rect 16212 3884 16264 3893
rect 16580 3927 16632 3936
rect 16580 3893 16589 3927
rect 16589 3893 16623 3927
rect 16623 3893 16632 3927
rect 16580 3884 16632 3893
rect 16764 3884 16816 3936
rect 18328 3884 18380 3936
rect 3106 3782 3158 3834
rect 3170 3782 3222 3834
rect 3234 3782 3286 3834
rect 3298 3782 3350 3834
rect 3362 3782 3414 3834
rect 6206 3782 6258 3834
rect 6270 3782 6322 3834
rect 6334 3782 6386 3834
rect 6398 3782 6450 3834
rect 6462 3782 6514 3834
rect 9306 3782 9358 3834
rect 9370 3782 9422 3834
rect 9434 3782 9486 3834
rect 9498 3782 9550 3834
rect 9562 3782 9614 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 12534 3782 12586 3834
rect 12598 3782 12650 3834
rect 12662 3782 12714 3834
rect 15506 3782 15558 3834
rect 15570 3782 15622 3834
rect 15634 3782 15686 3834
rect 15698 3782 15750 3834
rect 15762 3782 15814 3834
rect 18606 3782 18658 3834
rect 18670 3782 18722 3834
rect 18734 3782 18786 3834
rect 18798 3782 18850 3834
rect 18862 3782 18914 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 3608 3680 3660 3732
rect 4252 3680 4304 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 11336 3680 11388 3732
rect 11520 3680 11572 3732
rect 2688 3544 2740 3596
rect 2964 3587 3016 3596
rect 2964 3553 2973 3587
rect 2973 3553 3007 3587
rect 3007 3553 3016 3587
rect 2964 3544 3016 3553
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 3700 3544 3752 3596
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 12532 3612 12584 3664
rect 12992 3680 13044 3732
rect 13084 3680 13136 3732
rect 16580 3680 16632 3732
rect 18052 3680 18104 3732
rect 12808 3612 12860 3664
rect 5264 3544 5316 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 11428 3544 11480 3596
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 12900 3476 12952 3528
rect 13820 3544 13872 3596
rect 14372 3544 14424 3596
rect 14924 3612 14976 3664
rect 16028 3612 16080 3664
rect 17684 3612 17736 3664
rect 13544 3476 13596 3528
rect 14280 3476 14332 3528
rect 15384 3476 15436 3528
rect 17868 3544 17920 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 18328 3587 18380 3596
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 4344 3451 4396 3460
rect 4344 3417 4353 3451
rect 4353 3417 4387 3451
rect 4387 3417 4396 3451
rect 4344 3408 4396 3417
rect 14740 3408 14792 3460
rect 16856 3408 16908 3460
rect 5724 3340 5776 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 1556 3238 1608 3290
rect 1620 3238 1672 3290
rect 1684 3238 1736 3290
rect 1748 3238 1800 3290
rect 1812 3238 1864 3290
rect 4656 3238 4708 3290
rect 4720 3238 4772 3290
rect 4784 3238 4836 3290
rect 4848 3238 4900 3290
rect 4912 3238 4964 3290
rect 7756 3238 7808 3290
rect 7820 3238 7872 3290
rect 7884 3238 7936 3290
rect 7948 3238 8000 3290
rect 8012 3238 8064 3290
rect 10856 3238 10908 3290
rect 10920 3238 10972 3290
rect 10984 3238 11036 3290
rect 11048 3238 11100 3290
rect 11112 3238 11164 3290
rect 13956 3238 14008 3290
rect 14020 3238 14072 3290
rect 14084 3238 14136 3290
rect 14148 3238 14200 3290
rect 14212 3238 14264 3290
rect 17056 3238 17108 3290
rect 17120 3238 17172 3290
rect 17184 3238 17236 3290
rect 17248 3238 17300 3290
rect 17312 3238 17364 3290
rect 1032 3136 1084 3188
rect 1952 3136 2004 3188
rect 4160 3136 4212 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 9128 3136 9180 3188
rect 12532 3136 12584 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 17592 3136 17644 3188
rect 17868 3136 17920 3188
rect 6368 3068 6420 3120
rect 8944 3068 8996 3120
rect 2780 3000 2832 3052
rect 5632 3000 5684 3052
rect 6828 3000 6880 3052
rect 1032 2975 1084 2984
rect 1032 2941 1041 2975
rect 1041 2941 1075 2975
rect 1075 2941 1084 2975
rect 1032 2932 1084 2941
rect 2044 2932 2096 2984
rect 2964 2932 3016 2984
rect 3700 2932 3752 2984
rect 5356 2932 5408 2984
rect 5816 2932 5868 2984
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 13728 3068 13780 3120
rect 9220 3000 9272 3052
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 13636 3000 13688 3052
rect 16580 3068 16632 3120
rect 17500 3068 17552 3120
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 19064 2932 19116 2984
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 5632 2839 5684 2848
rect 1952 2796 2004 2805
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 12440 2796 12492 2848
rect 12992 2796 13044 2848
rect 13544 2796 13596 2848
rect 13912 2796 13964 2848
rect 14372 2796 14424 2848
rect 15200 2796 15252 2848
rect 16212 2839 16264 2848
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 16304 2796 16356 2805
rect 3106 2694 3158 2746
rect 3170 2694 3222 2746
rect 3234 2694 3286 2746
rect 3298 2694 3350 2746
rect 3362 2694 3414 2746
rect 6206 2694 6258 2746
rect 6270 2694 6322 2746
rect 6334 2694 6386 2746
rect 6398 2694 6450 2746
rect 6462 2694 6514 2746
rect 9306 2694 9358 2746
rect 9370 2694 9422 2746
rect 9434 2694 9486 2746
rect 9498 2694 9550 2746
rect 9562 2694 9614 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 12534 2694 12586 2746
rect 12598 2694 12650 2746
rect 12662 2694 12714 2746
rect 15506 2694 15558 2746
rect 15570 2694 15622 2746
rect 15634 2694 15686 2746
rect 15698 2694 15750 2746
rect 15762 2694 15814 2746
rect 18606 2694 18658 2746
rect 18670 2694 18722 2746
rect 18734 2694 18786 2746
rect 18798 2694 18850 2746
rect 18862 2694 18914 2746
rect 1032 2592 1084 2644
rect 5540 2592 5592 2644
rect 6000 2592 6052 2644
rect 8024 2592 8076 2644
rect 9220 2592 9272 2644
rect 13820 2592 13872 2644
rect 3332 2524 3384 2576
rect 3884 2524 3936 2576
rect 7288 2524 7340 2576
rect 2872 2456 2924 2508
rect 4068 2456 4120 2508
rect 5356 2499 5408 2508
rect 5356 2465 5365 2499
rect 5365 2465 5399 2499
rect 5399 2465 5408 2499
rect 5356 2456 5408 2465
rect 7104 2456 7156 2508
rect 7656 2524 7708 2576
rect 8024 2456 8076 2508
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 5724 2388 5776 2440
rect 8668 2524 8720 2576
rect 9864 2524 9916 2576
rect 9680 2456 9732 2508
rect 10600 2524 10652 2576
rect 13912 2524 13964 2576
rect 14832 2524 14884 2576
rect 15384 2592 15436 2644
rect 16580 2592 16632 2644
rect 17776 2592 17828 2644
rect 13728 2499 13780 2508
rect 9864 2388 9916 2440
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 16764 2524 16816 2576
rect 17408 2456 17460 2508
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17868 2499 17920 2508
rect 17500 2456 17552 2465
rect 17868 2465 17877 2499
rect 17877 2465 17911 2499
rect 17911 2465 17920 2499
rect 17868 2456 17920 2465
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 15016 2388 15068 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16488 2388 16540 2440
rect 9220 2320 9272 2372
rect 9036 2252 9088 2304
rect 16764 2320 16816 2372
rect 17684 2320 17736 2372
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 10324 2252 10376 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 1556 2150 1608 2202
rect 1620 2150 1672 2202
rect 1684 2150 1736 2202
rect 1748 2150 1800 2202
rect 1812 2150 1864 2202
rect 4656 2150 4708 2202
rect 4720 2150 4772 2202
rect 4784 2150 4836 2202
rect 4848 2150 4900 2202
rect 4912 2150 4964 2202
rect 7756 2150 7808 2202
rect 7820 2150 7872 2202
rect 7884 2150 7936 2202
rect 7948 2150 8000 2202
rect 8012 2150 8064 2202
rect 10856 2150 10908 2202
rect 10920 2150 10972 2202
rect 10984 2150 11036 2202
rect 11048 2150 11100 2202
rect 11112 2150 11164 2202
rect 13956 2150 14008 2202
rect 14020 2150 14072 2202
rect 14084 2150 14136 2202
rect 14148 2150 14200 2202
rect 14212 2150 14264 2202
rect 17056 2150 17108 2202
rect 17120 2150 17172 2202
rect 17184 2150 17236 2202
rect 17248 2150 17300 2202
rect 17312 2150 17364 2202
rect 1952 2048 2004 2100
rect 2872 2091 2924 2100
rect 2872 2057 2881 2091
rect 2881 2057 2915 2091
rect 2915 2057 2924 2091
rect 2872 2048 2924 2057
rect 5632 2048 5684 2100
rect 5816 2048 5868 2100
rect 7012 2048 7064 2100
rect 9220 2091 9272 2100
rect 9220 2057 9229 2091
rect 9229 2057 9263 2091
rect 9263 2057 9272 2091
rect 9220 2048 9272 2057
rect 9772 1980 9824 2032
rect 12808 1980 12860 2032
rect 14556 2048 14608 2100
rect 15016 2048 15068 2100
rect 16304 2048 16356 2100
rect 2780 1912 2832 1964
rect 4528 1912 4580 1964
rect 6920 1912 6972 1964
rect 3608 1844 3660 1896
rect 3976 1887 4028 1896
rect 3976 1853 3985 1887
rect 3985 1853 4019 1887
rect 4019 1853 4028 1887
rect 3976 1844 4028 1853
rect 4068 1844 4120 1896
rect 4344 1887 4396 1896
rect 4344 1853 4353 1887
rect 4353 1853 4387 1887
rect 4387 1853 4396 1887
rect 4344 1844 4396 1853
rect 5356 1844 5408 1896
rect 8300 1844 8352 1896
rect 9036 1887 9088 1896
rect 9036 1853 9045 1887
rect 9045 1853 9079 1887
rect 9079 1853 9088 1887
rect 12072 1912 12124 1964
rect 13820 1980 13872 2032
rect 9036 1844 9088 1853
rect 10600 1887 10652 1896
rect 10600 1853 10609 1887
rect 10609 1853 10643 1887
rect 10643 1853 10652 1887
rect 10600 1844 10652 1853
rect 12992 1844 13044 1896
rect 13636 1912 13688 1964
rect 3332 1819 3384 1828
rect 3332 1785 3341 1819
rect 3341 1785 3375 1819
rect 3375 1785 3384 1819
rect 3332 1776 3384 1785
rect 5816 1776 5868 1828
rect 14832 1980 14884 2032
rect 15200 1912 15252 1964
rect 16856 1912 16908 1964
rect 16948 1912 17000 1964
rect 15384 1887 15436 1896
rect 15384 1853 15393 1887
rect 15393 1853 15427 1887
rect 15427 1853 15436 1887
rect 15384 1844 15436 1853
rect 15936 1844 15988 1896
rect 16212 1776 16264 1828
rect 17408 1776 17460 1828
rect 2964 1708 3016 1760
rect 4528 1751 4580 1760
rect 4528 1717 4537 1751
rect 4537 1717 4571 1751
rect 4571 1717 4580 1751
rect 4528 1708 4580 1717
rect 5632 1751 5684 1760
rect 5632 1717 5641 1751
rect 5641 1717 5675 1751
rect 5675 1717 5684 1751
rect 5632 1708 5684 1717
rect 7288 1751 7340 1760
rect 7288 1717 7297 1751
rect 7297 1717 7331 1751
rect 7331 1717 7340 1751
rect 7288 1708 7340 1717
rect 13084 1751 13136 1760
rect 13084 1717 13093 1751
rect 13093 1717 13127 1751
rect 13127 1717 13136 1751
rect 13084 1708 13136 1717
rect 13544 1751 13596 1760
rect 13544 1717 13553 1751
rect 13553 1717 13587 1751
rect 13587 1717 13596 1751
rect 13544 1708 13596 1717
rect 15016 1751 15068 1760
rect 15016 1717 15025 1751
rect 15025 1717 15059 1751
rect 15059 1717 15068 1751
rect 15016 1708 15068 1717
rect 16488 1751 16540 1760
rect 16488 1717 16497 1751
rect 16497 1717 16531 1751
rect 16531 1717 16540 1751
rect 16488 1708 16540 1717
rect 18420 1751 18472 1760
rect 18420 1717 18429 1751
rect 18429 1717 18463 1751
rect 18463 1717 18472 1751
rect 18420 1708 18472 1717
rect 3106 1606 3158 1658
rect 3170 1606 3222 1658
rect 3234 1606 3286 1658
rect 3298 1606 3350 1658
rect 3362 1606 3414 1658
rect 6206 1606 6258 1658
rect 6270 1606 6322 1658
rect 6334 1606 6386 1658
rect 6398 1606 6450 1658
rect 6462 1606 6514 1658
rect 9306 1606 9358 1658
rect 9370 1606 9422 1658
rect 9434 1606 9486 1658
rect 9498 1606 9550 1658
rect 9562 1606 9614 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 12534 1606 12586 1658
rect 12598 1606 12650 1658
rect 12662 1606 12714 1658
rect 15506 1606 15558 1658
rect 15570 1606 15622 1658
rect 15634 1606 15686 1658
rect 15698 1606 15750 1658
rect 15762 1606 15814 1658
rect 18606 1606 18658 1658
rect 18670 1606 18722 1658
rect 18734 1606 18786 1658
rect 18798 1606 18850 1658
rect 18862 1606 18914 1658
rect 2964 1504 3016 1556
rect 5632 1504 5684 1556
rect 7288 1504 7340 1556
rect 8300 1504 8352 1556
rect 13728 1504 13780 1556
rect 15384 1504 15436 1556
rect 15936 1547 15988 1556
rect 15936 1513 15945 1547
rect 15945 1513 15979 1547
rect 15979 1513 15988 1547
rect 15936 1504 15988 1513
rect 16856 1504 16908 1556
rect 3976 1411 4028 1420
rect 3976 1377 3985 1411
rect 3985 1377 4019 1411
rect 4019 1377 4028 1411
rect 3976 1368 4028 1377
rect 4344 1411 4396 1420
rect 4344 1377 4353 1411
rect 4353 1377 4387 1411
rect 4387 1377 4396 1411
rect 4344 1368 4396 1377
rect 14924 1436 14976 1488
rect 5356 1368 5408 1420
rect 8668 1343 8720 1352
rect 8668 1309 8677 1343
rect 8677 1309 8711 1343
rect 8711 1309 8720 1343
rect 8668 1300 8720 1309
rect 10048 1368 10100 1420
rect 10324 1411 10376 1420
rect 10324 1377 10333 1411
rect 10333 1377 10367 1411
rect 10367 1377 10376 1411
rect 13084 1411 13136 1420
rect 10324 1368 10376 1377
rect 13084 1377 13093 1411
rect 13093 1377 13127 1411
rect 13127 1377 13136 1411
rect 13084 1368 13136 1377
rect 13544 1368 13596 1420
rect 15016 1411 15068 1420
rect 15016 1377 15024 1411
rect 15024 1377 15058 1411
rect 15058 1377 15068 1411
rect 15016 1368 15068 1377
rect 16488 1436 16540 1488
rect 16396 1368 16448 1420
rect 14740 1343 14792 1352
rect 14740 1309 14749 1343
rect 14749 1309 14783 1343
rect 14783 1309 14792 1343
rect 14740 1300 14792 1309
rect 16764 1411 16816 1420
rect 16764 1377 16773 1411
rect 16773 1377 16807 1411
rect 16807 1377 16816 1411
rect 16764 1368 16816 1377
rect 17408 1368 17460 1420
rect 17868 1300 17920 1352
rect 3976 1164 4028 1216
rect 17408 1164 17460 1216
rect 1556 1062 1608 1114
rect 1620 1062 1672 1114
rect 1684 1062 1736 1114
rect 1748 1062 1800 1114
rect 1812 1062 1864 1114
rect 4656 1062 4708 1114
rect 4720 1062 4772 1114
rect 4784 1062 4836 1114
rect 4848 1062 4900 1114
rect 4912 1062 4964 1114
rect 7756 1062 7808 1114
rect 7820 1062 7872 1114
rect 7884 1062 7936 1114
rect 7948 1062 8000 1114
rect 8012 1062 8064 1114
rect 10856 1062 10908 1114
rect 10920 1062 10972 1114
rect 10984 1062 11036 1114
rect 11048 1062 11100 1114
rect 11112 1062 11164 1114
rect 13956 1062 14008 1114
rect 14020 1062 14072 1114
rect 14084 1062 14136 1114
rect 14148 1062 14200 1114
rect 14212 1062 14264 1114
rect 17056 1062 17108 1114
rect 17120 1062 17172 1114
rect 17184 1062 17236 1114
rect 17248 1062 17300 1114
rect 17312 1062 17364 1114
rect 3106 518 3158 570
rect 3170 518 3222 570
rect 3234 518 3286 570
rect 3298 518 3350 570
rect 3362 518 3414 570
rect 6206 518 6258 570
rect 6270 518 6322 570
rect 6334 518 6386 570
rect 6398 518 6450 570
rect 6462 518 6514 570
rect 9306 518 9358 570
rect 9370 518 9422 570
rect 9434 518 9486 570
rect 9498 518 9550 570
rect 9562 518 9614 570
rect 12406 518 12458 570
rect 12470 518 12522 570
rect 12534 518 12586 570
rect 12598 518 12650 570
rect 12662 518 12714 570
rect 15506 518 15558 570
rect 15570 518 15622 570
rect 15634 518 15686 570
rect 15698 518 15750 570
rect 15762 518 15814 570
rect 18606 518 18658 570
rect 18670 518 18722 570
rect 18734 518 18786 570
rect 18798 518 18850 570
rect 18862 518 18914 570
<< metal2 >>
rect 1398 19200 1454 20000
rect 4250 19200 4306 20000
rect 7102 19200 7158 20000
rect 9954 19200 10010 20000
rect 12806 19200 12862 20000
rect 15304 19230 15608 19258
rect 1412 18222 1440 19200
rect 1556 18524 1864 18533
rect 1556 18522 1562 18524
rect 1618 18522 1642 18524
rect 1698 18522 1722 18524
rect 1778 18522 1802 18524
rect 1858 18522 1864 18524
rect 1618 18470 1620 18522
rect 1800 18470 1802 18522
rect 1556 18468 1562 18470
rect 1618 18468 1642 18470
rect 1698 18468 1722 18470
rect 1778 18468 1802 18470
rect 1858 18468 1864 18470
rect 1556 18459 1864 18468
rect 4264 18426 4292 19200
rect 4656 18524 4964 18533
rect 4656 18522 4662 18524
rect 4718 18522 4742 18524
rect 4798 18522 4822 18524
rect 4878 18522 4902 18524
rect 4958 18522 4964 18524
rect 4718 18470 4720 18522
rect 4900 18470 4902 18522
rect 4656 18468 4662 18470
rect 4718 18468 4742 18470
rect 4798 18468 4822 18470
rect 4878 18468 4902 18470
rect 4958 18468 4964 18470
rect 4656 18459 4964 18468
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 3106 17980 3414 17989
rect 3106 17978 3112 17980
rect 3168 17978 3192 17980
rect 3248 17978 3272 17980
rect 3328 17978 3352 17980
rect 3408 17978 3414 17980
rect 3168 17926 3170 17978
rect 3350 17926 3352 17978
rect 3106 17924 3112 17926
rect 3168 17924 3192 17926
rect 3248 17924 3272 17926
rect 3328 17924 3352 17926
rect 3408 17924 3414 17926
rect 3106 17915 3414 17924
rect 4264 17814 4292 18362
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 1556 17436 1864 17445
rect 1556 17434 1562 17436
rect 1618 17434 1642 17436
rect 1698 17434 1722 17436
rect 1778 17434 1802 17436
rect 1858 17434 1864 17436
rect 1618 17382 1620 17434
rect 1800 17382 1802 17434
rect 1556 17380 1562 17382
rect 1618 17380 1642 17382
rect 1698 17380 1722 17382
rect 1778 17380 1802 17382
rect 1858 17380 1864 17382
rect 1556 17371 1864 17380
rect 1964 17338 1992 17682
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1124 16992 1176 16998
rect 1124 16934 1176 16940
rect 940 16040 992 16046
rect 940 15982 992 15988
rect 952 15570 980 15982
rect 1136 15706 1164 16934
rect 1556 16348 1864 16357
rect 1556 16346 1562 16348
rect 1618 16346 1642 16348
rect 1698 16346 1722 16348
rect 1778 16346 1802 16348
rect 1858 16346 1864 16348
rect 1618 16294 1620 16346
rect 1800 16294 1802 16346
rect 1556 16292 1562 16294
rect 1618 16292 1642 16294
rect 1698 16292 1722 16294
rect 1778 16292 1802 16294
rect 1858 16292 1864 16294
rect 1556 16283 1864 16292
rect 1400 16176 1452 16182
rect 1400 16118 1452 16124
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 940 15564 992 15570
rect 940 15506 992 15512
rect 952 14550 980 15506
rect 1412 15502 1440 16118
rect 1964 16046 1992 17138
rect 2424 16998 2452 17682
rect 4356 17610 4384 18362
rect 6000 18352 6052 18358
rect 6000 18294 6052 18300
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2608 16574 2636 16934
rect 2516 16546 2636 16574
rect 2516 16114 2544 16546
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15706 1992 15846
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 940 14544 992 14550
rect 940 14486 992 14492
rect 1216 14476 1268 14482
rect 1216 14418 1268 14424
rect 1228 13530 1256 14418
rect 1320 13530 1348 15302
rect 1216 13524 1268 13530
rect 1216 13466 1268 13472
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1412 13326 1440 15438
rect 1556 15260 1864 15269
rect 1556 15258 1562 15260
rect 1618 15258 1642 15260
rect 1698 15258 1722 15260
rect 1778 15258 1802 15260
rect 1858 15258 1864 15260
rect 1618 15206 1620 15258
rect 1800 15206 1802 15258
rect 1556 15204 1562 15206
rect 1618 15204 1642 15206
rect 1698 15204 1722 15206
rect 1778 15204 1802 15206
rect 1858 15204 1864 15206
rect 1556 15195 1864 15204
rect 2056 15162 2084 15914
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1556 14172 1864 14181
rect 1556 14170 1562 14172
rect 1618 14170 1642 14172
rect 1698 14170 1722 14172
rect 1778 14170 1802 14172
rect 1858 14170 1864 14172
rect 1618 14118 1620 14170
rect 1800 14118 1802 14170
rect 1556 14116 1562 14118
rect 1618 14116 1642 14118
rect 1698 14116 1722 14118
rect 1778 14116 1802 14118
rect 1858 14116 1864 14118
rect 1556 14107 1864 14116
rect 2056 13870 2084 14962
rect 2148 14414 2176 16050
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 14890 2360 15846
rect 2700 15162 2728 17274
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2792 16046 2820 16934
rect 2884 16590 2912 17478
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16794 3004 17070
rect 3106 16892 3414 16901
rect 3106 16890 3112 16892
rect 3168 16890 3192 16892
rect 3248 16890 3272 16892
rect 3328 16890 3352 16892
rect 3408 16890 3414 16892
rect 3168 16838 3170 16890
rect 3350 16838 3352 16890
rect 3106 16836 3112 16838
rect 3168 16836 3192 16838
rect 3248 16836 3272 16838
rect 3328 16836 3352 16838
rect 3408 16836 3414 16838
rect 3106 16827 3414 16836
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 2792 14550 2820 15982
rect 3106 15804 3414 15813
rect 3106 15802 3112 15804
rect 3168 15802 3192 15804
rect 3248 15802 3272 15804
rect 3328 15802 3352 15804
rect 3408 15802 3414 15804
rect 3168 15750 3170 15802
rect 3350 15750 3352 15802
rect 3106 15748 3112 15750
rect 3168 15748 3192 15750
rect 3248 15748 3272 15750
rect 3328 15748 3352 15750
rect 3408 15748 3414 15750
rect 3106 15739 3414 15748
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2148 13938 2176 14214
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1556 13084 1864 13093
rect 1556 13082 1562 13084
rect 1618 13082 1642 13084
rect 1698 13082 1722 13084
rect 1778 13082 1802 13084
rect 1858 13082 1864 13084
rect 1618 13030 1620 13082
rect 1800 13030 1802 13082
rect 1556 13028 1562 13030
rect 1618 13028 1642 13030
rect 1698 13028 1722 13030
rect 1778 13028 1802 13030
rect 1858 13028 1864 13030
rect 1556 13019 1864 13028
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12306 1532 12582
rect 1688 12374 1716 12718
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1032 12096 1084 12102
rect 1032 12038 1084 12044
rect 1044 11694 1072 12038
rect 1032 11688 1084 11694
rect 1032 11630 1084 11636
rect 1412 10810 1440 12174
rect 1556 11996 1864 12005
rect 1556 11994 1562 11996
rect 1618 11994 1642 11996
rect 1698 11994 1722 11996
rect 1778 11994 1802 11996
rect 1858 11994 1864 11996
rect 1618 11942 1620 11994
rect 1800 11942 1802 11994
rect 1556 11940 1562 11942
rect 1618 11940 1642 11942
rect 1698 11940 1722 11942
rect 1778 11940 1802 11942
rect 1858 11940 1864 11942
rect 1556 11931 1864 11940
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11354 1624 11494
rect 1964 11354 1992 12718
rect 2056 12306 2084 13806
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1556 10908 1864 10917
rect 1556 10906 1562 10908
rect 1618 10906 1642 10908
rect 1698 10906 1722 10908
rect 1778 10906 1802 10908
rect 1858 10906 1864 10908
rect 1618 10854 1620 10906
rect 1800 10854 1802 10906
rect 1556 10852 1562 10854
rect 1618 10852 1642 10854
rect 1698 10852 1722 10854
rect 1778 10852 1802 10854
rect 1858 10852 1864 10854
rect 1556 10843 1864 10852
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 952 10033 980 10066
rect 938 10024 994 10033
rect 938 9959 994 9968
rect 1412 9654 1440 10746
rect 1556 9820 1864 9829
rect 1556 9818 1562 9820
rect 1618 9818 1642 9820
rect 1698 9818 1722 9820
rect 1778 9818 1802 9820
rect 1858 9818 1864 9820
rect 1618 9766 1620 9818
rect 1800 9766 1802 9818
rect 1556 9764 1562 9766
rect 1618 9764 1642 9766
rect 1698 9764 1722 9766
rect 1778 9764 1802 9766
rect 1858 9764 1864 9766
rect 1556 9755 1864 9764
rect 1400 9648 1452 9654
rect 1964 9602 1992 11154
rect 1400 9590 1452 9596
rect 1412 9450 1440 9590
rect 1780 9586 1992 9602
rect 2056 9586 2084 11494
rect 2148 11286 2176 12582
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10266 2176 11018
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1768 9580 1992 9586
rect 1820 9574 1992 9580
rect 1768 9522 1820 9528
rect 1964 9466 1992 9574
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2148 9518 2176 10202
rect 2240 9994 2268 11086
rect 2424 10130 2452 11698
rect 2884 10826 2912 15506
rect 3804 14890 3832 16662
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3106 14716 3414 14725
rect 3106 14714 3112 14716
rect 3168 14714 3192 14716
rect 3248 14714 3272 14716
rect 3328 14714 3352 14716
rect 3408 14714 3414 14716
rect 3168 14662 3170 14714
rect 3350 14662 3352 14714
rect 3106 14660 3112 14662
rect 3168 14660 3192 14662
rect 3248 14660 3272 14662
rect 3328 14660 3352 14662
rect 3408 14660 3414 14662
rect 3106 14651 3414 14660
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 2976 13394 3004 14350
rect 3528 14074 3556 14350
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3620 14074 3648 14282
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3106 13628 3414 13637
rect 3106 13626 3112 13628
rect 3168 13626 3192 13628
rect 3248 13626 3272 13628
rect 3328 13626 3352 13628
rect 3408 13626 3414 13628
rect 3168 13574 3170 13626
rect 3350 13574 3352 13626
rect 3106 13572 3112 13574
rect 3168 13572 3192 13574
rect 3248 13572 3272 13574
rect 3328 13572 3352 13574
rect 3408 13572 3414 13574
rect 3106 13563 3414 13572
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3620 13326 3648 14010
rect 3804 13802 3832 14826
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 2976 12714 3096 12730
rect 3804 12714 3832 13738
rect 3988 13530 4016 14894
rect 4172 14618 4200 14894
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 2976 12708 3108 12714
rect 2976 12702 3056 12708
rect 2976 11286 3004 12702
rect 3056 12650 3108 12656
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3106 12540 3414 12549
rect 3106 12538 3112 12540
rect 3168 12538 3192 12540
rect 3248 12538 3272 12540
rect 3328 12538 3352 12540
rect 3408 12538 3414 12540
rect 3168 12486 3170 12538
rect 3350 12486 3352 12538
rect 3106 12484 3112 12486
rect 3168 12484 3192 12486
rect 3248 12484 3272 12486
rect 3328 12484 3352 12486
rect 3408 12484 3414 12486
rect 3106 12475 3414 12484
rect 4172 12306 4200 12718
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3106 11452 3414 11461
rect 3106 11450 3112 11452
rect 3168 11450 3192 11452
rect 3248 11450 3272 11452
rect 3328 11450 3352 11452
rect 3408 11450 3414 11452
rect 3168 11398 3170 11450
rect 3350 11398 3352 11450
rect 3106 11396 3112 11398
rect 3168 11396 3192 11398
rect 3248 11396 3272 11398
rect 3328 11396 3352 11398
rect 3408 11396 3414 11398
rect 3106 11387 3414 11396
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2792 10798 2912 10826
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 9654 2268 9930
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 9512 2188 9518
rect 1400 9444 1452 9450
rect 1964 9438 2084 9466
rect 2136 9454 2188 9460
rect 1400 9386 1452 9392
rect 1032 9376 1084 9382
rect 1032 9318 1084 9324
rect 1044 7954 1072 9318
rect 1412 8430 1440 9386
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1556 8732 1864 8741
rect 1556 8730 1562 8732
rect 1618 8730 1642 8732
rect 1698 8730 1722 8732
rect 1778 8730 1802 8732
rect 1858 8730 1864 8732
rect 1618 8678 1620 8730
rect 1800 8678 1802 8730
rect 1556 8676 1562 8678
rect 1618 8676 1642 8678
rect 1698 8676 1722 8678
rect 1778 8676 1802 8678
rect 1858 8676 1864 8678
rect 1556 8667 1864 8676
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1124 8356 1176 8362
rect 1124 8298 1176 8304
rect 1136 8022 1164 8298
rect 1216 8288 1268 8294
rect 1216 8230 1268 8236
rect 1228 8090 1256 8230
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 1124 8016 1176 8022
rect 1124 7958 1176 7964
rect 1032 7948 1084 7954
rect 1032 7890 1084 7896
rect 1228 7002 1256 8026
rect 1556 7644 1864 7653
rect 1556 7642 1562 7644
rect 1618 7642 1642 7644
rect 1698 7642 1722 7644
rect 1778 7642 1802 7644
rect 1858 7642 1864 7644
rect 1618 7590 1620 7642
rect 1800 7590 1802 7642
rect 1556 7588 1562 7590
rect 1618 7588 1642 7590
rect 1698 7588 1722 7590
rect 1778 7588 1802 7590
rect 1858 7588 1864 7590
rect 1556 7579 1864 7588
rect 1216 6996 1268 7002
rect 1216 6938 1268 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6458 1440 6734
rect 1964 6730 1992 9318
rect 2056 9042 2084 9438
rect 2148 9110 2176 9454
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2056 7954 2084 8842
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1556 6556 1864 6565
rect 1556 6554 1562 6556
rect 1618 6554 1642 6556
rect 1698 6554 1722 6556
rect 1778 6554 1802 6556
rect 1858 6554 1864 6556
rect 1618 6502 1620 6554
rect 1800 6502 1802 6554
rect 1556 6500 1562 6502
rect 1618 6500 1642 6502
rect 1698 6500 1722 6502
rect 1778 6500 1802 6502
rect 1858 6500 1864 6502
rect 1556 6491 1864 6500
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 2056 5914 2084 7890
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1556 5468 1864 5477
rect 1556 5466 1562 5468
rect 1618 5466 1642 5468
rect 1698 5466 1722 5468
rect 1778 5466 1802 5468
rect 1858 5466 1864 5468
rect 1618 5414 1620 5466
rect 1800 5414 1802 5466
rect 1556 5412 1562 5414
rect 1618 5412 1642 5414
rect 1698 5412 1722 5414
rect 1778 5412 1802 5414
rect 1858 5412 1864 5414
rect 1556 5403 1864 5412
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 848 5160 900 5166
rect 848 5102 900 5108
rect 860 4826 888 5102
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 1596 4690 1624 5306
rect 940 4684 992 4690
rect 940 4626 992 4632
rect 1032 4684 1084 4690
rect 1032 4626 1084 4632
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 952 3942 980 4626
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 1044 3194 1072 4626
rect 1556 4380 1864 4389
rect 1556 4378 1562 4380
rect 1618 4378 1642 4380
rect 1698 4378 1722 4380
rect 1778 4378 1802 4380
rect 1858 4378 1864 4380
rect 1618 4326 1620 4378
rect 1800 4326 1802 4378
rect 1556 4324 1562 4326
rect 1618 4324 1642 4326
rect 1698 4324 1722 4326
rect 1778 4324 1802 4326
rect 1858 4324 1864 4326
rect 1556 4315 1864 4324
rect 1964 4146 1992 5714
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5370 2084 5510
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2148 5302 2176 7210
rect 2240 6458 2268 9590
rect 2332 8634 2360 9998
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2424 8430 2452 10066
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 8498 2728 9454
rect 2792 9450 2820 10798
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2884 9654 2912 10610
rect 2976 10470 3004 11222
rect 4172 11014 4200 12242
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3620 10606 3648 10950
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3106 10364 3414 10373
rect 3106 10362 3112 10364
rect 3168 10362 3192 10364
rect 3248 10362 3272 10364
rect 3328 10362 3352 10364
rect 3408 10362 3414 10364
rect 3168 10310 3170 10362
rect 3350 10310 3352 10362
rect 3106 10308 3112 10310
rect 3168 10308 3192 10310
rect 3248 10308 3272 10310
rect 3328 10308 3352 10310
rect 3408 10308 3414 10310
rect 3106 10299 3414 10308
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4264 10198 4292 11086
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4356 9926 4384 17546
rect 4656 17436 4964 17445
rect 4656 17434 4662 17436
rect 4718 17434 4742 17436
rect 4798 17434 4822 17436
rect 4878 17434 4902 17436
rect 4958 17434 4964 17436
rect 4718 17382 4720 17434
rect 4900 17382 4902 17434
rect 4656 17380 4662 17382
rect 4718 17380 4742 17382
rect 4798 17380 4822 17382
rect 4878 17380 4902 17382
rect 4958 17380 4964 17382
rect 4656 17371 4964 17380
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4448 17134 4476 17274
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4448 16794 4476 17070
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16114 4476 16390
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4448 15026 4476 16050
rect 4540 16046 4568 16934
rect 4656 16348 4964 16357
rect 4656 16346 4662 16348
rect 4718 16346 4742 16348
rect 4798 16346 4822 16348
rect 4878 16346 4902 16348
rect 4958 16346 4964 16348
rect 4718 16294 4720 16346
rect 4900 16294 4902 16346
rect 4656 16292 4662 16294
rect 4718 16292 4742 16294
rect 4798 16292 4822 16294
rect 4878 16292 4902 16294
rect 4958 16292 4964 16294
rect 4656 16283 4964 16292
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4656 15260 4964 15269
rect 4656 15258 4662 15260
rect 4718 15258 4742 15260
rect 4798 15258 4822 15260
rect 4878 15258 4902 15260
rect 4958 15258 4964 15260
rect 4718 15206 4720 15258
rect 4900 15206 4902 15258
rect 4656 15204 4662 15206
rect 4718 15204 4742 15206
rect 4798 15204 4822 15206
rect 4878 15204 4902 15206
rect 4958 15204 4964 15206
rect 4656 15195 4964 15204
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4448 14482 4476 14962
rect 5000 14958 5028 18022
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5092 16794 5120 17002
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5184 16726 5212 17682
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17134 5304 17478
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5368 16998 5396 17546
rect 5460 16998 5488 18090
rect 5736 17338 5764 18090
rect 5724 17332 5776 17338
rect 5776 17292 5856 17320
rect 5724 17274 5776 17280
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5736 16250 5764 16730
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5736 14958 5764 16186
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 13938 4476 14418
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4448 13394 4476 13874
rect 4540 13870 4568 14758
rect 5552 14550 5580 14758
rect 5828 14550 5856 17292
rect 6012 17134 6040 18294
rect 6206 17980 6514 17989
rect 6206 17978 6212 17980
rect 6268 17978 6292 17980
rect 6348 17978 6372 17980
rect 6428 17978 6452 17980
rect 6508 17978 6514 17980
rect 6268 17926 6270 17978
rect 6450 17926 6452 17978
rect 6206 17924 6212 17926
rect 6268 17924 6292 17926
rect 6348 17924 6372 17926
rect 6428 17924 6452 17926
rect 6508 17924 6514 17926
rect 6206 17915 6514 17924
rect 7116 17218 7144 19200
rect 7756 18524 8064 18533
rect 7756 18522 7762 18524
rect 7818 18522 7842 18524
rect 7898 18522 7922 18524
rect 7978 18522 8002 18524
rect 8058 18522 8064 18524
rect 7818 18470 7820 18522
rect 8000 18470 8002 18522
rect 7756 18468 7762 18470
rect 7818 18468 7842 18470
rect 7898 18468 7922 18470
rect 7978 18468 8002 18470
rect 8058 18468 8064 18470
rect 7756 18459 8064 18468
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 7852 17746 7880 18090
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7756 17436 8064 17445
rect 7756 17434 7762 17436
rect 7818 17434 7842 17436
rect 7898 17434 7922 17436
rect 7978 17434 8002 17436
rect 8058 17434 8064 17436
rect 7818 17382 7820 17434
rect 8000 17382 8002 17434
rect 7756 17380 7762 17382
rect 7818 17380 7842 17382
rect 7898 17380 7922 17382
rect 7978 17380 8002 17382
rect 8058 17380 8064 17382
rect 7756 17371 8064 17380
rect 7116 17190 7236 17218
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6206 16892 6514 16901
rect 6206 16890 6212 16892
rect 6268 16890 6292 16892
rect 6348 16890 6372 16892
rect 6428 16890 6452 16892
rect 6508 16890 6514 16892
rect 6268 16838 6270 16890
rect 6450 16838 6452 16890
rect 6206 16836 6212 16838
rect 6268 16836 6292 16838
rect 6348 16836 6372 16838
rect 6428 16836 6452 16838
rect 6508 16836 6514 16838
rect 6206 16827 6514 16836
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16046 6868 16390
rect 7208 16046 7236 17190
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7484 16114 7512 17138
rect 8128 17082 8156 18090
rect 8036 17066 8156 17082
rect 8024 17060 8156 17066
rect 8076 17054 8156 17060
rect 8024 17002 8076 17008
rect 8128 16726 8156 17054
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 7756 16348 8064 16357
rect 7756 16346 7762 16348
rect 7818 16346 7842 16348
rect 7898 16346 7922 16348
rect 7978 16346 8002 16348
rect 8058 16346 8064 16348
rect 7818 16294 7820 16346
rect 8000 16294 8002 16346
rect 7756 16292 7762 16294
rect 7818 16292 7842 16294
rect 7898 16292 7922 16294
rect 7978 16292 8002 16294
rect 8058 16292 8064 16294
rect 7756 16283 8064 16292
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6206 15804 6514 15813
rect 6206 15802 6212 15804
rect 6268 15802 6292 15804
rect 6348 15802 6372 15804
rect 6428 15802 6452 15804
rect 6508 15802 6514 15804
rect 6268 15750 6270 15802
rect 6450 15750 6452 15802
rect 6206 15748 6212 15750
rect 6268 15748 6292 15750
rect 6348 15748 6372 15750
rect 6428 15748 6452 15750
rect 6508 15748 6514 15750
rect 6206 15739 6514 15748
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6206 14716 6514 14725
rect 6206 14714 6212 14716
rect 6268 14714 6292 14716
rect 6348 14714 6372 14716
rect 6428 14714 6452 14716
rect 6508 14714 6514 14716
rect 6268 14662 6270 14714
rect 6450 14662 6452 14714
rect 6206 14660 6212 14662
rect 6268 14660 6292 14662
rect 6348 14660 6372 14662
rect 6428 14660 6452 14662
rect 6508 14660 6514 14662
rect 6206 14651 6514 14660
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 4656 14172 4964 14181
rect 4656 14170 4662 14172
rect 4718 14170 4742 14172
rect 4798 14170 4822 14172
rect 4878 14170 4902 14172
rect 4958 14170 4964 14172
rect 4718 14118 4720 14170
rect 4900 14118 4902 14170
rect 4656 14116 4662 14118
rect 4718 14116 4742 14118
rect 4798 14116 4822 14118
rect 4878 14116 4902 14118
rect 4958 14116 4964 14118
rect 4656 14107 4964 14116
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 5828 13802 5856 14486
rect 6932 14074 6960 14826
rect 7024 14618 7052 15846
rect 7208 15706 7236 15982
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7300 13938 7328 16050
rect 7756 15260 8064 15269
rect 7756 15258 7762 15260
rect 7818 15258 7842 15260
rect 7898 15258 7922 15260
rect 7978 15258 8002 15260
rect 8058 15258 8064 15260
rect 7818 15206 7820 15258
rect 8000 15206 8002 15258
rect 7756 15204 7762 15206
rect 7818 15204 7842 15206
rect 7898 15204 7922 15206
rect 7978 15204 8002 15206
rect 8058 15204 8064 15206
rect 7756 15195 8064 15204
rect 8128 14890 8156 16662
rect 8220 15978 8248 18158
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17678 8340 18022
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8404 16794 8432 18158
rect 8680 17814 8708 18226
rect 9680 18216 9732 18222
rect 9968 18170 9996 19200
rect 10856 18524 11164 18533
rect 10856 18522 10862 18524
rect 10918 18522 10942 18524
rect 10998 18522 11022 18524
rect 11078 18522 11102 18524
rect 11158 18522 11164 18524
rect 10918 18470 10920 18522
rect 11100 18470 11102 18522
rect 10856 18468 10862 18470
rect 10918 18468 10942 18470
rect 10998 18468 11022 18470
rect 11078 18468 11102 18470
rect 11158 18468 11164 18470
rect 10856 18459 11164 18468
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 9680 18158 9732 18164
rect 9306 17980 9614 17989
rect 9306 17978 9312 17980
rect 9368 17978 9392 17980
rect 9448 17978 9472 17980
rect 9528 17978 9552 17980
rect 9608 17978 9614 17980
rect 9368 17926 9370 17978
rect 9550 17926 9552 17978
rect 9306 17924 9312 17926
rect 9368 17924 9392 17926
rect 9448 17924 9472 17926
rect 9528 17924 9552 17926
rect 9608 17924 9614 17926
rect 9306 17915 9614 17924
rect 9692 17882 9720 18158
rect 9876 18142 9996 18170
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8220 15706 8248 15914
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8128 14550 8156 14826
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7756 14172 8064 14181
rect 7756 14170 7762 14172
rect 7818 14170 7842 14172
rect 7898 14170 7922 14172
rect 7978 14170 8002 14172
rect 8058 14170 8064 14172
rect 7818 14118 7820 14170
rect 8000 14118 8002 14170
rect 7756 14116 7762 14118
rect 7818 14116 7842 14118
rect 7898 14116 7922 14118
rect 7978 14116 8002 14118
rect 8058 14116 8064 14118
rect 7756 14107 8064 14116
rect 8312 14074 8340 14350
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 4448 12986 4476 13330
rect 4656 13084 4964 13093
rect 4656 13082 4662 13084
rect 4718 13082 4742 13084
rect 4798 13082 4822 13084
rect 4878 13082 4902 13084
rect 4958 13082 4964 13084
rect 4718 13030 4720 13082
rect 4900 13030 4902 13082
rect 4656 13028 4662 13030
rect 4718 13028 4742 13030
rect 4798 13028 4822 13030
rect 4878 13028 4902 13030
rect 4958 13028 4964 13030
rect 4656 13019 4964 13028
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 5276 12442 5304 13330
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5368 12374 5396 13398
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4656 11996 4964 12005
rect 4656 11994 4662 11996
rect 4718 11994 4742 11996
rect 4798 11994 4822 11996
rect 4878 11994 4902 11996
rect 4958 11994 4964 11996
rect 4718 11942 4720 11994
rect 4900 11942 4902 11994
rect 4656 11940 4662 11942
rect 4718 11940 4742 11942
rect 4798 11940 4822 11942
rect 4878 11940 4902 11942
rect 4958 11940 4964 11942
rect 4656 11931 4964 11940
rect 5368 11778 5396 12310
rect 5460 12306 5488 12582
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5276 11750 5396 11778
rect 5276 11694 5304 11750
rect 5460 11694 5488 12242
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 4656 10908 4964 10917
rect 4656 10906 4662 10908
rect 4718 10906 4742 10908
rect 4798 10906 4822 10908
rect 4878 10906 4902 10908
rect 4958 10906 4964 10908
rect 4718 10854 4720 10906
rect 4900 10854 4902 10906
rect 4656 10852 4662 10854
rect 4718 10852 4742 10854
rect 4798 10852 4822 10854
rect 4878 10852 4902 10854
rect 4958 10852 4964 10854
rect 4656 10843 4964 10852
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 9110 2820 9386
rect 2884 9178 2912 9454
rect 3106 9276 3414 9285
rect 3106 9274 3112 9276
rect 3168 9274 3192 9276
rect 3248 9274 3272 9276
rect 3328 9274 3352 9276
rect 3408 9274 3414 9276
rect 3168 9222 3170 9274
rect 3350 9222 3352 9274
rect 3106 9220 3112 9222
rect 3168 9220 3192 9222
rect 3248 9220 3272 9222
rect 3328 9220 3352 9222
rect 3408 9220 3414 9222
rect 3106 9211 3414 9220
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 3436 8430 3464 8842
rect 4172 8498 4200 8978
rect 4448 8974 4476 9862
rect 4656 9820 4964 9829
rect 4656 9818 4662 9820
rect 4718 9818 4742 9820
rect 4798 9818 4822 9820
rect 4878 9818 4902 9820
rect 4958 9818 4964 9820
rect 4718 9766 4720 9818
rect 4900 9766 4902 9818
rect 4656 9764 4662 9766
rect 4718 9764 4742 9766
rect 4798 9764 4822 9766
rect 4878 9764 4902 9766
rect 4958 9764 4964 9766
rect 4656 9755 4964 9764
rect 5000 9518 5028 10406
rect 5460 10266 5488 11086
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 10130 5580 12038
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4632 9042 4660 9318
rect 4724 9042 4752 9318
rect 5460 9178 5488 10066
rect 5644 9178 5672 12650
rect 5828 12434 5856 13738
rect 6206 13628 6514 13637
rect 6206 13626 6212 13628
rect 6268 13626 6292 13628
rect 6348 13626 6372 13628
rect 6428 13626 6452 13628
rect 6508 13626 6514 13628
rect 6268 13574 6270 13626
rect 6450 13574 6452 13626
rect 6206 13572 6212 13574
rect 6268 13572 6292 13574
rect 6348 13572 6372 13574
rect 6428 13572 6452 13574
rect 6508 13572 6514 13574
rect 6206 13563 6514 13572
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6206 12540 6514 12549
rect 6206 12538 6212 12540
rect 6268 12538 6292 12540
rect 6348 12538 6372 12540
rect 6428 12538 6452 12540
rect 6508 12538 6514 12540
rect 6268 12486 6270 12538
rect 6450 12486 6452 12538
rect 6206 12484 6212 12486
rect 6268 12484 6292 12486
rect 6348 12484 6372 12486
rect 6428 12484 6452 12486
rect 6508 12484 6514 12486
rect 6206 12475 6514 12484
rect 5736 12406 5856 12434
rect 5736 12170 5764 12406
rect 6656 12374 6684 13126
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11286 5764 12106
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 2424 6866 2452 8366
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3106 8188 3414 8197
rect 3106 8186 3112 8188
rect 3168 8186 3192 8188
rect 3248 8186 3272 8188
rect 3328 8186 3352 8188
rect 3408 8186 3414 8188
rect 3168 8134 3170 8186
rect 3350 8134 3352 8186
rect 3106 8132 3112 8134
rect 3168 8132 3192 8134
rect 3248 8132 3272 8134
rect 3328 8132 3352 8134
rect 3408 8132 3414 8134
rect 3106 8123 3414 8132
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 6866 2912 7346
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3106 7100 3414 7109
rect 3106 7098 3112 7100
rect 3168 7098 3192 7100
rect 3248 7098 3272 7100
rect 3328 7098 3352 7100
rect 3408 7098 3414 7100
rect 3168 7046 3170 7098
rect 3350 7046 3352 7098
rect 3106 7044 3112 7046
rect 3168 7044 3192 7046
rect 3248 7044 3272 7046
rect 3328 7044 3352 7046
rect 3408 7044 3414 7046
rect 3106 7035 3414 7044
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 5710 2268 6258
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2240 5148 2268 5646
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5166 2728 5578
rect 2792 5352 2820 6734
rect 2884 6662 2912 6802
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 3106 6012 3414 6021
rect 3106 6010 3112 6012
rect 3168 6010 3192 6012
rect 3248 6010 3272 6012
rect 3328 6010 3352 6012
rect 3408 6010 3414 6012
rect 3168 5958 3170 6010
rect 3350 5958 3352 6010
rect 3106 5956 3112 5958
rect 3168 5956 3192 5958
rect 3248 5956 3272 5958
rect 3328 5956 3352 5958
rect 3408 5956 3414 5958
rect 3106 5947 3414 5956
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3252 5642 3280 5714
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 2792 5324 2912 5352
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2056 5120 2268 5148
rect 2688 5160 2740 5166
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2056 3942 2084 5120
rect 2688 5102 2740 5108
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2608 4282 2636 4558
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1556 3292 1864 3301
rect 1556 3290 1562 3292
rect 1618 3290 1642 3292
rect 1698 3290 1722 3292
rect 1778 3290 1802 3292
rect 1858 3290 1864 3292
rect 1618 3238 1620 3290
rect 1800 3238 1802 3290
rect 1556 3236 1562 3238
rect 1618 3236 1642 3238
rect 1698 3236 1722 3238
rect 1778 3236 1802 3238
rect 1858 3236 1864 3238
rect 1556 3227 1864 3236
rect 1964 3194 1992 3878
rect 1032 3188 1084 3194
rect 1032 3130 1084 3136
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2056 2990 2084 3878
rect 1032 2984 1084 2990
rect 1032 2926 1084 2932
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1044 2650 1072 2926
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1032 2644 1084 2650
rect 1032 2586 1084 2592
rect 1556 2204 1864 2213
rect 1556 2202 1562 2204
rect 1618 2202 1642 2204
rect 1698 2202 1722 2204
rect 1778 2202 1802 2204
rect 1858 2202 1864 2204
rect 1618 2150 1620 2202
rect 1800 2150 1802 2202
rect 1556 2148 1562 2150
rect 1618 2148 1642 2150
rect 1698 2148 1722 2150
rect 1778 2148 1802 2150
rect 1858 2148 1864 2150
rect 1556 2139 1864 2148
rect 1964 2106 1992 2790
rect 2332 2446 2360 4082
rect 2700 4078 2728 5102
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3602 2728 4014
rect 2792 3738 2820 5170
rect 2884 4826 2912 5324
rect 3106 4924 3414 4933
rect 3106 4922 3112 4924
rect 3168 4922 3192 4924
rect 3248 4922 3272 4924
rect 3328 4922 3352 4924
rect 3408 4922 3414 4924
rect 3168 4870 3170 4922
rect 3350 4870 3352 4922
rect 3106 4868 3112 4870
rect 3168 4868 3192 4870
rect 3248 4868 3272 4870
rect 3328 4868 3352 4870
rect 3408 4868 3414 4870
rect 3106 4859 3414 4868
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2884 3942 2912 4150
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3106 3836 3414 3845
rect 3106 3834 3112 3836
rect 3168 3834 3192 3836
rect 3248 3834 3272 3836
rect 3328 3834 3352 3836
rect 3408 3834 3414 3836
rect 3168 3782 3170 3834
rect 3350 3782 3352 3834
rect 3106 3780 3112 3782
rect 3168 3780 3192 3782
rect 3248 3780 3272 3782
rect 3328 3780 3352 3782
rect 3408 3780 3414 3782
rect 3106 3771 3414 3780
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3528 3602 3556 4014
rect 3620 3738 3648 7142
rect 3804 6118 3832 8298
rect 4448 7546 4476 8910
rect 4656 8732 4964 8741
rect 4656 8730 4662 8732
rect 4718 8730 4742 8732
rect 4798 8730 4822 8732
rect 4878 8730 4902 8732
rect 4958 8730 4964 8732
rect 4718 8678 4720 8730
rect 4900 8678 4902 8730
rect 4656 8676 4662 8678
rect 4718 8676 4742 8678
rect 4798 8676 4822 8678
rect 4878 8676 4902 8678
rect 4958 8676 4964 8678
rect 4656 8667 4964 8676
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5184 7834 5212 8434
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 7954 5304 8298
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4656 7644 4964 7653
rect 4656 7642 4662 7644
rect 4718 7642 4742 7644
rect 4798 7642 4822 7644
rect 4878 7642 4902 7644
rect 4958 7642 4964 7644
rect 4718 7590 4720 7642
rect 4900 7590 4902 7642
rect 4656 7588 4662 7590
rect 4718 7588 4742 7590
rect 4798 7588 4822 7590
rect 4878 7588 4902 7590
rect 4958 7588 4964 7590
rect 4656 7579 4964 7588
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6934 4200 7210
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5710 3832 6054
rect 3896 5778 3924 6190
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3804 5148 3832 5646
rect 3896 5302 3924 5714
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3884 5160 3936 5166
rect 3804 5120 3884 5148
rect 3884 5102 3936 5108
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 1952 2100 2004 2106
rect 1952 2042 2004 2048
rect 2792 1970 2820 2994
rect 2976 2990 3004 3538
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3106 2748 3414 2757
rect 3106 2746 3112 2748
rect 3168 2746 3192 2748
rect 3248 2746 3272 2748
rect 3328 2746 3352 2748
rect 3408 2746 3414 2748
rect 3168 2694 3170 2746
rect 3350 2694 3352 2746
rect 3106 2692 3112 2694
rect 3168 2692 3192 2694
rect 3248 2692 3272 2694
rect 3328 2692 3352 2694
rect 3408 2692 3414 2694
rect 3106 2683 3414 2692
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2884 2106 2912 2450
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 3344 1834 3372 2518
rect 3620 1902 3648 3674
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3712 2990 3740 3538
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3896 2582 3924 5102
rect 4172 4214 4200 6666
rect 4656 6556 4964 6565
rect 4656 6554 4662 6556
rect 4718 6554 4742 6556
rect 4798 6554 4822 6556
rect 4878 6554 4902 6556
rect 4958 6554 4964 6556
rect 4718 6502 4720 6554
rect 4900 6502 4902 6554
rect 4656 6500 4662 6502
rect 4718 6500 4742 6502
rect 4798 6500 4822 6502
rect 4878 6500 4902 6502
rect 4958 6500 4964 6502
rect 4656 6491 4964 6500
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5166 4292 5510
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4160 4208 4212 4214
rect 4080 4168 4160 4196
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 4080 2514 4108 4168
rect 4160 4150 4212 4156
rect 4264 3738 4292 4626
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3194 4200 3538
rect 4356 3466 4384 5714
rect 4448 5166 4476 5782
rect 4540 5370 4568 6258
rect 4656 5468 4964 5477
rect 4656 5466 4662 5468
rect 4718 5466 4742 5468
rect 4798 5466 4822 5468
rect 4878 5466 4902 5468
rect 4958 5466 4964 5468
rect 4718 5414 4720 5466
rect 4900 5414 4902 5466
rect 4656 5412 4662 5414
rect 4718 5412 4742 5414
rect 4798 5412 4822 5414
rect 4878 5412 4902 5414
rect 4958 5412 4964 5414
rect 4656 5403 4964 5412
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4080 1902 4108 2450
rect 4540 1970 4568 4966
rect 4724 4690 4752 4966
rect 4816 4690 4844 5034
rect 5000 4826 5028 7822
rect 5184 7806 5304 7834
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5092 5642 5120 7482
rect 5276 7342 5304 7806
rect 5644 7546 5672 9114
rect 5736 8430 5764 9454
rect 5828 8906 5856 12242
rect 6380 11830 6408 12242
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6206 11452 6514 11461
rect 6206 11450 6212 11452
rect 6268 11450 6292 11452
rect 6348 11450 6372 11452
rect 6428 11450 6452 11452
rect 6508 11450 6514 11452
rect 6268 11398 6270 11450
rect 6450 11398 6452 11450
rect 6206 11396 6212 11398
rect 6268 11396 6292 11398
rect 6348 11396 6372 11398
rect 6428 11396 6452 11398
rect 6508 11396 6514 11398
rect 6206 11387 6514 11396
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6564 10606 6592 10950
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5920 9042 5948 10474
rect 6206 10364 6514 10373
rect 6206 10362 6212 10364
rect 6268 10362 6292 10364
rect 6348 10362 6372 10364
rect 6428 10362 6452 10364
rect 6508 10362 6514 10364
rect 6268 10310 6270 10362
rect 6450 10310 6452 10362
rect 6206 10308 6212 10310
rect 6268 10308 6292 10310
rect 6348 10308 6372 10310
rect 6428 10308 6452 10310
rect 6508 10308 6514 10310
rect 6206 10299 6514 10308
rect 6564 9518 6592 10542
rect 6932 10130 6960 10950
rect 7024 10198 7052 11494
rect 7116 10470 7144 13806
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6206 9276 6514 9285
rect 6206 9274 6212 9276
rect 6268 9274 6292 9276
rect 6348 9274 6372 9276
rect 6428 9274 6452 9276
rect 6508 9274 6514 9276
rect 6268 9222 6270 9274
rect 6450 9222 6452 9274
rect 6206 9220 6212 9222
rect 6268 9220 6292 9222
rect 6348 9220 6372 9222
rect 6428 9220 6452 9222
rect 6508 9220 6514 9222
rect 6206 9211 6514 9220
rect 6656 9042 6684 9386
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5828 8566 5856 8842
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5276 6322 5304 7278
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4656 4380 4964 4389
rect 4656 4378 4662 4380
rect 4718 4378 4742 4380
rect 4798 4378 4822 4380
rect 4878 4378 4902 4380
rect 4958 4378 4964 4380
rect 4718 4326 4720 4378
rect 4900 4326 4902 4378
rect 4656 4324 4662 4326
rect 4718 4324 4742 4326
rect 4798 4324 4822 4326
rect 4878 4324 4902 4326
rect 4958 4324 4964 4326
rect 4656 4315 4964 4324
rect 5092 4282 5120 5578
rect 5184 5370 5212 5646
rect 5276 5556 5304 6258
rect 5368 6254 5396 7482
rect 5736 6662 5764 8366
rect 5920 7426 5948 8978
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5828 7410 5948 7426
rect 5828 7404 5960 7410
rect 5828 7398 5908 7404
rect 5828 6662 5856 7398
rect 5908 7346 5960 7352
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 5658 5396 6190
rect 5552 6118 5580 6326
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5368 5630 5488 5658
rect 5356 5568 5408 5574
rect 5276 5528 5356 5556
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5276 5234 5304 5528
rect 5356 5510 5408 5516
rect 5264 5228 5316 5234
rect 5460 5216 5488 5630
rect 5264 5170 5316 5176
rect 5368 5188 5488 5216
rect 5368 4826 5396 5188
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5184 3738 5212 4694
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5460 3602 5488 5034
rect 5644 5012 5672 6394
rect 5736 6186 5764 6598
rect 5828 6390 5856 6598
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5828 6254 5856 6326
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5736 5166 5764 6122
rect 5920 5846 5948 7210
rect 6012 6390 6040 8842
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6206 8188 6514 8197
rect 6206 8186 6212 8188
rect 6268 8186 6292 8188
rect 6348 8186 6372 8188
rect 6428 8186 6452 8188
rect 6508 8186 6514 8188
rect 6268 8134 6270 8186
rect 6450 8134 6452 8186
rect 6206 8132 6212 8134
rect 6268 8132 6292 8134
rect 6348 8132 6372 8134
rect 6428 8132 6452 8134
rect 6508 8132 6514 8134
rect 6206 8123 6514 8132
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6564 7274 6592 7958
rect 6932 7886 6960 8366
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6206 7100 6514 7109
rect 6206 7098 6212 7100
rect 6268 7098 6292 7100
rect 6348 7098 6372 7100
rect 6428 7098 6452 7100
rect 6508 7098 6514 7100
rect 6268 7046 6270 7098
rect 6450 7046 6452 7098
rect 6206 7044 6212 7046
rect 6268 7044 6292 7046
rect 6348 7044 6372 7046
rect 6428 7044 6452 7046
rect 6508 7044 6514 7046
rect 6206 7035 6514 7044
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5644 4984 5764 5012
rect 5736 4486 5764 4984
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4078 5764 4422
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 4656 3292 4964 3301
rect 4656 3290 4662 3292
rect 4718 3290 4742 3292
rect 4798 3290 4822 3292
rect 4878 3290 4902 3292
rect 4958 3290 4964 3292
rect 4718 3238 4720 3290
rect 4900 3238 4902 3290
rect 4656 3236 4662 3238
rect 4718 3236 4742 3238
rect 4798 3236 4822 3238
rect 4878 3236 4902 3238
rect 4958 3236 4964 3238
rect 4656 3227 4964 3236
rect 5276 3194 5304 3538
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5368 2514 5396 2926
rect 5552 2650 5580 3470
rect 5644 3058 5672 3538
rect 5736 3398 5764 4014
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 4656 2204 4964 2213
rect 4656 2202 4662 2204
rect 4718 2202 4742 2204
rect 4798 2202 4822 2204
rect 4878 2202 4902 2204
rect 4958 2202 4964 2204
rect 4718 2150 4720 2202
rect 4900 2150 4902 2202
rect 4656 2148 4662 2150
rect 4718 2148 4742 2150
rect 4798 2148 4822 2150
rect 4878 2148 4902 2150
rect 4958 2148 4964 2150
rect 4656 2139 4964 2148
rect 4528 1964 4580 1970
rect 4528 1906 4580 1912
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3976 1896 4028 1902
rect 3976 1838 4028 1844
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4344 1896 4396 1902
rect 4344 1838 4396 1844
rect 3332 1828 3384 1834
rect 3332 1770 3384 1776
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2976 1562 3004 1702
rect 3106 1660 3414 1669
rect 3106 1658 3112 1660
rect 3168 1658 3192 1660
rect 3248 1658 3272 1660
rect 3328 1658 3352 1660
rect 3408 1658 3414 1660
rect 3168 1606 3170 1658
rect 3350 1606 3352 1658
rect 3106 1604 3112 1606
rect 3168 1604 3192 1606
rect 3248 1604 3272 1606
rect 3328 1604 3352 1606
rect 3408 1604 3414 1606
rect 3106 1595 3414 1604
rect 2964 1556 3016 1562
rect 2964 1498 3016 1504
rect 3988 1426 4016 1838
rect 4356 1426 4384 1838
rect 4540 1766 4568 1906
rect 5368 1902 5396 2450
rect 5644 2106 5672 2790
rect 5736 2446 5764 3334
rect 5828 2990 5856 4762
rect 6012 4758 6040 6326
rect 6656 6322 6684 6598
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6206 6012 6514 6021
rect 6206 6010 6212 6012
rect 6268 6010 6292 6012
rect 6348 6010 6372 6012
rect 6428 6010 6452 6012
rect 6508 6010 6514 6012
rect 6268 5958 6270 6010
rect 6450 5958 6452 6010
rect 6206 5956 6212 5958
rect 6268 5956 6292 5958
rect 6348 5956 6372 5958
rect 6428 5956 6452 5958
rect 6508 5956 6514 5958
rect 6206 5947 6514 5956
rect 6206 4924 6514 4933
rect 6206 4922 6212 4924
rect 6268 4922 6292 4924
rect 6348 4922 6372 4924
rect 6428 4922 6452 4924
rect 6508 4922 6514 4924
rect 6268 4870 6270 4922
rect 6450 4870 6452 4922
rect 6206 4868 6212 4870
rect 6268 4868 6292 4870
rect 6348 4868 6372 4870
rect 6428 4868 6452 4870
rect 6508 4868 6514 4870
rect 6206 4859 6514 4868
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5828 2106 5856 2926
rect 6012 2650 6040 4082
rect 6656 3942 6684 6122
rect 6840 5710 6868 6666
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6932 5166 6960 7822
rect 7024 6866 7052 10134
rect 7208 9178 7236 10610
rect 7300 10606 7328 13330
rect 7668 12170 7696 13874
rect 7756 13084 8064 13093
rect 7756 13082 7762 13084
rect 7818 13082 7842 13084
rect 7898 13082 7922 13084
rect 7978 13082 8002 13084
rect 8058 13082 8064 13084
rect 7818 13030 7820 13082
rect 8000 13030 8002 13082
rect 7756 13028 7762 13030
rect 7818 13028 7842 13030
rect 7898 13028 7922 13030
rect 7978 13028 8002 13030
rect 8058 13028 8064 13030
rect 7756 13019 8064 13028
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8588 12238 8616 12310
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7756 11996 8064 12005
rect 7756 11994 7762 11996
rect 7818 11994 7842 11996
rect 7898 11994 7922 11996
rect 7978 11994 8002 11996
rect 8058 11994 8064 11996
rect 7818 11942 7820 11994
rect 8000 11942 8002 11994
rect 7756 11940 7762 11942
rect 7818 11940 7842 11942
rect 7898 11940 7922 11942
rect 7978 11940 8002 11942
rect 8058 11940 8064 11942
rect 7756 11931 8064 11940
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8220 11354 8248 11562
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8588 11286 8616 12174
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 7756 10908 8064 10917
rect 7756 10906 7762 10908
rect 7818 10906 7842 10908
rect 7898 10906 7922 10908
rect 7978 10906 8002 10908
rect 8058 10906 8064 10908
rect 7818 10854 7820 10906
rect 8000 10854 8002 10906
rect 7756 10852 7762 10854
rect 7818 10852 7842 10854
rect 7898 10852 7922 10854
rect 7978 10852 8002 10854
rect 8058 10852 8064 10854
rect 7756 10843 8064 10852
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7300 9994 7328 10542
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7576 7546 7604 8026
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7576 7274 7604 7482
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7668 6866 7696 9998
rect 7756 9820 8064 9829
rect 7756 9818 7762 9820
rect 7818 9818 7842 9820
rect 7898 9818 7922 9820
rect 7978 9818 8002 9820
rect 8058 9818 8064 9820
rect 7818 9766 7820 9818
rect 8000 9766 8002 9818
rect 7756 9764 7762 9766
rect 7818 9764 7842 9766
rect 7898 9764 7922 9766
rect 7978 9764 8002 9766
rect 8058 9764 8064 9766
rect 7756 9755 8064 9764
rect 8128 9042 8156 10474
rect 8680 9450 8708 17750
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 16114 8800 16934
rect 9048 16250 9076 17002
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16250 9168 16526
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 9232 15162 9260 17614
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9306 16892 9614 16901
rect 9306 16890 9312 16892
rect 9368 16890 9392 16892
rect 9448 16890 9472 16892
rect 9528 16890 9552 16892
rect 9608 16890 9614 16892
rect 9368 16838 9370 16890
rect 9550 16838 9552 16890
rect 9306 16836 9312 16838
rect 9368 16836 9392 16838
rect 9448 16836 9472 16838
rect 9528 16836 9552 16838
rect 9608 16836 9614 16838
rect 9306 16827 9614 16836
rect 9306 15804 9614 15813
rect 9306 15802 9312 15804
rect 9368 15802 9392 15804
rect 9448 15802 9472 15804
rect 9528 15802 9552 15804
rect 9608 15802 9614 15804
rect 9368 15750 9370 15802
rect 9550 15750 9552 15802
rect 9306 15748 9312 15750
rect 9368 15748 9392 15750
rect 9448 15748 9472 15750
rect 9528 15748 9552 15750
rect 9608 15748 9614 15750
rect 9306 15739 9614 15748
rect 9692 15638 9720 17478
rect 9876 16522 9904 18142
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 9968 16726 9996 18022
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 10060 16250 10088 16594
rect 10336 16250 10364 18022
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 12850 8800 13806
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8772 12714 8800 12786
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 11354 8892 12582
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 9048 10266 9076 14758
rect 9140 13530 9168 14758
rect 9306 14716 9614 14725
rect 9306 14714 9312 14716
rect 9368 14714 9392 14716
rect 9448 14714 9472 14716
rect 9528 14714 9552 14716
rect 9608 14714 9614 14716
rect 9368 14662 9370 14714
rect 9550 14662 9552 14714
rect 9306 14660 9312 14662
rect 9368 14660 9392 14662
rect 9448 14660 9472 14662
rect 9528 14660 9552 14662
rect 9608 14660 9614 14662
rect 9306 14651 9614 14660
rect 9784 14278 9812 14758
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9306 13628 9614 13637
rect 9306 13626 9312 13628
rect 9368 13626 9392 13628
rect 9448 13626 9472 13628
rect 9528 13626 9552 13628
rect 9608 13626 9614 13628
rect 9368 13574 9370 13626
rect 9550 13574 9552 13626
rect 9306 13572 9312 13574
rect 9368 13572 9392 13574
rect 9448 13572 9472 13574
rect 9528 13572 9552 13574
rect 9608 13572 9614 13574
rect 9306 13563 9614 13572
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 12986 9720 13262
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 11694 9260 12718
rect 9306 12540 9614 12549
rect 9306 12538 9312 12540
rect 9368 12538 9392 12540
rect 9448 12538 9472 12540
rect 9528 12538 9552 12540
rect 9608 12538 9614 12540
rect 9368 12486 9370 12538
rect 9550 12486 9552 12538
rect 9306 12484 9312 12486
rect 9368 12484 9392 12486
rect 9448 12484 9472 12486
rect 9528 12484 9552 12486
rect 9608 12484 9614 12486
rect 9306 12475 9614 12484
rect 9784 11830 9812 14214
rect 9876 13462 9904 15846
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10060 15162 10088 15506
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10336 15094 10364 15506
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10336 14958 10364 15030
rect 10520 15026 10548 18226
rect 12406 17980 12714 17989
rect 12406 17978 12412 17980
rect 12468 17978 12492 17980
rect 12548 17978 12572 17980
rect 12628 17978 12652 17980
rect 12708 17978 12714 17980
rect 12468 17926 12470 17978
rect 12650 17926 12652 17978
rect 12406 17924 12412 17926
rect 12468 17924 12492 17926
rect 12548 17924 12572 17926
rect 12628 17924 12652 17926
rect 12708 17924 12714 17926
rect 12406 17915 12714 17924
rect 12820 17678 12848 19200
rect 13956 18524 14264 18533
rect 13956 18522 13962 18524
rect 14018 18522 14042 18524
rect 14098 18522 14122 18524
rect 14178 18522 14202 18524
rect 14258 18522 14264 18524
rect 14018 18470 14020 18522
rect 14200 18470 14202 18522
rect 13956 18468 13962 18470
rect 14018 18468 14042 18470
rect 14098 18468 14122 18470
rect 14178 18468 14202 18470
rect 14258 18468 14264 18470
rect 13956 18459 14264 18468
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12912 17746 12940 18158
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 10856 17436 11164 17445
rect 10856 17434 10862 17436
rect 10918 17434 10942 17436
rect 10998 17434 11022 17436
rect 11078 17434 11102 17436
rect 11158 17434 11164 17436
rect 10918 17382 10920 17434
rect 11100 17382 11102 17434
rect 10856 17380 10862 17382
rect 10918 17380 10942 17382
rect 10998 17380 11022 17382
rect 11078 17380 11102 17382
rect 11158 17380 11164 17382
rect 10856 17371 11164 17380
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12176 17066 12204 17138
rect 12348 17128 12400 17134
rect 12268 17088 12348 17116
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 10612 15910 10640 17002
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 10856 16348 11164 16357
rect 10856 16346 10862 16348
rect 10918 16346 10942 16348
rect 10998 16346 11022 16348
rect 11078 16346 11102 16348
rect 11158 16346 11164 16348
rect 10918 16294 10920 16346
rect 11100 16294 11102 16346
rect 10856 16292 10862 16294
rect 10918 16292 10942 16294
rect 10998 16292 11022 16294
rect 11078 16292 11102 16294
rect 11158 16292 11164 16294
rect 10856 16283 11164 16292
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 11716 15706 11744 16934
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 12084 15570 12112 16662
rect 12176 16454 12204 17002
rect 12268 16658 12296 17088
rect 12348 17070 12400 17076
rect 12544 16998 12572 17206
rect 13464 17134 13492 18158
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12406 16892 12714 16901
rect 12406 16890 12412 16892
rect 12468 16890 12492 16892
rect 12548 16890 12572 16892
rect 12628 16890 12652 16892
rect 12708 16890 12714 16892
rect 12468 16838 12470 16890
rect 12650 16838 12652 16890
rect 12406 16836 12412 16838
rect 12468 16836 12492 16838
rect 12548 16836 12572 16838
rect 12628 16836 12652 16838
rect 12708 16836 12714 16838
rect 12406 16827 12714 16836
rect 12820 16794 12848 17070
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13096 16658 13124 16934
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 10856 15260 11164 15269
rect 10856 15258 10862 15260
rect 10918 15258 10942 15260
rect 10998 15258 11022 15260
rect 11078 15258 11102 15260
rect 11158 15258 11164 15260
rect 10918 15206 10920 15258
rect 11100 15206 11102 15258
rect 10856 15204 10862 15206
rect 10918 15204 10942 15206
rect 10998 15204 11022 15206
rect 11078 15204 11102 15206
rect 11158 15204 11164 15206
rect 10856 15195 11164 15204
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 11256 14958 11284 15302
rect 11348 15162 11376 15438
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10336 14822 10364 14894
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 10060 13870 10088 14418
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10060 13530 10088 13806
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 10152 12850 10180 14282
rect 10856 14172 11164 14181
rect 10856 14170 10862 14172
rect 10918 14170 10942 14172
rect 10998 14170 11022 14172
rect 11078 14170 11102 14172
rect 11158 14170 11164 14172
rect 10918 14118 10920 14170
rect 11100 14118 11102 14170
rect 10856 14116 10862 14118
rect 10918 14116 10942 14118
rect 10998 14116 11022 14118
rect 11078 14116 11102 14118
rect 11158 14116 11164 14118
rect 10856 14107 11164 14116
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11354 9168 11494
rect 9306 11452 9614 11461
rect 9306 11450 9312 11452
rect 9368 11450 9392 11452
rect 9448 11450 9472 11452
rect 9528 11450 9552 11452
rect 9608 11450 9614 11452
rect 9368 11398 9370 11450
rect 9550 11398 9552 11450
rect 9306 11396 9312 11398
rect 9368 11396 9392 11398
rect 9448 11396 9472 11398
rect 9528 11396 9552 11398
rect 9608 11396 9614 11398
rect 9306 11387 9614 11396
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9784 11218 9812 11766
rect 9968 11218 9996 12038
rect 10060 11762 10088 12786
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10428 11694 10456 13126
rect 10520 12918 10548 13126
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10704 11898 10732 12242
rect 10796 12238 10824 13126
rect 10856 13084 11164 13093
rect 10856 13082 10862 13084
rect 10918 13082 10942 13084
rect 10998 13082 11022 13084
rect 11078 13082 11102 13084
rect 11158 13082 11164 13084
rect 10918 13030 10920 13082
rect 11100 13030 11102 13082
rect 10856 13028 10862 13030
rect 10918 13028 10942 13030
rect 10998 13028 11022 13030
rect 11078 13028 11102 13030
rect 11158 13028 11164 13030
rect 10856 13019 11164 13028
rect 11256 12374 11284 14418
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 13938 11376 14214
rect 11532 13938 11560 15370
rect 11624 15026 11652 15370
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 12176 14958 12204 15506
rect 12268 15094 12296 16594
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12406 15804 12714 15813
rect 12406 15802 12412 15804
rect 12468 15802 12492 15804
rect 12548 15802 12572 15804
rect 12628 15802 12652 15804
rect 12708 15802 12714 15804
rect 12468 15750 12470 15802
rect 12650 15750 12652 15802
rect 12406 15748 12412 15750
rect 12468 15748 12492 15750
rect 12548 15748 12572 15750
rect 12628 15748 12652 15750
rect 12708 15748 12714 15750
rect 12406 15739 12714 15748
rect 12820 15706 12848 16390
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12164 14952 12216 14958
rect 12084 14912 12164 14940
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11808 13394 11836 14826
rect 12084 13462 12112 14912
rect 12164 14894 12216 14900
rect 12406 14716 12714 14725
rect 12406 14714 12412 14716
rect 12468 14714 12492 14716
rect 12548 14714 12572 14716
rect 12628 14714 12652 14716
rect 12708 14714 12714 14716
rect 12468 14662 12470 14714
rect 12650 14662 12652 14714
rect 12406 14660 12412 14662
rect 12468 14660 12492 14662
rect 12548 14660 12572 14662
rect 12628 14660 12652 14662
rect 12708 14660 12714 14662
rect 12406 14651 12714 14660
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12636 13802 12664 14486
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12782 11468 13262
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11440 12306 11468 12718
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10856 11996 11164 12005
rect 10856 11994 10862 11996
rect 10918 11994 10942 11996
rect 10998 11994 11022 11996
rect 11078 11994 11102 11996
rect 11158 11994 11164 11996
rect 10918 11942 10920 11994
rect 11100 11942 11102 11994
rect 10856 11940 10862 11942
rect 10918 11940 10942 11942
rect 10998 11940 11022 11942
rect 11078 11940 11102 11942
rect 11158 11940 11164 11942
rect 10856 11931 11164 11940
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10244 11218 10272 11494
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 10810 10640 11086
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10704 10606 10732 11494
rect 10856 10908 11164 10917
rect 10856 10906 10862 10908
rect 10918 10906 10942 10908
rect 10998 10906 11022 10908
rect 11078 10906 11102 10908
rect 11158 10906 11164 10908
rect 10918 10854 10920 10906
rect 11100 10854 11102 10906
rect 10856 10852 10862 10854
rect 10918 10852 10942 10854
rect 10998 10852 11022 10854
rect 11078 10852 11102 10854
rect 11158 10852 11164 10854
rect 10856 10843 11164 10852
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 9306 10364 9614 10373
rect 9306 10362 9312 10364
rect 9368 10362 9392 10364
rect 9448 10362 9472 10364
rect 9528 10362 9552 10364
rect 9608 10362 9614 10364
rect 9368 10310 9370 10362
rect 9550 10310 9552 10362
rect 9306 10308 9312 10310
rect 9368 10308 9392 10310
rect 9448 10308 9472 10310
rect 9528 10308 9552 10310
rect 9608 10308 9614 10310
rect 9306 10299 9614 10308
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7756 8732 8064 8741
rect 7756 8730 7762 8732
rect 7818 8730 7842 8732
rect 7898 8730 7922 8732
rect 7978 8730 8002 8732
rect 8058 8730 8064 8732
rect 7818 8678 7820 8730
rect 8000 8678 8002 8730
rect 7756 8676 7762 8678
rect 7818 8676 7842 8678
rect 7898 8676 7922 8678
rect 7978 8676 8002 8678
rect 8058 8676 8064 8678
rect 7756 8667 8064 8676
rect 8128 8634 8156 8774
rect 8312 8634 8340 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8514 8432 9318
rect 8680 9042 8708 9386
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8312 8486 8432 8514
rect 8312 8430 8340 8486
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7756 7644 8064 7653
rect 7756 7642 7762 7644
rect 7818 7642 7842 7644
rect 7898 7642 7922 7644
rect 7978 7642 8002 7644
rect 8058 7642 8064 7644
rect 7818 7590 7820 7642
rect 8000 7590 8002 7642
rect 7756 7588 7762 7590
rect 7818 7588 7842 7590
rect 7898 7588 7922 7590
rect 7978 7588 8002 7590
rect 8058 7588 8064 7590
rect 7756 7579 8064 7588
rect 8312 7342 8340 8366
rect 8680 8362 8708 8978
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8680 8090 8708 8298
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8680 6934 8708 8026
rect 8956 7546 8984 9522
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 9110 9076 9318
rect 9306 9276 9614 9285
rect 9306 9274 9312 9276
rect 9368 9274 9392 9276
rect 9448 9274 9472 9276
rect 9528 9274 9552 9276
rect 9608 9274 9614 9276
rect 9368 9222 9370 9274
rect 9550 9222 9552 9274
rect 9306 9220 9312 9222
rect 9368 9220 9392 9222
rect 9448 9220 9472 9222
rect 9528 9220 9552 9222
rect 9608 9220 9614 9222
rect 9306 9211 9614 9220
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 9876 8974 9904 9998
rect 10704 9722 10732 10542
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9586 10824 10202
rect 11256 10130 11284 11494
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10856 9820 11164 9829
rect 10856 9818 10862 9820
rect 10918 9818 10942 9820
rect 10998 9818 11022 9820
rect 11078 9818 11102 9820
rect 11158 9818 11164 9820
rect 10918 9766 10920 9818
rect 11100 9766 11102 9818
rect 10856 9764 10862 9766
rect 10918 9764 10942 9766
rect 10998 9764 11022 9766
rect 11078 9764 11102 9766
rect 11158 9764 11164 9766
rect 10856 9755 11164 9764
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10796 9110 10824 9386
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9306 8188 9614 8197
rect 9306 8186 9312 8188
rect 9368 8186 9392 8188
rect 9448 8186 9472 8188
rect 9528 8186 9552 8188
rect 9608 8186 9614 8188
rect 9368 8134 9370 8186
rect 9550 8134 9552 8186
rect 9306 8132 9312 8134
rect 9368 8132 9392 8134
rect 9448 8132 9472 8134
rect 9528 8132 9552 8134
rect 9608 8132 9614 8134
rect 9306 8123 9614 8132
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7756 6556 8064 6565
rect 7756 6554 7762 6556
rect 7818 6554 7842 6556
rect 7898 6554 7922 6556
rect 7978 6554 8002 6556
rect 8058 6554 8064 6556
rect 7818 6502 7820 6554
rect 8000 6502 8002 6554
rect 7756 6500 7762 6502
rect 7818 6500 7842 6502
rect 7898 6500 7922 6502
rect 7978 6500 8002 6502
rect 8058 6500 8064 6502
rect 7756 6491 8064 6500
rect 8220 6186 8248 6802
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4554 6868 4966
rect 7024 4826 7052 6054
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6840 4214 6868 4490
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6840 4010 6868 4150
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6206 3836 6514 3845
rect 6206 3834 6212 3836
rect 6268 3834 6292 3836
rect 6348 3834 6372 3836
rect 6428 3834 6452 3836
rect 6508 3834 6514 3836
rect 6268 3782 6270 3834
rect 6450 3782 6452 3834
rect 6206 3780 6212 3782
rect 6268 3780 6292 3782
rect 6348 3780 6372 3782
rect 6428 3780 6452 3782
rect 6508 3780 6514 3782
rect 6206 3771 6514 3780
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6380 2990 6408 3062
rect 6840 3058 6868 3946
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6840 2802 6868 2994
rect 6840 2774 6960 2802
rect 6206 2748 6514 2757
rect 6206 2746 6212 2748
rect 6268 2746 6292 2748
rect 6348 2746 6372 2748
rect 6428 2746 6452 2748
rect 6508 2746 6514 2748
rect 6268 2694 6270 2746
rect 6450 2694 6452 2746
rect 6206 2692 6212 2694
rect 6268 2692 6292 2694
rect 6348 2692 6372 2694
rect 6428 2692 6452 2694
rect 6508 2692 6514 2694
rect 6206 2683 6514 2692
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 4528 1760 4580 1766
rect 4528 1702 4580 1708
rect 5368 1426 5396 1838
rect 5828 1834 5856 2042
rect 6932 1970 6960 2774
rect 7024 2106 7052 3946
rect 7116 2514 7144 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7208 4282 7236 4762
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7208 4010 7236 4218
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7300 2582 7328 5170
rect 7392 4010 7420 5782
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7484 4486 7512 4626
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4010 7512 4422
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7576 3942 7604 6054
rect 8036 5914 8064 6122
rect 8024 5908 8076 5914
rect 8076 5868 8156 5896
rect 8024 5850 8076 5856
rect 7756 5468 8064 5477
rect 7756 5466 7762 5468
rect 7818 5466 7842 5468
rect 7898 5466 7922 5468
rect 7978 5466 8002 5468
rect 8058 5466 8064 5468
rect 7818 5414 7820 5466
rect 8000 5414 8002 5466
rect 7756 5412 7762 5414
rect 7818 5412 7842 5414
rect 7898 5412 7922 5414
rect 7978 5412 8002 5414
rect 8058 5412 8064 5414
rect 7756 5403 8064 5412
rect 8128 5370 8156 5868
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8220 5166 8248 6122
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 7756 4380 8064 4389
rect 7756 4378 7762 4380
rect 7818 4378 7842 4380
rect 7898 4378 7922 4380
rect 7978 4378 8002 4380
rect 8058 4378 8064 4380
rect 7818 4326 7820 4378
rect 8000 4326 8002 4378
rect 7756 4324 7762 4326
rect 7818 4324 7842 4326
rect 7898 4324 7922 4326
rect 7978 4324 8002 4326
rect 8058 4324 8064 4326
rect 7756 4315 8064 4324
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7668 2582 7696 4014
rect 7756 3292 8064 3301
rect 7756 3290 7762 3292
rect 7818 3290 7842 3292
rect 7898 3290 7922 3292
rect 7978 3290 8002 3292
rect 8058 3290 8064 3292
rect 7818 3238 7820 3290
rect 8000 3238 8002 3290
rect 7756 3236 7762 3238
rect 7818 3236 7842 3238
rect 7898 3236 7922 3238
rect 7978 3236 8002 3238
rect 8058 3236 8064 3238
rect 7756 3227 8064 3236
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7288 2576 7340 2582
rect 7288 2518 7340 2524
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 8036 2514 8064 2586
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 7756 2204 8064 2213
rect 7756 2202 7762 2204
rect 7818 2202 7842 2204
rect 7898 2202 7922 2204
rect 7978 2202 8002 2204
rect 8058 2202 8064 2204
rect 7818 2150 7820 2202
rect 8000 2150 8002 2202
rect 7756 2148 7762 2150
rect 7818 2148 7842 2150
rect 7898 2148 7922 2150
rect 7978 2148 8002 2150
rect 8058 2148 8064 2150
rect 7756 2139 8064 2148
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 8312 1902 8340 5102
rect 8404 4826 8432 6734
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4622 8524 6258
rect 8772 5166 8800 6326
rect 8864 5302 8892 7278
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4282 8800 4490
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 3992 8892 5102
rect 8956 4690 8984 6598
rect 9232 6390 9260 7210
rect 9306 7100 9614 7109
rect 9306 7098 9312 7100
rect 9368 7098 9392 7100
rect 9448 7098 9472 7100
rect 9528 7098 9552 7100
rect 9608 7098 9614 7100
rect 9368 7046 9370 7098
rect 9550 7046 9552 7098
rect 9306 7044 9312 7046
rect 9368 7044 9392 7046
rect 9448 7044 9472 7046
rect 9528 7044 9552 7046
rect 9608 7044 9614 7046
rect 9306 7035 9614 7044
rect 9876 6914 9904 8910
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10428 8090 10456 8366
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 9876 6886 9996 6914
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5846 9260 6054
rect 9306 6012 9614 6021
rect 9306 6010 9312 6012
rect 9368 6010 9392 6012
rect 9448 6010 9472 6012
rect 9528 6010 9552 6012
rect 9608 6010 9614 6012
rect 9368 5958 9370 6010
rect 9550 5958 9552 6010
rect 9306 5956 9312 5958
rect 9368 5956 9392 5958
rect 9448 5956 9472 5958
rect 9528 5956 9552 5958
rect 9608 5956 9614 5958
rect 9306 5947 9614 5956
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5166 9628 5646
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4282 8984 4626
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8944 4004 8996 4010
rect 8864 3964 8944 3992
rect 8944 3946 8996 3952
rect 8956 3126 8984 3946
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 5816 1828 5868 1834
rect 5816 1770 5868 1776
rect 5632 1760 5684 1766
rect 5632 1702 5684 1708
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 5644 1562 5672 1702
rect 6206 1660 6514 1669
rect 6206 1658 6212 1660
rect 6268 1658 6292 1660
rect 6348 1658 6372 1660
rect 6428 1658 6452 1660
rect 6508 1658 6514 1660
rect 6268 1606 6270 1658
rect 6450 1606 6452 1658
rect 6206 1604 6212 1606
rect 6268 1604 6292 1606
rect 6348 1604 6372 1606
rect 6428 1604 6452 1606
rect 6508 1604 6514 1606
rect 6206 1595 6514 1604
rect 7300 1562 7328 1702
rect 8312 1562 8340 1838
rect 5632 1556 5684 1562
rect 5632 1498 5684 1504
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 4344 1420 4396 1426
rect 4344 1362 4396 1368
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 3988 1222 4016 1362
rect 8680 1358 8708 2518
rect 9048 2310 9076 5034
rect 9232 4758 9260 5102
rect 9306 4924 9614 4933
rect 9306 4922 9312 4924
rect 9368 4922 9392 4924
rect 9448 4922 9472 4924
rect 9528 4922 9552 4924
rect 9608 4922 9614 4924
rect 9368 4870 9370 4922
rect 9550 4870 9552 4922
rect 9306 4868 9312 4870
rect 9368 4868 9392 4870
rect 9448 4868 9472 4870
rect 9528 4868 9552 4870
rect 9608 4868 9614 4870
rect 9306 4859 9614 4868
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9784 4282 9812 5102
rect 9968 4690 9996 6886
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5098 10272 5510
rect 10520 5166 10548 8434
rect 10796 8378 10824 9046
rect 10856 8732 11164 8741
rect 10856 8730 10862 8732
rect 10918 8730 10942 8732
rect 10998 8730 11022 8732
rect 11078 8730 11102 8732
rect 11158 8730 11164 8732
rect 10918 8678 10920 8730
rect 11100 8678 11102 8730
rect 10856 8676 10862 8678
rect 10918 8676 10942 8678
rect 10998 8676 11022 8678
rect 11078 8676 11102 8678
rect 11158 8676 11164 8678
rect 10856 8667 11164 8676
rect 10796 8362 10916 8378
rect 10796 8356 10928 8362
rect 10796 8350 10876 8356
rect 10876 8298 10928 8304
rect 10888 8022 10916 8298
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10856 7644 11164 7653
rect 10856 7642 10862 7644
rect 10918 7642 10942 7644
rect 10998 7642 11022 7644
rect 11078 7642 11102 7644
rect 11158 7642 11164 7644
rect 10918 7590 10920 7642
rect 11100 7590 11102 7642
rect 10856 7588 10862 7590
rect 10918 7588 10942 7590
rect 10998 7588 11022 7590
rect 11078 7588 11102 7590
rect 11158 7588 11164 7590
rect 10856 7579 11164 7588
rect 11256 7342 11284 10066
rect 11348 9178 11376 11630
rect 11440 10810 11468 12242
rect 11532 11762 11560 13330
rect 11808 12238 11836 13330
rect 12176 12714 12204 13670
rect 12406 13628 12714 13637
rect 12406 13626 12412 13628
rect 12468 13626 12492 13628
rect 12548 13626 12572 13628
rect 12628 13626 12652 13628
rect 12708 13626 12714 13628
rect 12468 13574 12470 13626
rect 12650 13574 12652 13626
rect 12406 13572 12412 13574
rect 12468 13572 12492 13574
rect 12548 13572 12572 13574
rect 12628 13572 12652 13574
rect 12708 13572 12714 13574
rect 12406 13563 12714 13572
rect 12820 12986 12848 15642
rect 12912 15570 12940 16594
rect 13096 16266 13124 16594
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13004 16238 13124 16266
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 14958 12940 15506
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12912 14414 12940 14758
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11354 11560 11698
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 9178 11468 10542
rect 12176 10538 12204 12650
rect 12406 12540 12714 12549
rect 12406 12538 12412 12540
rect 12468 12538 12492 12540
rect 12548 12538 12572 12540
rect 12628 12538 12652 12540
rect 12708 12538 12714 12540
rect 12468 12486 12470 12538
rect 12650 12486 12652 12538
rect 12406 12484 12412 12486
rect 12468 12484 12492 12486
rect 12548 12484 12572 12486
rect 12628 12484 12652 12486
rect 12708 12484 12714 12486
rect 12406 12475 12714 12484
rect 12912 12434 12940 14010
rect 13004 13938 13032 16238
rect 13372 15706 13400 16526
rect 13464 16454 13492 17070
rect 13648 16998 13676 17070
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14482 13124 14758
rect 13556 14482 13584 16390
rect 13832 16250 13860 18090
rect 13956 17436 14264 17445
rect 13956 17434 13962 17436
rect 14018 17434 14042 17436
rect 14098 17434 14122 17436
rect 14178 17434 14202 17436
rect 14258 17434 14264 17436
rect 14018 17382 14020 17434
rect 14200 17382 14202 17434
rect 13956 17380 13962 17382
rect 14018 17380 14042 17382
rect 14098 17380 14122 17382
rect 14178 17380 14202 17382
rect 14258 17380 14264 17382
rect 13956 17371 14264 17380
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 13956 16348 14264 16357
rect 13956 16346 13962 16348
rect 14018 16346 14042 16348
rect 14098 16346 14122 16348
rect 14178 16346 14202 16348
rect 14258 16346 14264 16348
rect 14018 16294 14020 16346
rect 14200 16294 14202 16346
rect 13956 16292 13962 16294
rect 14018 16292 14042 16294
rect 14098 16292 14122 16294
rect 14178 16292 14202 16294
rect 14258 16292 14264 16294
rect 13956 16283 14264 16292
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14292 15706 14320 17138
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 16658 14504 16934
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14384 15586 14412 16390
rect 14292 15558 14412 15586
rect 14292 15502 14320 15558
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 13956 15260 14264 15269
rect 13956 15258 13962 15260
rect 14018 15258 14042 15260
rect 14098 15258 14122 15260
rect 14178 15258 14202 15260
rect 14258 15258 14264 15260
rect 14018 15206 14020 15258
rect 14200 15206 14202 15258
rect 13956 15204 13962 15206
rect 14018 15204 14042 15206
rect 14098 15204 14122 15206
rect 14178 15204 14202 15206
rect 14258 15204 14264 15206
rect 13956 15195 14264 15204
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13464 13462 13492 14350
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 12912 12406 13032 12434
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12406 11452 12714 11461
rect 12406 11450 12412 11452
rect 12468 11450 12492 11452
rect 12548 11450 12572 11452
rect 12628 11450 12652 11452
rect 12708 11450 12714 11452
rect 12468 11398 12470 11450
rect 12650 11398 12652 11450
rect 12406 11396 12412 11398
rect 12468 11396 12492 11398
rect 12548 11396 12572 11398
rect 12628 11396 12652 11398
rect 12708 11396 12714 11398
rect 12406 11387 12714 11396
rect 12820 10554 12848 12106
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 10674 12940 12038
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12164 10532 12216 10538
rect 12820 10526 12940 10554
rect 12164 10474 12216 10480
rect 12176 9674 12204 10474
rect 12406 10364 12714 10373
rect 12406 10362 12412 10364
rect 12468 10362 12492 10364
rect 12548 10362 12572 10364
rect 12628 10362 12652 10364
rect 12708 10362 12714 10364
rect 12468 10310 12470 10362
rect 12650 10310 12652 10362
rect 12406 10308 12412 10310
rect 12468 10308 12492 10310
rect 12548 10308 12572 10310
rect 12628 10308 12652 10310
rect 12708 10308 12714 10310
rect 12406 10299 12714 10308
rect 11612 9648 11664 9654
rect 12176 9646 12296 9674
rect 11612 9590 11664 9596
rect 11624 9382 11652 9590
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11900 9042 11928 9522
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10856 6556 11164 6565
rect 10856 6554 10862 6556
rect 10918 6554 10942 6556
rect 10998 6554 11022 6556
rect 11078 6554 11102 6556
rect 11158 6554 11164 6556
rect 10918 6502 10920 6554
rect 11100 6502 11102 6554
rect 10856 6500 10862 6502
rect 10918 6500 10942 6502
rect 10998 6500 11022 6502
rect 11078 6500 11102 6502
rect 11158 6500 11164 6502
rect 10856 6491 11164 6500
rect 11256 5794 11284 6734
rect 11348 6458 11376 8910
rect 11900 8498 11928 8978
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 7954 11928 8434
rect 12268 8430 12296 9646
rect 12406 9276 12714 9285
rect 12406 9274 12412 9276
rect 12468 9274 12492 9276
rect 12548 9274 12572 9276
rect 12628 9274 12652 9276
rect 12708 9274 12714 9276
rect 12468 9222 12470 9274
rect 12650 9222 12652 9274
rect 12406 9220 12412 9222
rect 12468 9220 12492 9222
rect 12548 9220 12572 9222
rect 12628 9220 12652 9222
rect 12708 9220 12714 9222
rect 12406 9211 12714 9220
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7478 11928 7890
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 6322 11468 7414
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11256 5766 11376 5794
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 10856 5468 11164 5477
rect 10856 5466 10862 5468
rect 10918 5466 10942 5468
rect 10998 5466 11022 5468
rect 11078 5466 11102 5468
rect 11158 5466 11164 5468
rect 10918 5414 10920 5466
rect 11100 5414 11102 5466
rect 10856 5412 10862 5414
rect 10918 5412 10942 5414
rect 10998 5412 11022 5414
rect 11078 5412 11102 5414
rect 11158 5412 11164 5414
rect 10856 5403 11164 5412
rect 11256 5370 11284 5578
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3194 9168 3878
rect 9306 3836 9614 3845
rect 9306 3834 9312 3836
rect 9368 3834 9392 3836
rect 9448 3834 9472 3836
rect 9528 3834 9552 3836
rect 9608 3834 9614 3836
rect 9368 3782 9370 3834
rect 9550 3782 9552 3834
rect 9306 3780 9312 3782
rect 9368 3780 9392 3782
rect 9448 3780 9472 3782
rect 9528 3780 9552 3782
rect 9608 3780 9614 3782
rect 9306 3771 9614 3780
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9232 2650 9260 2994
rect 9306 2748 9614 2757
rect 9306 2746 9312 2748
rect 9368 2746 9392 2748
rect 9448 2746 9472 2748
rect 9528 2746 9552 2748
rect 9608 2746 9614 2748
rect 9368 2694 9370 2746
rect 9550 2694 9552 2746
rect 9306 2692 9312 2694
rect 9368 2692 9392 2694
rect 9448 2692 9472 2694
rect 9528 2692 9552 2694
rect 9608 2692 9614 2694
rect 9306 2683 9614 2692
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9692 2514 9720 4082
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 1902 9076 2246
rect 9232 2106 9260 2314
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9784 2038 9812 2790
rect 9876 2582 9904 4014
rect 10244 4010 10272 5034
rect 11348 4826 11376 5766
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 5658 11468 5714
rect 11532 5658 11560 6802
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11624 5778 11652 6734
rect 12176 6662 12204 8298
rect 12406 8188 12714 8197
rect 12406 8186 12412 8188
rect 12468 8186 12492 8188
rect 12548 8186 12572 8188
rect 12628 8186 12652 8188
rect 12708 8186 12714 8188
rect 12468 8134 12470 8186
rect 12650 8134 12652 8186
rect 12406 8132 12412 8134
rect 12468 8132 12492 8134
rect 12548 8132 12572 8134
rect 12628 8132 12652 8134
rect 12708 8132 12714 8134
rect 12406 8123 12714 8132
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7546 12572 7686
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12406 7100 12714 7109
rect 12406 7098 12412 7100
rect 12468 7098 12492 7100
rect 12548 7098 12572 7100
rect 12628 7098 12652 7100
rect 12708 7098 12714 7100
rect 12468 7046 12470 7098
rect 12650 7046 12652 7098
rect 12406 7044 12412 7046
rect 12468 7044 12492 7046
rect 12548 7044 12572 7046
rect 12628 7044 12652 7046
rect 12708 7044 12714 7046
rect 12406 7035 12714 7044
rect 12820 6730 12848 7822
rect 12912 6866 12940 10526
rect 13004 9110 13032 12406
rect 13188 12374 13216 12786
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11694 13216 12310
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 10674 13216 11630
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13188 10062 13216 10610
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13280 9994 13308 13330
rect 13556 13258 13584 14418
rect 14016 14414 14044 14962
rect 14188 14816 14240 14822
rect 14292 14804 14320 15438
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14958 14412 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14476 14822 14504 16594
rect 14464 14816 14516 14822
rect 14292 14776 14412 14804
rect 14188 14758 14240 14764
rect 14200 14634 14228 14758
rect 14200 14606 14320 14634
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13648 13530 13676 13942
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13648 12434 13676 13466
rect 13556 12406 13676 12434
rect 13556 12374 13584 12406
rect 13740 12374 13768 14282
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13832 11626 13860 14214
rect 13956 14172 14264 14181
rect 13956 14170 13962 14172
rect 14018 14170 14042 14172
rect 14098 14170 14122 14172
rect 14178 14170 14202 14172
rect 14258 14170 14264 14172
rect 14018 14118 14020 14170
rect 14200 14118 14202 14170
rect 13956 14116 13962 14118
rect 14018 14116 14042 14118
rect 14098 14116 14122 14118
rect 14178 14116 14202 14118
rect 14258 14116 14264 14118
rect 13956 14107 14264 14116
rect 13956 13084 14264 13093
rect 13956 13082 13962 13084
rect 14018 13082 14042 13084
rect 14098 13082 14122 13084
rect 14178 13082 14202 13084
rect 14258 13082 14264 13084
rect 14018 13030 14020 13082
rect 14200 13030 14202 13082
rect 13956 13028 13962 13030
rect 14018 13028 14042 13030
rect 14098 13028 14122 13030
rect 14178 13028 14202 13030
rect 14258 13028 14264 13030
rect 13956 13019 14264 13028
rect 14292 12306 14320 14606
rect 14384 13870 14412 14776
rect 14464 14758 14516 14764
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14384 12442 14412 13806
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 13956 11996 14264 12005
rect 13956 11994 13962 11996
rect 14018 11994 14042 11996
rect 14098 11994 14122 11996
rect 14178 11994 14202 11996
rect 14258 11994 14264 11996
rect 14018 11942 14020 11994
rect 14200 11942 14202 11994
rect 13956 11940 13962 11942
rect 14018 11940 14042 11942
rect 14098 11940 14122 11942
rect 14178 11940 14202 11942
rect 14258 11940 14264 11942
rect 13956 11931 14264 11940
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 14188 11552 14240 11558
rect 14240 11512 14320 11540
rect 14188 11494 14240 11500
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13832 10130 13860 11290
rect 13956 10908 14264 10917
rect 13956 10906 13962 10908
rect 14018 10906 14042 10908
rect 14098 10906 14122 10908
rect 14178 10906 14202 10908
rect 14258 10906 14264 10908
rect 14018 10854 14020 10906
rect 14200 10854 14202 10906
rect 13956 10852 13962 10854
rect 14018 10852 14042 10854
rect 14098 10852 14122 10854
rect 14178 10852 14202 10854
rect 14258 10852 14264 10854
rect 13956 10843 14264 10852
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13004 8634 13032 9046
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6186 12204 6598
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5846 12204 6122
rect 12406 6012 12714 6021
rect 12406 6010 12412 6012
rect 12468 6010 12492 6012
rect 12548 6010 12572 6012
rect 12628 6010 12652 6012
rect 12708 6010 12714 6012
rect 12468 5958 12470 6010
rect 12650 5958 12652 6010
rect 12406 5956 12412 5958
rect 12468 5956 12492 5958
rect 12548 5956 12572 5958
rect 12628 5956 12652 5958
rect 12708 5956 12714 5958
rect 12406 5947 12714 5956
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11808 5658 11836 5714
rect 11440 5630 11836 5658
rect 11808 5234 11836 5630
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10856 4380 11164 4389
rect 10856 4378 10862 4380
rect 10918 4378 10942 4380
rect 10998 4378 11022 4380
rect 11078 4378 11102 4380
rect 11158 4378 11164 4380
rect 10918 4326 10920 4378
rect 11100 4326 11102 4378
rect 10856 4324 10862 4326
rect 10918 4324 10942 4326
rect 10998 4324 11022 4326
rect 11078 4324 11102 4326
rect 11158 4324 11164 4326
rect 10856 4315 11164 4324
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 11348 3738 11376 4626
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 4282 11468 4558
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11440 3602 11468 4218
rect 11532 3738 11560 4966
rect 11808 4690 11836 5170
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 10856 3292 11164 3301
rect 10856 3290 10862 3292
rect 10918 3290 10942 3292
rect 10998 3290 11022 3292
rect 11078 3290 11102 3292
rect 11158 3290 11164 3292
rect 10918 3238 10920 3290
rect 11100 3238 11102 3290
rect 10856 3236 10862 3238
rect 10918 3236 10942 3238
rect 10998 3236 11022 3238
rect 11078 3236 11102 3238
rect 11158 3236 11164 3238
rect 10856 3227 11164 3236
rect 12268 3108 12296 5578
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12406 4924 12714 4933
rect 12406 4922 12412 4924
rect 12468 4922 12492 4924
rect 12548 4922 12572 4924
rect 12628 4922 12652 4924
rect 12708 4922 12714 4924
rect 12468 4870 12470 4922
rect 12650 4870 12652 4922
rect 12406 4868 12412 4870
rect 12468 4868 12492 4870
rect 12548 4868 12572 4870
rect 12628 4868 12652 4870
rect 12708 4868 12714 4870
rect 12406 4859 12714 4868
rect 12912 3942 12940 4966
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12406 3836 12714 3845
rect 12406 3834 12412 3836
rect 12468 3834 12492 3836
rect 12548 3834 12572 3836
rect 12628 3834 12652 3836
rect 12708 3834 12714 3836
rect 12468 3782 12470 3834
rect 12650 3782 12652 3834
rect 12406 3780 12412 3782
rect 12468 3780 12492 3782
rect 12548 3780 12572 3782
rect 12628 3780 12652 3782
rect 12708 3780 12714 3782
rect 12406 3771 12714 3780
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12544 3194 12572 3606
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12268 3080 12480 3108
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 9876 2446 9904 2518
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 9306 1660 9614 1669
rect 9306 1658 9312 1660
rect 9368 1658 9392 1660
rect 9448 1658 9472 1660
rect 9528 1658 9552 1660
rect 9608 1658 9614 1660
rect 9368 1606 9370 1658
rect 9550 1606 9552 1658
rect 9306 1604 9312 1606
rect 9368 1604 9392 1606
rect 9448 1604 9472 1606
rect 9528 1604 9552 1606
rect 9608 1604 9614 1606
rect 9306 1595 9614 1604
rect 10060 1426 10088 2246
rect 10336 1426 10364 2246
rect 10612 1902 10640 2518
rect 10856 2204 11164 2213
rect 10856 2202 10862 2204
rect 10918 2202 10942 2204
rect 10998 2202 11022 2204
rect 11078 2202 11102 2204
rect 11158 2202 11164 2204
rect 10918 2150 10920 2202
rect 11100 2150 11102 2202
rect 10856 2148 10862 2150
rect 10918 2148 10942 2150
rect 10998 2148 11022 2150
rect 11078 2148 11102 2150
rect 11158 2148 11164 2150
rect 10856 2139 11164 2148
rect 12084 1970 12112 2926
rect 12452 2854 12480 3080
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12406 2748 12714 2757
rect 12406 2746 12412 2748
rect 12468 2746 12492 2748
rect 12548 2746 12572 2748
rect 12628 2746 12652 2748
rect 12708 2746 12714 2748
rect 12468 2694 12470 2746
rect 12650 2694 12652 2746
rect 12406 2692 12412 2694
rect 12468 2692 12492 2694
rect 12548 2692 12572 2694
rect 12628 2692 12652 2694
rect 12708 2692 12714 2694
rect 12406 2683 12714 2692
rect 12820 2038 12848 3606
rect 12912 3534 12940 3878
rect 13004 3738 13032 7890
rect 13556 7818 13584 9930
rect 13956 9820 14264 9829
rect 13956 9818 13962 9820
rect 14018 9818 14042 9820
rect 14098 9818 14122 9820
rect 14178 9818 14202 9820
rect 14258 9818 14264 9820
rect 14018 9766 14020 9818
rect 14200 9766 14202 9818
rect 13956 9764 13962 9766
rect 14018 9764 14042 9766
rect 14098 9764 14122 9766
rect 14178 9764 14202 9766
rect 14258 9764 14264 9766
rect 13956 9755 14264 9764
rect 13956 8732 14264 8741
rect 13956 8730 13962 8732
rect 14018 8730 14042 8732
rect 14098 8730 14122 8732
rect 14178 8730 14202 8732
rect 14258 8730 14264 8732
rect 14018 8678 14020 8730
rect 14200 8678 14202 8730
rect 13956 8676 13962 8678
rect 14018 8676 14042 8678
rect 14098 8676 14122 8678
rect 14178 8676 14202 8678
rect 14258 8676 14264 8678
rect 13956 8667 14264 8676
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13832 6798 13860 8434
rect 14292 8294 14320 11512
rect 14476 10130 14504 14418
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9722 14504 10066
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14384 9382 14412 9454
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8906 14412 9318
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14568 8498 14596 13330
rect 14660 9042 14688 18226
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16590 14780 17002
rect 14844 16794 14872 18022
rect 14936 17746 14964 18090
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15028 16674 15056 18022
rect 15212 16794 15240 18022
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 14936 16646 15056 16674
rect 15200 16652 15252 16658
rect 14936 16590 14964 16646
rect 15200 16594 15252 16600
rect 14740 16584 14792 16590
rect 14924 16584 14976 16590
rect 14740 16526 14792 16532
rect 14844 16532 14924 16538
rect 14844 16526 14976 16532
rect 14752 15570 14780 16526
rect 14844 16510 14964 16526
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 14890 14780 15506
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14752 13938 14780 14826
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14844 12434 14872 16510
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 15028 15366 15056 15914
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14936 13870 14964 14962
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 13394 14964 13806
rect 15028 13462 15056 15302
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15120 13938 15148 14894
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14936 12702 15148 12730
rect 15212 12714 15240 16594
rect 14936 12646 14964 12702
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 12434 15056 12582
rect 14752 12406 14872 12434
rect 14936 12406 15056 12434
rect 14752 12238 14780 12406
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11150 14780 12174
rect 14844 12102 14872 12310
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11150 14872 12038
rect 14936 11354 14964 12406
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15028 11218 15056 12242
rect 15120 11626 15148 12702
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15212 11286 15240 12378
rect 15304 11762 15332 19230
rect 15580 19122 15608 19230
rect 15658 19200 15714 20000
rect 18510 19200 18566 20000
rect 15672 19122 15700 19200
rect 15580 19094 15700 19122
rect 18418 18592 18474 18601
rect 17056 18524 17364 18533
rect 18418 18527 18474 18536
rect 17056 18522 17062 18524
rect 17118 18522 17142 18524
rect 17198 18522 17222 18524
rect 17278 18522 17302 18524
rect 17358 18522 17364 18524
rect 17118 18470 17120 18522
rect 17300 18470 17302 18522
rect 17056 18468 17062 18470
rect 17118 18468 17142 18470
rect 17198 18468 17222 18470
rect 17278 18468 17302 18470
rect 17358 18468 17364 18470
rect 17056 18459 17364 18468
rect 18432 18426 18460 18527
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18432 18222 18460 18362
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 16658 15424 18022
rect 15506 17980 15814 17989
rect 15506 17978 15512 17980
rect 15568 17978 15592 17980
rect 15648 17978 15672 17980
rect 15728 17978 15752 17980
rect 15808 17978 15814 17980
rect 15568 17926 15570 17978
rect 15750 17926 15752 17978
rect 15506 17924 15512 17926
rect 15568 17924 15592 17926
rect 15648 17924 15672 17926
rect 15728 17924 15752 17926
rect 15808 17924 15814 17926
rect 15506 17915 15814 17924
rect 15506 16892 15814 16901
rect 15506 16890 15512 16892
rect 15568 16890 15592 16892
rect 15648 16890 15672 16892
rect 15728 16890 15752 16892
rect 15808 16890 15814 16892
rect 15568 16838 15570 16890
rect 15750 16838 15752 16890
rect 15506 16836 15512 16838
rect 15568 16836 15592 16838
rect 15648 16836 15672 16838
rect 15728 16836 15752 16838
rect 15808 16836 15814 16838
rect 15506 16827 15814 16836
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15506 15804 15814 15813
rect 15506 15802 15512 15804
rect 15568 15802 15592 15804
rect 15648 15802 15672 15804
rect 15728 15802 15752 15804
rect 15808 15802 15814 15804
rect 15568 15750 15570 15802
rect 15750 15750 15752 15802
rect 15506 15748 15512 15750
rect 15568 15748 15592 15750
rect 15648 15748 15672 15750
rect 15728 15748 15752 15750
rect 15808 15748 15814 15750
rect 15506 15739 15814 15748
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 14498 15424 14758
rect 15506 14716 15814 14725
rect 15506 14714 15512 14716
rect 15568 14714 15592 14716
rect 15648 14714 15672 14716
rect 15728 14714 15752 14716
rect 15808 14714 15814 14716
rect 15568 14662 15570 14714
rect 15750 14662 15752 14714
rect 15506 14660 15512 14662
rect 15568 14660 15592 14662
rect 15648 14660 15672 14662
rect 15728 14660 15752 14662
rect 15808 14660 15814 14662
rect 15506 14651 15814 14660
rect 15396 14470 15516 14498
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 13938 15424 14282
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15488 13784 15516 14470
rect 15856 14074 15884 14894
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16040 14414 16068 14486
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16132 14278 16160 18158
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15706 16344 15982
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15396 13756 15516 13784
rect 15396 11898 15424 13756
rect 15506 13628 15814 13637
rect 15506 13626 15512 13628
rect 15568 13626 15592 13628
rect 15648 13626 15672 13628
rect 15728 13626 15752 13628
rect 15808 13626 15814 13628
rect 15568 13574 15570 13626
rect 15750 13574 15752 13626
rect 15506 13572 15512 13574
rect 15568 13572 15592 13574
rect 15648 13572 15672 13574
rect 15728 13572 15752 13574
rect 15808 13572 15814 13574
rect 15506 13563 15814 13572
rect 16316 12918 16344 15506
rect 16500 15162 16528 17002
rect 16684 16794 16712 17614
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16868 15978 16896 17750
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17056 17436 17364 17445
rect 17056 17434 17062 17436
rect 17118 17434 17142 17436
rect 17198 17434 17222 17436
rect 17278 17434 17302 17436
rect 17358 17434 17364 17436
rect 17118 17382 17120 17434
rect 17300 17382 17302 17434
rect 17056 17380 17062 17382
rect 17118 17380 17142 17382
rect 17198 17380 17222 17382
rect 17278 17380 17302 17382
rect 17358 17380 17364 17382
rect 17056 17371 17364 17380
rect 17512 17202 17540 17478
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17056 16348 17364 16357
rect 17056 16346 17062 16348
rect 17118 16346 17142 16348
rect 17198 16346 17222 16348
rect 17278 16346 17302 16348
rect 17358 16346 17364 16348
rect 17118 16294 17120 16346
rect 17300 16294 17302 16346
rect 17056 16292 17062 16294
rect 17118 16292 17142 16294
rect 17198 16292 17222 16294
rect 17278 16292 17302 16294
rect 17358 16292 17364 16294
rect 17056 16283 17364 16292
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16592 14958 16620 15370
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16776 14482 16804 14962
rect 16868 14890 16896 15914
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15502 17724 15846
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17056 15260 17364 15269
rect 17056 15258 17062 15260
rect 17118 15258 17142 15260
rect 17198 15258 17222 15260
rect 17278 15258 17302 15260
rect 17358 15258 17364 15260
rect 17118 15206 17120 15258
rect 17300 15206 17302 15258
rect 17056 15204 17062 15206
rect 17118 15204 17142 15206
rect 17198 15204 17222 15206
rect 17278 15204 17302 15206
rect 17358 15204 17364 15206
rect 17056 15195 17364 15204
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 14550 16896 14826
rect 16960 14618 16988 15098
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16776 13954 16804 14418
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16592 13938 16804 13954
rect 16580 13932 16804 13938
rect 16632 13926 16804 13932
rect 16580 13874 16632 13880
rect 16592 13818 16620 13874
rect 16500 13790 16620 13818
rect 16764 13796 16816 13802
rect 16500 13530 16528 13790
rect 16764 13738 16816 13744
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16776 13462 16804 13738
rect 16868 13734 16896 14282
rect 16960 13802 16988 14554
rect 17696 14362 17724 15438
rect 17788 14482 17816 17070
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16153 18460 16594
rect 18418 16144 18474 16153
rect 18418 16079 18474 16088
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17880 15162 17908 15438
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 18432 14822 18460 15506
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18064 14482 18092 14758
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17960 14408 18012 14414
rect 17696 14334 17816 14362
rect 17960 14350 18012 14356
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17056 14172 17364 14181
rect 17056 14170 17062 14172
rect 17118 14170 17142 14172
rect 17198 14170 17222 14172
rect 17278 14170 17302 14172
rect 17358 14170 17364 14172
rect 17118 14118 17120 14170
rect 17300 14118 17302 14170
rect 17056 14116 17062 14118
rect 17118 14116 17142 14118
rect 17198 14116 17222 14118
rect 17278 14116 17302 14118
rect 17358 14116 17364 14118
rect 17056 14107 17364 14116
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17056 13084 17364 13093
rect 17056 13082 17062 13084
rect 17118 13082 17142 13084
rect 17198 13082 17222 13084
rect 17278 13082 17302 13084
rect 17358 13082 17364 13084
rect 17118 13030 17120 13082
rect 17300 13030 17302 13082
rect 17056 13028 17062 13030
rect 17118 13028 17142 13030
rect 17198 13028 17222 13030
rect 17278 13028 17302 13030
rect 17358 13028 17364 13030
rect 17056 13019 17364 13028
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 17604 12850 17632 13330
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 15506 12540 15814 12549
rect 15506 12538 15512 12540
rect 15568 12538 15592 12540
rect 15648 12538 15672 12540
rect 15728 12538 15752 12540
rect 15808 12538 15814 12540
rect 15568 12486 15570 12538
rect 15750 12486 15752 12538
rect 15506 12484 15512 12486
rect 15568 12484 15592 12486
rect 15648 12484 15672 12486
rect 15728 12484 15752 12486
rect 15808 12484 15814 12486
rect 15506 12475 15814 12484
rect 16132 12374 16160 12718
rect 16776 12442 16804 12718
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 17144 12306 17172 12718
rect 17604 12696 17632 12786
rect 17420 12668 17632 12696
rect 17420 12306 17448 12668
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15506 11452 15814 11461
rect 15506 11450 15512 11452
rect 15568 11450 15592 11452
rect 15648 11450 15672 11452
rect 15728 11450 15752 11452
rect 15808 11450 15814 11452
rect 15568 11398 15570 11450
rect 15750 11398 15752 11450
rect 15506 11396 15512 11398
rect 15568 11396 15592 11398
rect 15648 11396 15672 11398
rect 15728 11396 15752 11398
rect 15808 11396 15814 11398
rect 15506 11387 15814 11396
rect 16040 11354 16068 12174
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14752 9654 14780 11086
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 13956 7644 14264 7653
rect 13956 7642 13962 7644
rect 14018 7642 14042 7644
rect 14098 7642 14122 7644
rect 14178 7642 14202 7644
rect 14258 7642 14264 7644
rect 14018 7590 14020 7642
rect 14200 7590 14202 7642
rect 13956 7588 13962 7590
rect 14018 7588 14042 7590
rect 14098 7588 14122 7590
rect 14178 7588 14202 7590
rect 14258 7588 14264 7590
rect 13956 7579 14264 7588
rect 14292 7274 14320 8230
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14476 6798 14504 8366
rect 14568 7750 14596 8434
rect 14660 8090 14688 8978
rect 14844 8974 14872 11086
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14936 10826 14964 11018
rect 14936 10798 15056 10826
rect 16132 10810 16160 11630
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 15028 10266 15056 10798
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15028 9586 15056 10202
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8430 14872 8910
rect 15028 8430 15056 9318
rect 15212 8498 15240 9590
rect 15304 8838 15332 10474
rect 15506 10364 15814 10373
rect 15506 10362 15512 10364
rect 15568 10362 15592 10364
rect 15648 10362 15672 10364
rect 15728 10362 15752 10364
rect 15808 10362 15814 10364
rect 15568 10310 15570 10362
rect 15750 10310 15752 10362
rect 15506 10308 15512 10310
rect 15568 10308 15592 10310
rect 15648 10308 15672 10310
rect 15728 10308 15752 10310
rect 15808 10308 15814 10310
rect 15506 10299 15814 10308
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14844 7818 14872 8366
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 3738 13124 4422
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 13188 3194 13216 6190
rect 13832 4758 13860 6734
rect 13956 6556 14264 6565
rect 13956 6554 13962 6556
rect 14018 6554 14042 6556
rect 14098 6554 14122 6556
rect 14178 6554 14202 6556
rect 14258 6554 14264 6556
rect 14018 6502 14020 6554
rect 14200 6502 14202 6554
rect 13956 6500 13962 6502
rect 14018 6500 14042 6502
rect 14098 6500 14122 6502
rect 14178 6500 14202 6502
rect 14258 6500 14264 6502
rect 13956 6491 14264 6500
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 13956 5468 14264 5477
rect 13956 5466 13962 5468
rect 14018 5466 14042 5468
rect 14098 5466 14122 5468
rect 14178 5466 14202 5468
rect 14258 5466 14264 5468
rect 14018 5414 14020 5466
rect 14200 5414 14202 5466
rect 13956 5412 13962 5414
rect 14018 5412 14042 5414
rect 14098 5412 14122 5414
rect 14178 5412 14202 5414
rect 14258 5412 14264 5414
rect 13956 5403 14264 5412
rect 14292 5370 14320 5646
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13648 4146 13676 4490
rect 13956 4380 14264 4389
rect 13956 4378 13962 4380
rect 14018 4378 14042 4380
rect 14098 4378 14122 4380
rect 14178 4378 14202 4380
rect 14258 4378 14264 4380
rect 14018 4326 14020 4378
rect 14200 4326 14202 4378
rect 13956 4324 13962 4326
rect 14018 4324 14042 4326
rect 14098 4324 14122 4326
rect 14178 4324 14202 4326
rect 14258 4324 14264 4326
rect 13956 4315 14264 4324
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13556 2854 13584 3470
rect 13648 3058 13676 4082
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 12808 2032 12860 2038
rect 12808 1974 12860 1980
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 13004 1902 13032 2790
rect 13556 2446 13584 2790
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13648 1970 13676 2994
rect 13740 2990 13768 3062
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13832 2650 13860 3538
rect 14292 3534 14320 4626
rect 14384 3602 14412 6258
rect 14476 6254 14504 6734
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14568 6186 14596 7142
rect 14844 6254 14872 7754
rect 15028 6390 15056 8366
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13956 3292 14264 3301
rect 13956 3290 13962 3292
rect 14018 3290 14042 3292
rect 14098 3290 14122 3292
rect 14178 3290 14202 3292
rect 14258 3290 14264 3292
rect 14018 3238 14020 3290
rect 14200 3238 14202 3290
rect 13956 3236 13962 3238
rect 14018 3236 14042 3238
rect 14098 3236 14122 3238
rect 14178 3236 14202 3238
rect 14258 3236 14264 3238
rect 13956 3227 14264 3236
rect 14384 2854 14412 3538
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13924 2582 13952 2790
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 10600 1896 10652 1902
rect 10600 1838 10652 1844
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 13084 1760 13136 1766
rect 13084 1702 13136 1708
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 12406 1660 12714 1669
rect 12406 1658 12412 1660
rect 12468 1658 12492 1660
rect 12548 1658 12572 1660
rect 12628 1658 12652 1660
rect 12708 1658 12714 1660
rect 12468 1606 12470 1658
rect 12650 1606 12652 1658
rect 12406 1604 12412 1606
rect 12468 1604 12492 1606
rect 12548 1604 12572 1606
rect 12628 1604 12652 1606
rect 12708 1604 12714 1606
rect 12406 1595 12714 1604
rect 13096 1426 13124 1702
rect 13556 1426 13584 1702
rect 13740 1562 13768 2450
rect 13924 2360 13952 2518
rect 13832 2332 13952 2360
rect 13832 2038 13860 2332
rect 13956 2204 14264 2213
rect 13956 2202 13962 2204
rect 14018 2202 14042 2204
rect 14098 2202 14122 2204
rect 14178 2202 14202 2204
rect 14258 2202 14264 2204
rect 14018 2150 14020 2202
rect 14200 2150 14202 2202
rect 13956 2148 13962 2150
rect 14018 2148 14042 2150
rect 14098 2148 14122 2150
rect 14178 2148 14202 2150
rect 14258 2148 14264 2150
rect 13956 2139 14264 2148
rect 14568 2106 14596 6122
rect 14660 4282 14688 6190
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 10048 1420 10100 1426
rect 10048 1362 10100 1368
rect 10324 1420 10376 1426
rect 10324 1362 10376 1368
rect 13084 1420 13136 1426
rect 13084 1362 13136 1368
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 14752 1358 14780 3402
rect 14844 2582 14872 5510
rect 15304 5166 15332 8774
rect 15396 8634 15424 9998
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15580 9518 15608 9862
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15506 9276 15814 9285
rect 15506 9274 15512 9276
rect 15568 9274 15592 9276
rect 15648 9274 15672 9276
rect 15728 9274 15752 9276
rect 15808 9274 15814 9276
rect 15568 9222 15570 9274
rect 15750 9222 15752 9274
rect 15506 9220 15512 9222
rect 15568 9220 15592 9222
rect 15648 9220 15672 9222
rect 15728 9220 15752 9222
rect 15808 9220 15814 9222
rect 15506 9211 15814 9220
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15580 8362 15608 8842
rect 15856 8430 15884 9862
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 8498 15976 9454
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15568 8356 15620 8362
rect 16040 8344 16068 10134
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16224 8974 16252 9386
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15568 8298 15620 8304
rect 15948 8316 16068 8344
rect 15506 8188 15814 8197
rect 15506 8186 15512 8188
rect 15568 8186 15592 8188
rect 15648 8186 15672 8188
rect 15728 8186 15752 8188
rect 15808 8186 15814 8188
rect 15568 8134 15570 8186
rect 15750 8134 15752 8186
rect 15506 8132 15512 8134
rect 15568 8132 15592 8134
rect 15648 8132 15672 8134
rect 15728 8132 15752 8134
rect 15808 8132 15814 8134
rect 15506 8123 15814 8132
rect 15948 8022 15976 8316
rect 16408 8294 16436 11290
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16500 10674 16528 11086
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16592 9926 16620 12242
rect 17056 11996 17364 12005
rect 17056 11994 17062 11996
rect 17118 11994 17142 11996
rect 17198 11994 17222 11996
rect 17278 11994 17302 11996
rect 17358 11994 17364 11996
rect 17118 11942 17120 11994
rect 17300 11942 17302 11994
rect 17056 11940 17062 11942
rect 17118 11940 17142 11942
rect 17198 11940 17222 11942
rect 17278 11940 17302 11942
rect 17358 11940 17364 11942
rect 17056 11931 17364 11940
rect 17420 11898 17448 12242
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16592 8412 16620 8774
rect 16672 8424 16724 8430
rect 16592 8384 16672 8412
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15506 7100 15814 7109
rect 15506 7098 15512 7100
rect 15568 7098 15592 7100
rect 15648 7098 15672 7100
rect 15728 7098 15752 7100
rect 15808 7098 15814 7100
rect 15568 7046 15570 7098
rect 15750 7046 15752 7098
rect 15506 7044 15512 7046
rect 15568 7044 15592 7046
rect 15648 7044 15672 7046
rect 15728 7044 15752 7046
rect 15808 7044 15814 7046
rect 15506 7035 15814 7044
rect 15948 6746 15976 7958
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 15764 6730 15976 6746
rect 15752 6724 15976 6730
rect 15804 6718 15976 6724
rect 15752 6666 15804 6672
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15396 6186 15424 6598
rect 15856 6322 15884 6598
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14936 3670 14964 4082
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 15028 2802 15056 4422
rect 15396 3942 15424 6122
rect 15948 6118 15976 6718
rect 16132 6322 16160 7346
rect 16408 7274 16436 8230
rect 16500 7954 16528 8366
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16500 7546 16528 7890
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16408 6730 16436 7210
rect 16592 6798 16620 8384
rect 16672 8366 16724 8372
rect 16868 7546 16896 9318
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15506 6012 15814 6021
rect 15506 6010 15512 6012
rect 15568 6010 15592 6012
rect 15648 6010 15672 6012
rect 15728 6010 15752 6012
rect 15808 6010 15814 6012
rect 15568 5958 15570 6010
rect 15750 5958 15752 6010
rect 15506 5956 15512 5958
rect 15568 5956 15592 5958
rect 15648 5956 15672 5958
rect 15728 5956 15752 5958
rect 15808 5956 15814 5958
rect 15506 5947 15814 5956
rect 15948 5846 15976 6054
rect 16132 5914 16160 6258
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15506 4924 15814 4933
rect 15506 4922 15512 4924
rect 15568 4922 15592 4924
rect 15648 4922 15672 4924
rect 15728 4922 15752 4924
rect 15808 4922 15814 4924
rect 15568 4870 15570 4922
rect 15750 4870 15752 4922
rect 15506 4868 15512 4870
rect 15568 4868 15592 4870
rect 15648 4868 15672 4870
rect 15728 4868 15752 4870
rect 15808 4868 15814 4870
rect 15506 4859 15814 4868
rect 15948 4758 15976 5782
rect 16132 5710 16160 5850
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15948 4026 15976 4694
rect 15948 4010 16068 4026
rect 15936 4004 16068 4010
rect 15988 3998 16068 4004
rect 15936 3946 15988 3952
rect 15384 3936 15436 3942
rect 15948 3915 15976 3946
rect 15384 3878 15436 3884
rect 15396 3534 15424 3878
rect 15506 3836 15814 3845
rect 15506 3834 15512 3836
rect 15568 3834 15592 3836
rect 15648 3834 15672 3836
rect 15728 3834 15752 3836
rect 15808 3834 15814 3836
rect 15568 3782 15570 3834
rect 15750 3782 15752 3834
rect 15506 3780 15512 3782
rect 15568 3780 15592 3782
rect 15648 3780 15672 3782
rect 15728 3780 15752 3782
rect 15808 3780 15814 3782
rect 15506 3771 15814 3780
rect 16040 3670 16068 3998
rect 16224 3942 16252 5646
rect 16592 4758 16620 6734
rect 16776 6066 16804 6802
rect 16960 6118 16988 11154
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17056 10908 17364 10917
rect 17056 10906 17062 10908
rect 17118 10906 17142 10908
rect 17198 10906 17222 10908
rect 17278 10906 17302 10908
rect 17358 10906 17364 10908
rect 17118 10854 17120 10906
rect 17300 10854 17302 10906
rect 17056 10852 17062 10854
rect 17118 10852 17142 10854
rect 17198 10852 17222 10854
rect 17278 10852 17302 10854
rect 17358 10852 17364 10854
rect 17056 10843 17364 10852
rect 17512 10606 17540 10950
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10062 17172 10406
rect 17420 10130 17448 10542
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17056 9820 17364 9829
rect 17056 9818 17062 9820
rect 17118 9818 17142 9820
rect 17198 9818 17222 9820
rect 17278 9818 17302 9820
rect 17358 9818 17364 9820
rect 17118 9766 17120 9818
rect 17300 9766 17302 9818
rect 17056 9764 17062 9766
rect 17118 9764 17142 9766
rect 17198 9764 17222 9766
rect 17278 9764 17302 9766
rect 17358 9764 17364 9766
rect 17056 9755 17364 9764
rect 17420 9722 17448 10066
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17328 9178 17356 9454
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17056 8732 17364 8741
rect 17056 8730 17062 8732
rect 17118 8730 17142 8732
rect 17198 8730 17222 8732
rect 17278 8730 17302 8732
rect 17358 8730 17364 8732
rect 17118 8678 17120 8730
rect 17300 8678 17302 8730
rect 17056 8676 17062 8678
rect 17118 8676 17142 8678
rect 17198 8676 17222 8678
rect 17278 8676 17302 8678
rect 17358 8676 17364 8678
rect 17056 8667 17364 8676
rect 17420 8514 17448 9318
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17328 8486 17448 8514
rect 17328 7954 17356 8486
rect 17512 7954 17540 9114
rect 17604 8634 17632 9386
rect 17696 9042 17724 14214
rect 17788 12434 17816 14334
rect 17972 14074 18000 14350
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17788 12406 17908 12434
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 9518 17816 10406
rect 17880 10198 17908 12406
rect 18156 11762 18184 14214
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18248 11354 18276 13942
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18418 11248 18474 11257
rect 18418 11183 18420 11192
rect 18472 11183 18474 11192
rect 18420 11154 18472 11160
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 18432 10130 18460 10406
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17880 9518 17908 9930
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17972 9382 18000 9998
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17972 8974 18000 9318
rect 18524 9110 18552 19200
rect 18606 17980 18914 17989
rect 18606 17978 18612 17980
rect 18668 17978 18692 17980
rect 18748 17978 18772 17980
rect 18828 17978 18852 17980
rect 18908 17978 18914 17980
rect 18668 17926 18670 17978
rect 18850 17926 18852 17978
rect 18606 17924 18612 17926
rect 18668 17924 18692 17926
rect 18748 17924 18772 17926
rect 18828 17924 18852 17926
rect 18908 17924 18914 17926
rect 18606 17915 18914 17924
rect 18606 16892 18914 16901
rect 18606 16890 18612 16892
rect 18668 16890 18692 16892
rect 18748 16890 18772 16892
rect 18828 16890 18852 16892
rect 18908 16890 18914 16892
rect 18668 16838 18670 16890
rect 18850 16838 18852 16890
rect 18606 16836 18612 16838
rect 18668 16836 18692 16838
rect 18748 16836 18772 16838
rect 18828 16836 18852 16838
rect 18908 16836 18914 16838
rect 18606 16827 18914 16836
rect 18606 15804 18914 15813
rect 18606 15802 18612 15804
rect 18668 15802 18692 15804
rect 18748 15802 18772 15804
rect 18828 15802 18852 15804
rect 18908 15802 18914 15804
rect 18668 15750 18670 15802
rect 18850 15750 18852 15802
rect 18606 15748 18612 15750
rect 18668 15748 18692 15750
rect 18748 15748 18772 15750
rect 18828 15748 18852 15750
rect 18908 15748 18914 15750
rect 18606 15739 18914 15748
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18606 14716 18914 14725
rect 18606 14714 18612 14716
rect 18668 14714 18692 14716
rect 18748 14714 18772 14716
rect 18828 14714 18852 14716
rect 18908 14714 18914 14716
rect 18668 14662 18670 14714
rect 18850 14662 18852 14714
rect 18606 14660 18612 14662
rect 18668 14660 18692 14662
rect 18748 14660 18772 14662
rect 18828 14660 18852 14662
rect 18908 14660 18914 14662
rect 18606 14651 18914 14660
rect 19076 13705 19104 14758
rect 19062 13696 19118 13705
rect 18606 13628 18914 13637
rect 19062 13631 19118 13640
rect 18606 13626 18612 13628
rect 18668 13626 18692 13628
rect 18748 13626 18772 13628
rect 18828 13626 18852 13628
rect 18908 13626 18914 13628
rect 18668 13574 18670 13626
rect 18850 13574 18852 13626
rect 18606 13572 18612 13574
rect 18668 13572 18692 13574
rect 18748 13572 18772 13574
rect 18828 13572 18852 13574
rect 18908 13572 18914 13574
rect 18606 13563 18914 13572
rect 18606 12540 18914 12549
rect 18606 12538 18612 12540
rect 18668 12538 18692 12540
rect 18748 12538 18772 12540
rect 18828 12538 18852 12540
rect 18908 12538 18914 12540
rect 18668 12486 18670 12538
rect 18850 12486 18852 12538
rect 18606 12484 18612 12486
rect 18668 12484 18692 12486
rect 18748 12484 18772 12486
rect 18828 12484 18852 12486
rect 18908 12484 18914 12486
rect 18606 12475 18914 12484
rect 18606 11452 18914 11461
rect 18606 11450 18612 11452
rect 18668 11450 18692 11452
rect 18748 11450 18772 11452
rect 18828 11450 18852 11452
rect 18908 11450 18914 11452
rect 18668 11398 18670 11450
rect 18850 11398 18852 11450
rect 18606 11396 18612 11398
rect 18668 11396 18692 11398
rect 18748 11396 18772 11398
rect 18828 11396 18852 11398
rect 18908 11396 18914 11398
rect 18606 11387 18914 11396
rect 18606 10364 18914 10373
rect 18606 10362 18612 10364
rect 18668 10362 18692 10364
rect 18748 10362 18772 10364
rect 18828 10362 18852 10364
rect 18908 10362 18914 10364
rect 18668 10310 18670 10362
rect 18850 10310 18852 10362
rect 18606 10308 18612 10310
rect 18668 10308 18692 10310
rect 18748 10308 18772 10310
rect 18828 10308 18852 10310
rect 18908 10308 18914 10310
rect 18606 10299 18914 10308
rect 18606 9276 18914 9285
rect 18606 9274 18612 9276
rect 18668 9274 18692 9276
rect 18748 9274 18772 9276
rect 18828 9274 18852 9276
rect 18908 9274 18914 9276
rect 18668 9222 18670 9274
rect 18850 9222 18852 9274
rect 18606 9220 18612 9222
rect 18668 9220 18692 9222
rect 18748 9220 18772 9222
rect 18828 9220 18852 9222
rect 18908 9220 18914 9222
rect 18606 9211 18914 9220
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18420 8832 18472 8838
rect 17958 8800 18014 8809
rect 18420 8774 18472 8780
rect 17958 8735 18014 8744
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17056 7644 17364 7653
rect 17056 7642 17062 7644
rect 17118 7642 17142 7644
rect 17198 7642 17222 7644
rect 17278 7642 17302 7644
rect 17358 7642 17364 7644
rect 17118 7590 17120 7642
rect 17300 7590 17302 7642
rect 17056 7588 17062 7590
rect 17118 7588 17142 7590
rect 17198 7588 17222 7590
rect 17278 7588 17302 7590
rect 17358 7588 17364 7590
rect 17056 7579 17364 7588
rect 17512 7290 17540 7890
rect 17972 7342 18000 8735
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 17420 7262 17540 7290
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17056 6556 17364 6565
rect 17056 6554 17062 6556
rect 17118 6554 17142 6556
rect 17198 6554 17222 6556
rect 17278 6554 17302 6556
rect 17358 6554 17364 6556
rect 17118 6502 17120 6554
rect 17300 6502 17302 6554
rect 17056 6500 17062 6502
rect 17118 6500 17142 6502
rect 17198 6500 17222 6502
rect 17278 6500 17302 6502
rect 17358 6500 17364 6502
rect 17056 6491 17364 6500
rect 16948 6112 17000 6118
rect 16776 6038 16896 6066
rect 16948 6054 17000 6060
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16592 4078 16620 4694
rect 16776 4690 16804 5714
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16580 4072 16632 4078
rect 16500 4020 16580 4026
rect 16500 4014 16632 4020
rect 16500 3998 16620 4014
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16500 3618 16528 3998
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3738 16620 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16500 3590 16620 3618
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15200 2848 15252 2854
rect 15028 2796 15200 2802
rect 15028 2790 15252 2796
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 15028 2774 15240 2790
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 14844 2038 14872 2518
rect 15028 2446 15056 2774
rect 15506 2748 15814 2757
rect 15506 2746 15512 2748
rect 15568 2746 15592 2748
rect 15648 2746 15672 2748
rect 15728 2746 15752 2748
rect 15808 2746 15814 2748
rect 15568 2694 15570 2746
rect 15750 2694 15752 2746
rect 15506 2692 15512 2694
rect 15568 2692 15592 2694
rect 15648 2692 15672 2694
rect 15728 2692 15752 2694
rect 15808 2692 15814 2694
rect 15506 2683 15814 2692
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14832 2032 14884 2038
rect 14832 1974 14884 1980
rect 14936 1494 14964 2246
rect 15028 2106 15056 2382
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 15212 1970 15240 2382
rect 15200 1964 15252 1970
rect 15200 1906 15252 1912
rect 15396 1902 15424 2586
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 15016 1760 15068 1766
rect 15016 1702 15068 1708
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 15028 1426 15056 1702
rect 15396 1562 15424 1838
rect 15506 1660 15814 1669
rect 15506 1658 15512 1660
rect 15568 1658 15592 1660
rect 15648 1658 15672 1660
rect 15728 1658 15752 1660
rect 15808 1658 15814 1660
rect 15568 1606 15570 1658
rect 15750 1606 15752 1658
rect 15506 1604 15512 1606
rect 15568 1604 15592 1606
rect 15648 1604 15672 1606
rect 15728 1604 15752 1606
rect 15808 1604 15814 1606
rect 15506 1595 15814 1604
rect 15948 1562 15976 1838
rect 16224 1834 16252 2790
rect 16316 2106 16344 2790
rect 16500 2446 16528 3334
rect 16592 3126 16620 3590
rect 16684 3194 16712 4422
rect 16776 4282 16804 4626
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16868 4026 16896 6038
rect 16960 4690 16988 6054
rect 17056 5468 17364 5477
rect 17056 5466 17062 5468
rect 17118 5466 17142 5468
rect 17198 5466 17222 5468
rect 17278 5466 17302 5468
rect 17358 5466 17364 5468
rect 17118 5414 17120 5466
rect 17300 5414 17302 5466
rect 17056 5412 17062 5414
rect 17118 5412 17142 5414
rect 17198 5412 17222 5414
rect 17278 5412 17302 5414
rect 17358 5412 17364 5414
rect 17056 5403 17364 5412
rect 17420 4826 17448 7262
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6866 17540 7142
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17972 6458 18000 7278
rect 18156 7002 18184 7686
rect 18248 7002 18276 7890
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16960 4146 16988 4626
rect 17056 4380 17364 4389
rect 17056 4378 17062 4380
rect 17118 4378 17142 4380
rect 17198 4378 17222 4380
rect 17278 4378 17302 4380
rect 17358 4378 17364 4380
rect 17118 4326 17120 4378
rect 17300 4326 17302 4378
rect 17056 4324 17062 4326
rect 17118 4324 17142 4326
rect 17198 4324 17222 4326
rect 17278 4324 17302 4326
rect 17358 4324 17364 4326
rect 17056 4315 17364 4324
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16868 3998 16988 4026
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16592 2650 16620 3062
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16776 2582 16804 3878
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16500 1850 16528 2382
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16212 1828 16264 1834
rect 16212 1770 16264 1776
rect 16408 1822 16528 1850
rect 15384 1556 15436 1562
rect 15384 1498 15436 1504
rect 15936 1556 15988 1562
rect 15936 1498 15988 1504
rect 16408 1426 16436 1822
rect 16488 1760 16540 1766
rect 16488 1702 16540 1708
rect 16500 1494 16528 1702
rect 16488 1488 16540 1494
rect 16488 1430 16540 1436
rect 16776 1426 16804 2314
rect 16868 1970 16896 3402
rect 16960 1970 16988 3998
rect 17056 3292 17364 3301
rect 17056 3290 17062 3292
rect 17118 3290 17142 3292
rect 17198 3290 17222 3292
rect 17278 3290 17302 3292
rect 17358 3290 17364 3292
rect 17118 3238 17120 3290
rect 17300 3238 17302 3290
rect 17056 3236 17062 3238
rect 17118 3236 17142 3238
rect 17198 3236 17222 3238
rect 17278 3236 17302 3238
rect 17358 3236 17364 3238
rect 17056 3227 17364 3236
rect 17604 3194 17632 6394
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17788 4078 17816 4490
rect 17880 4146 17908 4626
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17512 2514 17540 3062
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17056 2204 17364 2213
rect 17056 2202 17062 2204
rect 17118 2202 17142 2204
rect 17198 2202 17222 2204
rect 17278 2202 17302 2204
rect 17358 2202 17364 2204
rect 17118 2150 17120 2202
rect 17300 2150 17302 2202
rect 17056 2148 17062 2150
rect 17118 2148 17142 2150
rect 17198 2148 17222 2150
rect 17278 2148 17302 2150
rect 17358 2148 17364 2150
rect 17056 2139 17364 2148
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 16868 1562 16896 1906
rect 17420 1834 17448 2450
rect 17696 2378 17724 3606
rect 17788 2650 17816 4014
rect 18064 3738 18092 6258
rect 18340 5914 18368 8026
rect 18432 7546 18460 8774
rect 18524 8634 18552 9046
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18606 8188 18914 8197
rect 18606 8186 18612 8188
rect 18668 8186 18692 8188
rect 18748 8186 18772 8188
rect 18828 8186 18852 8188
rect 18908 8186 18914 8188
rect 18668 8134 18670 8186
rect 18850 8134 18852 8186
rect 18606 8132 18612 8134
rect 18668 8132 18692 8134
rect 18748 8132 18772 8134
rect 18828 8132 18852 8134
rect 18908 8132 18914 8134
rect 18606 8123 18914 8132
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18606 7100 18914 7109
rect 18606 7098 18612 7100
rect 18668 7098 18692 7100
rect 18748 7098 18772 7100
rect 18828 7098 18852 7100
rect 18908 7098 18914 7100
rect 18668 7046 18670 7098
rect 18850 7046 18852 7098
rect 18606 7044 18612 7046
rect 18668 7044 18692 7046
rect 18748 7044 18772 7046
rect 18828 7044 18852 7046
rect 18908 7044 18914 7046
rect 18606 7035 18914 7044
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18432 5778 18460 6287
rect 18606 6012 18914 6021
rect 18606 6010 18612 6012
rect 18668 6010 18692 6012
rect 18748 6010 18772 6012
rect 18828 6010 18852 6012
rect 18908 6010 18914 6012
rect 18668 5958 18670 6010
rect 18850 5958 18852 6010
rect 18606 5956 18612 5958
rect 18668 5956 18692 5958
rect 18748 5956 18772 5958
rect 18828 5956 18852 5958
rect 18908 5956 18914 5958
rect 18606 5947 18914 5956
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18606 4924 18914 4933
rect 18606 4922 18612 4924
rect 18668 4922 18692 4924
rect 18748 4922 18772 4924
rect 18828 4922 18852 4924
rect 18908 4922 18914 4924
rect 18668 4870 18670 4922
rect 18850 4870 18852 4922
rect 18606 4868 18612 4870
rect 18668 4868 18692 4870
rect 18748 4868 18772 4870
rect 18828 4868 18852 4870
rect 18908 4868 18914 4870
rect 18606 4859 18914 4868
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18156 3602 18184 4422
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 19062 3904 19118 3913
rect 18340 3602 18368 3878
rect 18606 3836 18914 3845
rect 19062 3839 19118 3848
rect 18606 3834 18612 3836
rect 18668 3834 18692 3836
rect 18748 3834 18772 3836
rect 18828 3834 18852 3836
rect 18908 3834 18914 3836
rect 18668 3782 18670 3834
rect 18850 3782 18852 3834
rect 18606 3780 18612 3782
rect 18668 3780 18692 3782
rect 18748 3780 18772 3782
rect 18828 3780 18852 3782
rect 18908 3780 18914 3782
rect 18606 3771 18914 3780
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 17880 3194 17908 3538
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 19076 2990 19104 3839
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18606 2748 18914 2757
rect 18606 2746 18612 2748
rect 18668 2746 18692 2748
rect 18748 2746 18772 2748
rect 18828 2746 18852 2748
rect 18908 2746 18914 2748
rect 18668 2694 18670 2746
rect 18850 2694 18852 2746
rect 18606 2692 18612 2694
rect 18668 2692 18692 2694
rect 18748 2692 18772 2694
rect 18828 2692 18852 2694
rect 18908 2692 18914 2694
rect 18606 2683 18914 2692
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17408 1828 17460 1834
rect 17408 1770 17460 1776
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 17420 1426 17448 1770
rect 15016 1420 15068 1426
rect 15016 1362 15068 1368
rect 16396 1420 16448 1426
rect 16396 1362 16448 1368
rect 16764 1420 16816 1426
rect 16764 1362 16816 1368
rect 17408 1420 17460 1426
rect 17408 1362 17460 1368
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 17420 1222 17448 1362
rect 17880 1358 17908 2450
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 18432 1465 18460 1702
rect 18606 1660 18914 1669
rect 18606 1658 18612 1660
rect 18668 1658 18692 1660
rect 18748 1658 18772 1660
rect 18828 1658 18852 1660
rect 18908 1658 18914 1660
rect 18668 1606 18670 1658
rect 18850 1606 18852 1658
rect 18606 1604 18612 1606
rect 18668 1604 18692 1606
rect 18748 1604 18772 1606
rect 18828 1604 18852 1606
rect 18908 1604 18914 1606
rect 18606 1595 18914 1604
rect 18418 1456 18474 1465
rect 18418 1391 18474 1400
rect 17868 1352 17920 1358
rect 17868 1294 17920 1300
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 17408 1216 17460 1222
rect 17408 1158 17460 1164
rect 1556 1116 1864 1125
rect 1556 1114 1562 1116
rect 1618 1114 1642 1116
rect 1698 1114 1722 1116
rect 1778 1114 1802 1116
rect 1858 1114 1864 1116
rect 1618 1062 1620 1114
rect 1800 1062 1802 1114
rect 1556 1060 1562 1062
rect 1618 1060 1642 1062
rect 1698 1060 1722 1062
rect 1778 1060 1802 1062
rect 1858 1060 1864 1062
rect 1556 1051 1864 1060
rect 4656 1116 4964 1125
rect 4656 1114 4662 1116
rect 4718 1114 4742 1116
rect 4798 1114 4822 1116
rect 4878 1114 4902 1116
rect 4958 1114 4964 1116
rect 4718 1062 4720 1114
rect 4900 1062 4902 1114
rect 4656 1060 4662 1062
rect 4718 1060 4742 1062
rect 4798 1060 4822 1062
rect 4878 1060 4902 1062
rect 4958 1060 4964 1062
rect 4656 1051 4964 1060
rect 7756 1116 8064 1125
rect 7756 1114 7762 1116
rect 7818 1114 7842 1116
rect 7898 1114 7922 1116
rect 7978 1114 8002 1116
rect 8058 1114 8064 1116
rect 7818 1062 7820 1114
rect 8000 1062 8002 1114
rect 7756 1060 7762 1062
rect 7818 1060 7842 1062
rect 7898 1060 7922 1062
rect 7978 1060 8002 1062
rect 8058 1060 8064 1062
rect 7756 1051 8064 1060
rect 10856 1116 11164 1125
rect 10856 1114 10862 1116
rect 10918 1114 10942 1116
rect 10998 1114 11022 1116
rect 11078 1114 11102 1116
rect 11158 1114 11164 1116
rect 10918 1062 10920 1114
rect 11100 1062 11102 1114
rect 10856 1060 10862 1062
rect 10918 1060 10942 1062
rect 10998 1060 11022 1062
rect 11078 1060 11102 1062
rect 11158 1060 11164 1062
rect 10856 1051 11164 1060
rect 13956 1116 14264 1125
rect 13956 1114 13962 1116
rect 14018 1114 14042 1116
rect 14098 1114 14122 1116
rect 14178 1114 14202 1116
rect 14258 1114 14264 1116
rect 14018 1062 14020 1114
rect 14200 1062 14202 1114
rect 13956 1060 13962 1062
rect 14018 1060 14042 1062
rect 14098 1060 14122 1062
rect 14178 1060 14202 1062
rect 14258 1060 14264 1062
rect 13956 1051 14264 1060
rect 17056 1116 17364 1125
rect 17056 1114 17062 1116
rect 17118 1114 17142 1116
rect 17198 1114 17222 1116
rect 17278 1114 17302 1116
rect 17358 1114 17364 1116
rect 17118 1062 17120 1114
rect 17300 1062 17302 1114
rect 17056 1060 17062 1062
rect 17118 1060 17142 1062
rect 17198 1060 17222 1062
rect 17278 1060 17302 1062
rect 17358 1060 17364 1062
rect 17056 1051 17364 1060
rect 3106 572 3414 581
rect 3106 570 3112 572
rect 3168 570 3192 572
rect 3248 570 3272 572
rect 3328 570 3352 572
rect 3408 570 3414 572
rect 3168 518 3170 570
rect 3350 518 3352 570
rect 3106 516 3112 518
rect 3168 516 3192 518
rect 3248 516 3272 518
rect 3328 516 3352 518
rect 3408 516 3414 518
rect 3106 507 3414 516
rect 6206 572 6514 581
rect 6206 570 6212 572
rect 6268 570 6292 572
rect 6348 570 6372 572
rect 6428 570 6452 572
rect 6508 570 6514 572
rect 6268 518 6270 570
rect 6450 518 6452 570
rect 6206 516 6212 518
rect 6268 516 6292 518
rect 6348 516 6372 518
rect 6428 516 6452 518
rect 6508 516 6514 518
rect 6206 507 6514 516
rect 9306 572 9614 581
rect 9306 570 9312 572
rect 9368 570 9392 572
rect 9448 570 9472 572
rect 9528 570 9552 572
rect 9608 570 9614 572
rect 9368 518 9370 570
rect 9550 518 9552 570
rect 9306 516 9312 518
rect 9368 516 9392 518
rect 9448 516 9472 518
rect 9528 516 9552 518
rect 9608 516 9614 518
rect 9306 507 9614 516
rect 12406 572 12714 581
rect 12406 570 12412 572
rect 12468 570 12492 572
rect 12548 570 12572 572
rect 12628 570 12652 572
rect 12708 570 12714 572
rect 12468 518 12470 570
rect 12650 518 12652 570
rect 12406 516 12412 518
rect 12468 516 12492 518
rect 12548 516 12572 518
rect 12628 516 12652 518
rect 12708 516 12714 518
rect 12406 507 12714 516
rect 15506 572 15814 581
rect 15506 570 15512 572
rect 15568 570 15592 572
rect 15648 570 15672 572
rect 15728 570 15752 572
rect 15808 570 15814 572
rect 15568 518 15570 570
rect 15750 518 15752 570
rect 15506 516 15512 518
rect 15568 516 15592 518
rect 15648 516 15672 518
rect 15728 516 15752 518
rect 15808 516 15814 518
rect 15506 507 15814 516
rect 18606 572 18914 581
rect 18606 570 18612 572
rect 18668 570 18692 572
rect 18748 570 18772 572
rect 18828 570 18852 572
rect 18908 570 18914 572
rect 18668 518 18670 570
rect 18850 518 18852 570
rect 18606 516 18612 518
rect 18668 516 18692 518
rect 18748 516 18772 518
rect 18828 516 18852 518
rect 18908 516 18914 518
rect 18606 507 18914 516
<< via2 >>
rect 1562 18522 1618 18524
rect 1642 18522 1698 18524
rect 1722 18522 1778 18524
rect 1802 18522 1858 18524
rect 1562 18470 1608 18522
rect 1608 18470 1618 18522
rect 1642 18470 1672 18522
rect 1672 18470 1684 18522
rect 1684 18470 1698 18522
rect 1722 18470 1736 18522
rect 1736 18470 1748 18522
rect 1748 18470 1778 18522
rect 1802 18470 1812 18522
rect 1812 18470 1858 18522
rect 1562 18468 1618 18470
rect 1642 18468 1698 18470
rect 1722 18468 1778 18470
rect 1802 18468 1858 18470
rect 4662 18522 4718 18524
rect 4742 18522 4798 18524
rect 4822 18522 4878 18524
rect 4902 18522 4958 18524
rect 4662 18470 4708 18522
rect 4708 18470 4718 18522
rect 4742 18470 4772 18522
rect 4772 18470 4784 18522
rect 4784 18470 4798 18522
rect 4822 18470 4836 18522
rect 4836 18470 4848 18522
rect 4848 18470 4878 18522
rect 4902 18470 4912 18522
rect 4912 18470 4958 18522
rect 4662 18468 4718 18470
rect 4742 18468 4798 18470
rect 4822 18468 4878 18470
rect 4902 18468 4958 18470
rect 3112 17978 3168 17980
rect 3192 17978 3248 17980
rect 3272 17978 3328 17980
rect 3352 17978 3408 17980
rect 3112 17926 3158 17978
rect 3158 17926 3168 17978
rect 3192 17926 3222 17978
rect 3222 17926 3234 17978
rect 3234 17926 3248 17978
rect 3272 17926 3286 17978
rect 3286 17926 3298 17978
rect 3298 17926 3328 17978
rect 3352 17926 3362 17978
rect 3362 17926 3408 17978
rect 3112 17924 3168 17926
rect 3192 17924 3248 17926
rect 3272 17924 3328 17926
rect 3352 17924 3408 17926
rect 1562 17434 1618 17436
rect 1642 17434 1698 17436
rect 1722 17434 1778 17436
rect 1802 17434 1858 17436
rect 1562 17382 1608 17434
rect 1608 17382 1618 17434
rect 1642 17382 1672 17434
rect 1672 17382 1684 17434
rect 1684 17382 1698 17434
rect 1722 17382 1736 17434
rect 1736 17382 1748 17434
rect 1748 17382 1778 17434
rect 1802 17382 1812 17434
rect 1812 17382 1858 17434
rect 1562 17380 1618 17382
rect 1642 17380 1698 17382
rect 1722 17380 1778 17382
rect 1802 17380 1858 17382
rect 1562 16346 1618 16348
rect 1642 16346 1698 16348
rect 1722 16346 1778 16348
rect 1802 16346 1858 16348
rect 1562 16294 1608 16346
rect 1608 16294 1618 16346
rect 1642 16294 1672 16346
rect 1672 16294 1684 16346
rect 1684 16294 1698 16346
rect 1722 16294 1736 16346
rect 1736 16294 1748 16346
rect 1748 16294 1778 16346
rect 1802 16294 1812 16346
rect 1812 16294 1858 16346
rect 1562 16292 1618 16294
rect 1642 16292 1698 16294
rect 1722 16292 1778 16294
rect 1802 16292 1858 16294
rect 1562 15258 1618 15260
rect 1642 15258 1698 15260
rect 1722 15258 1778 15260
rect 1802 15258 1858 15260
rect 1562 15206 1608 15258
rect 1608 15206 1618 15258
rect 1642 15206 1672 15258
rect 1672 15206 1684 15258
rect 1684 15206 1698 15258
rect 1722 15206 1736 15258
rect 1736 15206 1748 15258
rect 1748 15206 1778 15258
rect 1802 15206 1812 15258
rect 1812 15206 1858 15258
rect 1562 15204 1618 15206
rect 1642 15204 1698 15206
rect 1722 15204 1778 15206
rect 1802 15204 1858 15206
rect 1562 14170 1618 14172
rect 1642 14170 1698 14172
rect 1722 14170 1778 14172
rect 1802 14170 1858 14172
rect 1562 14118 1608 14170
rect 1608 14118 1618 14170
rect 1642 14118 1672 14170
rect 1672 14118 1684 14170
rect 1684 14118 1698 14170
rect 1722 14118 1736 14170
rect 1736 14118 1748 14170
rect 1748 14118 1778 14170
rect 1802 14118 1812 14170
rect 1812 14118 1858 14170
rect 1562 14116 1618 14118
rect 1642 14116 1698 14118
rect 1722 14116 1778 14118
rect 1802 14116 1858 14118
rect 3112 16890 3168 16892
rect 3192 16890 3248 16892
rect 3272 16890 3328 16892
rect 3352 16890 3408 16892
rect 3112 16838 3158 16890
rect 3158 16838 3168 16890
rect 3192 16838 3222 16890
rect 3222 16838 3234 16890
rect 3234 16838 3248 16890
rect 3272 16838 3286 16890
rect 3286 16838 3298 16890
rect 3298 16838 3328 16890
rect 3352 16838 3362 16890
rect 3362 16838 3408 16890
rect 3112 16836 3168 16838
rect 3192 16836 3248 16838
rect 3272 16836 3328 16838
rect 3352 16836 3408 16838
rect 3112 15802 3168 15804
rect 3192 15802 3248 15804
rect 3272 15802 3328 15804
rect 3352 15802 3408 15804
rect 3112 15750 3158 15802
rect 3158 15750 3168 15802
rect 3192 15750 3222 15802
rect 3222 15750 3234 15802
rect 3234 15750 3248 15802
rect 3272 15750 3286 15802
rect 3286 15750 3298 15802
rect 3298 15750 3328 15802
rect 3352 15750 3362 15802
rect 3362 15750 3408 15802
rect 3112 15748 3168 15750
rect 3192 15748 3248 15750
rect 3272 15748 3328 15750
rect 3352 15748 3408 15750
rect 1562 13082 1618 13084
rect 1642 13082 1698 13084
rect 1722 13082 1778 13084
rect 1802 13082 1858 13084
rect 1562 13030 1608 13082
rect 1608 13030 1618 13082
rect 1642 13030 1672 13082
rect 1672 13030 1684 13082
rect 1684 13030 1698 13082
rect 1722 13030 1736 13082
rect 1736 13030 1748 13082
rect 1748 13030 1778 13082
rect 1802 13030 1812 13082
rect 1812 13030 1858 13082
rect 1562 13028 1618 13030
rect 1642 13028 1698 13030
rect 1722 13028 1778 13030
rect 1802 13028 1858 13030
rect 1562 11994 1618 11996
rect 1642 11994 1698 11996
rect 1722 11994 1778 11996
rect 1802 11994 1858 11996
rect 1562 11942 1608 11994
rect 1608 11942 1618 11994
rect 1642 11942 1672 11994
rect 1672 11942 1684 11994
rect 1684 11942 1698 11994
rect 1722 11942 1736 11994
rect 1736 11942 1748 11994
rect 1748 11942 1778 11994
rect 1802 11942 1812 11994
rect 1812 11942 1858 11994
rect 1562 11940 1618 11942
rect 1642 11940 1698 11942
rect 1722 11940 1778 11942
rect 1802 11940 1858 11942
rect 1562 10906 1618 10908
rect 1642 10906 1698 10908
rect 1722 10906 1778 10908
rect 1802 10906 1858 10908
rect 1562 10854 1608 10906
rect 1608 10854 1618 10906
rect 1642 10854 1672 10906
rect 1672 10854 1684 10906
rect 1684 10854 1698 10906
rect 1722 10854 1736 10906
rect 1736 10854 1748 10906
rect 1748 10854 1778 10906
rect 1802 10854 1812 10906
rect 1812 10854 1858 10906
rect 1562 10852 1618 10854
rect 1642 10852 1698 10854
rect 1722 10852 1778 10854
rect 1802 10852 1858 10854
rect 938 9968 994 10024
rect 1562 9818 1618 9820
rect 1642 9818 1698 9820
rect 1722 9818 1778 9820
rect 1802 9818 1858 9820
rect 1562 9766 1608 9818
rect 1608 9766 1618 9818
rect 1642 9766 1672 9818
rect 1672 9766 1684 9818
rect 1684 9766 1698 9818
rect 1722 9766 1736 9818
rect 1736 9766 1748 9818
rect 1748 9766 1778 9818
rect 1802 9766 1812 9818
rect 1812 9766 1858 9818
rect 1562 9764 1618 9766
rect 1642 9764 1698 9766
rect 1722 9764 1778 9766
rect 1802 9764 1858 9766
rect 3112 14714 3168 14716
rect 3192 14714 3248 14716
rect 3272 14714 3328 14716
rect 3352 14714 3408 14716
rect 3112 14662 3158 14714
rect 3158 14662 3168 14714
rect 3192 14662 3222 14714
rect 3222 14662 3234 14714
rect 3234 14662 3248 14714
rect 3272 14662 3286 14714
rect 3286 14662 3298 14714
rect 3298 14662 3328 14714
rect 3352 14662 3362 14714
rect 3362 14662 3408 14714
rect 3112 14660 3168 14662
rect 3192 14660 3248 14662
rect 3272 14660 3328 14662
rect 3352 14660 3408 14662
rect 3112 13626 3168 13628
rect 3192 13626 3248 13628
rect 3272 13626 3328 13628
rect 3352 13626 3408 13628
rect 3112 13574 3158 13626
rect 3158 13574 3168 13626
rect 3192 13574 3222 13626
rect 3222 13574 3234 13626
rect 3234 13574 3248 13626
rect 3272 13574 3286 13626
rect 3286 13574 3298 13626
rect 3298 13574 3328 13626
rect 3352 13574 3362 13626
rect 3362 13574 3408 13626
rect 3112 13572 3168 13574
rect 3192 13572 3248 13574
rect 3272 13572 3328 13574
rect 3352 13572 3408 13574
rect 3112 12538 3168 12540
rect 3192 12538 3248 12540
rect 3272 12538 3328 12540
rect 3352 12538 3408 12540
rect 3112 12486 3158 12538
rect 3158 12486 3168 12538
rect 3192 12486 3222 12538
rect 3222 12486 3234 12538
rect 3234 12486 3248 12538
rect 3272 12486 3286 12538
rect 3286 12486 3298 12538
rect 3298 12486 3328 12538
rect 3352 12486 3362 12538
rect 3362 12486 3408 12538
rect 3112 12484 3168 12486
rect 3192 12484 3248 12486
rect 3272 12484 3328 12486
rect 3352 12484 3408 12486
rect 3112 11450 3168 11452
rect 3192 11450 3248 11452
rect 3272 11450 3328 11452
rect 3352 11450 3408 11452
rect 3112 11398 3158 11450
rect 3158 11398 3168 11450
rect 3192 11398 3222 11450
rect 3222 11398 3234 11450
rect 3234 11398 3248 11450
rect 3272 11398 3286 11450
rect 3286 11398 3298 11450
rect 3298 11398 3328 11450
rect 3352 11398 3362 11450
rect 3362 11398 3408 11450
rect 3112 11396 3168 11398
rect 3192 11396 3248 11398
rect 3272 11396 3328 11398
rect 3352 11396 3408 11398
rect 1562 8730 1618 8732
rect 1642 8730 1698 8732
rect 1722 8730 1778 8732
rect 1802 8730 1858 8732
rect 1562 8678 1608 8730
rect 1608 8678 1618 8730
rect 1642 8678 1672 8730
rect 1672 8678 1684 8730
rect 1684 8678 1698 8730
rect 1722 8678 1736 8730
rect 1736 8678 1748 8730
rect 1748 8678 1778 8730
rect 1802 8678 1812 8730
rect 1812 8678 1858 8730
rect 1562 8676 1618 8678
rect 1642 8676 1698 8678
rect 1722 8676 1778 8678
rect 1802 8676 1858 8678
rect 1562 7642 1618 7644
rect 1642 7642 1698 7644
rect 1722 7642 1778 7644
rect 1802 7642 1858 7644
rect 1562 7590 1608 7642
rect 1608 7590 1618 7642
rect 1642 7590 1672 7642
rect 1672 7590 1684 7642
rect 1684 7590 1698 7642
rect 1722 7590 1736 7642
rect 1736 7590 1748 7642
rect 1748 7590 1778 7642
rect 1802 7590 1812 7642
rect 1812 7590 1858 7642
rect 1562 7588 1618 7590
rect 1642 7588 1698 7590
rect 1722 7588 1778 7590
rect 1802 7588 1858 7590
rect 1562 6554 1618 6556
rect 1642 6554 1698 6556
rect 1722 6554 1778 6556
rect 1802 6554 1858 6556
rect 1562 6502 1608 6554
rect 1608 6502 1618 6554
rect 1642 6502 1672 6554
rect 1672 6502 1684 6554
rect 1684 6502 1698 6554
rect 1722 6502 1736 6554
rect 1736 6502 1748 6554
rect 1748 6502 1778 6554
rect 1802 6502 1812 6554
rect 1812 6502 1858 6554
rect 1562 6500 1618 6502
rect 1642 6500 1698 6502
rect 1722 6500 1778 6502
rect 1802 6500 1858 6502
rect 1562 5466 1618 5468
rect 1642 5466 1698 5468
rect 1722 5466 1778 5468
rect 1802 5466 1858 5468
rect 1562 5414 1608 5466
rect 1608 5414 1618 5466
rect 1642 5414 1672 5466
rect 1672 5414 1684 5466
rect 1684 5414 1698 5466
rect 1722 5414 1736 5466
rect 1736 5414 1748 5466
rect 1748 5414 1778 5466
rect 1802 5414 1812 5466
rect 1812 5414 1858 5466
rect 1562 5412 1618 5414
rect 1642 5412 1698 5414
rect 1722 5412 1778 5414
rect 1802 5412 1858 5414
rect 1562 4378 1618 4380
rect 1642 4378 1698 4380
rect 1722 4378 1778 4380
rect 1802 4378 1858 4380
rect 1562 4326 1608 4378
rect 1608 4326 1618 4378
rect 1642 4326 1672 4378
rect 1672 4326 1684 4378
rect 1684 4326 1698 4378
rect 1722 4326 1736 4378
rect 1736 4326 1748 4378
rect 1748 4326 1778 4378
rect 1802 4326 1812 4378
rect 1812 4326 1858 4378
rect 1562 4324 1618 4326
rect 1642 4324 1698 4326
rect 1722 4324 1778 4326
rect 1802 4324 1858 4326
rect 3112 10362 3168 10364
rect 3192 10362 3248 10364
rect 3272 10362 3328 10364
rect 3352 10362 3408 10364
rect 3112 10310 3158 10362
rect 3158 10310 3168 10362
rect 3192 10310 3222 10362
rect 3222 10310 3234 10362
rect 3234 10310 3248 10362
rect 3272 10310 3286 10362
rect 3286 10310 3298 10362
rect 3298 10310 3328 10362
rect 3352 10310 3362 10362
rect 3362 10310 3408 10362
rect 3112 10308 3168 10310
rect 3192 10308 3248 10310
rect 3272 10308 3328 10310
rect 3352 10308 3408 10310
rect 4662 17434 4718 17436
rect 4742 17434 4798 17436
rect 4822 17434 4878 17436
rect 4902 17434 4958 17436
rect 4662 17382 4708 17434
rect 4708 17382 4718 17434
rect 4742 17382 4772 17434
rect 4772 17382 4784 17434
rect 4784 17382 4798 17434
rect 4822 17382 4836 17434
rect 4836 17382 4848 17434
rect 4848 17382 4878 17434
rect 4902 17382 4912 17434
rect 4912 17382 4958 17434
rect 4662 17380 4718 17382
rect 4742 17380 4798 17382
rect 4822 17380 4878 17382
rect 4902 17380 4958 17382
rect 4662 16346 4718 16348
rect 4742 16346 4798 16348
rect 4822 16346 4878 16348
rect 4902 16346 4958 16348
rect 4662 16294 4708 16346
rect 4708 16294 4718 16346
rect 4742 16294 4772 16346
rect 4772 16294 4784 16346
rect 4784 16294 4798 16346
rect 4822 16294 4836 16346
rect 4836 16294 4848 16346
rect 4848 16294 4878 16346
rect 4902 16294 4912 16346
rect 4912 16294 4958 16346
rect 4662 16292 4718 16294
rect 4742 16292 4798 16294
rect 4822 16292 4878 16294
rect 4902 16292 4958 16294
rect 4662 15258 4718 15260
rect 4742 15258 4798 15260
rect 4822 15258 4878 15260
rect 4902 15258 4958 15260
rect 4662 15206 4708 15258
rect 4708 15206 4718 15258
rect 4742 15206 4772 15258
rect 4772 15206 4784 15258
rect 4784 15206 4798 15258
rect 4822 15206 4836 15258
rect 4836 15206 4848 15258
rect 4848 15206 4878 15258
rect 4902 15206 4912 15258
rect 4912 15206 4958 15258
rect 4662 15204 4718 15206
rect 4742 15204 4798 15206
rect 4822 15204 4878 15206
rect 4902 15204 4958 15206
rect 6212 17978 6268 17980
rect 6292 17978 6348 17980
rect 6372 17978 6428 17980
rect 6452 17978 6508 17980
rect 6212 17926 6258 17978
rect 6258 17926 6268 17978
rect 6292 17926 6322 17978
rect 6322 17926 6334 17978
rect 6334 17926 6348 17978
rect 6372 17926 6386 17978
rect 6386 17926 6398 17978
rect 6398 17926 6428 17978
rect 6452 17926 6462 17978
rect 6462 17926 6508 17978
rect 6212 17924 6268 17926
rect 6292 17924 6348 17926
rect 6372 17924 6428 17926
rect 6452 17924 6508 17926
rect 7762 18522 7818 18524
rect 7842 18522 7898 18524
rect 7922 18522 7978 18524
rect 8002 18522 8058 18524
rect 7762 18470 7808 18522
rect 7808 18470 7818 18522
rect 7842 18470 7872 18522
rect 7872 18470 7884 18522
rect 7884 18470 7898 18522
rect 7922 18470 7936 18522
rect 7936 18470 7948 18522
rect 7948 18470 7978 18522
rect 8002 18470 8012 18522
rect 8012 18470 8058 18522
rect 7762 18468 7818 18470
rect 7842 18468 7898 18470
rect 7922 18468 7978 18470
rect 8002 18468 8058 18470
rect 7762 17434 7818 17436
rect 7842 17434 7898 17436
rect 7922 17434 7978 17436
rect 8002 17434 8058 17436
rect 7762 17382 7808 17434
rect 7808 17382 7818 17434
rect 7842 17382 7872 17434
rect 7872 17382 7884 17434
rect 7884 17382 7898 17434
rect 7922 17382 7936 17434
rect 7936 17382 7948 17434
rect 7948 17382 7978 17434
rect 8002 17382 8012 17434
rect 8012 17382 8058 17434
rect 7762 17380 7818 17382
rect 7842 17380 7898 17382
rect 7922 17380 7978 17382
rect 8002 17380 8058 17382
rect 6212 16890 6268 16892
rect 6292 16890 6348 16892
rect 6372 16890 6428 16892
rect 6452 16890 6508 16892
rect 6212 16838 6258 16890
rect 6258 16838 6268 16890
rect 6292 16838 6322 16890
rect 6322 16838 6334 16890
rect 6334 16838 6348 16890
rect 6372 16838 6386 16890
rect 6386 16838 6398 16890
rect 6398 16838 6428 16890
rect 6452 16838 6462 16890
rect 6462 16838 6508 16890
rect 6212 16836 6268 16838
rect 6292 16836 6348 16838
rect 6372 16836 6428 16838
rect 6452 16836 6508 16838
rect 7762 16346 7818 16348
rect 7842 16346 7898 16348
rect 7922 16346 7978 16348
rect 8002 16346 8058 16348
rect 7762 16294 7808 16346
rect 7808 16294 7818 16346
rect 7842 16294 7872 16346
rect 7872 16294 7884 16346
rect 7884 16294 7898 16346
rect 7922 16294 7936 16346
rect 7936 16294 7948 16346
rect 7948 16294 7978 16346
rect 8002 16294 8012 16346
rect 8012 16294 8058 16346
rect 7762 16292 7818 16294
rect 7842 16292 7898 16294
rect 7922 16292 7978 16294
rect 8002 16292 8058 16294
rect 6212 15802 6268 15804
rect 6292 15802 6348 15804
rect 6372 15802 6428 15804
rect 6452 15802 6508 15804
rect 6212 15750 6258 15802
rect 6258 15750 6268 15802
rect 6292 15750 6322 15802
rect 6322 15750 6334 15802
rect 6334 15750 6348 15802
rect 6372 15750 6386 15802
rect 6386 15750 6398 15802
rect 6398 15750 6428 15802
rect 6452 15750 6462 15802
rect 6462 15750 6508 15802
rect 6212 15748 6268 15750
rect 6292 15748 6348 15750
rect 6372 15748 6428 15750
rect 6452 15748 6508 15750
rect 6212 14714 6268 14716
rect 6292 14714 6348 14716
rect 6372 14714 6428 14716
rect 6452 14714 6508 14716
rect 6212 14662 6258 14714
rect 6258 14662 6268 14714
rect 6292 14662 6322 14714
rect 6322 14662 6334 14714
rect 6334 14662 6348 14714
rect 6372 14662 6386 14714
rect 6386 14662 6398 14714
rect 6398 14662 6428 14714
rect 6452 14662 6462 14714
rect 6462 14662 6508 14714
rect 6212 14660 6268 14662
rect 6292 14660 6348 14662
rect 6372 14660 6428 14662
rect 6452 14660 6508 14662
rect 4662 14170 4718 14172
rect 4742 14170 4798 14172
rect 4822 14170 4878 14172
rect 4902 14170 4958 14172
rect 4662 14118 4708 14170
rect 4708 14118 4718 14170
rect 4742 14118 4772 14170
rect 4772 14118 4784 14170
rect 4784 14118 4798 14170
rect 4822 14118 4836 14170
rect 4836 14118 4848 14170
rect 4848 14118 4878 14170
rect 4902 14118 4912 14170
rect 4912 14118 4958 14170
rect 4662 14116 4718 14118
rect 4742 14116 4798 14118
rect 4822 14116 4878 14118
rect 4902 14116 4958 14118
rect 7762 15258 7818 15260
rect 7842 15258 7898 15260
rect 7922 15258 7978 15260
rect 8002 15258 8058 15260
rect 7762 15206 7808 15258
rect 7808 15206 7818 15258
rect 7842 15206 7872 15258
rect 7872 15206 7884 15258
rect 7884 15206 7898 15258
rect 7922 15206 7936 15258
rect 7936 15206 7948 15258
rect 7948 15206 7978 15258
rect 8002 15206 8012 15258
rect 8012 15206 8058 15258
rect 7762 15204 7818 15206
rect 7842 15204 7898 15206
rect 7922 15204 7978 15206
rect 8002 15204 8058 15206
rect 10862 18522 10918 18524
rect 10942 18522 10998 18524
rect 11022 18522 11078 18524
rect 11102 18522 11158 18524
rect 10862 18470 10908 18522
rect 10908 18470 10918 18522
rect 10942 18470 10972 18522
rect 10972 18470 10984 18522
rect 10984 18470 10998 18522
rect 11022 18470 11036 18522
rect 11036 18470 11048 18522
rect 11048 18470 11078 18522
rect 11102 18470 11112 18522
rect 11112 18470 11158 18522
rect 10862 18468 10918 18470
rect 10942 18468 10998 18470
rect 11022 18468 11078 18470
rect 11102 18468 11158 18470
rect 9312 17978 9368 17980
rect 9392 17978 9448 17980
rect 9472 17978 9528 17980
rect 9552 17978 9608 17980
rect 9312 17926 9358 17978
rect 9358 17926 9368 17978
rect 9392 17926 9422 17978
rect 9422 17926 9434 17978
rect 9434 17926 9448 17978
rect 9472 17926 9486 17978
rect 9486 17926 9498 17978
rect 9498 17926 9528 17978
rect 9552 17926 9562 17978
rect 9562 17926 9608 17978
rect 9312 17924 9368 17926
rect 9392 17924 9448 17926
rect 9472 17924 9528 17926
rect 9552 17924 9608 17926
rect 7762 14170 7818 14172
rect 7842 14170 7898 14172
rect 7922 14170 7978 14172
rect 8002 14170 8058 14172
rect 7762 14118 7808 14170
rect 7808 14118 7818 14170
rect 7842 14118 7872 14170
rect 7872 14118 7884 14170
rect 7884 14118 7898 14170
rect 7922 14118 7936 14170
rect 7936 14118 7948 14170
rect 7948 14118 7978 14170
rect 8002 14118 8012 14170
rect 8012 14118 8058 14170
rect 7762 14116 7818 14118
rect 7842 14116 7898 14118
rect 7922 14116 7978 14118
rect 8002 14116 8058 14118
rect 4662 13082 4718 13084
rect 4742 13082 4798 13084
rect 4822 13082 4878 13084
rect 4902 13082 4958 13084
rect 4662 13030 4708 13082
rect 4708 13030 4718 13082
rect 4742 13030 4772 13082
rect 4772 13030 4784 13082
rect 4784 13030 4798 13082
rect 4822 13030 4836 13082
rect 4836 13030 4848 13082
rect 4848 13030 4878 13082
rect 4902 13030 4912 13082
rect 4912 13030 4958 13082
rect 4662 13028 4718 13030
rect 4742 13028 4798 13030
rect 4822 13028 4878 13030
rect 4902 13028 4958 13030
rect 4662 11994 4718 11996
rect 4742 11994 4798 11996
rect 4822 11994 4878 11996
rect 4902 11994 4958 11996
rect 4662 11942 4708 11994
rect 4708 11942 4718 11994
rect 4742 11942 4772 11994
rect 4772 11942 4784 11994
rect 4784 11942 4798 11994
rect 4822 11942 4836 11994
rect 4836 11942 4848 11994
rect 4848 11942 4878 11994
rect 4902 11942 4912 11994
rect 4912 11942 4958 11994
rect 4662 11940 4718 11942
rect 4742 11940 4798 11942
rect 4822 11940 4878 11942
rect 4902 11940 4958 11942
rect 4662 10906 4718 10908
rect 4742 10906 4798 10908
rect 4822 10906 4878 10908
rect 4902 10906 4958 10908
rect 4662 10854 4708 10906
rect 4708 10854 4718 10906
rect 4742 10854 4772 10906
rect 4772 10854 4784 10906
rect 4784 10854 4798 10906
rect 4822 10854 4836 10906
rect 4836 10854 4848 10906
rect 4848 10854 4878 10906
rect 4902 10854 4912 10906
rect 4912 10854 4958 10906
rect 4662 10852 4718 10854
rect 4742 10852 4798 10854
rect 4822 10852 4878 10854
rect 4902 10852 4958 10854
rect 3112 9274 3168 9276
rect 3192 9274 3248 9276
rect 3272 9274 3328 9276
rect 3352 9274 3408 9276
rect 3112 9222 3158 9274
rect 3158 9222 3168 9274
rect 3192 9222 3222 9274
rect 3222 9222 3234 9274
rect 3234 9222 3248 9274
rect 3272 9222 3286 9274
rect 3286 9222 3298 9274
rect 3298 9222 3328 9274
rect 3352 9222 3362 9274
rect 3362 9222 3408 9274
rect 3112 9220 3168 9222
rect 3192 9220 3248 9222
rect 3272 9220 3328 9222
rect 3352 9220 3408 9222
rect 4662 9818 4718 9820
rect 4742 9818 4798 9820
rect 4822 9818 4878 9820
rect 4902 9818 4958 9820
rect 4662 9766 4708 9818
rect 4708 9766 4718 9818
rect 4742 9766 4772 9818
rect 4772 9766 4784 9818
rect 4784 9766 4798 9818
rect 4822 9766 4836 9818
rect 4836 9766 4848 9818
rect 4848 9766 4878 9818
rect 4902 9766 4912 9818
rect 4912 9766 4958 9818
rect 4662 9764 4718 9766
rect 4742 9764 4798 9766
rect 4822 9764 4878 9766
rect 4902 9764 4958 9766
rect 6212 13626 6268 13628
rect 6292 13626 6348 13628
rect 6372 13626 6428 13628
rect 6452 13626 6508 13628
rect 6212 13574 6258 13626
rect 6258 13574 6268 13626
rect 6292 13574 6322 13626
rect 6322 13574 6334 13626
rect 6334 13574 6348 13626
rect 6372 13574 6386 13626
rect 6386 13574 6398 13626
rect 6398 13574 6428 13626
rect 6452 13574 6462 13626
rect 6462 13574 6508 13626
rect 6212 13572 6268 13574
rect 6292 13572 6348 13574
rect 6372 13572 6428 13574
rect 6452 13572 6508 13574
rect 6212 12538 6268 12540
rect 6292 12538 6348 12540
rect 6372 12538 6428 12540
rect 6452 12538 6508 12540
rect 6212 12486 6258 12538
rect 6258 12486 6268 12538
rect 6292 12486 6322 12538
rect 6322 12486 6334 12538
rect 6334 12486 6348 12538
rect 6372 12486 6386 12538
rect 6386 12486 6398 12538
rect 6398 12486 6428 12538
rect 6452 12486 6462 12538
rect 6462 12486 6508 12538
rect 6212 12484 6268 12486
rect 6292 12484 6348 12486
rect 6372 12484 6428 12486
rect 6452 12484 6508 12486
rect 3112 8186 3168 8188
rect 3192 8186 3248 8188
rect 3272 8186 3328 8188
rect 3352 8186 3408 8188
rect 3112 8134 3158 8186
rect 3158 8134 3168 8186
rect 3192 8134 3222 8186
rect 3222 8134 3234 8186
rect 3234 8134 3248 8186
rect 3272 8134 3286 8186
rect 3286 8134 3298 8186
rect 3298 8134 3328 8186
rect 3352 8134 3362 8186
rect 3362 8134 3408 8186
rect 3112 8132 3168 8134
rect 3192 8132 3248 8134
rect 3272 8132 3328 8134
rect 3352 8132 3408 8134
rect 3112 7098 3168 7100
rect 3192 7098 3248 7100
rect 3272 7098 3328 7100
rect 3352 7098 3408 7100
rect 3112 7046 3158 7098
rect 3158 7046 3168 7098
rect 3192 7046 3222 7098
rect 3222 7046 3234 7098
rect 3234 7046 3248 7098
rect 3272 7046 3286 7098
rect 3286 7046 3298 7098
rect 3298 7046 3328 7098
rect 3352 7046 3362 7098
rect 3362 7046 3408 7098
rect 3112 7044 3168 7046
rect 3192 7044 3248 7046
rect 3272 7044 3328 7046
rect 3352 7044 3408 7046
rect 3112 6010 3168 6012
rect 3192 6010 3248 6012
rect 3272 6010 3328 6012
rect 3352 6010 3408 6012
rect 3112 5958 3158 6010
rect 3158 5958 3168 6010
rect 3192 5958 3222 6010
rect 3222 5958 3234 6010
rect 3234 5958 3248 6010
rect 3272 5958 3286 6010
rect 3286 5958 3298 6010
rect 3298 5958 3328 6010
rect 3352 5958 3362 6010
rect 3362 5958 3408 6010
rect 3112 5956 3168 5958
rect 3192 5956 3248 5958
rect 3272 5956 3328 5958
rect 3352 5956 3408 5958
rect 1562 3290 1618 3292
rect 1642 3290 1698 3292
rect 1722 3290 1778 3292
rect 1802 3290 1858 3292
rect 1562 3238 1608 3290
rect 1608 3238 1618 3290
rect 1642 3238 1672 3290
rect 1672 3238 1684 3290
rect 1684 3238 1698 3290
rect 1722 3238 1736 3290
rect 1736 3238 1748 3290
rect 1748 3238 1778 3290
rect 1802 3238 1812 3290
rect 1812 3238 1858 3290
rect 1562 3236 1618 3238
rect 1642 3236 1698 3238
rect 1722 3236 1778 3238
rect 1802 3236 1858 3238
rect 1562 2202 1618 2204
rect 1642 2202 1698 2204
rect 1722 2202 1778 2204
rect 1802 2202 1858 2204
rect 1562 2150 1608 2202
rect 1608 2150 1618 2202
rect 1642 2150 1672 2202
rect 1672 2150 1684 2202
rect 1684 2150 1698 2202
rect 1722 2150 1736 2202
rect 1736 2150 1748 2202
rect 1748 2150 1778 2202
rect 1802 2150 1812 2202
rect 1812 2150 1858 2202
rect 1562 2148 1618 2150
rect 1642 2148 1698 2150
rect 1722 2148 1778 2150
rect 1802 2148 1858 2150
rect 3112 4922 3168 4924
rect 3192 4922 3248 4924
rect 3272 4922 3328 4924
rect 3352 4922 3408 4924
rect 3112 4870 3158 4922
rect 3158 4870 3168 4922
rect 3192 4870 3222 4922
rect 3222 4870 3234 4922
rect 3234 4870 3248 4922
rect 3272 4870 3286 4922
rect 3286 4870 3298 4922
rect 3298 4870 3328 4922
rect 3352 4870 3362 4922
rect 3362 4870 3408 4922
rect 3112 4868 3168 4870
rect 3192 4868 3248 4870
rect 3272 4868 3328 4870
rect 3352 4868 3408 4870
rect 3112 3834 3168 3836
rect 3192 3834 3248 3836
rect 3272 3834 3328 3836
rect 3352 3834 3408 3836
rect 3112 3782 3158 3834
rect 3158 3782 3168 3834
rect 3192 3782 3222 3834
rect 3222 3782 3234 3834
rect 3234 3782 3248 3834
rect 3272 3782 3286 3834
rect 3286 3782 3298 3834
rect 3298 3782 3328 3834
rect 3352 3782 3362 3834
rect 3362 3782 3408 3834
rect 3112 3780 3168 3782
rect 3192 3780 3248 3782
rect 3272 3780 3328 3782
rect 3352 3780 3408 3782
rect 4662 8730 4718 8732
rect 4742 8730 4798 8732
rect 4822 8730 4878 8732
rect 4902 8730 4958 8732
rect 4662 8678 4708 8730
rect 4708 8678 4718 8730
rect 4742 8678 4772 8730
rect 4772 8678 4784 8730
rect 4784 8678 4798 8730
rect 4822 8678 4836 8730
rect 4836 8678 4848 8730
rect 4848 8678 4878 8730
rect 4902 8678 4912 8730
rect 4912 8678 4958 8730
rect 4662 8676 4718 8678
rect 4742 8676 4798 8678
rect 4822 8676 4878 8678
rect 4902 8676 4958 8678
rect 4662 7642 4718 7644
rect 4742 7642 4798 7644
rect 4822 7642 4878 7644
rect 4902 7642 4958 7644
rect 4662 7590 4708 7642
rect 4708 7590 4718 7642
rect 4742 7590 4772 7642
rect 4772 7590 4784 7642
rect 4784 7590 4798 7642
rect 4822 7590 4836 7642
rect 4836 7590 4848 7642
rect 4848 7590 4878 7642
rect 4902 7590 4912 7642
rect 4912 7590 4958 7642
rect 4662 7588 4718 7590
rect 4742 7588 4798 7590
rect 4822 7588 4878 7590
rect 4902 7588 4958 7590
rect 3112 2746 3168 2748
rect 3192 2746 3248 2748
rect 3272 2746 3328 2748
rect 3352 2746 3408 2748
rect 3112 2694 3158 2746
rect 3158 2694 3168 2746
rect 3192 2694 3222 2746
rect 3222 2694 3234 2746
rect 3234 2694 3248 2746
rect 3272 2694 3286 2746
rect 3286 2694 3298 2746
rect 3298 2694 3328 2746
rect 3352 2694 3362 2746
rect 3362 2694 3408 2746
rect 3112 2692 3168 2694
rect 3192 2692 3248 2694
rect 3272 2692 3328 2694
rect 3352 2692 3408 2694
rect 4662 6554 4718 6556
rect 4742 6554 4798 6556
rect 4822 6554 4878 6556
rect 4902 6554 4958 6556
rect 4662 6502 4708 6554
rect 4708 6502 4718 6554
rect 4742 6502 4772 6554
rect 4772 6502 4784 6554
rect 4784 6502 4798 6554
rect 4822 6502 4836 6554
rect 4836 6502 4848 6554
rect 4848 6502 4878 6554
rect 4902 6502 4912 6554
rect 4912 6502 4958 6554
rect 4662 6500 4718 6502
rect 4742 6500 4798 6502
rect 4822 6500 4878 6502
rect 4902 6500 4958 6502
rect 4662 5466 4718 5468
rect 4742 5466 4798 5468
rect 4822 5466 4878 5468
rect 4902 5466 4958 5468
rect 4662 5414 4708 5466
rect 4708 5414 4718 5466
rect 4742 5414 4772 5466
rect 4772 5414 4784 5466
rect 4784 5414 4798 5466
rect 4822 5414 4836 5466
rect 4836 5414 4848 5466
rect 4848 5414 4878 5466
rect 4902 5414 4912 5466
rect 4912 5414 4958 5466
rect 4662 5412 4718 5414
rect 4742 5412 4798 5414
rect 4822 5412 4878 5414
rect 4902 5412 4958 5414
rect 6212 11450 6268 11452
rect 6292 11450 6348 11452
rect 6372 11450 6428 11452
rect 6452 11450 6508 11452
rect 6212 11398 6258 11450
rect 6258 11398 6268 11450
rect 6292 11398 6322 11450
rect 6322 11398 6334 11450
rect 6334 11398 6348 11450
rect 6372 11398 6386 11450
rect 6386 11398 6398 11450
rect 6398 11398 6428 11450
rect 6452 11398 6462 11450
rect 6462 11398 6508 11450
rect 6212 11396 6268 11398
rect 6292 11396 6348 11398
rect 6372 11396 6428 11398
rect 6452 11396 6508 11398
rect 6212 10362 6268 10364
rect 6292 10362 6348 10364
rect 6372 10362 6428 10364
rect 6452 10362 6508 10364
rect 6212 10310 6258 10362
rect 6258 10310 6268 10362
rect 6292 10310 6322 10362
rect 6322 10310 6334 10362
rect 6334 10310 6348 10362
rect 6372 10310 6386 10362
rect 6386 10310 6398 10362
rect 6398 10310 6428 10362
rect 6452 10310 6462 10362
rect 6462 10310 6508 10362
rect 6212 10308 6268 10310
rect 6292 10308 6348 10310
rect 6372 10308 6428 10310
rect 6452 10308 6508 10310
rect 6212 9274 6268 9276
rect 6292 9274 6348 9276
rect 6372 9274 6428 9276
rect 6452 9274 6508 9276
rect 6212 9222 6258 9274
rect 6258 9222 6268 9274
rect 6292 9222 6322 9274
rect 6322 9222 6334 9274
rect 6334 9222 6348 9274
rect 6372 9222 6386 9274
rect 6386 9222 6398 9274
rect 6398 9222 6428 9274
rect 6452 9222 6462 9274
rect 6462 9222 6508 9274
rect 6212 9220 6268 9222
rect 6292 9220 6348 9222
rect 6372 9220 6428 9222
rect 6452 9220 6508 9222
rect 4662 4378 4718 4380
rect 4742 4378 4798 4380
rect 4822 4378 4878 4380
rect 4902 4378 4958 4380
rect 4662 4326 4708 4378
rect 4708 4326 4718 4378
rect 4742 4326 4772 4378
rect 4772 4326 4784 4378
rect 4784 4326 4798 4378
rect 4822 4326 4836 4378
rect 4836 4326 4848 4378
rect 4848 4326 4878 4378
rect 4902 4326 4912 4378
rect 4912 4326 4958 4378
rect 4662 4324 4718 4326
rect 4742 4324 4798 4326
rect 4822 4324 4878 4326
rect 4902 4324 4958 4326
rect 6212 8186 6268 8188
rect 6292 8186 6348 8188
rect 6372 8186 6428 8188
rect 6452 8186 6508 8188
rect 6212 8134 6258 8186
rect 6258 8134 6268 8186
rect 6292 8134 6322 8186
rect 6322 8134 6334 8186
rect 6334 8134 6348 8186
rect 6372 8134 6386 8186
rect 6386 8134 6398 8186
rect 6398 8134 6428 8186
rect 6452 8134 6462 8186
rect 6462 8134 6508 8186
rect 6212 8132 6268 8134
rect 6292 8132 6348 8134
rect 6372 8132 6428 8134
rect 6452 8132 6508 8134
rect 6212 7098 6268 7100
rect 6292 7098 6348 7100
rect 6372 7098 6428 7100
rect 6452 7098 6508 7100
rect 6212 7046 6258 7098
rect 6258 7046 6268 7098
rect 6292 7046 6322 7098
rect 6322 7046 6334 7098
rect 6334 7046 6348 7098
rect 6372 7046 6386 7098
rect 6386 7046 6398 7098
rect 6398 7046 6428 7098
rect 6452 7046 6462 7098
rect 6462 7046 6508 7098
rect 6212 7044 6268 7046
rect 6292 7044 6348 7046
rect 6372 7044 6428 7046
rect 6452 7044 6508 7046
rect 4662 3290 4718 3292
rect 4742 3290 4798 3292
rect 4822 3290 4878 3292
rect 4902 3290 4958 3292
rect 4662 3238 4708 3290
rect 4708 3238 4718 3290
rect 4742 3238 4772 3290
rect 4772 3238 4784 3290
rect 4784 3238 4798 3290
rect 4822 3238 4836 3290
rect 4836 3238 4848 3290
rect 4848 3238 4878 3290
rect 4902 3238 4912 3290
rect 4912 3238 4958 3290
rect 4662 3236 4718 3238
rect 4742 3236 4798 3238
rect 4822 3236 4878 3238
rect 4902 3236 4958 3238
rect 4662 2202 4718 2204
rect 4742 2202 4798 2204
rect 4822 2202 4878 2204
rect 4902 2202 4958 2204
rect 4662 2150 4708 2202
rect 4708 2150 4718 2202
rect 4742 2150 4772 2202
rect 4772 2150 4784 2202
rect 4784 2150 4798 2202
rect 4822 2150 4836 2202
rect 4836 2150 4848 2202
rect 4848 2150 4878 2202
rect 4902 2150 4912 2202
rect 4912 2150 4958 2202
rect 4662 2148 4718 2150
rect 4742 2148 4798 2150
rect 4822 2148 4878 2150
rect 4902 2148 4958 2150
rect 3112 1658 3168 1660
rect 3192 1658 3248 1660
rect 3272 1658 3328 1660
rect 3352 1658 3408 1660
rect 3112 1606 3158 1658
rect 3158 1606 3168 1658
rect 3192 1606 3222 1658
rect 3222 1606 3234 1658
rect 3234 1606 3248 1658
rect 3272 1606 3286 1658
rect 3286 1606 3298 1658
rect 3298 1606 3328 1658
rect 3352 1606 3362 1658
rect 3362 1606 3408 1658
rect 3112 1604 3168 1606
rect 3192 1604 3248 1606
rect 3272 1604 3328 1606
rect 3352 1604 3408 1606
rect 6212 6010 6268 6012
rect 6292 6010 6348 6012
rect 6372 6010 6428 6012
rect 6452 6010 6508 6012
rect 6212 5958 6258 6010
rect 6258 5958 6268 6010
rect 6292 5958 6322 6010
rect 6322 5958 6334 6010
rect 6334 5958 6348 6010
rect 6372 5958 6386 6010
rect 6386 5958 6398 6010
rect 6398 5958 6428 6010
rect 6452 5958 6462 6010
rect 6462 5958 6508 6010
rect 6212 5956 6268 5958
rect 6292 5956 6348 5958
rect 6372 5956 6428 5958
rect 6452 5956 6508 5958
rect 6212 4922 6268 4924
rect 6292 4922 6348 4924
rect 6372 4922 6428 4924
rect 6452 4922 6508 4924
rect 6212 4870 6258 4922
rect 6258 4870 6268 4922
rect 6292 4870 6322 4922
rect 6322 4870 6334 4922
rect 6334 4870 6348 4922
rect 6372 4870 6386 4922
rect 6386 4870 6398 4922
rect 6398 4870 6428 4922
rect 6452 4870 6462 4922
rect 6462 4870 6508 4922
rect 6212 4868 6268 4870
rect 6292 4868 6348 4870
rect 6372 4868 6428 4870
rect 6452 4868 6508 4870
rect 7762 13082 7818 13084
rect 7842 13082 7898 13084
rect 7922 13082 7978 13084
rect 8002 13082 8058 13084
rect 7762 13030 7808 13082
rect 7808 13030 7818 13082
rect 7842 13030 7872 13082
rect 7872 13030 7884 13082
rect 7884 13030 7898 13082
rect 7922 13030 7936 13082
rect 7936 13030 7948 13082
rect 7948 13030 7978 13082
rect 8002 13030 8012 13082
rect 8012 13030 8058 13082
rect 7762 13028 7818 13030
rect 7842 13028 7898 13030
rect 7922 13028 7978 13030
rect 8002 13028 8058 13030
rect 7762 11994 7818 11996
rect 7842 11994 7898 11996
rect 7922 11994 7978 11996
rect 8002 11994 8058 11996
rect 7762 11942 7808 11994
rect 7808 11942 7818 11994
rect 7842 11942 7872 11994
rect 7872 11942 7884 11994
rect 7884 11942 7898 11994
rect 7922 11942 7936 11994
rect 7936 11942 7948 11994
rect 7948 11942 7978 11994
rect 8002 11942 8012 11994
rect 8012 11942 8058 11994
rect 7762 11940 7818 11942
rect 7842 11940 7898 11942
rect 7922 11940 7978 11942
rect 8002 11940 8058 11942
rect 7762 10906 7818 10908
rect 7842 10906 7898 10908
rect 7922 10906 7978 10908
rect 8002 10906 8058 10908
rect 7762 10854 7808 10906
rect 7808 10854 7818 10906
rect 7842 10854 7872 10906
rect 7872 10854 7884 10906
rect 7884 10854 7898 10906
rect 7922 10854 7936 10906
rect 7936 10854 7948 10906
rect 7948 10854 7978 10906
rect 8002 10854 8012 10906
rect 8012 10854 8058 10906
rect 7762 10852 7818 10854
rect 7842 10852 7898 10854
rect 7922 10852 7978 10854
rect 8002 10852 8058 10854
rect 7762 9818 7818 9820
rect 7842 9818 7898 9820
rect 7922 9818 7978 9820
rect 8002 9818 8058 9820
rect 7762 9766 7808 9818
rect 7808 9766 7818 9818
rect 7842 9766 7872 9818
rect 7872 9766 7884 9818
rect 7884 9766 7898 9818
rect 7922 9766 7936 9818
rect 7936 9766 7948 9818
rect 7948 9766 7978 9818
rect 8002 9766 8012 9818
rect 8012 9766 8058 9818
rect 7762 9764 7818 9766
rect 7842 9764 7898 9766
rect 7922 9764 7978 9766
rect 8002 9764 8058 9766
rect 9312 16890 9368 16892
rect 9392 16890 9448 16892
rect 9472 16890 9528 16892
rect 9552 16890 9608 16892
rect 9312 16838 9358 16890
rect 9358 16838 9368 16890
rect 9392 16838 9422 16890
rect 9422 16838 9434 16890
rect 9434 16838 9448 16890
rect 9472 16838 9486 16890
rect 9486 16838 9498 16890
rect 9498 16838 9528 16890
rect 9552 16838 9562 16890
rect 9562 16838 9608 16890
rect 9312 16836 9368 16838
rect 9392 16836 9448 16838
rect 9472 16836 9528 16838
rect 9552 16836 9608 16838
rect 9312 15802 9368 15804
rect 9392 15802 9448 15804
rect 9472 15802 9528 15804
rect 9552 15802 9608 15804
rect 9312 15750 9358 15802
rect 9358 15750 9368 15802
rect 9392 15750 9422 15802
rect 9422 15750 9434 15802
rect 9434 15750 9448 15802
rect 9472 15750 9486 15802
rect 9486 15750 9498 15802
rect 9498 15750 9528 15802
rect 9552 15750 9562 15802
rect 9562 15750 9608 15802
rect 9312 15748 9368 15750
rect 9392 15748 9448 15750
rect 9472 15748 9528 15750
rect 9552 15748 9608 15750
rect 9312 14714 9368 14716
rect 9392 14714 9448 14716
rect 9472 14714 9528 14716
rect 9552 14714 9608 14716
rect 9312 14662 9358 14714
rect 9358 14662 9368 14714
rect 9392 14662 9422 14714
rect 9422 14662 9434 14714
rect 9434 14662 9448 14714
rect 9472 14662 9486 14714
rect 9486 14662 9498 14714
rect 9498 14662 9528 14714
rect 9552 14662 9562 14714
rect 9562 14662 9608 14714
rect 9312 14660 9368 14662
rect 9392 14660 9448 14662
rect 9472 14660 9528 14662
rect 9552 14660 9608 14662
rect 9312 13626 9368 13628
rect 9392 13626 9448 13628
rect 9472 13626 9528 13628
rect 9552 13626 9608 13628
rect 9312 13574 9358 13626
rect 9358 13574 9368 13626
rect 9392 13574 9422 13626
rect 9422 13574 9434 13626
rect 9434 13574 9448 13626
rect 9472 13574 9486 13626
rect 9486 13574 9498 13626
rect 9498 13574 9528 13626
rect 9552 13574 9562 13626
rect 9562 13574 9608 13626
rect 9312 13572 9368 13574
rect 9392 13572 9448 13574
rect 9472 13572 9528 13574
rect 9552 13572 9608 13574
rect 9312 12538 9368 12540
rect 9392 12538 9448 12540
rect 9472 12538 9528 12540
rect 9552 12538 9608 12540
rect 9312 12486 9358 12538
rect 9358 12486 9368 12538
rect 9392 12486 9422 12538
rect 9422 12486 9434 12538
rect 9434 12486 9448 12538
rect 9472 12486 9486 12538
rect 9486 12486 9498 12538
rect 9498 12486 9528 12538
rect 9552 12486 9562 12538
rect 9562 12486 9608 12538
rect 9312 12484 9368 12486
rect 9392 12484 9448 12486
rect 9472 12484 9528 12486
rect 9552 12484 9608 12486
rect 12412 17978 12468 17980
rect 12492 17978 12548 17980
rect 12572 17978 12628 17980
rect 12652 17978 12708 17980
rect 12412 17926 12458 17978
rect 12458 17926 12468 17978
rect 12492 17926 12522 17978
rect 12522 17926 12534 17978
rect 12534 17926 12548 17978
rect 12572 17926 12586 17978
rect 12586 17926 12598 17978
rect 12598 17926 12628 17978
rect 12652 17926 12662 17978
rect 12662 17926 12708 17978
rect 12412 17924 12468 17926
rect 12492 17924 12548 17926
rect 12572 17924 12628 17926
rect 12652 17924 12708 17926
rect 13962 18522 14018 18524
rect 14042 18522 14098 18524
rect 14122 18522 14178 18524
rect 14202 18522 14258 18524
rect 13962 18470 14008 18522
rect 14008 18470 14018 18522
rect 14042 18470 14072 18522
rect 14072 18470 14084 18522
rect 14084 18470 14098 18522
rect 14122 18470 14136 18522
rect 14136 18470 14148 18522
rect 14148 18470 14178 18522
rect 14202 18470 14212 18522
rect 14212 18470 14258 18522
rect 13962 18468 14018 18470
rect 14042 18468 14098 18470
rect 14122 18468 14178 18470
rect 14202 18468 14258 18470
rect 10862 17434 10918 17436
rect 10942 17434 10998 17436
rect 11022 17434 11078 17436
rect 11102 17434 11158 17436
rect 10862 17382 10908 17434
rect 10908 17382 10918 17434
rect 10942 17382 10972 17434
rect 10972 17382 10984 17434
rect 10984 17382 10998 17434
rect 11022 17382 11036 17434
rect 11036 17382 11048 17434
rect 11048 17382 11078 17434
rect 11102 17382 11112 17434
rect 11112 17382 11158 17434
rect 10862 17380 10918 17382
rect 10942 17380 10998 17382
rect 11022 17380 11078 17382
rect 11102 17380 11158 17382
rect 10862 16346 10918 16348
rect 10942 16346 10998 16348
rect 11022 16346 11078 16348
rect 11102 16346 11158 16348
rect 10862 16294 10908 16346
rect 10908 16294 10918 16346
rect 10942 16294 10972 16346
rect 10972 16294 10984 16346
rect 10984 16294 10998 16346
rect 11022 16294 11036 16346
rect 11036 16294 11048 16346
rect 11048 16294 11078 16346
rect 11102 16294 11112 16346
rect 11112 16294 11158 16346
rect 10862 16292 10918 16294
rect 10942 16292 10998 16294
rect 11022 16292 11078 16294
rect 11102 16292 11158 16294
rect 12412 16890 12468 16892
rect 12492 16890 12548 16892
rect 12572 16890 12628 16892
rect 12652 16890 12708 16892
rect 12412 16838 12458 16890
rect 12458 16838 12468 16890
rect 12492 16838 12522 16890
rect 12522 16838 12534 16890
rect 12534 16838 12548 16890
rect 12572 16838 12586 16890
rect 12586 16838 12598 16890
rect 12598 16838 12628 16890
rect 12652 16838 12662 16890
rect 12662 16838 12708 16890
rect 12412 16836 12468 16838
rect 12492 16836 12548 16838
rect 12572 16836 12628 16838
rect 12652 16836 12708 16838
rect 10862 15258 10918 15260
rect 10942 15258 10998 15260
rect 11022 15258 11078 15260
rect 11102 15258 11158 15260
rect 10862 15206 10908 15258
rect 10908 15206 10918 15258
rect 10942 15206 10972 15258
rect 10972 15206 10984 15258
rect 10984 15206 10998 15258
rect 11022 15206 11036 15258
rect 11036 15206 11048 15258
rect 11048 15206 11078 15258
rect 11102 15206 11112 15258
rect 11112 15206 11158 15258
rect 10862 15204 10918 15206
rect 10942 15204 10998 15206
rect 11022 15204 11078 15206
rect 11102 15204 11158 15206
rect 10862 14170 10918 14172
rect 10942 14170 10998 14172
rect 11022 14170 11078 14172
rect 11102 14170 11158 14172
rect 10862 14118 10908 14170
rect 10908 14118 10918 14170
rect 10942 14118 10972 14170
rect 10972 14118 10984 14170
rect 10984 14118 10998 14170
rect 11022 14118 11036 14170
rect 11036 14118 11048 14170
rect 11048 14118 11078 14170
rect 11102 14118 11112 14170
rect 11112 14118 11158 14170
rect 10862 14116 10918 14118
rect 10942 14116 10998 14118
rect 11022 14116 11078 14118
rect 11102 14116 11158 14118
rect 9312 11450 9368 11452
rect 9392 11450 9448 11452
rect 9472 11450 9528 11452
rect 9552 11450 9608 11452
rect 9312 11398 9358 11450
rect 9358 11398 9368 11450
rect 9392 11398 9422 11450
rect 9422 11398 9434 11450
rect 9434 11398 9448 11450
rect 9472 11398 9486 11450
rect 9486 11398 9498 11450
rect 9498 11398 9528 11450
rect 9552 11398 9562 11450
rect 9562 11398 9608 11450
rect 9312 11396 9368 11398
rect 9392 11396 9448 11398
rect 9472 11396 9528 11398
rect 9552 11396 9608 11398
rect 10862 13082 10918 13084
rect 10942 13082 10998 13084
rect 11022 13082 11078 13084
rect 11102 13082 11158 13084
rect 10862 13030 10908 13082
rect 10908 13030 10918 13082
rect 10942 13030 10972 13082
rect 10972 13030 10984 13082
rect 10984 13030 10998 13082
rect 11022 13030 11036 13082
rect 11036 13030 11048 13082
rect 11048 13030 11078 13082
rect 11102 13030 11112 13082
rect 11112 13030 11158 13082
rect 10862 13028 10918 13030
rect 10942 13028 10998 13030
rect 11022 13028 11078 13030
rect 11102 13028 11158 13030
rect 12412 15802 12468 15804
rect 12492 15802 12548 15804
rect 12572 15802 12628 15804
rect 12652 15802 12708 15804
rect 12412 15750 12458 15802
rect 12458 15750 12468 15802
rect 12492 15750 12522 15802
rect 12522 15750 12534 15802
rect 12534 15750 12548 15802
rect 12572 15750 12586 15802
rect 12586 15750 12598 15802
rect 12598 15750 12628 15802
rect 12652 15750 12662 15802
rect 12662 15750 12708 15802
rect 12412 15748 12468 15750
rect 12492 15748 12548 15750
rect 12572 15748 12628 15750
rect 12652 15748 12708 15750
rect 12412 14714 12468 14716
rect 12492 14714 12548 14716
rect 12572 14714 12628 14716
rect 12652 14714 12708 14716
rect 12412 14662 12458 14714
rect 12458 14662 12468 14714
rect 12492 14662 12522 14714
rect 12522 14662 12534 14714
rect 12534 14662 12548 14714
rect 12572 14662 12586 14714
rect 12586 14662 12598 14714
rect 12598 14662 12628 14714
rect 12652 14662 12662 14714
rect 12662 14662 12708 14714
rect 12412 14660 12468 14662
rect 12492 14660 12548 14662
rect 12572 14660 12628 14662
rect 12652 14660 12708 14662
rect 10862 11994 10918 11996
rect 10942 11994 10998 11996
rect 11022 11994 11078 11996
rect 11102 11994 11158 11996
rect 10862 11942 10908 11994
rect 10908 11942 10918 11994
rect 10942 11942 10972 11994
rect 10972 11942 10984 11994
rect 10984 11942 10998 11994
rect 11022 11942 11036 11994
rect 11036 11942 11048 11994
rect 11048 11942 11078 11994
rect 11102 11942 11112 11994
rect 11112 11942 11158 11994
rect 10862 11940 10918 11942
rect 10942 11940 10998 11942
rect 11022 11940 11078 11942
rect 11102 11940 11158 11942
rect 10862 10906 10918 10908
rect 10942 10906 10998 10908
rect 11022 10906 11078 10908
rect 11102 10906 11158 10908
rect 10862 10854 10908 10906
rect 10908 10854 10918 10906
rect 10942 10854 10972 10906
rect 10972 10854 10984 10906
rect 10984 10854 10998 10906
rect 11022 10854 11036 10906
rect 11036 10854 11048 10906
rect 11048 10854 11078 10906
rect 11102 10854 11112 10906
rect 11112 10854 11158 10906
rect 10862 10852 10918 10854
rect 10942 10852 10998 10854
rect 11022 10852 11078 10854
rect 11102 10852 11158 10854
rect 9312 10362 9368 10364
rect 9392 10362 9448 10364
rect 9472 10362 9528 10364
rect 9552 10362 9608 10364
rect 9312 10310 9358 10362
rect 9358 10310 9368 10362
rect 9392 10310 9422 10362
rect 9422 10310 9434 10362
rect 9434 10310 9448 10362
rect 9472 10310 9486 10362
rect 9486 10310 9498 10362
rect 9498 10310 9528 10362
rect 9552 10310 9562 10362
rect 9562 10310 9608 10362
rect 9312 10308 9368 10310
rect 9392 10308 9448 10310
rect 9472 10308 9528 10310
rect 9552 10308 9608 10310
rect 7762 8730 7818 8732
rect 7842 8730 7898 8732
rect 7922 8730 7978 8732
rect 8002 8730 8058 8732
rect 7762 8678 7808 8730
rect 7808 8678 7818 8730
rect 7842 8678 7872 8730
rect 7872 8678 7884 8730
rect 7884 8678 7898 8730
rect 7922 8678 7936 8730
rect 7936 8678 7948 8730
rect 7948 8678 7978 8730
rect 8002 8678 8012 8730
rect 8012 8678 8058 8730
rect 7762 8676 7818 8678
rect 7842 8676 7898 8678
rect 7922 8676 7978 8678
rect 8002 8676 8058 8678
rect 7762 7642 7818 7644
rect 7842 7642 7898 7644
rect 7922 7642 7978 7644
rect 8002 7642 8058 7644
rect 7762 7590 7808 7642
rect 7808 7590 7818 7642
rect 7842 7590 7872 7642
rect 7872 7590 7884 7642
rect 7884 7590 7898 7642
rect 7922 7590 7936 7642
rect 7936 7590 7948 7642
rect 7948 7590 7978 7642
rect 8002 7590 8012 7642
rect 8012 7590 8058 7642
rect 7762 7588 7818 7590
rect 7842 7588 7898 7590
rect 7922 7588 7978 7590
rect 8002 7588 8058 7590
rect 9312 9274 9368 9276
rect 9392 9274 9448 9276
rect 9472 9274 9528 9276
rect 9552 9274 9608 9276
rect 9312 9222 9358 9274
rect 9358 9222 9368 9274
rect 9392 9222 9422 9274
rect 9422 9222 9434 9274
rect 9434 9222 9448 9274
rect 9472 9222 9486 9274
rect 9486 9222 9498 9274
rect 9498 9222 9528 9274
rect 9552 9222 9562 9274
rect 9562 9222 9608 9274
rect 9312 9220 9368 9222
rect 9392 9220 9448 9222
rect 9472 9220 9528 9222
rect 9552 9220 9608 9222
rect 10862 9818 10918 9820
rect 10942 9818 10998 9820
rect 11022 9818 11078 9820
rect 11102 9818 11158 9820
rect 10862 9766 10908 9818
rect 10908 9766 10918 9818
rect 10942 9766 10972 9818
rect 10972 9766 10984 9818
rect 10984 9766 10998 9818
rect 11022 9766 11036 9818
rect 11036 9766 11048 9818
rect 11048 9766 11078 9818
rect 11102 9766 11112 9818
rect 11112 9766 11158 9818
rect 10862 9764 10918 9766
rect 10942 9764 10998 9766
rect 11022 9764 11078 9766
rect 11102 9764 11158 9766
rect 9312 8186 9368 8188
rect 9392 8186 9448 8188
rect 9472 8186 9528 8188
rect 9552 8186 9608 8188
rect 9312 8134 9358 8186
rect 9358 8134 9368 8186
rect 9392 8134 9422 8186
rect 9422 8134 9434 8186
rect 9434 8134 9448 8186
rect 9472 8134 9486 8186
rect 9486 8134 9498 8186
rect 9498 8134 9528 8186
rect 9552 8134 9562 8186
rect 9562 8134 9608 8186
rect 9312 8132 9368 8134
rect 9392 8132 9448 8134
rect 9472 8132 9528 8134
rect 9552 8132 9608 8134
rect 7762 6554 7818 6556
rect 7842 6554 7898 6556
rect 7922 6554 7978 6556
rect 8002 6554 8058 6556
rect 7762 6502 7808 6554
rect 7808 6502 7818 6554
rect 7842 6502 7872 6554
rect 7872 6502 7884 6554
rect 7884 6502 7898 6554
rect 7922 6502 7936 6554
rect 7936 6502 7948 6554
rect 7948 6502 7978 6554
rect 8002 6502 8012 6554
rect 8012 6502 8058 6554
rect 7762 6500 7818 6502
rect 7842 6500 7898 6502
rect 7922 6500 7978 6502
rect 8002 6500 8058 6502
rect 6212 3834 6268 3836
rect 6292 3834 6348 3836
rect 6372 3834 6428 3836
rect 6452 3834 6508 3836
rect 6212 3782 6258 3834
rect 6258 3782 6268 3834
rect 6292 3782 6322 3834
rect 6322 3782 6334 3834
rect 6334 3782 6348 3834
rect 6372 3782 6386 3834
rect 6386 3782 6398 3834
rect 6398 3782 6428 3834
rect 6452 3782 6462 3834
rect 6462 3782 6508 3834
rect 6212 3780 6268 3782
rect 6292 3780 6348 3782
rect 6372 3780 6428 3782
rect 6452 3780 6508 3782
rect 6212 2746 6268 2748
rect 6292 2746 6348 2748
rect 6372 2746 6428 2748
rect 6452 2746 6508 2748
rect 6212 2694 6258 2746
rect 6258 2694 6268 2746
rect 6292 2694 6322 2746
rect 6322 2694 6334 2746
rect 6334 2694 6348 2746
rect 6372 2694 6386 2746
rect 6386 2694 6398 2746
rect 6398 2694 6428 2746
rect 6452 2694 6462 2746
rect 6462 2694 6508 2746
rect 6212 2692 6268 2694
rect 6292 2692 6348 2694
rect 6372 2692 6428 2694
rect 6452 2692 6508 2694
rect 7762 5466 7818 5468
rect 7842 5466 7898 5468
rect 7922 5466 7978 5468
rect 8002 5466 8058 5468
rect 7762 5414 7808 5466
rect 7808 5414 7818 5466
rect 7842 5414 7872 5466
rect 7872 5414 7884 5466
rect 7884 5414 7898 5466
rect 7922 5414 7936 5466
rect 7936 5414 7948 5466
rect 7948 5414 7978 5466
rect 8002 5414 8012 5466
rect 8012 5414 8058 5466
rect 7762 5412 7818 5414
rect 7842 5412 7898 5414
rect 7922 5412 7978 5414
rect 8002 5412 8058 5414
rect 7762 4378 7818 4380
rect 7842 4378 7898 4380
rect 7922 4378 7978 4380
rect 8002 4378 8058 4380
rect 7762 4326 7808 4378
rect 7808 4326 7818 4378
rect 7842 4326 7872 4378
rect 7872 4326 7884 4378
rect 7884 4326 7898 4378
rect 7922 4326 7936 4378
rect 7936 4326 7948 4378
rect 7948 4326 7978 4378
rect 8002 4326 8012 4378
rect 8012 4326 8058 4378
rect 7762 4324 7818 4326
rect 7842 4324 7898 4326
rect 7922 4324 7978 4326
rect 8002 4324 8058 4326
rect 7762 3290 7818 3292
rect 7842 3290 7898 3292
rect 7922 3290 7978 3292
rect 8002 3290 8058 3292
rect 7762 3238 7808 3290
rect 7808 3238 7818 3290
rect 7842 3238 7872 3290
rect 7872 3238 7884 3290
rect 7884 3238 7898 3290
rect 7922 3238 7936 3290
rect 7936 3238 7948 3290
rect 7948 3238 7978 3290
rect 8002 3238 8012 3290
rect 8012 3238 8058 3290
rect 7762 3236 7818 3238
rect 7842 3236 7898 3238
rect 7922 3236 7978 3238
rect 8002 3236 8058 3238
rect 7762 2202 7818 2204
rect 7842 2202 7898 2204
rect 7922 2202 7978 2204
rect 8002 2202 8058 2204
rect 7762 2150 7808 2202
rect 7808 2150 7818 2202
rect 7842 2150 7872 2202
rect 7872 2150 7884 2202
rect 7884 2150 7898 2202
rect 7922 2150 7936 2202
rect 7936 2150 7948 2202
rect 7948 2150 7978 2202
rect 8002 2150 8012 2202
rect 8012 2150 8058 2202
rect 7762 2148 7818 2150
rect 7842 2148 7898 2150
rect 7922 2148 7978 2150
rect 8002 2148 8058 2150
rect 9312 7098 9368 7100
rect 9392 7098 9448 7100
rect 9472 7098 9528 7100
rect 9552 7098 9608 7100
rect 9312 7046 9358 7098
rect 9358 7046 9368 7098
rect 9392 7046 9422 7098
rect 9422 7046 9434 7098
rect 9434 7046 9448 7098
rect 9472 7046 9486 7098
rect 9486 7046 9498 7098
rect 9498 7046 9528 7098
rect 9552 7046 9562 7098
rect 9562 7046 9608 7098
rect 9312 7044 9368 7046
rect 9392 7044 9448 7046
rect 9472 7044 9528 7046
rect 9552 7044 9608 7046
rect 9312 6010 9368 6012
rect 9392 6010 9448 6012
rect 9472 6010 9528 6012
rect 9552 6010 9608 6012
rect 9312 5958 9358 6010
rect 9358 5958 9368 6010
rect 9392 5958 9422 6010
rect 9422 5958 9434 6010
rect 9434 5958 9448 6010
rect 9472 5958 9486 6010
rect 9486 5958 9498 6010
rect 9498 5958 9528 6010
rect 9552 5958 9562 6010
rect 9562 5958 9608 6010
rect 9312 5956 9368 5958
rect 9392 5956 9448 5958
rect 9472 5956 9528 5958
rect 9552 5956 9608 5958
rect 6212 1658 6268 1660
rect 6292 1658 6348 1660
rect 6372 1658 6428 1660
rect 6452 1658 6508 1660
rect 6212 1606 6258 1658
rect 6258 1606 6268 1658
rect 6292 1606 6322 1658
rect 6322 1606 6334 1658
rect 6334 1606 6348 1658
rect 6372 1606 6386 1658
rect 6386 1606 6398 1658
rect 6398 1606 6428 1658
rect 6452 1606 6462 1658
rect 6462 1606 6508 1658
rect 6212 1604 6268 1606
rect 6292 1604 6348 1606
rect 6372 1604 6428 1606
rect 6452 1604 6508 1606
rect 9312 4922 9368 4924
rect 9392 4922 9448 4924
rect 9472 4922 9528 4924
rect 9552 4922 9608 4924
rect 9312 4870 9358 4922
rect 9358 4870 9368 4922
rect 9392 4870 9422 4922
rect 9422 4870 9434 4922
rect 9434 4870 9448 4922
rect 9472 4870 9486 4922
rect 9486 4870 9498 4922
rect 9498 4870 9528 4922
rect 9552 4870 9562 4922
rect 9562 4870 9608 4922
rect 9312 4868 9368 4870
rect 9392 4868 9448 4870
rect 9472 4868 9528 4870
rect 9552 4868 9608 4870
rect 10862 8730 10918 8732
rect 10942 8730 10998 8732
rect 11022 8730 11078 8732
rect 11102 8730 11158 8732
rect 10862 8678 10908 8730
rect 10908 8678 10918 8730
rect 10942 8678 10972 8730
rect 10972 8678 10984 8730
rect 10984 8678 10998 8730
rect 11022 8678 11036 8730
rect 11036 8678 11048 8730
rect 11048 8678 11078 8730
rect 11102 8678 11112 8730
rect 11112 8678 11158 8730
rect 10862 8676 10918 8678
rect 10942 8676 10998 8678
rect 11022 8676 11078 8678
rect 11102 8676 11158 8678
rect 10862 7642 10918 7644
rect 10942 7642 10998 7644
rect 11022 7642 11078 7644
rect 11102 7642 11158 7644
rect 10862 7590 10908 7642
rect 10908 7590 10918 7642
rect 10942 7590 10972 7642
rect 10972 7590 10984 7642
rect 10984 7590 10998 7642
rect 11022 7590 11036 7642
rect 11036 7590 11048 7642
rect 11048 7590 11078 7642
rect 11102 7590 11112 7642
rect 11112 7590 11158 7642
rect 10862 7588 10918 7590
rect 10942 7588 10998 7590
rect 11022 7588 11078 7590
rect 11102 7588 11158 7590
rect 12412 13626 12468 13628
rect 12492 13626 12548 13628
rect 12572 13626 12628 13628
rect 12652 13626 12708 13628
rect 12412 13574 12458 13626
rect 12458 13574 12468 13626
rect 12492 13574 12522 13626
rect 12522 13574 12534 13626
rect 12534 13574 12548 13626
rect 12572 13574 12586 13626
rect 12586 13574 12598 13626
rect 12598 13574 12628 13626
rect 12652 13574 12662 13626
rect 12662 13574 12708 13626
rect 12412 13572 12468 13574
rect 12492 13572 12548 13574
rect 12572 13572 12628 13574
rect 12652 13572 12708 13574
rect 12412 12538 12468 12540
rect 12492 12538 12548 12540
rect 12572 12538 12628 12540
rect 12652 12538 12708 12540
rect 12412 12486 12458 12538
rect 12458 12486 12468 12538
rect 12492 12486 12522 12538
rect 12522 12486 12534 12538
rect 12534 12486 12548 12538
rect 12572 12486 12586 12538
rect 12586 12486 12598 12538
rect 12598 12486 12628 12538
rect 12652 12486 12662 12538
rect 12662 12486 12708 12538
rect 12412 12484 12468 12486
rect 12492 12484 12548 12486
rect 12572 12484 12628 12486
rect 12652 12484 12708 12486
rect 13962 17434 14018 17436
rect 14042 17434 14098 17436
rect 14122 17434 14178 17436
rect 14202 17434 14258 17436
rect 13962 17382 14008 17434
rect 14008 17382 14018 17434
rect 14042 17382 14072 17434
rect 14072 17382 14084 17434
rect 14084 17382 14098 17434
rect 14122 17382 14136 17434
rect 14136 17382 14148 17434
rect 14148 17382 14178 17434
rect 14202 17382 14212 17434
rect 14212 17382 14258 17434
rect 13962 17380 14018 17382
rect 14042 17380 14098 17382
rect 14122 17380 14178 17382
rect 14202 17380 14258 17382
rect 13962 16346 14018 16348
rect 14042 16346 14098 16348
rect 14122 16346 14178 16348
rect 14202 16346 14258 16348
rect 13962 16294 14008 16346
rect 14008 16294 14018 16346
rect 14042 16294 14072 16346
rect 14072 16294 14084 16346
rect 14084 16294 14098 16346
rect 14122 16294 14136 16346
rect 14136 16294 14148 16346
rect 14148 16294 14178 16346
rect 14202 16294 14212 16346
rect 14212 16294 14258 16346
rect 13962 16292 14018 16294
rect 14042 16292 14098 16294
rect 14122 16292 14178 16294
rect 14202 16292 14258 16294
rect 13962 15258 14018 15260
rect 14042 15258 14098 15260
rect 14122 15258 14178 15260
rect 14202 15258 14258 15260
rect 13962 15206 14008 15258
rect 14008 15206 14018 15258
rect 14042 15206 14072 15258
rect 14072 15206 14084 15258
rect 14084 15206 14098 15258
rect 14122 15206 14136 15258
rect 14136 15206 14148 15258
rect 14148 15206 14178 15258
rect 14202 15206 14212 15258
rect 14212 15206 14258 15258
rect 13962 15204 14018 15206
rect 14042 15204 14098 15206
rect 14122 15204 14178 15206
rect 14202 15204 14258 15206
rect 12412 11450 12468 11452
rect 12492 11450 12548 11452
rect 12572 11450 12628 11452
rect 12652 11450 12708 11452
rect 12412 11398 12458 11450
rect 12458 11398 12468 11450
rect 12492 11398 12522 11450
rect 12522 11398 12534 11450
rect 12534 11398 12548 11450
rect 12572 11398 12586 11450
rect 12586 11398 12598 11450
rect 12598 11398 12628 11450
rect 12652 11398 12662 11450
rect 12662 11398 12708 11450
rect 12412 11396 12468 11398
rect 12492 11396 12548 11398
rect 12572 11396 12628 11398
rect 12652 11396 12708 11398
rect 12412 10362 12468 10364
rect 12492 10362 12548 10364
rect 12572 10362 12628 10364
rect 12652 10362 12708 10364
rect 12412 10310 12458 10362
rect 12458 10310 12468 10362
rect 12492 10310 12522 10362
rect 12522 10310 12534 10362
rect 12534 10310 12548 10362
rect 12572 10310 12586 10362
rect 12586 10310 12598 10362
rect 12598 10310 12628 10362
rect 12652 10310 12662 10362
rect 12662 10310 12708 10362
rect 12412 10308 12468 10310
rect 12492 10308 12548 10310
rect 12572 10308 12628 10310
rect 12652 10308 12708 10310
rect 10862 6554 10918 6556
rect 10942 6554 10998 6556
rect 11022 6554 11078 6556
rect 11102 6554 11158 6556
rect 10862 6502 10908 6554
rect 10908 6502 10918 6554
rect 10942 6502 10972 6554
rect 10972 6502 10984 6554
rect 10984 6502 10998 6554
rect 11022 6502 11036 6554
rect 11036 6502 11048 6554
rect 11048 6502 11078 6554
rect 11102 6502 11112 6554
rect 11112 6502 11158 6554
rect 10862 6500 10918 6502
rect 10942 6500 10998 6502
rect 11022 6500 11078 6502
rect 11102 6500 11158 6502
rect 12412 9274 12468 9276
rect 12492 9274 12548 9276
rect 12572 9274 12628 9276
rect 12652 9274 12708 9276
rect 12412 9222 12458 9274
rect 12458 9222 12468 9274
rect 12492 9222 12522 9274
rect 12522 9222 12534 9274
rect 12534 9222 12548 9274
rect 12572 9222 12586 9274
rect 12586 9222 12598 9274
rect 12598 9222 12628 9274
rect 12652 9222 12662 9274
rect 12662 9222 12708 9274
rect 12412 9220 12468 9222
rect 12492 9220 12548 9222
rect 12572 9220 12628 9222
rect 12652 9220 12708 9222
rect 10862 5466 10918 5468
rect 10942 5466 10998 5468
rect 11022 5466 11078 5468
rect 11102 5466 11158 5468
rect 10862 5414 10908 5466
rect 10908 5414 10918 5466
rect 10942 5414 10972 5466
rect 10972 5414 10984 5466
rect 10984 5414 10998 5466
rect 11022 5414 11036 5466
rect 11036 5414 11048 5466
rect 11048 5414 11078 5466
rect 11102 5414 11112 5466
rect 11112 5414 11158 5466
rect 10862 5412 10918 5414
rect 10942 5412 10998 5414
rect 11022 5412 11078 5414
rect 11102 5412 11158 5414
rect 9312 3834 9368 3836
rect 9392 3834 9448 3836
rect 9472 3834 9528 3836
rect 9552 3834 9608 3836
rect 9312 3782 9358 3834
rect 9358 3782 9368 3834
rect 9392 3782 9422 3834
rect 9422 3782 9434 3834
rect 9434 3782 9448 3834
rect 9472 3782 9486 3834
rect 9486 3782 9498 3834
rect 9498 3782 9528 3834
rect 9552 3782 9562 3834
rect 9562 3782 9608 3834
rect 9312 3780 9368 3782
rect 9392 3780 9448 3782
rect 9472 3780 9528 3782
rect 9552 3780 9608 3782
rect 9312 2746 9368 2748
rect 9392 2746 9448 2748
rect 9472 2746 9528 2748
rect 9552 2746 9608 2748
rect 9312 2694 9358 2746
rect 9358 2694 9368 2746
rect 9392 2694 9422 2746
rect 9422 2694 9434 2746
rect 9434 2694 9448 2746
rect 9472 2694 9486 2746
rect 9486 2694 9498 2746
rect 9498 2694 9528 2746
rect 9552 2694 9562 2746
rect 9562 2694 9608 2746
rect 9312 2692 9368 2694
rect 9392 2692 9448 2694
rect 9472 2692 9528 2694
rect 9552 2692 9608 2694
rect 12412 8186 12468 8188
rect 12492 8186 12548 8188
rect 12572 8186 12628 8188
rect 12652 8186 12708 8188
rect 12412 8134 12458 8186
rect 12458 8134 12468 8186
rect 12492 8134 12522 8186
rect 12522 8134 12534 8186
rect 12534 8134 12548 8186
rect 12572 8134 12586 8186
rect 12586 8134 12598 8186
rect 12598 8134 12628 8186
rect 12652 8134 12662 8186
rect 12662 8134 12708 8186
rect 12412 8132 12468 8134
rect 12492 8132 12548 8134
rect 12572 8132 12628 8134
rect 12652 8132 12708 8134
rect 12412 7098 12468 7100
rect 12492 7098 12548 7100
rect 12572 7098 12628 7100
rect 12652 7098 12708 7100
rect 12412 7046 12458 7098
rect 12458 7046 12468 7098
rect 12492 7046 12522 7098
rect 12522 7046 12534 7098
rect 12534 7046 12548 7098
rect 12572 7046 12586 7098
rect 12586 7046 12598 7098
rect 12598 7046 12628 7098
rect 12652 7046 12662 7098
rect 12662 7046 12708 7098
rect 12412 7044 12468 7046
rect 12492 7044 12548 7046
rect 12572 7044 12628 7046
rect 12652 7044 12708 7046
rect 13962 14170 14018 14172
rect 14042 14170 14098 14172
rect 14122 14170 14178 14172
rect 14202 14170 14258 14172
rect 13962 14118 14008 14170
rect 14008 14118 14018 14170
rect 14042 14118 14072 14170
rect 14072 14118 14084 14170
rect 14084 14118 14098 14170
rect 14122 14118 14136 14170
rect 14136 14118 14148 14170
rect 14148 14118 14178 14170
rect 14202 14118 14212 14170
rect 14212 14118 14258 14170
rect 13962 14116 14018 14118
rect 14042 14116 14098 14118
rect 14122 14116 14178 14118
rect 14202 14116 14258 14118
rect 13962 13082 14018 13084
rect 14042 13082 14098 13084
rect 14122 13082 14178 13084
rect 14202 13082 14258 13084
rect 13962 13030 14008 13082
rect 14008 13030 14018 13082
rect 14042 13030 14072 13082
rect 14072 13030 14084 13082
rect 14084 13030 14098 13082
rect 14122 13030 14136 13082
rect 14136 13030 14148 13082
rect 14148 13030 14178 13082
rect 14202 13030 14212 13082
rect 14212 13030 14258 13082
rect 13962 13028 14018 13030
rect 14042 13028 14098 13030
rect 14122 13028 14178 13030
rect 14202 13028 14258 13030
rect 13962 11994 14018 11996
rect 14042 11994 14098 11996
rect 14122 11994 14178 11996
rect 14202 11994 14258 11996
rect 13962 11942 14008 11994
rect 14008 11942 14018 11994
rect 14042 11942 14072 11994
rect 14072 11942 14084 11994
rect 14084 11942 14098 11994
rect 14122 11942 14136 11994
rect 14136 11942 14148 11994
rect 14148 11942 14178 11994
rect 14202 11942 14212 11994
rect 14212 11942 14258 11994
rect 13962 11940 14018 11942
rect 14042 11940 14098 11942
rect 14122 11940 14178 11942
rect 14202 11940 14258 11942
rect 13962 10906 14018 10908
rect 14042 10906 14098 10908
rect 14122 10906 14178 10908
rect 14202 10906 14258 10908
rect 13962 10854 14008 10906
rect 14008 10854 14018 10906
rect 14042 10854 14072 10906
rect 14072 10854 14084 10906
rect 14084 10854 14098 10906
rect 14122 10854 14136 10906
rect 14136 10854 14148 10906
rect 14148 10854 14178 10906
rect 14202 10854 14212 10906
rect 14212 10854 14258 10906
rect 13962 10852 14018 10854
rect 14042 10852 14098 10854
rect 14122 10852 14178 10854
rect 14202 10852 14258 10854
rect 12412 6010 12468 6012
rect 12492 6010 12548 6012
rect 12572 6010 12628 6012
rect 12652 6010 12708 6012
rect 12412 5958 12458 6010
rect 12458 5958 12468 6010
rect 12492 5958 12522 6010
rect 12522 5958 12534 6010
rect 12534 5958 12548 6010
rect 12572 5958 12586 6010
rect 12586 5958 12598 6010
rect 12598 5958 12628 6010
rect 12652 5958 12662 6010
rect 12662 5958 12708 6010
rect 12412 5956 12468 5958
rect 12492 5956 12548 5958
rect 12572 5956 12628 5958
rect 12652 5956 12708 5958
rect 10862 4378 10918 4380
rect 10942 4378 10998 4380
rect 11022 4378 11078 4380
rect 11102 4378 11158 4380
rect 10862 4326 10908 4378
rect 10908 4326 10918 4378
rect 10942 4326 10972 4378
rect 10972 4326 10984 4378
rect 10984 4326 10998 4378
rect 11022 4326 11036 4378
rect 11036 4326 11048 4378
rect 11048 4326 11078 4378
rect 11102 4326 11112 4378
rect 11112 4326 11158 4378
rect 10862 4324 10918 4326
rect 10942 4324 10998 4326
rect 11022 4324 11078 4326
rect 11102 4324 11158 4326
rect 10862 3290 10918 3292
rect 10942 3290 10998 3292
rect 11022 3290 11078 3292
rect 11102 3290 11158 3292
rect 10862 3238 10908 3290
rect 10908 3238 10918 3290
rect 10942 3238 10972 3290
rect 10972 3238 10984 3290
rect 10984 3238 10998 3290
rect 11022 3238 11036 3290
rect 11036 3238 11048 3290
rect 11048 3238 11078 3290
rect 11102 3238 11112 3290
rect 11112 3238 11158 3290
rect 10862 3236 10918 3238
rect 10942 3236 10998 3238
rect 11022 3236 11078 3238
rect 11102 3236 11158 3238
rect 12412 4922 12468 4924
rect 12492 4922 12548 4924
rect 12572 4922 12628 4924
rect 12652 4922 12708 4924
rect 12412 4870 12458 4922
rect 12458 4870 12468 4922
rect 12492 4870 12522 4922
rect 12522 4870 12534 4922
rect 12534 4870 12548 4922
rect 12572 4870 12586 4922
rect 12586 4870 12598 4922
rect 12598 4870 12628 4922
rect 12652 4870 12662 4922
rect 12662 4870 12708 4922
rect 12412 4868 12468 4870
rect 12492 4868 12548 4870
rect 12572 4868 12628 4870
rect 12652 4868 12708 4870
rect 12412 3834 12468 3836
rect 12492 3834 12548 3836
rect 12572 3834 12628 3836
rect 12652 3834 12708 3836
rect 12412 3782 12458 3834
rect 12458 3782 12468 3834
rect 12492 3782 12522 3834
rect 12522 3782 12534 3834
rect 12534 3782 12548 3834
rect 12572 3782 12586 3834
rect 12586 3782 12598 3834
rect 12598 3782 12628 3834
rect 12652 3782 12662 3834
rect 12662 3782 12708 3834
rect 12412 3780 12468 3782
rect 12492 3780 12548 3782
rect 12572 3780 12628 3782
rect 12652 3780 12708 3782
rect 9312 1658 9368 1660
rect 9392 1658 9448 1660
rect 9472 1658 9528 1660
rect 9552 1658 9608 1660
rect 9312 1606 9358 1658
rect 9358 1606 9368 1658
rect 9392 1606 9422 1658
rect 9422 1606 9434 1658
rect 9434 1606 9448 1658
rect 9472 1606 9486 1658
rect 9486 1606 9498 1658
rect 9498 1606 9528 1658
rect 9552 1606 9562 1658
rect 9562 1606 9608 1658
rect 9312 1604 9368 1606
rect 9392 1604 9448 1606
rect 9472 1604 9528 1606
rect 9552 1604 9608 1606
rect 10862 2202 10918 2204
rect 10942 2202 10998 2204
rect 11022 2202 11078 2204
rect 11102 2202 11158 2204
rect 10862 2150 10908 2202
rect 10908 2150 10918 2202
rect 10942 2150 10972 2202
rect 10972 2150 10984 2202
rect 10984 2150 10998 2202
rect 11022 2150 11036 2202
rect 11036 2150 11048 2202
rect 11048 2150 11078 2202
rect 11102 2150 11112 2202
rect 11112 2150 11158 2202
rect 10862 2148 10918 2150
rect 10942 2148 10998 2150
rect 11022 2148 11078 2150
rect 11102 2148 11158 2150
rect 12412 2746 12468 2748
rect 12492 2746 12548 2748
rect 12572 2746 12628 2748
rect 12652 2746 12708 2748
rect 12412 2694 12458 2746
rect 12458 2694 12468 2746
rect 12492 2694 12522 2746
rect 12522 2694 12534 2746
rect 12534 2694 12548 2746
rect 12572 2694 12586 2746
rect 12586 2694 12598 2746
rect 12598 2694 12628 2746
rect 12652 2694 12662 2746
rect 12662 2694 12708 2746
rect 12412 2692 12468 2694
rect 12492 2692 12548 2694
rect 12572 2692 12628 2694
rect 12652 2692 12708 2694
rect 13962 9818 14018 9820
rect 14042 9818 14098 9820
rect 14122 9818 14178 9820
rect 14202 9818 14258 9820
rect 13962 9766 14008 9818
rect 14008 9766 14018 9818
rect 14042 9766 14072 9818
rect 14072 9766 14084 9818
rect 14084 9766 14098 9818
rect 14122 9766 14136 9818
rect 14136 9766 14148 9818
rect 14148 9766 14178 9818
rect 14202 9766 14212 9818
rect 14212 9766 14258 9818
rect 13962 9764 14018 9766
rect 14042 9764 14098 9766
rect 14122 9764 14178 9766
rect 14202 9764 14258 9766
rect 13962 8730 14018 8732
rect 14042 8730 14098 8732
rect 14122 8730 14178 8732
rect 14202 8730 14258 8732
rect 13962 8678 14008 8730
rect 14008 8678 14018 8730
rect 14042 8678 14072 8730
rect 14072 8678 14084 8730
rect 14084 8678 14098 8730
rect 14122 8678 14136 8730
rect 14136 8678 14148 8730
rect 14148 8678 14178 8730
rect 14202 8678 14212 8730
rect 14212 8678 14258 8730
rect 13962 8676 14018 8678
rect 14042 8676 14098 8678
rect 14122 8676 14178 8678
rect 14202 8676 14258 8678
rect 18418 18536 18474 18592
rect 17062 18522 17118 18524
rect 17142 18522 17198 18524
rect 17222 18522 17278 18524
rect 17302 18522 17358 18524
rect 17062 18470 17108 18522
rect 17108 18470 17118 18522
rect 17142 18470 17172 18522
rect 17172 18470 17184 18522
rect 17184 18470 17198 18522
rect 17222 18470 17236 18522
rect 17236 18470 17248 18522
rect 17248 18470 17278 18522
rect 17302 18470 17312 18522
rect 17312 18470 17358 18522
rect 17062 18468 17118 18470
rect 17142 18468 17198 18470
rect 17222 18468 17278 18470
rect 17302 18468 17358 18470
rect 15512 17978 15568 17980
rect 15592 17978 15648 17980
rect 15672 17978 15728 17980
rect 15752 17978 15808 17980
rect 15512 17926 15558 17978
rect 15558 17926 15568 17978
rect 15592 17926 15622 17978
rect 15622 17926 15634 17978
rect 15634 17926 15648 17978
rect 15672 17926 15686 17978
rect 15686 17926 15698 17978
rect 15698 17926 15728 17978
rect 15752 17926 15762 17978
rect 15762 17926 15808 17978
rect 15512 17924 15568 17926
rect 15592 17924 15648 17926
rect 15672 17924 15728 17926
rect 15752 17924 15808 17926
rect 15512 16890 15568 16892
rect 15592 16890 15648 16892
rect 15672 16890 15728 16892
rect 15752 16890 15808 16892
rect 15512 16838 15558 16890
rect 15558 16838 15568 16890
rect 15592 16838 15622 16890
rect 15622 16838 15634 16890
rect 15634 16838 15648 16890
rect 15672 16838 15686 16890
rect 15686 16838 15698 16890
rect 15698 16838 15728 16890
rect 15752 16838 15762 16890
rect 15762 16838 15808 16890
rect 15512 16836 15568 16838
rect 15592 16836 15648 16838
rect 15672 16836 15728 16838
rect 15752 16836 15808 16838
rect 15512 15802 15568 15804
rect 15592 15802 15648 15804
rect 15672 15802 15728 15804
rect 15752 15802 15808 15804
rect 15512 15750 15558 15802
rect 15558 15750 15568 15802
rect 15592 15750 15622 15802
rect 15622 15750 15634 15802
rect 15634 15750 15648 15802
rect 15672 15750 15686 15802
rect 15686 15750 15698 15802
rect 15698 15750 15728 15802
rect 15752 15750 15762 15802
rect 15762 15750 15808 15802
rect 15512 15748 15568 15750
rect 15592 15748 15648 15750
rect 15672 15748 15728 15750
rect 15752 15748 15808 15750
rect 15512 14714 15568 14716
rect 15592 14714 15648 14716
rect 15672 14714 15728 14716
rect 15752 14714 15808 14716
rect 15512 14662 15558 14714
rect 15558 14662 15568 14714
rect 15592 14662 15622 14714
rect 15622 14662 15634 14714
rect 15634 14662 15648 14714
rect 15672 14662 15686 14714
rect 15686 14662 15698 14714
rect 15698 14662 15728 14714
rect 15752 14662 15762 14714
rect 15762 14662 15808 14714
rect 15512 14660 15568 14662
rect 15592 14660 15648 14662
rect 15672 14660 15728 14662
rect 15752 14660 15808 14662
rect 15512 13626 15568 13628
rect 15592 13626 15648 13628
rect 15672 13626 15728 13628
rect 15752 13626 15808 13628
rect 15512 13574 15558 13626
rect 15558 13574 15568 13626
rect 15592 13574 15622 13626
rect 15622 13574 15634 13626
rect 15634 13574 15648 13626
rect 15672 13574 15686 13626
rect 15686 13574 15698 13626
rect 15698 13574 15728 13626
rect 15752 13574 15762 13626
rect 15762 13574 15808 13626
rect 15512 13572 15568 13574
rect 15592 13572 15648 13574
rect 15672 13572 15728 13574
rect 15752 13572 15808 13574
rect 17062 17434 17118 17436
rect 17142 17434 17198 17436
rect 17222 17434 17278 17436
rect 17302 17434 17358 17436
rect 17062 17382 17108 17434
rect 17108 17382 17118 17434
rect 17142 17382 17172 17434
rect 17172 17382 17184 17434
rect 17184 17382 17198 17434
rect 17222 17382 17236 17434
rect 17236 17382 17248 17434
rect 17248 17382 17278 17434
rect 17302 17382 17312 17434
rect 17312 17382 17358 17434
rect 17062 17380 17118 17382
rect 17142 17380 17198 17382
rect 17222 17380 17278 17382
rect 17302 17380 17358 17382
rect 17062 16346 17118 16348
rect 17142 16346 17198 16348
rect 17222 16346 17278 16348
rect 17302 16346 17358 16348
rect 17062 16294 17108 16346
rect 17108 16294 17118 16346
rect 17142 16294 17172 16346
rect 17172 16294 17184 16346
rect 17184 16294 17198 16346
rect 17222 16294 17236 16346
rect 17236 16294 17248 16346
rect 17248 16294 17278 16346
rect 17302 16294 17312 16346
rect 17312 16294 17358 16346
rect 17062 16292 17118 16294
rect 17142 16292 17198 16294
rect 17222 16292 17278 16294
rect 17302 16292 17358 16294
rect 17062 15258 17118 15260
rect 17142 15258 17198 15260
rect 17222 15258 17278 15260
rect 17302 15258 17358 15260
rect 17062 15206 17108 15258
rect 17108 15206 17118 15258
rect 17142 15206 17172 15258
rect 17172 15206 17184 15258
rect 17184 15206 17198 15258
rect 17222 15206 17236 15258
rect 17236 15206 17248 15258
rect 17248 15206 17278 15258
rect 17302 15206 17312 15258
rect 17312 15206 17358 15258
rect 17062 15204 17118 15206
rect 17142 15204 17198 15206
rect 17222 15204 17278 15206
rect 17302 15204 17358 15206
rect 18418 16088 18474 16144
rect 17062 14170 17118 14172
rect 17142 14170 17198 14172
rect 17222 14170 17278 14172
rect 17302 14170 17358 14172
rect 17062 14118 17108 14170
rect 17108 14118 17118 14170
rect 17142 14118 17172 14170
rect 17172 14118 17184 14170
rect 17184 14118 17198 14170
rect 17222 14118 17236 14170
rect 17236 14118 17248 14170
rect 17248 14118 17278 14170
rect 17302 14118 17312 14170
rect 17312 14118 17358 14170
rect 17062 14116 17118 14118
rect 17142 14116 17198 14118
rect 17222 14116 17278 14118
rect 17302 14116 17358 14118
rect 17062 13082 17118 13084
rect 17142 13082 17198 13084
rect 17222 13082 17278 13084
rect 17302 13082 17358 13084
rect 17062 13030 17108 13082
rect 17108 13030 17118 13082
rect 17142 13030 17172 13082
rect 17172 13030 17184 13082
rect 17184 13030 17198 13082
rect 17222 13030 17236 13082
rect 17236 13030 17248 13082
rect 17248 13030 17278 13082
rect 17302 13030 17312 13082
rect 17312 13030 17358 13082
rect 17062 13028 17118 13030
rect 17142 13028 17198 13030
rect 17222 13028 17278 13030
rect 17302 13028 17358 13030
rect 15512 12538 15568 12540
rect 15592 12538 15648 12540
rect 15672 12538 15728 12540
rect 15752 12538 15808 12540
rect 15512 12486 15558 12538
rect 15558 12486 15568 12538
rect 15592 12486 15622 12538
rect 15622 12486 15634 12538
rect 15634 12486 15648 12538
rect 15672 12486 15686 12538
rect 15686 12486 15698 12538
rect 15698 12486 15728 12538
rect 15752 12486 15762 12538
rect 15762 12486 15808 12538
rect 15512 12484 15568 12486
rect 15592 12484 15648 12486
rect 15672 12484 15728 12486
rect 15752 12484 15808 12486
rect 15512 11450 15568 11452
rect 15592 11450 15648 11452
rect 15672 11450 15728 11452
rect 15752 11450 15808 11452
rect 15512 11398 15558 11450
rect 15558 11398 15568 11450
rect 15592 11398 15622 11450
rect 15622 11398 15634 11450
rect 15634 11398 15648 11450
rect 15672 11398 15686 11450
rect 15686 11398 15698 11450
rect 15698 11398 15728 11450
rect 15752 11398 15762 11450
rect 15762 11398 15808 11450
rect 15512 11396 15568 11398
rect 15592 11396 15648 11398
rect 15672 11396 15728 11398
rect 15752 11396 15808 11398
rect 13962 7642 14018 7644
rect 14042 7642 14098 7644
rect 14122 7642 14178 7644
rect 14202 7642 14258 7644
rect 13962 7590 14008 7642
rect 14008 7590 14018 7642
rect 14042 7590 14072 7642
rect 14072 7590 14084 7642
rect 14084 7590 14098 7642
rect 14122 7590 14136 7642
rect 14136 7590 14148 7642
rect 14148 7590 14178 7642
rect 14202 7590 14212 7642
rect 14212 7590 14258 7642
rect 13962 7588 14018 7590
rect 14042 7588 14098 7590
rect 14122 7588 14178 7590
rect 14202 7588 14258 7590
rect 15512 10362 15568 10364
rect 15592 10362 15648 10364
rect 15672 10362 15728 10364
rect 15752 10362 15808 10364
rect 15512 10310 15558 10362
rect 15558 10310 15568 10362
rect 15592 10310 15622 10362
rect 15622 10310 15634 10362
rect 15634 10310 15648 10362
rect 15672 10310 15686 10362
rect 15686 10310 15698 10362
rect 15698 10310 15728 10362
rect 15752 10310 15762 10362
rect 15762 10310 15808 10362
rect 15512 10308 15568 10310
rect 15592 10308 15648 10310
rect 15672 10308 15728 10310
rect 15752 10308 15808 10310
rect 13962 6554 14018 6556
rect 14042 6554 14098 6556
rect 14122 6554 14178 6556
rect 14202 6554 14258 6556
rect 13962 6502 14008 6554
rect 14008 6502 14018 6554
rect 14042 6502 14072 6554
rect 14072 6502 14084 6554
rect 14084 6502 14098 6554
rect 14122 6502 14136 6554
rect 14136 6502 14148 6554
rect 14148 6502 14178 6554
rect 14202 6502 14212 6554
rect 14212 6502 14258 6554
rect 13962 6500 14018 6502
rect 14042 6500 14098 6502
rect 14122 6500 14178 6502
rect 14202 6500 14258 6502
rect 13962 5466 14018 5468
rect 14042 5466 14098 5468
rect 14122 5466 14178 5468
rect 14202 5466 14258 5468
rect 13962 5414 14008 5466
rect 14008 5414 14018 5466
rect 14042 5414 14072 5466
rect 14072 5414 14084 5466
rect 14084 5414 14098 5466
rect 14122 5414 14136 5466
rect 14136 5414 14148 5466
rect 14148 5414 14178 5466
rect 14202 5414 14212 5466
rect 14212 5414 14258 5466
rect 13962 5412 14018 5414
rect 14042 5412 14098 5414
rect 14122 5412 14178 5414
rect 14202 5412 14258 5414
rect 13962 4378 14018 4380
rect 14042 4378 14098 4380
rect 14122 4378 14178 4380
rect 14202 4378 14258 4380
rect 13962 4326 14008 4378
rect 14008 4326 14018 4378
rect 14042 4326 14072 4378
rect 14072 4326 14084 4378
rect 14084 4326 14098 4378
rect 14122 4326 14136 4378
rect 14136 4326 14148 4378
rect 14148 4326 14178 4378
rect 14202 4326 14212 4378
rect 14212 4326 14258 4378
rect 13962 4324 14018 4326
rect 14042 4324 14098 4326
rect 14122 4324 14178 4326
rect 14202 4324 14258 4326
rect 13962 3290 14018 3292
rect 14042 3290 14098 3292
rect 14122 3290 14178 3292
rect 14202 3290 14258 3292
rect 13962 3238 14008 3290
rect 14008 3238 14018 3290
rect 14042 3238 14072 3290
rect 14072 3238 14084 3290
rect 14084 3238 14098 3290
rect 14122 3238 14136 3290
rect 14136 3238 14148 3290
rect 14148 3238 14178 3290
rect 14202 3238 14212 3290
rect 14212 3238 14258 3290
rect 13962 3236 14018 3238
rect 14042 3236 14098 3238
rect 14122 3236 14178 3238
rect 14202 3236 14258 3238
rect 12412 1658 12468 1660
rect 12492 1658 12548 1660
rect 12572 1658 12628 1660
rect 12652 1658 12708 1660
rect 12412 1606 12458 1658
rect 12458 1606 12468 1658
rect 12492 1606 12522 1658
rect 12522 1606 12534 1658
rect 12534 1606 12548 1658
rect 12572 1606 12586 1658
rect 12586 1606 12598 1658
rect 12598 1606 12628 1658
rect 12652 1606 12662 1658
rect 12662 1606 12708 1658
rect 12412 1604 12468 1606
rect 12492 1604 12548 1606
rect 12572 1604 12628 1606
rect 12652 1604 12708 1606
rect 13962 2202 14018 2204
rect 14042 2202 14098 2204
rect 14122 2202 14178 2204
rect 14202 2202 14258 2204
rect 13962 2150 14008 2202
rect 14008 2150 14018 2202
rect 14042 2150 14072 2202
rect 14072 2150 14084 2202
rect 14084 2150 14098 2202
rect 14122 2150 14136 2202
rect 14136 2150 14148 2202
rect 14148 2150 14178 2202
rect 14202 2150 14212 2202
rect 14212 2150 14258 2202
rect 13962 2148 14018 2150
rect 14042 2148 14098 2150
rect 14122 2148 14178 2150
rect 14202 2148 14258 2150
rect 15512 9274 15568 9276
rect 15592 9274 15648 9276
rect 15672 9274 15728 9276
rect 15752 9274 15808 9276
rect 15512 9222 15558 9274
rect 15558 9222 15568 9274
rect 15592 9222 15622 9274
rect 15622 9222 15634 9274
rect 15634 9222 15648 9274
rect 15672 9222 15686 9274
rect 15686 9222 15698 9274
rect 15698 9222 15728 9274
rect 15752 9222 15762 9274
rect 15762 9222 15808 9274
rect 15512 9220 15568 9222
rect 15592 9220 15648 9222
rect 15672 9220 15728 9222
rect 15752 9220 15808 9222
rect 15512 8186 15568 8188
rect 15592 8186 15648 8188
rect 15672 8186 15728 8188
rect 15752 8186 15808 8188
rect 15512 8134 15558 8186
rect 15558 8134 15568 8186
rect 15592 8134 15622 8186
rect 15622 8134 15634 8186
rect 15634 8134 15648 8186
rect 15672 8134 15686 8186
rect 15686 8134 15698 8186
rect 15698 8134 15728 8186
rect 15752 8134 15762 8186
rect 15762 8134 15808 8186
rect 15512 8132 15568 8134
rect 15592 8132 15648 8134
rect 15672 8132 15728 8134
rect 15752 8132 15808 8134
rect 17062 11994 17118 11996
rect 17142 11994 17198 11996
rect 17222 11994 17278 11996
rect 17302 11994 17358 11996
rect 17062 11942 17108 11994
rect 17108 11942 17118 11994
rect 17142 11942 17172 11994
rect 17172 11942 17184 11994
rect 17184 11942 17198 11994
rect 17222 11942 17236 11994
rect 17236 11942 17248 11994
rect 17248 11942 17278 11994
rect 17302 11942 17312 11994
rect 17312 11942 17358 11994
rect 17062 11940 17118 11942
rect 17142 11940 17198 11942
rect 17222 11940 17278 11942
rect 17302 11940 17358 11942
rect 15512 7098 15568 7100
rect 15592 7098 15648 7100
rect 15672 7098 15728 7100
rect 15752 7098 15808 7100
rect 15512 7046 15558 7098
rect 15558 7046 15568 7098
rect 15592 7046 15622 7098
rect 15622 7046 15634 7098
rect 15634 7046 15648 7098
rect 15672 7046 15686 7098
rect 15686 7046 15698 7098
rect 15698 7046 15728 7098
rect 15752 7046 15762 7098
rect 15762 7046 15808 7098
rect 15512 7044 15568 7046
rect 15592 7044 15648 7046
rect 15672 7044 15728 7046
rect 15752 7044 15808 7046
rect 15512 6010 15568 6012
rect 15592 6010 15648 6012
rect 15672 6010 15728 6012
rect 15752 6010 15808 6012
rect 15512 5958 15558 6010
rect 15558 5958 15568 6010
rect 15592 5958 15622 6010
rect 15622 5958 15634 6010
rect 15634 5958 15648 6010
rect 15672 5958 15686 6010
rect 15686 5958 15698 6010
rect 15698 5958 15728 6010
rect 15752 5958 15762 6010
rect 15762 5958 15808 6010
rect 15512 5956 15568 5958
rect 15592 5956 15648 5958
rect 15672 5956 15728 5958
rect 15752 5956 15808 5958
rect 15512 4922 15568 4924
rect 15592 4922 15648 4924
rect 15672 4922 15728 4924
rect 15752 4922 15808 4924
rect 15512 4870 15558 4922
rect 15558 4870 15568 4922
rect 15592 4870 15622 4922
rect 15622 4870 15634 4922
rect 15634 4870 15648 4922
rect 15672 4870 15686 4922
rect 15686 4870 15698 4922
rect 15698 4870 15728 4922
rect 15752 4870 15762 4922
rect 15762 4870 15808 4922
rect 15512 4868 15568 4870
rect 15592 4868 15648 4870
rect 15672 4868 15728 4870
rect 15752 4868 15808 4870
rect 15512 3834 15568 3836
rect 15592 3834 15648 3836
rect 15672 3834 15728 3836
rect 15752 3834 15808 3836
rect 15512 3782 15558 3834
rect 15558 3782 15568 3834
rect 15592 3782 15622 3834
rect 15622 3782 15634 3834
rect 15634 3782 15648 3834
rect 15672 3782 15686 3834
rect 15686 3782 15698 3834
rect 15698 3782 15728 3834
rect 15752 3782 15762 3834
rect 15762 3782 15808 3834
rect 15512 3780 15568 3782
rect 15592 3780 15648 3782
rect 15672 3780 15728 3782
rect 15752 3780 15808 3782
rect 17062 10906 17118 10908
rect 17142 10906 17198 10908
rect 17222 10906 17278 10908
rect 17302 10906 17358 10908
rect 17062 10854 17108 10906
rect 17108 10854 17118 10906
rect 17142 10854 17172 10906
rect 17172 10854 17184 10906
rect 17184 10854 17198 10906
rect 17222 10854 17236 10906
rect 17236 10854 17248 10906
rect 17248 10854 17278 10906
rect 17302 10854 17312 10906
rect 17312 10854 17358 10906
rect 17062 10852 17118 10854
rect 17142 10852 17198 10854
rect 17222 10852 17278 10854
rect 17302 10852 17358 10854
rect 17062 9818 17118 9820
rect 17142 9818 17198 9820
rect 17222 9818 17278 9820
rect 17302 9818 17358 9820
rect 17062 9766 17108 9818
rect 17108 9766 17118 9818
rect 17142 9766 17172 9818
rect 17172 9766 17184 9818
rect 17184 9766 17198 9818
rect 17222 9766 17236 9818
rect 17236 9766 17248 9818
rect 17248 9766 17278 9818
rect 17302 9766 17312 9818
rect 17312 9766 17358 9818
rect 17062 9764 17118 9766
rect 17142 9764 17198 9766
rect 17222 9764 17278 9766
rect 17302 9764 17358 9766
rect 17062 8730 17118 8732
rect 17142 8730 17198 8732
rect 17222 8730 17278 8732
rect 17302 8730 17358 8732
rect 17062 8678 17108 8730
rect 17108 8678 17118 8730
rect 17142 8678 17172 8730
rect 17172 8678 17184 8730
rect 17184 8678 17198 8730
rect 17222 8678 17236 8730
rect 17236 8678 17248 8730
rect 17248 8678 17278 8730
rect 17302 8678 17312 8730
rect 17312 8678 17358 8730
rect 17062 8676 17118 8678
rect 17142 8676 17198 8678
rect 17222 8676 17278 8678
rect 17302 8676 17358 8678
rect 18418 11212 18474 11248
rect 18418 11192 18420 11212
rect 18420 11192 18472 11212
rect 18472 11192 18474 11212
rect 18612 17978 18668 17980
rect 18692 17978 18748 17980
rect 18772 17978 18828 17980
rect 18852 17978 18908 17980
rect 18612 17926 18658 17978
rect 18658 17926 18668 17978
rect 18692 17926 18722 17978
rect 18722 17926 18734 17978
rect 18734 17926 18748 17978
rect 18772 17926 18786 17978
rect 18786 17926 18798 17978
rect 18798 17926 18828 17978
rect 18852 17926 18862 17978
rect 18862 17926 18908 17978
rect 18612 17924 18668 17926
rect 18692 17924 18748 17926
rect 18772 17924 18828 17926
rect 18852 17924 18908 17926
rect 18612 16890 18668 16892
rect 18692 16890 18748 16892
rect 18772 16890 18828 16892
rect 18852 16890 18908 16892
rect 18612 16838 18658 16890
rect 18658 16838 18668 16890
rect 18692 16838 18722 16890
rect 18722 16838 18734 16890
rect 18734 16838 18748 16890
rect 18772 16838 18786 16890
rect 18786 16838 18798 16890
rect 18798 16838 18828 16890
rect 18852 16838 18862 16890
rect 18862 16838 18908 16890
rect 18612 16836 18668 16838
rect 18692 16836 18748 16838
rect 18772 16836 18828 16838
rect 18852 16836 18908 16838
rect 18612 15802 18668 15804
rect 18692 15802 18748 15804
rect 18772 15802 18828 15804
rect 18852 15802 18908 15804
rect 18612 15750 18658 15802
rect 18658 15750 18668 15802
rect 18692 15750 18722 15802
rect 18722 15750 18734 15802
rect 18734 15750 18748 15802
rect 18772 15750 18786 15802
rect 18786 15750 18798 15802
rect 18798 15750 18828 15802
rect 18852 15750 18862 15802
rect 18862 15750 18908 15802
rect 18612 15748 18668 15750
rect 18692 15748 18748 15750
rect 18772 15748 18828 15750
rect 18852 15748 18908 15750
rect 18612 14714 18668 14716
rect 18692 14714 18748 14716
rect 18772 14714 18828 14716
rect 18852 14714 18908 14716
rect 18612 14662 18658 14714
rect 18658 14662 18668 14714
rect 18692 14662 18722 14714
rect 18722 14662 18734 14714
rect 18734 14662 18748 14714
rect 18772 14662 18786 14714
rect 18786 14662 18798 14714
rect 18798 14662 18828 14714
rect 18852 14662 18862 14714
rect 18862 14662 18908 14714
rect 18612 14660 18668 14662
rect 18692 14660 18748 14662
rect 18772 14660 18828 14662
rect 18852 14660 18908 14662
rect 19062 13640 19118 13696
rect 18612 13626 18668 13628
rect 18692 13626 18748 13628
rect 18772 13626 18828 13628
rect 18852 13626 18908 13628
rect 18612 13574 18658 13626
rect 18658 13574 18668 13626
rect 18692 13574 18722 13626
rect 18722 13574 18734 13626
rect 18734 13574 18748 13626
rect 18772 13574 18786 13626
rect 18786 13574 18798 13626
rect 18798 13574 18828 13626
rect 18852 13574 18862 13626
rect 18862 13574 18908 13626
rect 18612 13572 18668 13574
rect 18692 13572 18748 13574
rect 18772 13572 18828 13574
rect 18852 13572 18908 13574
rect 18612 12538 18668 12540
rect 18692 12538 18748 12540
rect 18772 12538 18828 12540
rect 18852 12538 18908 12540
rect 18612 12486 18658 12538
rect 18658 12486 18668 12538
rect 18692 12486 18722 12538
rect 18722 12486 18734 12538
rect 18734 12486 18748 12538
rect 18772 12486 18786 12538
rect 18786 12486 18798 12538
rect 18798 12486 18828 12538
rect 18852 12486 18862 12538
rect 18862 12486 18908 12538
rect 18612 12484 18668 12486
rect 18692 12484 18748 12486
rect 18772 12484 18828 12486
rect 18852 12484 18908 12486
rect 18612 11450 18668 11452
rect 18692 11450 18748 11452
rect 18772 11450 18828 11452
rect 18852 11450 18908 11452
rect 18612 11398 18658 11450
rect 18658 11398 18668 11450
rect 18692 11398 18722 11450
rect 18722 11398 18734 11450
rect 18734 11398 18748 11450
rect 18772 11398 18786 11450
rect 18786 11398 18798 11450
rect 18798 11398 18828 11450
rect 18852 11398 18862 11450
rect 18862 11398 18908 11450
rect 18612 11396 18668 11398
rect 18692 11396 18748 11398
rect 18772 11396 18828 11398
rect 18852 11396 18908 11398
rect 18612 10362 18668 10364
rect 18692 10362 18748 10364
rect 18772 10362 18828 10364
rect 18852 10362 18908 10364
rect 18612 10310 18658 10362
rect 18658 10310 18668 10362
rect 18692 10310 18722 10362
rect 18722 10310 18734 10362
rect 18734 10310 18748 10362
rect 18772 10310 18786 10362
rect 18786 10310 18798 10362
rect 18798 10310 18828 10362
rect 18852 10310 18862 10362
rect 18862 10310 18908 10362
rect 18612 10308 18668 10310
rect 18692 10308 18748 10310
rect 18772 10308 18828 10310
rect 18852 10308 18908 10310
rect 18612 9274 18668 9276
rect 18692 9274 18748 9276
rect 18772 9274 18828 9276
rect 18852 9274 18908 9276
rect 18612 9222 18658 9274
rect 18658 9222 18668 9274
rect 18692 9222 18722 9274
rect 18722 9222 18734 9274
rect 18734 9222 18748 9274
rect 18772 9222 18786 9274
rect 18786 9222 18798 9274
rect 18798 9222 18828 9274
rect 18852 9222 18862 9274
rect 18862 9222 18908 9274
rect 18612 9220 18668 9222
rect 18692 9220 18748 9222
rect 18772 9220 18828 9222
rect 18852 9220 18908 9222
rect 17958 8744 18014 8800
rect 17062 7642 17118 7644
rect 17142 7642 17198 7644
rect 17222 7642 17278 7644
rect 17302 7642 17358 7644
rect 17062 7590 17108 7642
rect 17108 7590 17118 7642
rect 17142 7590 17172 7642
rect 17172 7590 17184 7642
rect 17184 7590 17198 7642
rect 17222 7590 17236 7642
rect 17236 7590 17248 7642
rect 17248 7590 17278 7642
rect 17302 7590 17312 7642
rect 17312 7590 17358 7642
rect 17062 7588 17118 7590
rect 17142 7588 17198 7590
rect 17222 7588 17278 7590
rect 17302 7588 17358 7590
rect 17062 6554 17118 6556
rect 17142 6554 17198 6556
rect 17222 6554 17278 6556
rect 17302 6554 17358 6556
rect 17062 6502 17108 6554
rect 17108 6502 17118 6554
rect 17142 6502 17172 6554
rect 17172 6502 17184 6554
rect 17184 6502 17198 6554
rect 17222 6502 17236 6554
rect 17236 6502 17248 6554
rect 17248 6502 17278 6554
rect 17302 6502 17312 6554
rect 17312 6502 17358 6554
rect 17062 6500 17118 6502
rect 17142 6500 17198 6502
rect 17222 6500 17278 6502
rect 17302 6500 17358 6502
rect 15512 2746 15568 2748
rect 15592 2746 15648 2748
rect 15672 2746 15728 2748
rect 15752 2746 15808 2748
rect 15512 2694 15558 2746
rect 15558 2694 15568 2746
rect 15592 2694 15622 2746
rect 15622 2694 15634 2746
rect 15634 2694 15648 2746
rect 15672 2694 15686 2746
rect 15686 2694 15698 2746
rect 15698 2694 15728 2746
rect 15752 2694 15762 2746
rect 15762 2694 15808 2746
rect 15512 2692 15568 2694
rect 15592 2692 15648 2694
rect 15672 2692 15728 2694
rect 15752 2692 15808 2694
rect 15512 1658 15568 1660
rect 15592 1658 15648 1660
rect 15672 1658 15728 1660
rect 15752 1658 15808 1660
rect 15512 1606 15558 1658
rect 15558 1606 15568 1658
rect 15592 1606 15622 1658
rect 15622 1606 15634 1658
rect 15634 1606 15648 1658
rect 15672 1606 15686 1658
rect 15686 1606 15698 1658
rect 15698 1606 15728 1658
rect 15752 1606 15762 1658
rect 15762 1606 15808 1658
rect 15512 1604 15568 1606
rect 15592 1604 15648 1606
rect 15672 1604 15728 1606
rect 15752 1604 15808 1606
rect 17062 5466 17118 5468
rect 17142 5466 17198 5468
rect 17222 5466 17278 5468
rect 17302 5466 17358 5468
rect 17062 5414 17108 5466
rect 17108 5414 17118 5466
rect 17142 5414 17172 5466
rect 17172 5414 17184 5466
rect 17184 5414 17198 5466
rect 17222 5414 17236 5466
rect 17236 5414 17248 5466
rect 17248 5414 17278 5466
rect 17302 5414 17312 5466
rect 17312 5414 17358 5466
rect 17062 5412 17118 5414
rect 17142 5412 17198 5414
rect 17222 5412 17278 5414
rect 17302 5412 17358 5414
rect 17062 4378 17118 4380
rect 17142 4378 17198 4380
rect 17222 4378 17278 4380
rect 17302 4378 17358 4380
rect 17062 4326 17108 4378
rect 17108 4326 17118 4378
rect 17142 4326 17172 4378
rect 17172 4326 17184 4378
rect 17184 4326 17198 4378
rect 17222 4326 17236 4378
rect 17236 4326 17248 4378
rect 17248 4326 17278 4378
rect 17302 4326 17312 4378
rect 17312 4326 17358 4378
rect 17062 4324 17118 4326
rect 17142 4324 17198 4326
rect 17222 4324 17278 4326
rect 17302 4324 17358 4326
rect 17062 3290 17118 3292
rect 17142 3290 17198 3292
rect 17222 3290 17278 3292
rect 17302 3290 17358 3292
rect 17062 3238 17108 3290
rect 17108 3238 17118 3290
rect 17142 3238 17172 3290
rect 17172 3238 17184 3290
rect 17184 3238 17198 3290
rect 17222 3238 17236 3290
rect 17236 3238 17248 3290
rect 17248 3238 17278 3290
rect 17302 3238 17312 3290
rect 17312 3238 17358 3290
rect 17062 3236 17118 3238
rect 17142 3236 17198 3238
rect 17222 3236 17278 3238
rect 17302 3236 17358 3238
rect 17062 2202 17118 2204
rect 17142 2202 17198 2204
rect 17222 2202 17278 2204
rect 17302 2202 17358 2204
rect 17062 2150 17108 2202
rect 17108 2150 17118 2202
rect 17142 2150 17172 2202
rect 17172 2150 17184 2202
rect 17184 2150 17198 2202
rect 17222 2150 17236 2202
rect 17236 2150 17248 2202
rect 17248 2150 17278 2202
rect 17302 2150 17312 2202
rect 17312 2150 17358 2202
rect 17062 2148 17118 2150
rect 17142 2148 17198 2150
rect 17222 2148 17278 2150
rect 17302 2148 17358 2150
rect 18612 8186 18668 8188
rect 18692 8186 18748 8188
rect 18772 8186 18828 8188
rect 18852 8186 18908 8188
rect 18612 8134 18658 8186
rect 18658 8134 18668 8186
rect 18692 8134 18722 8186
rect 18722 8134 18734 8186
rect 18734 8134 18748 8186
rect 18772 8134 18786 8186
rect 18786 8134 18798 8186
rect 18798 8134 18828 8186
rect 18852 8134 18862 8186
rect 18862 8134 18908 8186
rect 18612 8132 18668 8134
rect 18692 8132 18748 8134
rect 18772 8132 18828 8134
rect 18852 8132 18908 8134
rect 18612 7098 18668 7100
rect 18692 7098 18748 7100
rect 18772 7098 18828 7100
rect 18852 7098 18908 7100
rect 18612 7046 18658 7098
rect 18658 7046 18668 7098
rect 18692 7046 18722 7098
rect 18722 7046 18734 7098
rect 18734 7046 18748 7098
rect 18772 7046 18786 7098
rect 18786 7046 18798 7098
rect 18798 7046 18828 7098
rect 18852 7046 18862 7098
rect 18862 7046 18908 7098
rect 18612 7044 18668 7046
rect 18692 7044 18748 7046
rect 18772 7044 18828 7046
rect 18852 7044 18908 7046
rect 18418 6296 18474 6352
rect 18612 6010 18668 6012
rect 18692 6010 18748 6012
rect 18772 6010 18828 6012
rect 18852 6010 18908 6012
rect 18612 5958 18658 6010
rect 18658 5958 18668 6010
rect 18692 5958 18722 6010
rect 18722 5958 18734 6010
rect 18734 5958 18748 6010
rect 18772 5958 18786 6010
rect 18786 5958 18798 6010
rect 18798 5958 18828 6010
rect 18852 5958 18862 6010
rect 18862 5958 18908 6010
rect 18612 5956 18668 5958
rect 18692 5956 18748 5958
rect 18772 5956 18828 5958
rect 18852 5956 18908 5958
rect 18612 4922 18668 4924
rect 18692 4922 18748 4924
rect 18772 4922 18828 4924
rect 18852 4922 18908 4924
rect 18612 4870 18658 4922
rect 18658 4870 18668 4922
rect 18692 4870 18722 4922
rect 18722 4870 18734 4922
rect 18734 4870 18748 4922
rect 18772 4870 18786 4922
rect 18786 4870 18798 4922
rect 18798 4870 18828 4922
rect 18852 4870 18862 4922
rect 18862 4870 18908 4922
rect 18612 4868 18668 4870
rect 18692 4868 18748 4870
rect 18772 4868 18828 4870
rect 18852 4868 18908 4870
rect 19062 3848 19118 3904
rect 18612 3834 18668 3836
rect 18692 3834 18748 3836
rect 18772 3834 18828 3836
rect 18852 3834 18908 3836
rect 18612 3782 18658 3834
rect 18658 3782 18668 3834
rect 18692 3782 18722 3834
rect 18722 3782 18734 3834
rect 18734 3782 18748 3834
rect 18772 3782 18786 3834
rect 18786 3782 18798 3834
rect 18798 3782 18828 3834
rect 18852 3782 18862 3834
rect 18862 3782 18908 3834
rect 18612 3780 18668 3782
rect 18692 3780 18748 3782
rect 18772 3780 18828 3782
rect 18852 3780 18908 3782
rect 18612 2746 18668 2748
rect 18692 2746 18748 2748
rect 18772 2746 18828 2748
rect 18852 2746 18908 2748
rect 18612 2694 18658 2746
rect 18658 2694 18668 2746
rect 18692 2694 18722 2746
rect 18722 2694 18734 2746
rect 18734 2694 18748 2746
rect 18772 2694 18786 2746
rect 18786 2694 18798 2746
rect 18798 2694 18828 2746
rect 18852 2694 18862 2746
rect 18862 2694 18908 2746
rect 18612 2692 18668 2694
rect 18692 2692 18748 2694
rect 18772 2692 18828 2694
rect 18852 2692 18908 2694
rect 18612 1658 18668 1660
rect 18692 1658 18748 1660
rect 18772 1658 18828 1660
rect 18852 1658 18908 1660
rect 18612 1606 18658 1658
rect 18658 1606 18668 1658
rect 18692 1606 18722 1658
rect 18722 1606 18734 1658
rect 18734 1606 18748 1658
rect 18772 1606 18786 1658
rect 18786 1606 18798 1658
rect 18798 1606 18828 1658
rect 18852 1606 18862 1658
rect 18862 1606 18908 1658
rect 18612 1604 18668 1606
rect 18692 1604 18748 1606
rect 18772 1604 18828 1606
rect 18852 1604 18908 1606
rect 18418 1400 18474 1456
rect 1562 1114 1618 1116
rect 1642 1114 1698 1116
rect 1722 1114 1778 1116
rect 1802 1114 1858 1116
rect 1562 1062 1608 1114
rect 1608 1062 1618 1114
rect 1642 1062 1672 1114
rect 1672 1062 1684 1114
rect 1684 1062 1698 1114
rect 1722 1062 1736 1114
rect 1736 1062 1748 1114
rect 1748 1062 1778 1114
rect 1802 1062 1812 1114
rect 1812 1062 1858 1114
rect 1562 1060 1618 1062
rect 1642 1060 1698 1062
rect 1722 1060 1778 1062
rect 1802 1060 1858 1062
rect 4662 1114 4718 1116
rect 4742 1114 4798 1116
rect 4822 1114 4878 1116
rect 4902 1114 4958 1116
rect 4662 1062 4708 1114
rect 4708 1062 4718 1114
rect 4742 1062 4772 1114
rect 4772 1062 4784 1114
rect 4784 1062 4798 1114
rect 4822 1062 4836 1114
rect 4836 1062 4848 1114
rect 4848 1062 4878 1114
rect 4902 1062 4912 1114
rect 4912 1062 4958 1114
rect 4662 1060 4718 1062
rect 4742 1060 4798 1062
rect 4822 1060 4878 1062
rect 4902 1060 4958 1062
rect 7762 1114 7818 1116
rect 7842 1114 7898 1116
rect 7922 1114 7978 1116
rect 8002 1114 8058 1116
rect 7762 1062 7808 1114
rect 7808 1062 7818 1114
rect 7842 1062 7872 1114
rect 7872 1062 7884 1114
rect 7884 1062 7898 1114
rect 7922 1062 7936 1114
rect 7936 1062 7948 1114
rect 7948 1062 7978 1114
rect 8002 1062 8012 1114
rect 8012 1062 8058 1114
rect 7762 1060 7818 1062
rect 7842 1060 7898 1062
rect 7922 1060 7978 1062
rect 8002 1060 8058 1062
rect 10862 1114 10918 1116
rect 10942 1114 10998 1116
rect 11022 1114 11078 1116
rect 11102 1114 11158 1116
rect 10862 1062 10908 1114
rect 10908 1062 10918 1114
rect 10942 1062 10972 1114
rect 10972 1062 10984 1114
rect 10984 1062 10998 1114
rect 11022 1062 11036 1114
rect 11036 1062 11048 1114
rect 11048 1062 11078 1114
rect 11102 1062 11112 1114
rect 11112 1062 11158 1114
rect 10862 1060 10918 1062
rect 10942 1060 10998 1062
rect 11022 1060 11078 1062
rect 11102 1060 11158 1062
rect 13962 1114 14018 1116
rect 14042 1114 14098 1116
rect 14122 1114 14178 1116
rect 14202 1114 14258 1116
rect 13962 1062 14008 1114
rect 14008 1062 14018 1114
rect 14042 1062 14072 1114
rect 14072 1062 14084 1114
rect 14084 1062 14098 1114
rect 14122 1062 14136 1114
rect 14136 1062 14148 1114
rect 14148 1062 14178 1114
rect 14202 1062 14212 1114
rect 14212 1062 14258 1114
rect 13962 1060 14018 1062
rect 14042 1060 14098 1062
rect 14122 1060 14178 1062
rect 14202 1060 14258 1062
rect 17062 1114 17118 1116
rect 17142 1114 17198 1116
rect 17222 1114 17278 1116
rect 17302 1114 17358 1116
rect 17062 1062 17108 1114
rect 17108 1062 17118 1114
rect 17142 1062 17172 1114
rect 17172 1062 17184 1114
rect 17184 1062 17198 1114
rect 17222 1062 17236 1114
rect 17236 1062 17248 1114
rect 17248 1062 17278 1114
rect 17302 1062 17312 1114
rect 17312 1062 17358 1114
rect 17062 1060 17118 1062
rect 17142 1060 17198 1062
rect 17222 1060 17278 1062
rect 17302 1060 17358 1062
rect 3112 570 3168 572
rect 3192 570 3248 572
rect 3272 570 3328 572
rect 3352 570 3408 572
rect 3112 518 3158 570
rect 3158 518 3168 570
rect 3192 518 3222 570
rect 3222 518 3234 570
rect 3234 518 3248 570
rect 3272 518 3286 570
rect 3286 518 3298 570
rect 3298 518 3328 570
rect 3352 518 3362 570
rect 3362 518 3408 570
rect 3112 516 3168 518
rect 3192 516 3248 518
rect 3272 516 3328 518
rect 3352 516 3408 518
rect 6212 570 6268 572
rect 6292 570 6348 572
rect 6372 570 6428 572
rect 6452 570 6508 572
rect 6212 518 6258 570
rect 6258 518 6268 570
rect 6292 518 6322 570
rect 6322 518 6334 570
rect 6334 518 6348 570
rect 6372 518 6386 570
rect 6386 518 6398 570
rect 6398 518 6428 570
rect 6452 518 6462 570
rect 6462 518 6508 570
rect 6212 516 6268 518
rect 6292 516 6348 518
rect 6372 516 6428 518
rect 6452 516 6508 518
rect 9312 570 9368 572
rect 9392 570 9448 572
rect 9472 570 9528 572
rect 9552 570 9608 572
rect 9312 518 9358 570
rect 9358 518 9368 570
rect 9392 518 9422 570
rect 9422 518 9434 570
rect 9434 518 9448 570
rect 9472 518 9486 570
rect 9486 518 9498 570
rect 9498 518 9528 570
rect 9552 518 9562 570
rect 9562 518 9608 570
rect 9312 516 9368 518
rect 9392 516 9448 518
rect 9472 516 9528 518
rect 9552 516 9608 518
rect 12412 570 12468 572
rect 12492 570 12548 572
rect 12572 570 12628 572
rect 12652 570 12708 572
rect 12412 518 12458 570
rect 12458 518 12468 570
rect 12492 518 12522 570
rect 12522 518 12534 570
rect 12534 518 12548 570
rect 12572 518 12586 570
rect 12586 518 12598 570
rect 12598 518 12628 570
rect 12652 518 12662 570
rect 12662 518 12708 570
rect 12412 516 12468 518
rect 12492 516 12548 518
rect 12572 516 12628 518
rect 12652 516 12708 518
rect 15512 570 15568 572
rect 15592 570 15648 572
rect 15672 570 15728 572
rect 15752 570 15808 572
rect 15512 518 15558 570
rect 15558 518 15568 570
rect 15592 518 15622 570
rect 15622 518 15634 570
rect 15634 518 15648 570
rect 15672 518 15686 570
rect 15686 518 15698 570
rect 15698 518 15728 570
rect 15752 518 15762 570
rect 15762 518 15808 570
rect 15512 516 15568 518
rect 15592 516 15648 518
rect 15672 516 15728 518
rect 15752 516 15808 518
rect 18612 570 18668 572
rect 18692 570 18748 572
rect 18772 570 18828 572
rect 18852 570 18908 572
rect 18612 518 18658 570
rect 18658 518 18668 570
rect 18692 518 18722 570
rect 18722 518 18734 570
rect 18734 518 18748 570
rect 18772 518 18786 570
rect 18786 518 18798 570
rect 18798 518 18828 570
rect 18852 518 18862 570
rect 18862 518 18908 570
rect 18612 516 18668 518
rect 18692 516 18748 518
rect 18772 516 18828 518
rect 18852 516 18908 518
<< metal3 >>
rect 18413 18594 18479 18597
rect 19200 18594 20000 18624
rect 18413 18592 20000 18594
rect 18413 18536 18418 18592
rect 18474 18536 20000 18592
rect 18413 18534 20000 18536
rect 18413 18531 18479 18534
rect 1552 18528 1868 18529
rect 1552 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1868 18528
rect 1552 18463 1868 18464
rect 4652 18528 4968 18529
rect 4652 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4968 18528
rect 4652 18463 4968 18464
rect 7752 18528 8068 18529
rect 7752 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8068 18528
rect 7752 18463 8068 18464
rect 10852 18528 11168 18529
rect 10852 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11168 18528
rect 10852 18463 11168 18464
rect 13952 18528 14268 18529
rect 13952 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14268 18528
rect 13952 18463 14268 18464
rect 17052 18528 17368 18529
rect 17052 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17368 18528
rect 19200 18504 20000 18534
rect 17052 18463 17368 18464
rect 3102 17984 3418 17985
rect 3102 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3418 17984
rect 3102 17919 3418 17920
rect 6202 17984 6518 17985
rect 6202 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6518 17984
rect 6202 17919 6518 17920
rect 9302 17984 9618 17985
rect 9302 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9618 17984
rect 9302 17919 9618 17920
rect 12402 17984 12718 17985
rect 12402 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12718 17984
rect 12402 17919 12718 17920
rect 15502 17984 15818 17985
rect 15502 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15818 17984
rect 15502 17919 15818 17920
rect 18602 17984 18918 17985
rect 18602 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18918 17984
rect 18602 17919 18918 17920
rect 1552 17440 1868 17441
rect 1552 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1868 17440
rect 1552 17375 1868 17376
rect 4652 17440 4968 17441
rect 4652 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4968 17440
rect 4652 17375 4968 17376
rect 7752 17440 8068 17441
rect 7752 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8068 17440
rect 7752 17375 8068 17376
rect 10852 17440 11168 17441
rect 10852 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11168 17440
rect 10852 17375 11168 17376
rect 13952 17440 14268 17441
rect 13952 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14268 17440
rect 13952 17375 14268 17376
rect 17052 17440 17368 17441
rect 17052 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17368 17440
rect 17052 17375 17368 17376
rect 3102 16896 3418 16897
rect 3102 16832 3108 16896
rect 3172 16832 3188 16896
rect 3252 16832 3268 16896
rect 3332 16832 3348 16896
rect 3412 16832 3418 16896
rect 3102 16831 3418 16832
rect 6202 16896 6518 16897
rect 6202 16832 6208 16896
rect 6272 16832 6288 16896
rect 6352 16832 6368 16896
rect 6432 16832 6448 16896
rect 6512 16832 6518 16896
rect 6202 16831 6518 16832
rect 9302 16896 9618 16897
rect 9302 16832 9308 16896
rect 9372 16832 9388 16896
rect 9452 16832 9468 16896
rect 9532 16832 9548 16896
rect 9612 16832 9618 16896
rect 9302 16831 9618 16832
rect 12402 16896 12718 16897
rect 12402 16832 12408 16896
rect 12472 16832 12488 16896
rect 12552 16832 12568 16896
rect 12632 16832 12648 16896
rect 12712 16832 12718 16896
rect 12402 16831 12718 16832
rect 15502 16896 15818 16897
rect 15502 16832 15508 16896
rect 15572 16832 15588 16896
rect 15652 16832 15668 16896
rect 15732 16832 15748 16896
rect 15812 16832 15818 16896
rect 15502 16831 15818 16832
rect 18602 16896 18918 16897
rect 18602 16832 18608 16896
rect 18672 16832 18688 16896
rect 18752 16832 18768 16896
rect 18832 16832 18848 16896
rect 18912 16832 18918 16896
rect 18602 16831 18918 16832
rect 1552 16352 1868 16353
rect 1552 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1868 16352
rect 1552 16287 1868 16288
rect 4652 16352 4968 16353
rect 4652 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4968 16352
rect 4652 16287 4968 16288
rect 7752 16352 8068 16353
rect 7752 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8068 16352
rect 7752 16287 8068 16288
rect 10852 16352 11168 16353
rect 10852 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11168 16352
rect 10852 16287 11168 16288
rect 13952 16352 14268 16353
rect 13952 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14268 16352
rect 13952 16287 14268 16288
rect 17052 16352 17368 16353
rect 17052 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17368 16352
rect 17052 16287 17368 16288
rect 18413 16146 18479 16149
rect 19200 16146 20000 16176
rect 18413 16144 20000 16146
rect 18413 16088 18418 16144
rect 18474 16088 20000 16144
rect 18413 16086 20000 16088
rect 18413 16083 18479 16086
rect 19200 16056 20000 16086
rect 3102 15808 3418 15809
rect 3102 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3418 15808
rect 3102 15743 3418 15744
rect 6202 15808 6518 15809
rect 6202 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6518 15808
rect 6202 15743 6518 15744
rect 9302 15808 9618 15809
rect 9302 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9618 15808
rect 9302 15743 9618 15744
rect 12402 15808 12718 15809
rect 12402 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12718 15808
rect 12402 15743 12718 15744
rect 15502 15808 15818 15809
rect 15502 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15818 15808
rect 15502 15743 15818 15744
rect 18602 15808 18918 15809
rect 18602 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18918 15808
rect 18602 15743 18918 15744
rect 1552 15264 1868 15265
rect 1552 15200 1558 15264
rect 1622 15200 1638 15264
rect 1702 15200 1718 15264
rect 1782 15200 1798 15264
rect 1862 15200 1868 15264
rect 1552 15199 1868 15200
rect 4652 15264 4968 15265
rect 4652 15200 4658 15264
rect 4722 15200 4738 15264
rect 4802 15200 4818 15264
rect 4882 15200 4898 15264
rect 4962 15200 4968 15264
rect 4652 15199 4968 15200
rect 7752 15264 8068 15265
rect 7752 15200 7758 15264
rect 7822 15200 7838 15264
rect 7902 15200 7918 15264
rect 7982 15200 7998 15264
rect 8062 15200 8068 15264
rect 7752 15199 8068 15200
rect 10852 15264 11168 15265
rect 10852 15200 10858 15264
rect 10922 15200 10938 15264
rect 11002 15200 11018 15264
rect 11082 15200 11098 15264
rect 11162 15200 11168 15264
rect 10852 15199 11168 15200
rect 13952 15264 14268 15265
rect 13952 15200 13958 15264
rect 14022 15200 14038 15264
rect 14102 15200 14118 15264
rect 14182 15200 14198 15264
rect 14262 15200 14268 15264
rect 13952 15199 14268 15200
rect 17052 15264 17368 15265
rect 17052 15200 17058 15264
rect 17122 15200 17138 15264
rect 17202 15200 17218 15264
rect 17282 15200 17298 15264
rect 17362 15200 17368 15264
rect 17052 15199 17368 15200
rect 3102 14720 3418 14721
rect 3102 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3418 14720
rect 3102 14655 3418 14656
rect 6202 14720 6518 14721
rect 6202 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6518 14720
rect 6202 14655 6518 14656
rect 9302 14720 9618 14721
rect 9302 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9618 14720
rect 9302 14655 9618 14656
rect 12402 14720 12718 14721
rect 12402 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12718 14720
rect 12402 14655 12718 14656
rect 15502 14720 15818 14721
rect 15502 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15818 14720
rect 15502 14655 15818 14656
rect 18602 14720 18918 14721
rect 18602 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18918 14720
rect 18602 14655 18918 14656
rect 1552 14176 1868 14177
rect 1552 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1868 14176
rect 1552 14111 1868 14112
rect 4652 14176 4968 14177
rect 4652 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4968 14176
rect 4652 14111 4968 14112
rect 7752 14176 8068 14177
rect 7752 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8068 14176
rect 7752 14111 8068 14112
rect 10852 14176 11168 14177
rect 10852 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11168 14176
rect 10852 14111 11168 14112
rect 13952 14176 14268 14177
rect 13952 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14268 14176
rect 13952 14111 14268 14112
rect 17052 14176 17368 14177
rect 17052 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17368 14176
rect 17052 14111 17368 14112
rect 19057 13698 19123 13701
rect 19200 13698 20000 13728
rect 19057 13696 20000 13698
rect 19057 13640 19062 13696
rect 19118 13640 20000 13696
rect 19057 13638 20000 13640
rect 19057 13635 19123 13638
rect 3102 13632 3418 13633
rect 3102 13568 3108 13632
rect 3172 13568 3188 13632
rect 3252 13568 3268 13632
rect 3332 13568 3348 13632
rect 3412 13568 3418 13632
rect 3102 13567 3418 13568
rect 6202 13632 6518 13633
rect 6202 13568 6208 13632
rect 6272 13568 6288 13632
rect 6352 13568 6368 13632
rect 6432 13568 6448 13632
rect 6512 13568 6518 13632
rect 6202 13567 6518 13568
rect 9302 13632 9618 13633
rect 9302 13568 9308 13632
rect 9372 13568 9388 13632
rect 9452 13568 9468 13632
rect 9532 13568 9548 13632
rect 9612 13568 9618 13632
rect 9302 13567 9618 13568
rect 12402 13632 12718 13633
rect 12402 13568 12408 13632
rect 12472 13568 12488 13632
rect 12552 13568 12568 13632
rect 12632 13568 12648 13632
rect 12712 13568 12718 13632
rect 12402 13567 12718 13568
rect 15502 13632 15818 13633
rect 15502 13568 15508 13632
rect 15572 13568 15588 13632
rect 15652 13568 15668 13632
rect 15732 13568 15748 13632
rect 15812 13568 15818 13632
rect 15502 13567 15818 13568
rect 18602 13632 18918 13633
rect 18602 13568 18608 13632
rect 18672 13568 18688 13632
rect 18752 13568 18768 13632
rect 18832 13568 18848 13632
rect 18912 13568 18918 13632
rect 19200 13608 20000 13638
rect 18602 13567 18918 13568
rect 1552 13088 1868 13089
rect 1552 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1868 13088
rect 1552 13023 1868 13024
rect 4652 13088 4968 13089
rect 4652 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4968 13088
rect 4652 13023 4968 13024
rect 7752 13088 8068 13089
rect 7752 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8068 13088
rect 7752 13023 8068 13024
rect 10852 13088 11168 13089
rect 10852 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11168 13088
rect 10852 13023 11168 13024
rect 13952 13088 14268 13089
rect 13952 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14268 13088
rect 13952 13023 14268 13024
rect 17052 13088 17368 13089
rect 17052 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17368 13088
rect 17052 13023 17368 13024
rect 3102 12544 3418 12545
rect 3102 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3418 12544
rect 3102 12479 3418 12480
rect 6202 12544 6518 12545
rect 6202 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6518 12544
rect 6202 12479 6518 12480
rect 9302 12544 9618 12545
rect 9302 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9618 12544
rect 9302 12479 9618 12480
rect 12402 12544 12718 12545
rect 12402 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12718 12544
rect 12402 12479 12718 12480
rect 15502 12544 15818 12545
rect 15502 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15818 12544
rect 15502 12479 15818 12480
rect 18602 12544 18918 12545
rect 18602 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18918 12544
rect 18602 12479 18918 12480
rect 1552 12000 1868 12001
rect 1552 11936 1558 12000
rect 1622 11936 1638 12000
rect 1702 11936 1718 12000
rect 1782 11936 1798 12000
rect 1862 11936 1868 12000
rect 1552 11935 1868 11936
rect 4652 12000 4968 12001
rect 4652 11936 4658 12000
rect 4722 11936 4738 12000
rect 4802 11936 4818 12000
rect 4882 11936 4898 12000
rect 4962 11936 4968 12000
rect 4652 11935 4968 11936
rect 7752 12000 8068 12001
rect 7752 11936 7758 12000
rect 7822 11936 7838 12000
rect 7902 11936 7918 12000
rect 7982 11936 7998 12000
rect 8062 11936 8068 12000
rect 7752 11935 8068 11936
rect 10852 12000 11168 12001
rect 10852 11936 10858 12000
rect 10922 11936 10938 12000
rect 11002 11936 11018 12000
rect 11082 11936 11098 12000
rect 11162 11936 11168 12000
rect 10852 11935 11168 11936
rect 13952 12000 14268 12001
rect 13952 11936 13958 12000
rect 14022 11936 14038 12000
rect 14102 11936 14118 12000
rect 14182 11936 14198 12000
rect 14262 11936 14268 12000
rect 13952 11935 14268 11936
rect 17052 12000 17368 12001
rect 17052 11936 17058 12000
rect 17122 11936 17138 12000
rect 17202 11936 17218 12000
rect 17282 11936 17298 12000
rect 17362 11936 17368 12000
rect 17052 11935 17368 11936
rect 3102 11456 3418 11457
rect 3102 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3418 11456
rect 3102 11391 3418 11392
rect 6202 11456 6518 11457
rect 6202 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6518 11456
rect 6202 11391 6518 11392
rect 9302 11456 9618 11457
rect 9302 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9618 11456
rect 9302 11391 9618 11392
rect 12402 11456 12718 11457
rect 12402 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12718 11456
rect 12402 11391 12718 11392
rect 15502 11456 15818 11457
rect 15502 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15818 11456
rect 15502 11391 15818 11392
rect 18602 11456 18918 11457
rect 18602 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18918 11456
rect 18602 11391 18918 11392
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 1552 10912 1868 10913
rect 1552 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1868 10912
rect 1552 10847 1868 10848
rect 4652 10912 4968 10913
rect 4652 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4968 10912
rect 4652 10847 4968 10848
rect 7752 10912 8068 10913
rect 7752 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8068 10912
rect 7752 10847 8068 10848
rect 10852 10912 11168 10913
rect 10852 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11168 10912
rect 10852 10847 11168 10848
rect 13952 10912 14268 10913
rect 13952 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14268 10912
rect 13952 10847 14268 10848
rect 17052 10912 17368 10913
rect 17052 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17368 10912
rect 17052 10847 17368 10848
rect 3102 10368 3418 10369
rect 3102 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3418 10368
rect 3102 10303 3418 10304
rect 6202 10368 6518 10369
rect 6202 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6518 10368
rect 6202 10303 6518 10304
rect 9302 10368 9618 10369
rect 9302 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9618 10368
rect 9302 10303 9618 10304
rect 12402 10368 12718 10369
rect 12402 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12718 10368
rect 12402 10303 12718 10304
rect 15502 10368 15818 10369
rect 15502 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15818 10368
rect 15502 10303 15818 10304
rect 18602 10368 18918 10369
rect 18602 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18918 10368
rect 18602 10303 18918 10304
rect 0 10026 800 10056
rect 933 10026 999 10029
rect 0 10024 999 10026
rect 0 9968 938 10024
rect 994 9968 999 10024
rect 0 9966 999 9968
rect 0 9936 800 9966
rect 933 9963 999 9966
rect 1552 9824 1868 9825
rect 1552 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1868 9824
rect 1552 9759 1868 9760
rect 4652 9824 4968 9825
rect 4652 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4968 9824
rect 4652 9759 4968 9760
rect 7752 9824 8068 9825
rect 7752 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8068 9824
rect 7752 9759 8068 9760
rect 10852 9824 11168 9825
rect 10852 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11168 9824
rect 10852 9759 11168 9760
rect 13952 9824 14268 9825
rect 13952 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14268 9824
rect 13952 9759 14268 9760
rect 17052 9824 17368 9825
rect 17052 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17368 9824
rect 17052 9759 17368 9760
rect 3102 9280 3418 9281
rect 3102 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3418 9280
rect 3102 9215 3418 9216
rect 6202 9280 6518 9281
rect 6202 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6518 9280
rect 6202 9215 6518 9216
rect 9302 9280 9618 9281
rect 9302 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9618 9280
rect 9302 9215 9618 9216
rect 12402 9280 12718 9281
rect 12402 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12718 9280
rect 12402 9215 12718 9216
rect 15502 9280 15818 9281
rect 15502 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15818 9280
rect 15502 9215 15818 9216
rect 18602 9280 18918 9281
rect 18602 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18918 9280
rect 18602 9215 18918 9216
rect 17953 8802 18019 8805
rect 19200 8802 20000 8832
rect 17953 8800 20000 8802
rect 17953 8744 17958 8800
rect 18014 8744 20000 8800
rect 17953 8742 20000 8744
rect 17953 8739 18019 8742
rect 1552 8736 1868 8737
rect 1552 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1868 8736
rect 1552 8671 1868 8672
rect 4652 8736 4968 8737
rect 4652 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4968 8736
rect 4652 8671 4968 8672
rect 7752 8736 8068 8737
rect 7752 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8068 8736
rect 7752 8671 8068 8672
rect 10852 8736 11168 8737
rect 10852 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11168 8736
rect 10852 8671 11168 8672
rect 13952 8736 14268 8737
rect 13952 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14268 8736
rect 13952 8671 14268 8672
rect 17052 8736 17368 8737
rect 17052 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17368 8736
rect 19200 8712 20000 8742
rect 17052 8671 17368 8672
rect 3102 8192 3418 8193
rect 3102 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3418 8192
rect 3102 8127 3418 8128
rect 6202 8192 6518 8193
rect 6202 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6518 8192
rect 6202 8127 6518 8128
rect 9302 8192 9618 8193
rect 9302 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9618 8192
rect 9302 8127 9618 8128
rect 12402 8192 12718 8193
rect 12402 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12718 8192
rect 12402 8127 12718 8128
rect 15502 8192 15818 8193
rect 15502 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15818 8192
rect 15502 8127 15818 8128
rect 18602 8192 18918 8193
rect 18602 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18918 8192
rect 18602 8127 18918 8128
rect 1552 7648 1868 7649
rect 1552 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1868 7648
rect 1552 7583 1868 7584
rect 4652 7648 4968 7649
rect 4652 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4968 7648
rect 4652 7583 4968 7584
rect 7752 7648 8068 7649
rect 7752 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8068 7648
rect 7752 7583 8068 7584
rect 10852 7648 11168 7649
rect 10852 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11168 7648
rect 10852 7583 11168 7584
rect 13952 7648 14268 7649
rect 13952 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14268 7648
rect 13952 7583 14268 7584
rect 17052 7648 17368 7649
rect 17052 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17368 7648
rect 17052 7583 17368 7584
rect 3102 7104 3418 7105
rect 3102 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3418 7104
rect 3102 7039 3418 7040
rect 6202 7104 6518 7105
rect 6202 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6518 7104
rect 6202 7039 6518 7040
rect 9302 7104 9618 7105
rect 9302 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9618 7104
rect 9302 7039 9618 7040
rect 12402 7104 12718 7105
rect 12402 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12718 7104
rect 12402 7039 12718 7040
rect 15502 7104 15818 7105
rect 15502 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15818 7104
rect 15502 7039 15818 7040
rect 18602 7104 18918 7105
rect 18602 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18918 7104
rect 18602 7039 18918 7040
rect 1552 6560 1868 6561
rect 1552 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1868 6560
rect 1552 6495 1868 6496
rect 4652 6560 4968 6561
rect 4652 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4968 6560
rect 4652 6495 4968 6496
rect 7752 6560 8068 6561
rect 7752 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8068 6560
rect 7752 6495 8068 6496
rect 10852 6560 11168 6561
rect 10852 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11168 6560
rect 10852 6495 11168 6496
rect 13952 6560 14268 6561
rect 13952 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14268 6560
rect 13952 6495 14268 6496
rect 17052 6560 17368 6561
rect 17052 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17368 6560
rect 17052 6495 17368 6496
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 3102 6016 3418 6017
rect 3102 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3418 6016
rect 3102 5951 3418 5952
rect 6202 6016 6518 6017
rect 6202 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6518 6016
rect 6202 5951 6518 5952
rect 9302 6016 9618 6017
rect 9302 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9618 6016
rect 9302 5951 9618 5952
rect 12402 6016 12718 6017
rect 12402 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12718 6016
rect 12402 5951 12718 5952
rect 15502 6016 15818 6017
rect 15502 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15818 6016
rect 15502 5951 15818 5952
rect 18602 6016 18918 6017
rect 18602 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18918 6016
rect 18602 5951 18918 5952
rect 1552 5472 1868 5473
rect 1552 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1868 5472
rect 1552 5407 1868 5408
rect 4652 5472 4968 5473
rect 4652 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4968 5472
rect 4652 5407 4968 5408
rect 7752 5472 8068 5473
rect 7752 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8068 5472
rect 7752 5407 8068 5408
rect 10852 5472 11168 5473
rect 10852 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11168 5472
rect 10852 5407 11168 5408
rect 13952 5472 14268 5473
rect 13952 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14268 5472
rect 13952 5407 14268 5408
rect 17052 5472 17368 5473
rect 17052 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17368 5472
rect 17052 5407 17368 5408
rect 3102 4928 3418 4929
rect 3102 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3418 4928
rect 3102 4863 3418 4864
rect 6202 4928 6518 4929
rect 6202 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6518 4928
rect 6202 4863 6518 4864
rect 9302 4928 9618 4929
rect 9302 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9618 4928
rect 9302 4863 9618 4864
rect 12402 4928 12718 4929
rect 12402 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12718 4928
rect 12402 4863 12718 4864
rect 15502 4928 15818 4929
rect 15502 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15818 4928
rect 15502 4863 15818 4864
rect 18602 4928 18918 4929
rect 18602 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18918 4928
rect 18602 4863 18918 4864
rect 1552 4384 1868 4385
rect 1552 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1868 4384
rect 1552 4319 1868 4320
rect 4652 4384 4968 4385
rect 4652 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4968 4384
rect 4652 4319 4968 4320
rect 7752 4384 8068 4385
rect 7752 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8068 4384
rect 7752 4319 8068 4320
rect 10852 4384 11168 4385
rect 10852 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11168 4384
rect 10852 4319 11168 4320
rect 13952 4384 14268 4385
rect 13952 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14268 4384
rect 13952 4319 14268 4320
rect 17052 4384 17368 4385
rect 17052 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17368 4384
rect 17052 4319 17368 4320
rect 19057 3906 19123 3909
rect 19200 3906 20000 3936
rect 19057 3904 20000 3906
rect 19057 3848 19062 3904
rect 19118 3848 20000 3904
rect 19057 3846 20000 3848
rect 19057 3843 19123 3846
rect 3102 3840 3418 3841
rect 3102 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3418 3840
rect 3102 3775 3418 3776
rect 6202 3840 6518 3841
rect 6202 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6518 3840
rect 6202 3775 6518 3776
rect 9302 3840 9618 3841
rect 9302 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9618 3840
rect 9302 3775 9618 3776
rect 12402 3840 12718 3841
rect 12402 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12718 3840
rect 12402 3775 12718 3776
rect 15502 3840 15818 3841
rect 15502 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15818 3840
rect 15502 3775 15818 3776
rect 18602 3840 18918 3841
rect 18602 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18918 3840
rect 19200 3816 20000 3846
rect 18602 3775 18918 3776
rect 1552 3296 1868 3297
rect 1552 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1868 3296
rect 1552 3231 1868 3232
rect 4652 3296 4968 3297
rect 4652 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4968 3296
rect 4652 3231 4968 3232
rect 7752 3296 8068 3297
rect 7752 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8068 3296
rect 7752 3231 8068 3232
rect 10852 3296 11168 3297
rect 10852 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11168 3296
rect 10852 3231 11168 3232
rect 13952 3296 14268 3297
rect 13952 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14268 3296
rect 13952 3231 14268 3232
rect 17052 3296 17368 3297
rect 17052 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17368 3296
rect 17052 3231 17368 3232
rect 3102 2752 3418 2753
rect 3102 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3418 2752
rect 3102 2687 3418 2688
rect 6202 2752 6518 2753
rect 6202 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6518 2752
rect 6202 2687 6518 2688
rect 9302 2752 9618 2753
rect 9302 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9618 2752
rect 9302 2687 9618 2688
rect 12402 2752 12718 2753
rect 12402 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12718 2752
rect 12402 2687 12718 2688
rect 15502 2752 15818 2753
rect 15502 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15818 2752
rect 15502 2687 15818 2688
rect 18602 2752 18918 2753
rect 18602 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18918 2752
rect 18602 2687 18918 2688
rect 1552 2208 1868 2209
rect 1552 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1868 2208
rect 1552 2143 1868 2144
rect 4652 2208 4968 2209
rect 4652 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4968 2208
rect 4652 2143 4968 2144
rect 7752 2208 8068 2209
rect 7752 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8068 2208
rect 7752 2143 8068 2144
rect 10852 2208 11168 2209
rect 10852 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11168 2208
rect 10852 2143 11168 2144
rect 13952 2208 14268 2209
rect 13952 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14268 2208
rect 13952 2143 14268 2144
rect 17052 2208 17368 2209
rect 17052 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17368 2208
rect 17052 2143 17368 2144
rect 3102 1664 3418 1665
rect 3102 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3418 1664
rect 3102 1599 3418 1600
rect 6202 1664 6518 1665
rect 6202 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6518 1664
rect 6202 1599 6518 1600
rect 9302 1664 9618 1665
rect 9302 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9618 1664
rect 9302 1599 9618 1600
rect 12402 1664 12718 1665
rect 12402 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12718 1664
rect 12402 1599 12718 1600
rect 15502 1664 15818 1665
rect 15502 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15818 1664
rect 15502 1599 15818 1600
rect 18602 1664 18918 1665
rect 18602 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18918 1664
rect 18602 1599 18918 1600
rect 18413 1458 18479 1461
rect 19200 1458 20000 1488
rect 18413 1456 20000 1458
rect 18413 1400 18418 1456
rect 18474 1400 20000 1456
rect 18413 1398 20000 1400
rect 18413 1395 18479 1398
rect 19200 1368 20000 1398
rect 1552 1120 1868 1121
rect 1552 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1868 1120
rect 1552 1055 1868 1056
rect 4652 1120 4968 1121
rect 4652 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4968 1120
rect 4652 1055 4968 1056
rect 7752 1120 8068 1121
rect 7752 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8068 1120
rect 7752 1055 8068 1056
rect 10852 1120 11168 1121
rect 10852 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11168 1120
rect 10852 1055 11168 1056
rect 13952 1120 14268 1121
rect 13952 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14268 1120
rect 13952 1055 14268 1056
rect 17052 1120 17368 1121
rect 17052 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17368 1120
rect 17052 1055 17368 1056
rect 3102 576 3418 577
rect 3102 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3418 576
rect 3102 511 3418 512
rect 6202 576 6518 577
rect 6202 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6518 576
rect 6202 511 6518 512
rect 9302 576 9618 577
rect 9302 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9618 576
rect 9302 511 9618 512
rect 12402 576 12718 577
rect 12402 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12718 576
rect 12402 511 12718 512
rect 15502 576 15818 577
rect 15502 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15818 576
rect 15502 511 15818 512
rect 18602 576 18918 577
rect 18602 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18918 576
rect 18602 511 18918 512
<< via3 >>
rect 1558 18524 1622 18528
rect 1558 18468 1562 18524
rect 1562 18468 1618 18524
rect 1618 18468 1622 18524
rect 1558 18464 1622 18468
rect 1638 18524 1702 18528
rect 1638 18468 1642 18524
rect 1642 18468 1698 18524
rect 1698 18468 1702 18524
rect 1638 18464 1702 18468
rect 1718 18524 1782 18528
rect 1718 18468 1722 18524
rect 1722 18468 1778 18524
rect 1778 18468 1782 18524
rect 1718 18464 1782 18468
rect 1798 18524 1862 18528
rect 1798 18468 1802 18524
rect 1802 18468 1858 18524
rect 1858 18468 1862 18524
rect 1798 18464 1862 18468
rect 4658 18524 4722 18528
rect 4658 18468 4662 18524
rect 4662 18468 4718 18524
rect 4718 18468 4722 18524
rect 4658 18464 4722 18468
rect 4738 18524 4802 18528
rect 4738 18468 4742 18524
rect 4742 18468 4798 18524
rect 4798 18468 4802 18524
rect 4738 18464 4802 18468
rect 4818 18524 4882 18528
rect 4818 18468 4822 18524
rect 4822 18468 4878 18524
rect 4878 18468 4882 18524
rect 4818 18464 4882 18468
rect 4898 18524 4962 18528
rect 4898 18468 4902 18524
rect 4902 18468 4958 18524
rect 4958 18468 4962 18524
rect 4898 18464 4962 18468
rect 7758 18524 7822 18528
rect 7758 18468 7762 18524
rect 7762 18468 7818 18524
rect 7818 18468 7822 18524
rect 7758 18464 7822 18468
rect 7838 18524 7902 18528
rect 7838 18468 7842 18524
rect 7842 18468 7898 18524
rect 7898 18468 7902 18524
rect 7838 18464 7902 18468
rect 7918 18524 7982 18528
rect 7918 18468 7922 18524
rect 7922 18468 7978 18524
rect 7978 18468 7982 18524
rect 7918 18464 7982 18468
rect 7998 18524 8062 18528
rect 7998 18468 8002 18524
rect 8002 18468 8058 18524
rect 8058 18468 8062 18524
rect 7998 18464 8062 18468
rect 10858 18524 10922 18528
rect 10858 18468 10862 18524
rect 10862 18468 10918 18524
rect 10918 18468 10922 18524
rect 10858 18464 10922 18468
rect 10938 18524 11002 18528
rect 10938 18468 10942 18524
rect 10942 18468 10998 18524
rect 10998 18468 11002 18524
rect 10938 18464 11002 18468
rect 11018 18524 11082 18528
rect 11018 18468 11022 18524
rect 11022 18468 11078 18524
rect 11078 18468 11082 18524
rect 11018 18464 11082 18468
rect 11098 18524 11162 18528
rect 11098 18468 11102 18524
rect 11102 18468 11158 18524
rect 11158 18468 11162 18524
rect 11098 18464 11162 18468
rect 13958 18524 14022 18528
rect 13958 18468 13962 18524
rect 13962 18468 14018 18524
rect 14018 18468 14022 18524
rect 13958 18464 14022 18468
rect 14038 18524 14102 18528
rect 14038 18468 14042 18524
rect 14042 18468 14098 18524
rect 14098 18468 14102 18524
rect 14038 18464 14102 18468
rect 14118 18524 14182 18528
rect 14118 18468 14122 18524
rect 14122 18468 14178 18524
rect 14178 18468 14182 18524
rect 14118 18464 14182 18468
rect 14198 18524 14262 18528
rect 14198 18468 14202 18524
rect 14202 18468 14258 18524
rect 14258 18468 14262 18524
rect 14198 18464 14262 18468
rect 17058 18524 17122 18528
rect 17058 18468 17062 18524
rect 17062 18468 17118 18524
rect 17118 18468 17122 18524
rect 17058 18464 17122 18468
rect 17138 18524 17202 18528
rect 17138 18468 17142 18524
rect 17142 18468 17198 18524
rect 17198 18468 17202 18524
rect 17138 18464 17202 18468
rect 17218 18524 17282 18528
rect 17218 18468 17222 18524
rect 17222 18468 17278 18524
rect 17278 18468 17282 18524
rect 17218 18464 17282 18468
rect 17298 18524 17362 18528
rect 17298 18468 17302 18524
rect 17302 18468 17358 18524
rect 17358 18468 17362 18524
rect 17298 18464 17362 18468
rect 3108 17980 3172 17984
rect 3108 17924 3112 17980
rect 3112 17924 3168 17980
rect 3168 17924 3172 17980
rect 3108 17920 3172 17924
rect 3188 17980 3252 17984
rect 3188 17924 3192 17980
rect 3192 17924 3248 17980
rect 3248 17924 3252 17980
rect 3188 17920 3252 17924
rect 3268 17980 3332 17984
rect 3268 17924 3272 17980
rect 3272 17924 3328 17980
rect 3328 17924 3332 17980
rect 3268 17920 3332 17924
rect 3348 17980 3412 17984
rect 3348 17924 3352 17980
rect 3352 17924 3408 17980
rect 3408 17924 3412 17980
rect 3348 17920 3412 17924
rect 6208 17980 6272 17984
rect 6208 17924 6212 17980
rect 6212 17924 6268 17980
rect 6268 17924 6272 17980
rect 6208 17920 6272 17924
rect 6288 17980 6352 17984
rect 6288 17924 6292 17980
rect 6292 17924 6348 17980
rect 6348 17924 6352 17980
rect 6288 17920 6352 17924
rect 6368 17980 6432 17984
rect 6368 17924 6372 17980
rect 6372 17924 6428 17980
rect 6428 17924 6432 17980
rect 6368 17920 6432 17924
rect 6448 17980 6512 17984
rect 6448 17924 6452 17980
rect 6452 17924 6508 17980
rect 6508 17924 6512 17980
rect 6448 17920 6512 17924
rect 9308 17980 9372 17984
rect 9308 17924 9312 17980
rect 9312 17924 9368 17980
rect 9368 17924 9372 17980
rect 9308 17920 9372 17924
rect 9388 17980 9452 17984
rect 9388 17924 9392 17980
rect 9392 17924 9448 17980
rect 9448 17924 9452 17980
rect 9388 17920 9452 17924
rect 9468 17980 9532 17984
rect 9468 17924 9472 17980
rect 9472 17924 9528 17980
rect 9528 17924 9532 17980
rect 9468 17920 9532 17924
rect 9548 17980 9612 17984
rect 9548 17924 9552 17980
rect 9552 17924 9608 17980
rect 9608 17924 9612 17980
rect 9548 17920 9612 17924
rect 12408 17980 12472 17984
rect 12408 17924 12412 17980
rect 12412 17924 12468 17980
rect 12468 17924 12472 17980
rect 12408 17920 12472 17924
rect 12488 17980 12552 17984
rect 12488 17924 12492 17980
rect 12492 17924 12548 17980
rect 12548 17924 12552 17980
rect 12488 17920 12552 17924
rect 12568 17980 12632 17984
rect 12568 17924 12572 17980
rect 12572 17924 12628 17980
rect 12628 17924 12632 17980
rect 12568 17920 12632 17924
rect 12648 17980 12712 17984
rect 12648 17924 12652 17980
rect 12652 17924 12708 17980
rect 12708 17924 12712 17980
rect 12648 17920 12712 17924
rect 15508 17980 15572 17984
rect 15508 17924 15512 17980
rect 15512 17924 15568 17980
rect 15568 17924 15572 17980
rect 15508 17920 15572 17924
rect 15588 17980 15652 17984
rect 15588 17924 15592 17980
rect 15592 17924 15648 17980
rect 15648 17924 15652 17980
rect 15588 17920 15652 17924
rect 15668 17980 15732 17984
rect 15668 17924 15672 17980
rect 15672 17924 15728 17980
rect 15728 17924 15732 17980
rect 15668 17920 15732 17924
rect 15748 17980 15812 17984
rect 15748 17924 15752 17980
rect 15752 17924 15808 17980
rect 15808 17924 15812 17980
rect 15748 17920 15812 17924
rect 18608 17980 18672 17984
rect 18608 17924 18612 17980
rect 18612 17924 18668 17980
rect 18668 17924 18672 17980
rect 18608 17920 18672 17924
rect 18688 17980 18752 17984
rect 18688 17924 18692 17980
rect 18692 17924 18748 17980
rect 18748 17924 18752 17980
rect 18688 17920 18752 17924
rect 18768 17980 18832 17984
rect 18768 17924 18772 17980
rect 18772 17924 18828 17980
rect 18828 17924 18832 17980
rect 18768 17920 18832 17924
rect 18848 17980 18912 17984
rect 18848 17924 18852 17980
rect 18852 17924 18908 17980
rect 18908 17924 18912 17980
rect 18848 17920 18912 17924
rect 1558 17436 1622 17440
rect 1558 17380 1562 17436
rect 1562 17380 1618 17436
rect 1618 17380 1622 17436
rect 1558 17376 1622 17380
rect 1638 17436 1702 17440
rect 1638 17380 1642 17436
rect 1642 17380 1698 17436
rect 1698 17380 1702 17436
rect 1638 17376 1702 17380
rect 1718 17436 1782 17440
rect 1718 17380 1722 17436
rect 1722 17380 1778 17436
rect 1778 17380 1782 17436
rect 1718 17376 1782 17380
rect 1798 17436 1862 17440
rect 1798 17380 1802 17436
rect 1802 17380 1858 17436
rect 1858 17380 1862 17436
rect 1798 17376 1862 17380
rect 4658 17436 4722 17440
rect 4658 17380 4662 17436
rect 4662 17380 4718 17436
rect 4718 17380 4722 17436
rect 4658 17376 4722 17380
rect 4738 17436 4802 17440
rect 4738 17380 4742 17436
rect 4742 17380 4798 17436
rect 4798 17380 4802 17436
rect 4738 17376 4802 17380
rect 4818 17436 4882 17440
rect 4818 17380 4822 17436
rect 4822 17380 4878 17436
rect 4878 17380 4882 17436
rect 4818 17376 4882 17380
rect 4898 17436 4962 17440
rect 4898 17380 4902 17436
rect 4902 17380 4958 17436
rect 4958 17380 4962 17436
rect 4898 17376 4962 17380
rect 7758 17436 7822 17440
rect 7758 17380 7762 17436
rect 7762 17380 7818 17436
rect 7818 17380 7822 17436
rect 7758 17376 7822 17380
rect 7838 17436 7902 17440
rect 7838 17380 7842 17436
rect 7842 17380 7898 17436
rect 7898 17380 7902 17436
rect 7838 17376 7902 17380
rect 7918 17436 7982 17440
rect 7918 17380 7922 17436
rect 7922 17380 7978 17436
rect 7978 17380 7982 17436
rect 7918 17376 7982 17380
rect 7998 17436 8062 17440
rect 7998 17380 8002 17436
rect 8002 17380 8058 17436
rect 8058 17380 8062 17436
rect 7998 17376 8062 17380
rect 10858 17436 10922 17440
rect 10858 17380 10862 17436
rect 10862 17380 10918 17436
rect 10918 17380 10922 17436
rect 10858 17376 10922 17380
rect 10938 17436 11002 17440
rect 10938 17380 10942 17436
rect 10942 17380 10998 17436
rect 10998 17380 11002 17436
rect 10938 17376 11002 17380
rect 11018 17436 11082 17440
rect 11018 17380 11022 17436
rect 11022 17380 11078 17436
rect 11078 17380 11082 17436
rect 11018 17376 11082 17380
rect 11098 17436 11162 17440
rect 11098 17380 11102 17436
rect 11102 17380 11158 17436
rect 11158 17380 11162 17436
rect 11098 17376 11162 17380
rect 13958 17436 14022 17440
rect 13958 17380 13962 17436
rect 13962 17380 14018 17436
rect 14018 17380 14022 17436
rect 13958 17376 14022 17380
rect 14038 17436 14102 17440
rect 14038 17380 14042 17436
rect 14042 17380 14098 17436
rect 14098 17380 14102 17436
rect 14038 17376 14102 17380
rect 14118 17436 14182 17440
rect 14118 17380 14122 17436
rect 14122 17380 14178 17436
rect 14178 17380 14182 17436
rect 14118 17376 14182 17380
rect 14198 17436 14262 17440
rect 14198 17380 14202 17436
rect 14202 17380 14258 17436
rect 14258 17380 14262 17436
rect 14198 17376 14262 17380
rect 17058 17436 17122 17440
rect 17058 17380 17062 17436
rect 17062 17380 17118 17436
rect 17118 17380 17122 17436
rect 17058 17376 17122 17380
rect 17138 17436 17202 17440
rect 17138 17380 17142 17436
rect 17142 17380 17198 17436
rect 17198 17380 17202 17436
rect 17138 17376 17202 17380
rect 17218 17436 17282 17440
rect 17218 17380 17222 17436
rect 17222 17380 17278 17436
rect 17278 17380 17282 17436
rect 17218 17376 17282 17380
rect 17298 17436 17362 17440
rect 17298 17380 17302 17436
rect 17302 17380 17358 17436
rect 17358 17380 17362 17436
rect 17298 17376 17362 17380
rect 3108 16892 3172 16896
rect 3108 16836 3112 16892
rect 3112 16836 3168 16892
rect 3168 16836 3172 16892
rect 3108 16832 3172 16836
rect 3188 16892 3252 16896
rect 3188 16836 3192 16892
rect 3192 16836 3248 16892
rect 3248 16836 3252 16892
rect 3188 16832 3252 16836
rect 3268 16892 3332 16896
rect 3268 16836 3272 16892
rect 3272 16836 3328 16892
rect 3328 16836 3332 16892
rect 3268 16832 3332 16836
rect 3348 16892 3412 16896
rect 3348 16836 3352 16892
rect 3352 16836 3408 16892
rect 3408 16836 3412 16892
rect 3348 16832 3412 16836
rect 6208 16892 6272 16896
rect 6208 16836 6212 16892
rect 6212 16836 6268 16892
rect 6268 16836 6272 16892
rect 6208 16832 6272 16836
rect 6288 16892 6352 16896
rect 6288 16836 6292 16892
rect 6292 16836 6348 16892
rect 6348 16836 6352 16892
rect 6288 16832 6352 16836
rect 6368 16892 6432 16896
rect 6368 16836 6372 16892
rect 6372 16836 6428 16892
rect 6428 16836 6432 16892
rect 6368 16832 6432 16836
rect 6448 16892 6512 16896
rect 6448 16836 6452 16892
rect 6452 16836 6508 16892
rect 6508 16836 6512 16892
rect 6448 16832 6512 16836
rect 9308 16892 9372 16896
rect 9308 16836 9312 16892
rect 9312 16836 9368 16892
rect 9368 16836 9372 16892
rect 9308 16832 9372 16836
rect 9388 16892 9452 16896
rect 9388 16836 9392 16892
rect 9392 16836 9448 16892
rect 9448 16836 9452 16892
rect 9388 16832 9452 16836
rect 9468 16892 9532 16896
rect 9468 16836 9472 16892
rect 9472 16836 9528 16892
rect 9528 16836 9532 16892
rect 9468 16832 9532 16836
rect 9548 16892 9612 16896
rect 9548 16836 9552 16892
rect 9552 16836 9608 16892
rect 9608 16836 9612 16892
rect 9548 16832 9612 16836
rect 12408 16892 12472 16896
rect 12408 16836 12412 16892
rect 12412 16836 12468 16892
rect 12468 16836 12472 16892
rect 12408 16832 12472 16836
rect 12488 16892 12552 16896
rect 12488 16836 12492 16892
rect 12492 16836 12548 16892
rect 12548 16836 12552 16892
rect 12488 16832 12552 16836
rect 12568 16892 12632 16896
rect 12568 16836 12572 16892
rect 12572 16836 12628 16892
rect 12628 16836 12632 16892
rect 12568 16832 12632 16836
rect 12648 16892 12712 16896
rect 12648 16836 12652 16892
rect 12652 16836 12708 16892
rect 12708 16836 12712 16892
rect 12648 16832 12712 16836
rect 15508 16892 15572 16896
rect 15508 16836 15512 16892
rect 15512 16836 15568 16892
rect 15568 16836 15572 16892
rect 15508 16832 15572 16836
rect 15588 16892 15652 16896
rect 15588 16836 15592 16892
rect 15592 16836 15648 16892
rect 15648 16836 15652 16892
rect 15588 16832 15652 16836
rect 15668 16892 15732 16896
rect 15668 16836 15672 16892
rect 15672 16836 15728 16892
rect 15728 16836 15732 16892
rect 15668 16832 15732 16836
rect 15748 16892 15812 16896
rect 15748 16836 15752 16892
rect 15752 16836 15808 16892
rect 15808 16836 15812 16892
rect 15748 16832 15812 16836
rect 18608 16892 18672 16896
rect 18608 16836 18612 16892
rect 18612 16836 18668 16892
rect 18668 16836 18672 16892
rect 18608 16832 18672 16836
rect 18688 16892 18752 16896
rect 18688 16836 18692 16892
rect 18692 16836 18748 16892
rect 18748 16836 18752 16892
rect 18688 16832 18752 16836
rect 18768 16892 18832 16896
rect 18768 16836 18772 16892
rect 18772 16836 18828 16892
rect 18828 16836 18832 16892
rect 18768 16832 18832 16836
rect 18848 16892 18912 16896
rect 18848 16836 18852 16892
rect 18852 16836 18908 16892
rect 18908 16836 18912 16892
rect 18848 16832 18912 16836
rect 1558 16348 1622 16352
rect 1558 16292 1562 16348
rect 1562 16292 1618 16348
rect 1618 16292 1622 16348
rect 1558 16288 1622 16292
rect 1638 16348 1702 16352
rect 1638 16292 1642 16348
rect 1642 16292 1698 16348
rect 1698 16292 1702 16348
rect 1638 16288 1702 16292
rect 1718 16348 1782 16352
rect 1718 16292 1722 16348
rect 1722 16292 1778 16348
rect 1778 16292 1782 16348
rect 1718 16288 1782 16292
rect 1798 16348 1862 16352
rect 1798 16292 1802 16348
rect 1802 16292 1858 16348
rect 1858 16292 1862 16348
rect 1798 16288 1862 16292
rect 4658 16348 4722 16352
rect 4658 16292 4662 16348
rect 4662 16292 4718 16348
rect 4718 16292 4722 16348
rect 4658 16288 4722 16292
rect 4738 16348 4802 16352
rect 4738 16292 4742 16348
rect 4742 16292 4798 16348
rect 4798 16292 4802 16348
rect 4738 16288 4802 16292
rect 4818 16348 4882 16352
rect 4818 16292 4822 16348
rect 4822 16292 4878 16348
rect 4878 16292 4882 16348
rect 4818 16288 4882 16292
rect 4898 16348 4962 16352
rect 4898 16292 4902 16348
rect 4902 16292 4958 16348
rect 4958 16292 4962 16348
rect 4898 16288 4962 16292
rect 7758 16348 7822 16352
rect 7758 16292 7762 16348
rect 7762 16292 7818 16348
rect 7818 16292 7822 16348
rect 7758 16288 7822 16292
rect 7838 16348 7902 16352
rect 7838 16292 7842 16348
rect 7842 16292 7898 16348
rect 7898 16292 7902 16348
rect 7838 16288 7902 16292
rect 7918 16348 7982 16352
rect 7918 16292 7922 16348
rect 7922 16292 7978 16348
rect 7978 16292 7982 16348
rect 7918 16288 7982 16292
rect 7998 16348 8062 16352
rect 7998 16292 8002 16348
rect 8002 16292 8058 16348
rect 8058 16292 8062 16348
rect 7998 16288 8062 16292
rect 10858 16348 10922 16352
rect 10858 16292 10862 16348
rect 10862 16292 10918 16348
rect 10918 16292 10922 16348
rect 10858 16288 10922 16292
rect 10938 16348 11002 16352
rect 10938 16292 10942 16348
rect 10942 16292 10998 16348
rect 10998 16292 11002 16348
rect 10938 16288 11002 16292
rect 11018 16348 11082 16352
rect 11018 16292 11022 16348
rect 11022 16292 11078 16348
rect 11078 16292 11082 16348
rect 11018 16288 11082 16292
rect 11098 16348 11162 16352
rect 11098 16292 11102 16348
rect 11102 16292 11158 16348
rect 11158 16292 11162 16348
rect 11098 16288 11162 16292
rect 13958 16348 14022 16352
rect 13958 16292 13962 16348
rect 13962 16292 14018 16348
rect 14018 16292 14022 16348
rect 13958 16288 14022 16292
rect 14038 16348 14102 16352
rect 14038 16292 14042 16348
rect 14042 16292 14098 16348
rect 14098 16292 14102 16348
rect 14038 16288 14102 16292
rect 14118 16348 14182 16352
rect 14118 16292 14122 16348
rect 14122 16292 14178 16348
rect 14178 16292 14182 16348
rect 14118 16288 14182 16292
rect 14198 16348 14262 16352
rect 14198 16292 14202 16348
rect 14202 16292 14258 16348
rect 14258 16292 14262 16348
rect 14198 16288 14262 16292
rect 17058 16348 17122 16352
rect 17058 16292 17062 16348
rect 17062 16292 17118 16348
rect 17118 16292 17122 16348
rect 17058 16288 17122 16292
rect 17138 16348 17202 16352
rect 17138 16292 17142 16348
rect 17142 16292 17198 16348
rect 17198 16292 17202 16348
rect 17138 16288 17202 16292
rect 17218 16348 17282 16352
rect 17218 16292 17222 16348
rect 17222 16292 17278 16348
rect 17278 16292 17282 16348
rect 17218 16288 17282 16292
rect 17298 16348 17362 16352
rect 17298 16292 17302 16348
rect 17302 16292 17358 16348
rect 17358 16292 17362 16348
rect 17298 16288 17362 16292
rect 3108 15804 3172 15808
rect 3108 15748 3112 15804
rect 3112 15748 3168 15804
rect 3168 15748 3172 15804
rect 3108 15744 3172 15748
rect 3188 15804 3252 15808
rect 3188 15748 3192 15804
rect 3192 15748 3248 15804
rect 3248 15748 3252 15804
rect 3188 15744 3252 15748
rect 3268 15804 3332 15808
rect 3268 15748 3272 15804
rect 3272 15748 3328 15804
rect 3328 15748 3332 15804
rect 3268 15744 3332 15748
rect 3348 15804 3412 15808
rect 3348 15748 3352 15804
rect 3352 15748 3408 15804
rect 3408 15748 3412 15804
rect 3348 15744 3412 15748
rect 6208 15804 6272 15808
rect 6208 15748 6212 15804
rect 6212 15748 6268 15804
rect 6268 15748 6272 15804
rect 6208 15744 6272 15748
rect 6288 15804 6352 15808
rect 6288 15748 6292 15804
rect 6292 15748 6348 15804
rect 6348 15748 6352 15804
rect 6288 15744 6352 15748
rect 6368 15804 6432 15808
rect 6368 15748 6372 15804
rect 6372 15748 6428 15804
rect 6428 15748 6432 15804
rect 6368 15744 6432 15748
rect 6448 15804 6512 15808
rect 6448 15748 6452 15804
rect 6452 15748 6508 15804
rect 6508 15748 6512 15804
rect 6448 15744 6512 15748
rect 9308 15804 9372 15808
rect 9308 15748 9312 15804
rect 9312 15748 9368 15804
rect 9368 15748 9372 15804
rect 9308 15744 9372 15748
rect 9388 15804 9452 15808
rect 9388 15748 9392 15804
rect 9392 15748 9448 15804
rect 9448 15748 9452 15804
rect 9388 15744 9452 15748
rect 9468 15804 9532 15808
rect 9468 15748 9472 15804
rect 9472 15748 9528 15804
rect 9528 15748 9532 15804
rect 9468 15744 9532 15748
rect 9548 15804 9612 15808
rect 9548 15748 9552 15804
rect 9552 15748 9608 15804
rect 9608 15748 9612 15804
rect 9548 15744 9612 15748
rect 12408 15804 12472 15808
rect 12408 15748 12412 15804
rect 12412 15748 12468 15804
rect 12468 15748 12472 15804
rect 12408 15744 12472 15748
rect 12488 15804 12552 15808
rect 12488 15748 12492 15804
rect 12492 15748 12548 15804
rect 12548 15748 12552 15804
rect 12488 15744 12552 15748
rect 12568 15804 12632 15808
rect 12568 15748 12572 15804
rect 12572 15748 12628 15804
rect 12628 15748 12632 15804
rect 12568 15744 12632 15748
rect 12648 15804 12712 15808
rect 12648 15748 12652 15804
rect 12652 15748 12708 15804
rect 12708 15748 12712 15804
rect 12648 15744 12712 15748
rect 15508 15804 15572 15808
rect 15508 15748 15512 15804
rect 15512 15748 15568 15804
rect 15568 15748 15572 15804
rect 15508 15744 15572 15748
rect 15588 15804 15652 15808
rect 15588 15748 15592 15804
rect 15592 15748 15648 15804
rect 15648 15748 15652 15804
rect 15588 15744 15652 15748
rect 15668 15804 15732 15808
rect 15668 15748 15672 15804
rect 15672 15748 15728 15804
rect 15728 15748 15732 15804
rect 15668 15744 15732 15748
rect 15748 15804 15812 15808
rect 15748 15748 15752 15804
rect 15752 15748 15808 15804
rect 15808 15748 15812 15804
rect 15748 15744 15812 15748
rect 18608 15804 18672 15808
rect 18608 15748 18612 15804
rect 18612 15748 18668 15804
rect 18668 15748 18672 15804
rect 18608 15744 18672 15748
rect 18688 15804 18752 15808
rect 18688 15748 18692 15804
rect 18692 15748 18748 15804
rect 18748 15748 18752 15804
rect 18688 15744 18752 15748
rect 18768 15804 18832 15808
rect 18768 15748 18772 15804
rect 18772 15748 18828 15804
rect 18828 15748 18832 15804
rect 18768 15744 18832 15748
rect 18848 15804 18912 15808
rect 18848 15748 18852 15804
rect 18852 15748 18908 15804
rect 18908 15748 18912 15804
rect 18848 15744 18912 15748
rect 1558 15260 1622 15264
rect 1558 15204 1562 15260
rect 1562 15204 1618 15260
rect 1618 15204 1622 15260
rect 1558 15200 1622 15204
rect 1638 15260 1702 15264
rect 1638 15204 1642 15260
rect 1642 15204 1698 15260
rect 1698 15204 1702 15260
rect 1638 15200 1702 15204
rect 1718 15260 1782 15264
rect 1718 15204 1722 15260
rect 1722 15204 1778 15260
rect 1778 15204 1782 15260
rect 1718 15200 1782 15204
rect 1798 15260 1862 15264
rect 1798 15204 1802 15260
rect 1802 15204 1858 15260
rect 1858 15204 1862 15260
rect 1798 15200 1862 15204
rect 4658 15260 4722 15264
rect 4658 15204 4662 15260
rect 4662 15204 4718 15260
rect 4718 15204 4722 15260
rect 4658 15200 4722 15204
rect 4738 15260 4802 15264
rect 4738 15204 4742 15260
rect 4742 15204 4798 15260
rect 4798 15204 4802 15260
rect 4738 15200 4802 15204
rect 4818 15260 4882 15264
rect 4818 15204 4822 15260
rect 4822 15204 4878 15260
rect 4878 15204 4882 15260
rect 4818 15200 4882 15204
rect 4898 15260 4962 15264
rect 4898 15204 4902 15260
rect 4902 15204 4958 15260
rect 4958 15204 4962 15260
rect 4898 15200 4962 15204
rect 7758 15260 7822 15264
rect 7758 15204 7762 15260
rect 7762 15204 7818 15260
rect 7818 15204 7822 15260
rect 7758 15200 7822 15204
rect 7838 15260 7902 15264
rect 7838 15204 7842 15260
rect 7842 15204 7898 15260
rect 7898 15204 7902 15260
rect 7838 15200 7902 15204
rect 7918 15260 7982 15264
rect 7918 15204 7922 15260
rect 7922 15204 7978 15260
rect 7978 15204 7982 15260
rect 7918 15200 7982 15204
rect 7998 15260 8062 15264
rect 7998 15204 8002 15260
rect 8002 15204 8058 15260
rect 8058 15204 8062 15260
rect 7998 15200 8062 15204
rect 10858 15260 10922 15264
rect 10858 15204 10862 15260
rect 10862 15204 10918 15260
rect 10918 15204 10922 15260
rect 10858 15200 10922 15204
rect 10938 15260 11002 15264
rect 10938 15204 10942 15260
rect 10942 15204 10998 15260
rect 10998 15204 11002 15260
rect 10938 15200 11002 15204
rect 11018 15260 11082 15264
rect 11018 15204 11022 15260
rect 11022 15204 11078 15260
rect 11078 15204 11082 15260
rect 11018 15200 11082 15204
rect 11098 15260 11162 15264
rect 11098 15204 11102 15260
rect 11102 15204 11158 15260
rect 11158 15204 11162 15260
rect 11098 15200 11162 15204
rect 13958 15260 14022 15264
rect 13958 15204 13962 15260
rect 13962 15204 14018 15260
rect 14018 15204 14022 15260
rect 13958 15200 14022 15204
rect 14038 15260 14102 15264
rect 14038 15204 14042 15260
rect 14042 15204 14098 15260
rect 14098 15204 14102 15260
rect 14038 15200 14102 15204
rect 14118 15260 14182 15264
rect 14118 15204 14122 15260
rect 14122 15204 14178 15260
rect 14178 15204 14182 15260
rect 14118 15200 14182 15204
rect 14198 15260 14262 15264
rect 14198 15204 14202 15260
rect 14202 15204 14258 15260
rect 14258 15204 14262 15260
rect 14198 15200 14262 15204
rect 17058 15260 17122 15264
rect 17058 15204 17062 15260
rect 17062 15204 17118 15260
rect 17118 15204 17122 15260
rect 17058 15200 17122 15204
rect 17138 15260 17202 15264
rect 17138 15204 17142 15260
rect 17142 15204 17198 15260
rect 17198 15204 17202 15260
rect 17138 15200 17202 15204
rect 17218 15260 17282 15264
rect 17218 15204 17222 15260
rect 17222 15204 17278 15260
rect 17278 15204 17282 15260
rect 17218 15200 17282 15204
rect 17298 15260 17362 15264
rect 17298 15204 17302 15260
rect 17302 15204 17358 15260
rect 17358 15204 17362 15260
rect 17298 15200 17362 15204
rect 3108 14716 3172 14720
rect 3108 14660 3112 14716
rect 3112 14660 3168 14716
rect 3168 14660 3172 14716
rect 3108 14656 3172 14660
rect 3188 14716 3252 14720
rect 3188 14660 3192 14716
rect 3192 14660 3248 14716
rect 3248 14660 3252 14716
rect 3188 14656 3252 14660
rect 3268 14716 3332 14720
rect 3268 14660 3272 14716
rect 3272 14660 3328 14716
rect 3328 14660 3332 14716
rect 3268 14656 3332 14660
rect 3348 14716 3412 14720
rect 3348 14660 3352 14716
rect 3352 14660 3408 14716
rect 3408 14660 3412 14716
rect 3348 14656 3412 14660
rect 6208 14716 6272 14720
rect 6208 14660 6212 14716
rect 6212 14660 6268 14716
rect 6268 14660 6272 14716
rect 6208 14656 6272 14660
rect 6288 14716 6352 14720
rect 6288 14660 6292 14716
rect 6292 14660 6348 14716
rect 6348 14660 6352 14716
rect 6288 14656 6352 14660
rect 6368 14716 6432 14720
rect 6368 14660 6372 14716
rect 6372 14660 6428 14716
rect 6428 14660 6432 14716
rect 6368 14656 6432 14660
rect 6448 14716 6512 14720
rect 6448 14660 6452 14716
rect 6452 14660 6508 14716
rect 6508 14660 6512 14716
rect 6448 14656 6512 14660
rect 9308 14716 9372 14720
rect 9308 14660 9312 14716
rect 9312 14660 9368 14716
rect 9368 14660 9372 14716
rect 9308 14656 9372 14660
rect 9388 14716 9452 14720
rect 9388 14660 9392 14716
rect 9392 14660 9448 14716
rect 9448 14660 9452 14716
rect 9388 14656 9452 14660
rect 9468 14716 9532 14720
rect 9468 14660 9472 14716
rect 9472 14660 9528 14716
rect 9528 14660 9532 14716
rect 9468 14656 9532 14660
rect 9548 14716 9612 14720
rect 9548 14660 9552 14716
rect 9552 14660 9608 14716
rect 9608 14660 9612 14716
rect 9548 14656 9612 14660
rect 12408 14716 12472 14720
rect 12408 14660 12412 14716
rect 12412 14660 12468 14716
rect 12468 14660 12472 14716
rect 12408 14656 12472 14660
rect 12488 14716 12552 14720
rect 12488 14660 12492 14716
rect 12492 14660 12548 14716
rect 12548 14660 12552 14716
rect 12488 14656 12552 14660
rect 12568 14716 12632 14720
rect 12568 14660 12572 14716
rect 12572 14660 12628 14716
rect 12628 14660 12632 14716
rect 12568 14656 12632 14660
rect 12648 14716 12712 14720
rect 12648 14660 12652 14716
rect 12652 14660 12708 14716
rect 12708 14660 12712 14716
rect 12648 14656 12712 14660
rect 15508 14716 15572 14720
rect 15508 14660 15512 14716
rect 15512 14660 15568 14716
rect 15568 14660 15572 14716
rect 15508 14656 15572 14660
rect 15588 14716 15652 14720
rect 15588 14660 15592 14716
rect 15592 14660 15648 14716
rect 15648 14660 15652 14716
rect 15588 14656 15652 14660
rect 15668 14716 15732 14720
rect 15668 14660 15672 14716
rect 15672 14660 15728 14716
rect 15728 14660 15732 14716
rect 15668 14656 15732 14660
rect 15748 14716 15812 14720
rect 15748 14660 15752 14716
rect 15752 14660 15808 14716
rect 15808 14660 15812 14716
rect 15748 14656 15812 14660
rect 18608 14716 18672 14720
rect 18608 14660 18612 14716
rect 18612 14660 18668 14716
rect 18668 14660 18672 14716
rect 18608 14656 18672 14660
rect 18688 14716 18752 14720
rect 18688 14660 18692 14716
rect 18692 14660 18748 14716
rect 18748 14660 18752 14716
rect 18688 14656 18752 14660
rect 18768 14716 18832 14720
rect 18768 14660 18772 14716
rect 18772 14660 18828 14716
rect 18828 14660 18832 14716
rect 18768 14656 18832 14660
rect 18848 14716 18912 14720
rect 18848 14660 18852 14716
rect 18852 14660 18908 14716
rect 18908 14660 18912 14716
rect 18848 14656 18912 14660
rect 1558 14172 1622 14176
rect 1558 14116 1562 14172
rect 1562 14116 1618 14172
rect 1618 14116 1622 14172
rect 1558 14112 1622 14116
rect 1638 14172 1702 14176
rect 1638 14116 1642 14172
rect 1642 14116 1698 14172
rect 1698 14116 1702 14172
rect 1638 14112 1702 14116
rect 1718 14172 1782 14176
rect 1718 14116 1722 14172
rect 1722 14116 1778 14172
rect 1778 14116 1782 14172
rect 1718 14112 1782 14116
rect 1798 14172 1862 14176
rect 1798 14116 1802 14172
rect 1802 14116 1858 14172
rect 1858 14116 1862 14172
rect 1798 14112 1862 14116
rect 4658 14172 4722 14176
rect 4658 14116 4662 14172
rect 4662 14116 4718 14172
rect 4718 14116 4722 14172
rect 4658 14112 4722 14116
rect 4738 14172 4802 14176
rect 4738 14116 4742 14172
rect 4742 14116 4798 14172
rect 4798 14116 4802 14172
rect 4738 14112 4802 14116
rect 4818 14172 4882 14176
rect 4818 14116 4822 14172
rect 4822 14116 4878 14172
rect 4878 14116 4882 14172
rect 4818 14112 4882 14116
rect 4898 14172 4962 14176
rect 4898 14116 4902 14172
rect 4902 14116 4958 14172
rect 4958 14116 4962 14172
rect 4898 14112 4962 14116
rect 7758 14172 7822 14176
rect 7758 14116 7762 14172
rect 7762 14116 7818 14172
rect 7818 14116 7822 14172
rect 7758 14112 7822 14116
rect 7838 14172 7902 14176
rect 7838 14116 7842 14172
rect 7842 14116 7898 14172
rect 7898 14116 7902 14172
rect 7838 14112 7902 14116
rect 7918 14172 7982 14176
rect 7918 14116 7922 14172
rect 7922 14116 7978 14172
rect 7978 14116 7982 14172
rect 7918 14112 7982 14116
rect 7998 14172 8062 14176
rect 7998 14116 8002 14172
rect 8002 14116 8058 14172
rect 8058 14116 8062 14172
rect 7998 14112 8062 14116
rect 10858 14172 10922 14176
rect 10858 14116 10862 14172
rect 10862 14116 10918 14172
rect 10918 14116 10922 14172
rect 10858 14112 10922 14116
rect 10938 14172 11002 14176
rect 10938 14116 10942 14172
rect 10942 14116 10998 14172
rect 10998 14116 11002 14172
rect 10938 14112 11002 14116
rect 11018 14172 11082 14176
rect 11018 14116 11022 14172
rect 11022 14116 11078 14172
rect 11078 14116 11082 14172
rect 11018 14112 11082 14116
rect 11098 14172 11162 14176
rect 11098 14116 11102 14172
rect 11102 14116 11158 14172
rect 11158 14116 11162 14172
rect 11098 14112 11162 14116
rect 13958 14172 14022 14176
rect 13958 14116 13962 14172
rect 13962 14116 14018 14172
rect 14018 14116 14022 14172
rect 13958 14112 14022 14116
rect 14038 14172 14102 14176
rect 14038 14116 14042 14172
rect 14042 14116 14098 14172
rect 14098 14116 14102 14172
rect 14038 14112 14102 14116
rect 14118 14172 14182 14176
rect 14118 14116 14122 14172
rect 14122 14116 14178 14172
rect 14178 14116 14182 14172
rect 14118 14112 14182 14116
rect 14198 14172 14262 14176
rect 14198 14116 14202 14172
rect 14202 14116 14258 14172
rect 14258 14116 14262 14172
rect 14198 14112 14262 14116
rect 17058 14172 17122 14176
rect 17058 14116 17062 14172
rect 17062 14116 17118 14172
rect 17118 14116 17122 14172
rect 17058 14112 17122 14116
rect 17138 14172 17202 14176
rect 17138 14116 17142 14172
rect 17142 14116 17198 14172
rect 17198 14116 17202 14172
rect 17138 14112 17202 14116
rect 17218 14172 17282 14176
rect 17218 14116 17222 14172
rect 17222 14116 17278 14172
rect 17278 14116 17282 14172
rect 17218 14112 17282 14116
rect 17298 14172 17362 14176
rect 17298 14116 17302 14172
rect 17302 14116 17358 14172
rect 17358 14116 17362 14172
rect 17298 14112 17362 14116
rect 3108 13628 3172 13632
rect 3108 13572 3112 13628
rect 3112 13572 3168 13628
rect 3168 13572 3172 13628
rect 3108 13568 3172 13572
rect 3188 13628 3252 13632
rect 3188 13572 3192 13628
rect 3192 13572 3248 13628
rect 3248 13572 3252 13628
rect 3188 13568 3252 13572
rect 3268 13628 3332 13632
rect 3268 13572 3272 13628
rect 3272 13572 3328 13628
rect 3328 13572 3332 13628
rect 3268 13568 3332 13572
rect 3348 13628 3412 13632
rect 3348 13572 3352 13628
rect 3352 13572 3408 13628
rect 3408 13572 3412 13628
rect 3348 13568 3412 13572
rect 6208 13628 6272 13632
rect 6208 13572 6212 13628
rect 6212 13572 6268 13628
rect 6268 13572 6272 13628
rect 6208 13568 6272 13572
rect 6288 13628 6352 13632
rect 6288 13572 6292 13628
rect 6292 13572 6348 13628
rect 6348 13572 6352 13628
rect 6288 13568 6352 13572
rect 6368 13628 6432 13632
rect 6368 13572 6372 13628
rect 6372 13572 6428 13628
rect 6428 13572 6432 13628
rect 6368 13568 6432 13572
rect 6448 13628 6512 13632
rect 6448 13572 6452 13628
rect 6452 13572 6508 13628
rect 6508 13572 6512 13628
rect 6448 13568 6512 13572
rect 9308 13628 9372 13632
rect 9308 13572 9312 13628
rect 9312 13572 9368 13628
rect 9368 13572 9372 13628
rect 9308 13568 9372 13572
rect 9388 13628 9452 13632
rect 9388 13572 9392 13628
rect 9392 13572 9448 13628
rect 9448 13572 9452 13628
rect 9388 13568 9452 13572
rect 9468 13628 9532 13632
rect 9468 13572 9472 13628
rect 9472 13572 9528 13628
rect 9528 13572 9532 13628
rect 9468 13568 9532 13572
rect 9548 13628 9612 13632
rect 9548 13572 9552 13628
rect 9552 13572 9608 13628
rect 9608 13572 9612 13628
rect 9548 13568 9612 13572
rect 12408 13628 12472 13632
rect 12408 13572 12412 13628
rect 12412 13572 12468 13628
rect 12468 13572 12472 13628
rect 12408 13568 12472 13572
rect 12488 13628 12552 13632
rect 12488 13572 12492 13628
rect 12492 13572 12548 13628
rect 12548 13572 12552 13628
rect 12488 13568 12552 13572
rect 12568 13628 12632 13632
rect 12568 13572 12572 13628
rect 12572 13572 12628 13628
rect 12628 13572 12632 13628
rect 12568 13568 12632 13572
rect 12648 13628 12712 13632
rect 12648 13572 12652 13628
rect 12652 13572 12708 13628
rect 12708 13572 12712 13628
rect 12648 13568 12712 13572
rect 15508 13628 15572 13632
rect 15508 13572 15512 13628
rect 15512 13572 15568 13628
rect 15568 13572 15572 13628
rect 15508 13568 15572 13572
rect 15588 13628 15652 13632
rect 15588 13572 15592 13628
rect 15592 13572 15648 13628
rect 15648 13572 15652 13628
rect 15588 13568 15652 13572
rect 15668 13628 15732 13632
rect 15668 13572 15672 13628
rect 15672 13572 15728 13628
rect 15728 13572 15732 13628
rect 15668 13568 15732 13572
rect 15748 13628 15812 13632
rect 15748 13572 15752 13628
rect 15752 13572 15808 13628
rect 15808 13572 15812 13628
rect 15748 13568 15812 13572
rect 18608 13628 18672 13632
rect 18608 13572 18612 13628
rect 18612 13572 18668 13628
rect 18668 13572 18672 13628
rect 18608 13568 18672 13572
rect 18688 13628 18752 13632
rect 18688 13572 18692 13628
rect 18692 13572 18748 13628
rect 18748 13572 18752 13628
rect 18688 13568 18752 13572
rect 18768 13628 18832 13632
rect 18768 13572 18772 13628
rect 18772 13572 18828 13628
rect 18828 13572 18832 13628
rect 18768 13568 18832 13572
rect 18848 13628 18912 13632
rect 18848 13572 18852 13628
rect 18852 13572 18908 13628
rect 18908 13572 18912 13628
rect 18848 13568 18912 13572
rect 1558 13084 1622 13088
rect 1558 13028 1562 13084
rect 1562 13028 1618 13084
rect 1618 13028 1622 13084
rect 1558 13024 1622 13028
rect 1638 13084 1702 13088
rect 1638 13028 1642 13084
rect 1642 13028 1698 13084
rect 1698 13028 1702 13084
rect 1638 13024 1702 13028
rect 1718 13084 1782 13088
rect 1718 13028 1722 13084
rect 1722 13028 1778 13084
rect 1778 13028 1782 13084
rect 1718 13024 1782 13028
rect 1798 13084 1862 13088
rect 1798 13028 1802 13084
rect 1802 13028 1858 13084
rect 1858 13028 1862 13084
rect 1798 13024 1862 13028
rect 4658 13084 4722 13088
rect 4658 13028 4662 13084
rect 4662 13028 4718 13084
rect 4718 13028 4722 13084
rect 4658 13024 4722 13028
rect 4738 13084 4802 13088
rect 4738 13028 4742 13084
rect 4742 13028 4798 13084
rect 4798 13028 4802 13084
rect 4738 13024 4802 13028
rect 4818 13084 4882 13088
rect 4818 13028 4822 13084
rect 4822 13028 4878 13084
rect 4878 13028 4882 13084
rect 4818 13024 4882 13028
rect 4898 13084 4962 13088
rect 4898 13028 4902 13084
rect 4902 13028 4958 13084
rect 4958 13028 4962 13084
rect 4898 13024 4962 13028
rect 7758 13084 7822 13088
rect 7758 13028 7762 13084
rect 7762 13028 7818 13084
rect 7818 13028 7822 13084
rect 7758 13024 7822 13028
rect 7838 13084 7902 13088
rect 7838 13028 7842 13084
rect 7842 13028 7898 13084
rect 7898 13028 7902 13084
rect 7838 13024 7902 13028
rect 7918 13084 7982 13088
rect 7918 13028 7922 13084
rect 7922 13028 7978 13084
rect 7978 13028 7982 13084
rect 7918 13024 7982 13028
rect 7998 13084 8062 13088
rect 7998 13028 8002 13084
rect 8002 13028 8058 13084
rect 8058 13028 8062 13084
rect 7998 13024 8062 13028
rect 10858 13084 10922 13088
rect 10858 13028 10862 13084
rect 10862 13028 10918 13084
rect 10918 13028 10922 13084
rect 10858 13024 10922 13028
rect 10938 13084 11002 13088
rect 10938 13028 10942 13084
rect 10942 13028 10998 13084
rect 10998 13028 11002 13084
rect 10938 13024 11002 13028
rect 11018 13084 11082 13088
rect 11018 13028 11022 13084
rect 11022 13028 11078 13084
rect 11078 13028 11082 13084
rect 11018 13024 11082 13028
rect 11098 13084 11162 13088
rect 11098 13028 11102 13084
rect 11102 13028 11158 13084
rect 11158 13028 11162 13084
rect 11098 13024 11162 13028
rect 13958 13084 14022 13088
rect 13958 13028 13962 13084
rect 13962 13028 14018 13084
rect 14018 13028 14022 13084
rect 13958 13024 14022 13028
rect 14038 13084 14102 13088
rect 14038 13028 14042 13084
rect 14042 13028 14098 13084
rect 14098 13028 14102 13084
rect 14038 13024 14102 13028
rect 14118 13084 14182 13088
rect 14118 13028 14122 13084
rect 14122 13028 14178 13084
rect 14178 13028 14182 13084
rect 14118 13024 14182 13028
rect 14198 13084 14262 13088
rect 14198 13028 14202 13084
rect 14202 13028 14258 13084
rect 14258 13028 14262 13084
rect 14198 13024 14262 13028
rect 17058 13084 17122 13088
rect 17058 13028 17062 13084
rect 17062 13028 17118 13084
rect 17118 13028 17122 13084
rect 17058 13024 17122 13028
rect 17138 13084 17202 13088
rect 17138 13028 17142 13084
rect 17142 13028 17198 13084
rect 17198 13028 17202 13084
rect 17138 13024 17202 13028
rect 17218 13084 17282 13088
rect 17218 13028 17222 13084
rect 17222 13028 17278 13084
rect 17278 13028 17282 13084
rect 17218 13024 17282 13028
rect 17298 13084 17362 13088
rect 17298 13028 17302 13084
rect 17302 13028 17358 13084
rect 17358 13028 17362 13084
rect 17298 13024 17362 13028
rect 3108 12540 3172 12544
rect 3108 12484 3112 12540
rect 3112 12484 3168 12540
rect 3168 12484 3172 12540
rect 3108 12480 3172 12484
rect 3188 12540 3252 12544
rect 3188 12484 3192 12540
rect 3192 12484 3248 12540
rect 3248 12484 3252 12540
rect 3188 12480 3252 12484
rect 3268 12540 3332 12544
rect 3268 12484 3272 12540
rect 3272 12484 3328 12540
rect 3328 12484 3332 12540
rect 3268 12480 3332 12484
rect 3348 12540 3412 12544
rect 3348 12484 3352 12540
rect 3352 12484 3408 12540
rect 3408 12484 3412 12540
rect 3348 12480 3412 12484
rect 6208 12540 6272 12544
rect 6208 12484 6212 12540
rect 6212 12484 6268 12540
rect 6268 12484 6272 12540
rect 6208 12480 6272 12484
rect 6288 12540 6352 12544
rect 6288 12484 6292 12540
rect 6292 12484 6348 12540
rect 6348 12484 6352 12540
rect 6288 12480 6352 12484
rect 6368 12540 6432 12544
rect 6368 12484 6372 12540
rect 6372 12484 6428 12540
rect 6428 12484 6432 12540
rect 6368 12480 6432 12484
rect 6448 12540 6512 12544
rect 6448 12484 6452 12540
rect 6452 12484 6508 12540
rect 6508 12484 6512 12540
rect 6448 12480 6512 12484
rect 9308 12540 9372 12544
rect 9308 12484 9312 12540
rect 9312 12484 9368 12540
rect 9368 12484 9372 12540
rect 9308 12480 9372 12484
rect 9388 12540 9452 12544
rect 9388 12484 9392 12540
rect 9392 12484 9448 12540
rect 9448 12484 9452 12540
rect 9388 12480 9452 12484
rect 9468 12540 9532 12544
rect 9468 12484 9472 12540
rect 9472 12484 9528 12540
rect 9528 12484 9532 12540
rect 9468 12480 9532 12484
rect 9548 12540 9612 12544
rect 9548 12484 9552 12540
rect 9552 12484 9608 12540
rect 9608 12484 9612 12540
rect 9548 12480 9612 12484
rect 12408 12540 12472 12544
rect 12408 12484 12412 12540
rect 12412 12484 12468 12540
rect 12468 12484 12472 12540
rect 12408 12480 12472 12484
rect 12488 12540 12552 12544
rect 12488 12484 12492 12540
rect 12492 12484 12548 12540
rect 12548 12484 12552 12540
rect 12488 12480 12552 12484
rect 12568 12540 12632 12544
rect 12568 12484 12572 12540
rect 12572 12484 12628 12540
rect 12628 12484 12632 12540
rect 12568 12480 12632 12484
rect 12648 12540 12712 12544
rect 12648 12484 12652 12540
rect 12652 12484 12708 12540
rect 12708 12484 12712 12540
rect 12648 12480 12712 12484
rect 15508 12540 15572 12544
rect 15508 12484 15512 12540
rect 15512 12484 15568 12540
rect 15568 12484 15572 12540
rect 15508 12480 15572 12484
rect 15588 12540 15652 12544
rect 15588 12484 15592 12540
rect 15592 12484 15648 12540
rect 15648 12484 15652 12540
rect 15588 12480 15652 12484
rect 15668 12540 15732 12544
rect 15668 12484 15672 12540
rect 15672 12484 15728 12540
rect 15728 12484 15732 12540
rect 15668 12480 15732 12484
rect 15748 12540 15812 12544
rect 15748 12484 15752 12540
rect 15752 12484 15808 12540
rect 15808 12484 15812 12540
rect 15748 12480 15812 12484
rect 18608 12540 18672 12544
rect 18608 12484 18612 12540
rect 18612 12484 18668 12540
rect 18668 12484 18672 12540
rect 18608 12480 18672 12484
rect 18688 12540 18752 12544
rect 18688 12484 18692 12540
rect 18692 12484 18748 12540
rect 18748 12484 18752 12540
rect 18688 12480 18752 12484
rect 18768 12540 18832 12544
rect 18768 12484 18772 12540
rect 18772 12484 18828 12540
rect 18828 12484 18832 12540
rect 18768 12480 18832 12484
rect 18848 12540 18912 12544
rect 18848 12484 18852 12540
rect 18852 12484 18908 12540
rect 18908 12484 18912 12540
rect 18848 12480 18912 12484
rect 1558 11996 1622 12000
rect 1558 11940 1562 11996
rect 1562 11940 1618 11996
rect 1618 11940 1622 11996
rect 1558 11936 1622 11940
rect 1638 11996 1702 12000
rect 1638 11940 1642 11996
rect 1642 11940 1698 11996
rect 1698 11940 1702 11996
rect 1638 11936 1702 11940
rect 1718 11996 1782 12000
rect 1718 11940 1722 11996
rect 1722 11940 1778 11996
rect 1778 11940 1782 11996
rect 1718 11936 1782 11940
rect 1798 11996 1862 12000
rect 1798 11940 1802 11996
rect 1802 11940 1858 11996
rect 1858 11940 1862 11996
rect 1798 11936 1862 11940
rect 4658 11996 4722 12000
rect 4658 11940 4662 11996
rect 4662 11940 4718 11996
rect 4718 11940 4722 11996
rect 4658 11936 4722 11940
rect 4738 11996 4802 12000
rect 4738 11940 4742 11996
rect 4742 11940 4798 11996
rect 4798 11940 4802 11996
rect 4738 11936 4802 11940
rect 4818 11996 4882 12000
rect 4818 11940 4822 11996
rect 4822 11940 4878 11996
rect 4878 11940 4882 11996
rect 4818 11936 4882 11940
rect 4898 11996 4962 12000
rect 4898 11940 4902 11996
rect 4902 11940 4958 11996
rect 4958 11940 4962 11996
rect 4898 11936 4962 11940
rect 7758 11996 7822 12000
rect 7758 11940 7762 11996
rect 7762 11940 7818 11996
rect 7818 11940 7822 11996
rect 7758 11936 7822 11940
rect 7838 11996 7902 12000
rect 7838 11940 7842 11996
rect 7842 11940 7898 11996
rect 7898 11940 7902 11996
rect 7838 11936 7902 11940
rect 7918 11996 7982 12000
rect 7918 11940 7922 11996
rect 7922 11940 7978 11996
rect 7978 11940 7982 11996
rect 7918 11936 7982 11940
rect 7998 11996 8062 12000
rect 7998 11940 8002 11996
rect 8002 11940 8058 11996
rect 8058 11940 8062 11996
rect 7998 11936 8062 11940
rect 10858 11996 10922 12000
rect 10858 11940 10862 11996
rect 10862 11940 10918 11996
rect 10918 11940 10922 11996
rect 10858 11936 10922 11940
rect 10938 11996 11002 12000
rect 10938 11940 10942 11996
rect 10942 11940 10998 11996
rect 10998 11940 11002 11996
rect 10938 11936 11002 11940
rect 11018 11996 11082 12000
rect 11018 11940 11022 11996
rect 11022 11940 11078 11996
rect 11078 11940 11082 11996
rect 11018 11936 11082 11940
rect 11098 11996 11162 12000
rect 11098 11940 11102 11996
rect 11102 11940 11158 11996
rect 11158 11940 11162 11996
rect 11098 11936 11162 11940
rect 13958 11996 14022 12000
rect 13958 11940 13962 11996
rect 13962 11940 14018 11996
rect 14018 11940 14022 11996
rect 13958 11936 14022 11940
rect 14038 11996 14102 12000
rect 14038 11940 14042 11996
rect 14042 11940 14098 11996
rect 14098 11940 14102 11996
rect 14038 11936 14102 11940
rect 14118 11996 14182 12000
rect 14118 11940 14122 11996
rect 14122 11940 14178 11996
rect 14178 11940 14182 11996
rect 14118 11936 14182 11940
rect 14198 11996 14262 12000
rect 14198 11940 14202 11996
rect 14202 11940 14258 11996
rect 14258 11940 14262 11996
rect 14198 11936 14262 11940
rect 17058 11996 17122 12000
rect 17058 11940 17062 11996
rect 17062 11940 17118 11996
rect 17118 11940 17122 11996
rect 17058 11936 17122 11940
rect 17138 11996 17202 12000
rect 17138 11940 17142 11996
rect 17142 11940 17198 11996
rect 17198 11940 17202 11996
rect 17138 11936 17202 11940
rect 17218 11996 17282 12000
rect 17218 11940 17222 11996
rect 17222 11940 17278 11996
rect 17278 11940 17282 11996
rect 17218 11936 17282 11940
rect 17298 11996 17362 12000
rect 17298 11940 17302 11996
rect 17302 11940 17358 11996
rect 17358 11940 17362 11996
rect 17298 11936 17362 11940
rect 3108 11452 3172 11456
rect 3108 11396 3112 11452
rect 3112 11396 3168 11452
rect 3168 11396 3172 11452
rect 3108 11392 3172 11396
rect 3188 11452 3252 11456
rect 3188 11396 3192 11452
rect 3192 11396 3248 11452
rect 3248 11396 3252 11452
rect 3188 11392 3252 11396
rect 3268 11452 3332 11456
rect 3268 11396 3272 11452
rect 3272 11396 3328 11452
rect 3328 11396 3332 11452
rect 3268 11392 3332 11396
rect 3348 11452 3412 11456
rect 3348 11396 3352 11452
rect 3352 11396 3408 11452
rect 3408 11396 3412 11452
rect 3348 11392 3412 11396
rect 6208 11452 6272 11456
rect 6208 11396 6212 11452
rect 6212 11396 6268 11452
rect 6268 11396 6272 11452
rect 6208 11392 6272 11396
rect 6288 11452 6352 11456
rect 6288 11396 6292 11452
rect 6292 11396 6348 11452
rect 6348 11396 6352 11452
rect 6288 11392 6352 11396
rect 6368 11452 6432 11456
rect 6368 11396 6372 11452
rect 6372 11396 6428 11452
rect 6428 11396 6432 11452
rect 6368 11392 6432 11396
rect 6448 11452 6512 11456
rect 6448 11396 6452 11452
rect 6452 11396 6508 11452
rect 6508 11396 6512 11452
rect 6448 11392 6512 11396
rect 9308 11452 9372 11456
rect 9308 11396 9312 11452
rect 9312 11396 9368 11452
rect 9368 11396 9372 11452
rect 9308 11392 9372 11396
rect 9388 11452 9452 11456
rect 9388 11396 9392 11452
rect 9392 11396 9448 11452
rect 9448 11396 9452 11452
rect 9388 11392 9452 11396
rect 9468 11452 9532 11456
rect 9468 11396 9472 11452
rect 9472 11396 9528 11452
rect 9528 11396 9532 11452
rect 9468 11392 9532 11396
rect 9548 11452 9612 11456
rect 9548 11396 9552 11452
rect 9552 11396 9608 11452
rect 9608 11396 9612 11452
rect 9548 11392 9612 11396
rect 12408 11452 12472 11456
rect 12408 11396 12412 11452
rect 12412 11396 12468 11452
rect 12468 11396 12472 11452
rect 12408 11392 12472 11396
rect 12488 11452 12552 11456
rect 12488 11396 12492 11452
rect 12492 11396 12548 11452
rect 12548 11396 12552 11452
rect 12488 11392 12552 11396
rect 12568 11452 12632 11456
rect 12568 11396 12572 11452
rect 12572 11396 12628 11452
rect 12628 11396 12632 11452
rect 12568 11392 12632 11396
rect 12648 11452 12712 11456
rect 12648 11396 12652 11452
rect 12652 11396 12708 11452
rect 12708 11396 12712 11452
rect 12648 11392 12712 11396
rect 15508 11452 15572 11456
rect 15508 11396 15512 11452
rect 15512 11396 15568 11452
rect 15568 11396 15572 11452
rect 15508 11392 15572 11396
rect 15588 11452 15652 11456
rect 15588 11396 15592 11452
rect 15592 11396 15648 11452
rect 15648 11396 15652 11452
rect 15588 11392 15652 11396
rect 15668 11452 15732 11456
rect 15668 11396 15672 11452
rect 15672 11396 15728 11452
rect 15728 11396 15732 11452
rect 15668 11392 15732 11396
rect 15748 11452 15812 11456
rect 15748 11396 15752 11452
rect 15752 11396 15808 11452
rect 15808 11396 15812 11452
rect 15748 11392 15812 11396
rect 18608 11452 18672 11456
rect 18608 11396 18612 11452
rect 18612 11396 18668 11452
rect 18668 11396 18672 11452
rect 18608 11392 18672 11396
rect 18688 11452 18752 11456
rect 18688 11396 18692 11452
rect 18692 11396 18748 11452
rect 18748 11396 18752 11452
rect 18688 11392 18752 11396
rect 18768 11452 18832 11456
rect 18768 11396 18772 11452
rect 18772 11396 18828 11452
rect 18828 11396 18832 11452
rect 18768 11392 18832 11396
rect 18848 11452 18912 11456
rect 18848 11396 18852 11452
rect 18852 11396 18908 11452
rect 18908 11396 18912 11452
rect 18848 11392 18912 11396
rect 1558 10908 1622 10912
rect 1558 10852 1562 10908
rect 1562 10852 1618 10908
rect 1618 10852 1622 10908
rect 1558 10848 1622 10852
rect 1638 10908 1702 10912
rect 1638 10852 1642 10908
rect 1642 10852 1698 10908
rect 1698 10852 1702 10908
rect 1638 10848 1702 10852
rect 1718 10908 1782 10912
rect 1718 10852 1722 10908
rect 1722 10852 1778 10908
rect 1778 10852 1782 10908
rect 1718 10848 1782 10852
rect 1798 10908 1862 10912
rect 1798 10852 1802 10908
rect 1802 10852 1858 10908
rect 1858 10852 1862 10908
rect 1798 10848 1862 10852
rect 4658 10908 4722 10912
rect 4658 10852 4662 10908
rect 4662 10852 4718 10908
rect 4718 10852 4722 10908
rect 4658 10848 4722 10852
rect 4738 10908 4802 10912
rect 4738 10852 4742 10908
rect 4742 10852 4798 10908
rect 4798 10852 4802 10908
rect 4738 10848 4802 10852
rect 4818 10908 4882 10912
rect 4818 10852 4822 10908
rect 4822 10852 4878 10908
rect 4878 10852 4882 10908
rect 4818 10848 4882 10852
rect 4898 10908 4962 10912
rect 4898 10852 4902 10908
rect 4902 10852 4958 10908
rect 4958 10852 4962 10908
rect 4898 10848 4962 10852
rect 7758 10908 7822 10912
rect 7758 10852 7762 10908
rect 7762 10852 7818 10908
rect 7818 10852 7822 10908
rect 7758 10848 7822 10852
rect 7838 10908 7902 10912
rect 7838 10852 7842 10908
rect 7842 10852 7898 10908
rect 7898 10852 7902 10908
rect 7838 10848 7902 10852
rect 7918 10908 7982 10912
rect 7918 10852 7922 10908
rect 7922 10852 7978 10908
rect 7978 10852 7982 10908
rect 7918 10848 7982 10852
rect 7998 10908 8062 10912
rect 7998 10852 8002 10908
rect 8002 10852 8058 10908
rect 8058 10852 8062 10908
rect 7998 10848 8062 10852
rect 10858 10908 10922 10912
rect 10858 10852 10862 10908
rect 10862 10852 10918 10908
rect 10918 10852 10922 10908
rect 10858 10848 10922 10852
rect 10938 10908 11002 10912
rect 10938 10852 10942 10908
rect 10942 10852 10998 10908
rect 10998 10852 11002 10908
rect 10938 10848 11002 10852
rect 11018 10908 11082 10912
rect 11018 10852 11022 10908
rect 11022 10852 11078 10908
rect 11078 10852 11082 10908
rect 11018 10848 11082 10852
rect 11098 10908 11162 10912
rect 11098 10852 11102 10908
rect 11102 10852 11158 10908
rect 11158 10852 11162 10908
rect 11098 10848 11162 10852
rect 13958 10908 14022 10912
rect 13958 10852 13962 10908
rect 13962 10852 14018 10908
rect 14018 10852 14022 10908
rect 13958 10848 14022 10852
rect 14038 10908 14102 10912
rect 14038 10852 14042 10908
rect 14042 10852 14098 10908
rect 14098 10852 14102 10908
rect 14038 10848 14102 10852
rect 14118 10908 14182 10912
rect 14118 10852 14122 10908
rect 14122 10852 14178 10908
rect 14178 10852 14182 10908
rect 14118 10848 14182 10852
rect 14198 10908 14262 10912
rect 14198 10852 14202 10908
rect 14202 10852 14258 10908
rect 14258 10852 14262 10908
rect 14198 10848 14262 10852
rect 17058 10908 17122 10912
rect 17058 10852 17062 10908
rect 17062 10852 17118 10908
rect 17118 10852 17122 10908
rect 17058 10848 17122 10852
rect 17138 10908 17202 10912
rect 17138 10852 17142 10908
rect 17142 10852 17198 10908
rect 17198 10852 17202 10908
rect 17138 10848 17202 10852
rect 17218 10908 17282 10912
rect 17218 10852 17222 10908
rect 17222 10852 17278 10908
rect 17278 10852 17282 10908
rect 17218 10848 17282 10852
rect 17298 10908 17362 10912
rect 17298 10852 17302 10908
rect 17302 10852 17358 10908
rect 17358 10852 17362 10908
rect 17298 10848 17362 10852
rect 3108 10364 3172 10368
rect 3108 10308 3112 10364
rect 3112 10308 3168 10364
rect 3168 10308 3172 10364
rect 3108 10304 3172 10308
rect 3188 10364 3252 10368
rect 3188 10308 3192 10364
rect 3192 10308 3248 10364
rect 3248 10308 3252 10364
rect 3188 10304 3252 10308
rect 3268 10364 3332 10368
rect 3268 10308 3272 10364
rect 3272 10308 3328 10364
rect 3328 10308 3332 10364
rect 3268 10304 3332 10308
rect 3348 10364 3412 10368
rect 3348 10308 3352 10364
rect 3352 10308 3408 10364
rect 3408 10308 3412 10364
rect 3348 10304 3412 10308
rect 6208 10364 6272 10368
rect 6208 10308 6212 10364
rect 6212 10308 6268 10364
rect 6268 10308 6272 10364
rect 6208 10304 6272 10308
rect 6288 10364 6352 10368
rect 6288 10308 6292 10364
rect 6292 10308 6348 10364
rect 6348 10308 6352 10364
rect 6288 10304 6352 10308
rect 6368 10364 6432 10368
rect 6368 10308 6372 10364
rect 6372 10308 6428 10364
rect 6428 10308 6432 10364
rect 6368 10304 6432 10308
rect 6448 10364 6512 10368
rect 6448 10308 6452 10364
rect 6452 10308 6508 10364
rect 6508 10308 6512 10364
rect 6448 10304 6512 10308
rect 9308 10364 9372 10368
rect 9308 10308 9312 10364
rect 9312 10308 9368 10364
rect 9368 10308 9372 10364
rect 9308 10304 9372 10308
rect 9388 10364 9452 10368
rect 9388 10308 9392 10364
rect 9392 10308 9448 10364
rect 9448 10308 9452 10364
rect 9388 10304 9452 10308
rect 9468 10364 9532 10368
rect 9468 10308 9472 10364
rect 9472 10308 9528 10364
rect 9528 10308 9532 10364
rect 9468 10304 9532 10308
rect 9548 10364 9612 10368
rect 9548 10308 9552 10364
rect 9552 10308 9608 10364
rect 9608 10308 9612 10364
rect 9548 10304 9612 10308
rect 12408 10364 12472 10368
rect 12408 10308 12412 10364
rect 12412 10308 12468 10364
rect 12468 10308 12472 10364
rect 12408 10304 12472 10308
rect 12488 10364 12552 10368
rect 12488 10308 12492 10364
rect 12492 10308 12548 10364
rect 12548 10308 12552 10364
rect 12488 10304 12552 10308
rect 12568 10364 12632 10368
rect 12568 10308 12572 10364
rect 12572 10308 12628 10364
rect 12628 10308 12632 10364
rect 12568 10304 12632 10308
rect 12648 10364 12712 10368
rect 12648 10308 12652 10364
rect 12652 10308 12708 10364
rect 12708 10308 12712 10364
rect 12648 10304 12712 10308
rect 15508 10364 15572 10368
rect 15508 10308 15512 10364
rect 15512 10308 15568 10364
rect 15568 10308 15572 10364
rect 15508 10304 15572 10308
rect 15588 10364 15652 10368
rect 15588 10308 15592 10364
rect 15592 10308 15648 10364
rect 15648 10308 15652 10364
rect 15588 10304 15652 10308
rect 15668 10364 15732 10368
rect 15668 10308 15672 10364
rect 15672 10308 15728 10364
rect 15728 10308 15732 10364
rect 15668 10304 15732 10308
rect 15748 10364 15812 10368
rect 15748 10308 15752 10364
rect 15752 10308 15808 10364
rect 15808 10308 15812 10364
rect 15748 10304 15812 10308
rect 18608 10364 18672 10368
rect 18608 10308 18612 10364
rect 18612 10308 18668 10364
rect 18668 10308 18672 10364
rect 18608 10304 18672 10308
rect 18688 10364 18752 10368
rect 18688 10308 18692 10364
rect 18692 10308 18748 10364
rect 18748 10308 18752 10364
rect 18688 10304 18752 10308
rect 18768 10364 18832 10368
rect 18768 10308 18772 10364
rect 18772 10308 18828 10364
rect 18828 10308 18832 10364
rect 18768 10304 18832 10308
rect 18848 10364 18912 10368
rect 18848 10308 18852 10364
rect 18852 10308 18908 10364
rect 18908 10308 18912 10364
rect 18848 10304 18912 10308
rect 1558 9820 1622 9824
rect 1558 9764 1562 9820
rect 1562 9764 1618 9820
rect 1618 9764 1622 9820
rect 1558 9760 1622 9764
rect 1638 9820 1702 9824
rect 1638 9764 1642 9820
rect 1642 9764 1698 9820
rect 1698 9764 1702 9820
rect 1638 9760 1702 9764
rect 1718 9820 1782 9824
rect 1718 9764 1722 9820
rect 1722 9764 1778 9820
rect 1778 9764 1782 9820
rect 1718 9760 1782 9764
rect 1798 9820 1862 9824
rect 1798 9764 1802 9820
rect 1802 9764 1858 9820
rect 1858 9764 1862 9820
rect 1798 9760 1862 9764
rect 4658 9820 4722 9824
rect 4658 9764 4662 9820
rect 4662 9764 4718 9820
rect 4718 9764 4722 9820
rect 4658 9760 4722 9764
rect 4738 9820 4802 9824
rect 4738 9764 4742 9820
rect 4742 9764 4798 9820
rect 4798 9764 4802 9820
rect 4738 9760 4802 9764
rect 4818 9820 4882 9824
rect 4818 9764 4822 9820
rect 4822 9764 4878 9820
rect 4878 9764 4882 9820
rect 4818 9760 4882 9764
rect 4898 9820 4962 9824
rect 4898 9764 4902 9820
rect 4902 9764 4958 9820
rect 4958 9764 4962 9820
rect 4898 9760 4962 9764
rect 7758 9820 7822 9824
rect 7758 9764 7762 9820
rect 7762 9764 7818 9820
rect 7818 9764 7822 9820
rect 7758 9760 7822 9764
rect 7838 9820 7902 9824
rect 7838 9764 7842 9820
rect 7842 9764 7898 9820
rect 7898 9764 7902 9820
rect 7838 9760 7902 9764
rect 7918 9820 7982 9824
rect 7918 9764 7922 9820
rect 7922 9764 7978 9820
rect 7978 9764 7982 9820
rect 7918 9760 7982 9764
rect 7998 9820 8062 9824
rect 7998 9764 8002 9820
rect 8002 9764 8058 9820
rect 8058 9764 8062 9820
rect 7998 9760 8062 9764
rect 10858 9820 10922 9824
rect 10858 9764 10862 9820
rect 10862 9764 10918 9820
rect 10918 9764 10922 9820
rect 10858 9760 10922 9764
rect 10938 9820 11002 9824
rect 10938 9764 10942 9820
rect 10942 9764 10998 9820
rect 10998 9764 11002 9820
rect 10938 9760 11002 9764
rect 11018 9820 11082 9824
rect 11018 9764 11022 9820
rect 11022 9764 11078 9820
rect 11078 9764 11082 9820
rect 11018 9760 11082 9764
rect 11098 9820 11162 9824
rect 11098 9764 11102 9820
rect 11102 9764 11158 9820
rect 11158 9764 11162 9820
rect 11098 9760 11162 9764
rect 13958 9820 14022 9824
rect 13958 9764 13962 9820
rect 13962 9764 14018 9820
rect 14018 9764 14022 9820
rect 13958 9760 14022 9764
rect 14038 9820 14102 9824
rect 14038 9764 14042 9820
rect 14042 9764 14098 9820
rect 14098 9764 14102 9820
rect 14038 9760 14102 9764
rect 14118 9820 14182 9824
rect 14118 9764 14122 9820
rect 14122 9764 14178 9820
rect 14178 9764 14182 9820
rect 14118 9760 14182 9764
rect 14198 9820 14262 9824
rect 14198 9764 14202 9820
rect 14202 9764 14258 9820
rect 14258 9764 14262 9820
rect 14198 9760 14262 9764
rect 17058 9820 17122 9824
rect 17058 9764 17062 9820
rect 17062 9764 17118 9820
rect 17118 9764 17122 9820
rect 17058 9760 17122 9764
rect 17138 9820 17202 9824
rect 17138 9764 17142 9820
rect 17142 9764 17198 9820
rect 17198 9764 17202 9820
rect 17138 9760 17202 9764
rect 17218 9820 17282 9824
rect 17218 9764 17222 9820
rect 17222 9764 17278 9820
rect 17278 9764 17282 9820
rect 17218 9760 17282 9764
rect 17298 9820 17362 9824
rect 17298 9764 17302 9820
rect 17302 9764 17358 9820
rect 17358 9764 17362 9820
rect 17298 9760 17362 9764
rect 3108 9276 3172 9280
rect 3108 9220 3112 9276
rect 3112 9220 3168 9276
rect 3168 9220 3172 9276
rect 3108 9216 3172 9220
rect 3188 9276 3252 9280
rect 3188 9220 3192 9276
rect 3192 9220 3248 9276
rect 3248 9220 3252 9276
rect 3188 9216 3252 9220
rect 3268 9276 3332 9280
rect 3268 9220 3272 9276
rect 3272 9220 3328 9276
rect 3328 9220 3332 9276
rect 3268 9216 3332 9220
rect 3348 9276 3412 9280
rect 3348 9220 3352 9276
rect 3352 9220 3408 9276
rect 3408 9220 3412 9276
rect 3348 9216 3412 9220
rect 6208 9276 6272 9280
rect 6208 9220 6212 9276
rect 6212 9220 6268 9276
rect 6268 9220 6272 9276
rect 6208 9216 6272 9220
rect 6288 9276 6352 9280
rect 6288 9220 6292 9276
rect 6292 9220 6348 9276
rect 6348 9220 6352 9276
rect 6288 9216 6352 9220
rect 6368 9276 6432 9280
rect 6368 9220 6372 9276
rect 6372 9220 6428 9276
rect 6428 9220 6432 9276
rect 6368 9216 6432 9220
rect 6448 9276 6512 9280
rect 6448 9220 6452 9276
rect 6452 9220 6508 9276
rect 6508 9220 6512 9276
rect 6448 9216 6512 9220
rect 9308 9276 9372 9280
rect 9308 9220 9312 9276
rect 9312 9220 9368 9276
rect 9368 9220 9372 9276
rect 9308 9216 9372 9220
rect 9388 9276 9452 9280
rect 9388 9220 9392 9276
rect 9392 9220 9448 9276
rect 9448 9220 9452 9276
rect 9388 9216 9452 9220
rect 9468 9276 9532 9280
rect 9468 9220 9472 9276
rect 9472 9220 9528 9276
rect 9528 9220 9532 9276
rect 9468 9216 9532 9220
rect 9548 9276 9612 9280
rect 9548 9220 9552 9276
rect 9552 9220 9608 9276
rect 9608 9220 9612 9276
rect 9548 9216 9612 9220
rect 12408 9276 12472 9280
rect 12408 9220 12412 9276
rect 12412 9220 12468 9276
rect 12468 9220 12472 9276
rect 12408 9216 12472 9220
rect 12488 9276 12552 9280
rect 12488 9220 12492 9276
rect 12492 9220 12548 9276
rect 12548 9220 12552 9276
rect 12488 9216 12552 9220
rect 12568 9276 12632 9280
rect 12568 9220 12572 9276
rect 12572 9220 12628 9276
rect 12628 9220 12632 9276
rect 12568 9216 12632 9220
rect 12648 9276 12712 9280
rect 12648 9220 12652 9276
rect 12652 9220 12708 9276
rect 12708 9220 12712 9276
rect 12648 9216 12712 9220
rect 15508 9276 15572 9280
rect 15508 9220 15512 9276
rect 15512 9220 15568 9276
rect 15568 9220 15572 9276
rect 15508 9216 15572 9220
rect 15588 9276 15652 9280
rect 15588 9220 15592 9276
rect 15592 9220 15648 9276
rect 15648 9220 15652 9276
rect 15588 9216 15652 9220
rect 15668 9276 15732 9280
rect 15668 9220 15672 9276
rect 15672 9220 15728 9276
rect 15728 9220 15732 9276
rect 15668 9216 15732 9220
rect 15748 9276 15812 9280
rect 15748 9220 15752 9276
rect 15752 9220 15808 9276
rect 15808 9220 15812 9276
rect 15748 9216 15812 9220
rect 18608 9276 18672 9280
rect 18608 9220 18612 9276
rect 18612 9220 18668 9276
rect 18668 9220 18672 9276
rect 18608 9216 18672 9220
rect 18688 9276 18752 9280
rect 18688 9220 18692 9276
rect 18692 9220 18748 9276
rect 18748 9220 18752 9276
rect 18688 9216 18752 9220
rect 18768 9276 18832 9280
rect 18768 9220 18772 9276
rect 18772 9220 18828 9276
rect 18828 9220 18832 9276
rect 18768 9216 18832 9220
rect 18848 9276 18912 9280
rect 18848 9220 18852 9276
rect 18852 9220 18908 9276
rect 18908 9220 18912 9276
rect 18848 9216 18912 9220
rect 1558 8732 1622 8736
rect 1558 8676 1562 8732
rect 1562 8676 1618 8732
rect 1618 8676 1622 8732
rect 1558 8672 1622 8676
rect 1638 8732 1702 8736
rect 1638 8676 1642 8732
rect 1642 8676 1698 8732
rect 1698 8676 1702 8732
rect 1638 8672 1702 8676
rect 1718 8732 1782 8736
rect 1718 8676 1722 8732
rect 1722 8676 1778 8732
rect 1778 8676 1782 8732
rect 1718 8672 1782 8676
rect 1798 8732 1862 8736
rect 1798 8676 1802 8732
rect 1802 8676 1858 8732
rect 1858 8676 1862 8732
rect 1798 8672 1862 8676
rect 4658 8732 4722 8736
rect 4658 8676 4662 8732
rect 4662 8676 4718 8732
rect 4718 8676 4722 8732
rect 4658 8672 4722 8676
rect 4738 8732 4802 8736
rect 4738 8676 4742 8732
rect 4742 8676 4798 8732
rect 4798 8676 4802 8732
rect 4738 8672 4802 8676
rect 4818 8732 4882 8736
rect 4818 8676 4822 8732
rect 4822 8676 4878 8732
rect 4878 8676 4882 8732
rect 4818 8672 4882 8676
rect 4898 8732 4962 8736
rect 4898 8676 4902 8732
rect 4902 8676 4958 8732
rect 4958 8676 4962 8732
rect 4898 8672 4962 8676
rect 7758 8732 7822 8736
rect 7758 8676 7762 8732
rect 7762 8676 7818 8732
rect 7818 8676 7822 8732
rect 7758 8672 7822 8676
rect 7838 8732 7902 8736
rect 7838 8676 7842 8732
rect 7842 8676 7898 8732
rect 7898 8676 7902 8732
rect 7838 8672 7902 8676
rect 7918 8732 7982 8736
rect 7918 8676 7922 8732
rect 7922 8676 7978 8732
rect 7978 8676 7982 8732
rect 7918 8672 7982 8676
rect 7998 8732 8062 8736
rect 7998 8676 8002 8732
rect 8002 8676 8058 8732
rect 8058 8676 8062 8732
rect 7998 8672 8062 8676
rect 10858 8732 10922 8736
rect 10858 8676 10862 8732
rect 10862 8676 10918 8732
rect 10918 8676 10922 8732
rect 10858 8672 10922 8676
rect 10938 8732 11002 8736
rect 10938 8676 10942 8732
rect 10942 8676 10998 8732
rect 10998 8676 11002 8732
rect 10938 8672 11002 8676
rect 11018 8732 11082 8736
rect 11018 8676 11022 8732
rect 11022 8676 11078 8732
rect 11078 8676 11082 8732
rect 11018 8672 11082 8676
rect 11098 8732 11162 8736
rect 11098 8676 11102 8732
rect 11102 8676 11158 8732
rect 11158 8676 11162 8732
rect 11098 8672 11162 8676
rect 13958 8732 14022 8736
rect 13958 8676 13962 8732
rect 13962 8676 14018 8732
rect 14018 8676 14022 8732
rect 13958 8672 14022 8676
rect 14038 8732 14102 8736
rect 14038 8676 14042 8732
rect 14042 8676 14098 8732
rect 14098 8676 14102 8732
rect 14038 8672 14102 8676
rect 14118 8732 14182 8736
rect 14118 8676 14122 8732
rect 14122 8676 14178 8732
rect 14178 8676 14182 8732
rect 14118 8672 14182 8676
rect 14198 8732 14262 8736
rect 14198 8676 14202 8732
rect 14202 8676 14258 8732
rect 14258 8676 14262 8732
rect 14198 8672 14262 8676
rect 17058 8732 17122 8736
rect 17058 8676 17062 8732
rect 17062 8676 17118 8732
rect 17118 8676 17122 8732
rect 17058 8672 17122 8676
rect 17138 8732 17202 8736
rect 17138 8676 17142 8732
rect 17142 8676 17198 8732
rect 17198 8676 17202 8732
rect 17138 8672 17202 8676
rect 17218 8732 17282 8736
rect 17218 8676 17222 8732
rect 17222 8676 17278 8732
rect 17278 8676 17282 8732
rect 17218 8672 17282 8676
rect 17298 8732 17362 8736
rect 17298 8676 17302 8732
rect 17302 8676 17358 8732
rect 17358 8676 17362 8732
rect 17298 8672 17362 8676
rect 3108 8188 3172 8192
rect 3108 8132 3112 8188
rect 3112 8132 3168 8188
rect 3168 8132 3172 8188
rect 3108 8128 3172 8132
rect 3188 8188 3252 8192
rect 3188 8132 3192 8188
rect 3192 8132 3248 8188
rect 3248 8132 3252 8188
rect 3188 8128 3252 8132
rect 3268 8188 3332 8192
rect 3268 8132 3272 8188
rect 3272 8132 3328 8188
rect 3328 8132 3332 8188
rect 3268 8128 3332 8132
rect 3348 8188 3412 8192
rect 3348 8132 3352 8188
rect 3352 8132 3408 8188
rect 3408 8132 3412 8188
rect 3348 8128 3412 8132
rect 6208 8188 6272 8192
rect 6208 8132 6212 8188
rect 6212 8132 6268 8188
rect 6268 8132 6272 8188
rect 6208 8128 6272 8132
rect 6288 8188 6352 8192
rect 6288 8132 6292 8188
rect 6292 8132 6348 8188
rect 6348 8132 6352 8188
rect 6288 8128 6352 8132
rect 6368 8188 6432 8192
rect 6368 8132 6372 8188
rect 6372 8132 6428 8188
rect 6428 8132 6432 8188
rect 6368 8128 6432 8132
rect 6448 8188 6512 8192
rect 6448 8132 6452 8188
rect 6452 8132 6508 8188
rect 6508 8132 6512 8188
rect 6448 8128 6512 8132
rect 9308 8188 9372 8192
rect 9308 8132 9312 8188
rect 9312 8132 9368 8188
rect 9368 8132 9372 8188
rect 9308 8128 9372 8132
rect 9388 8188 9452 8192
rect 9388 8132 9392 8188
rect 9392 8132 9448 8188
rect 9448 8132 9452 8188
rect 9388 8128 9452 8132
rect 9468 8188 9532 8192
rect 9468 8132 9472 8188
rect 9472 8132 9528 8188
rect 9528 8132 9532 8188
rect 9468 8128 9532 8132
rect 9548 8188 9612 8192
rect 9548 8132 9552 8188
rect 9552 8132 9608 8188
rect 9608 8132 9612 8188
rect 9548 8128 9612 8132
rect 12408 8188 12472 8192
rect 12408 8132 12412 8188
rect 12412 8132 12468 8188
rect 12468 8132 12472 8188
rect 12408 8128 12472 8132
rect 12488 8188 12552 8192
rect 12488 8132 12492 8188
rect 12492 8132 12548 8188
rect 12548 8132 12552 8188
rect 12488 8128 12552 8132
rect 12568 8188 12632 8192
rect 12568 8132 12572 8188
rect 12572 8132 12628 8188
rect 12628 8132 12632 8188
rect 12568 8128 12632 8132
rect 12648 8188 12712 8192
rect 12648 8132 12652 8188
rect 12652 8132 12708 8188
rect 12708 8132 12712 8188
rect 12648 8128 12712 8132
rect 15508 8188 15572 8192
rect 15508 8132 15512 8188
rect 15512 8132 15568 8188
rect 15568 8132 15572 8188
rect 15508 8128 15572 8132
rect 15588 8188 15652 8192
rect 15588 8132 15592 8188
rect 15592 8132 15648 8188
rect 15648 8132 15652 8188
rect 15588 8128 15652 8132
rect 15668 8188 15732 8192
rect 15668 8132 15672 8188
rect 15672 8132 15728 8188
rect 15728 8132 15732 8188
rect 15668 8128 15732 8132
rect 15748 8188 15812 8192
rect 15748 8132 15752 8188
rect 15752 8132 15808 8188
rect 15808 8132 15812 8188
rect 15748 8128 15812 8132
rect 18608 8188 18672 8192
rect 18608 8132 18612 8188
rect 18612 8132 18668 8188
rect 18668 8132 18672 8188
rect 18608 8128 18672 8132
rect 18688 8188 18752 8192
rect 18688 8132 18692 8188
rect 18692 8132 18748 8188
rect 18748 8132 18752 8188
rect 18688 8128 18752 8132
rect 18768 8188 18832 8192
rect 18768 8132 18772 8188
rect 18772 8132 18828 8188
rect 18828 8132 18832 8188
rect 18768 8128 18832 8132
rect 18848 8188 18912 8192
rect 18848 8132 18852 8188
rect 18852 8132 18908 8188
rect 18908 8132 18912 8188
rect 18848 8128 18912 8132
rect 1558 7644 1622 7648
rect 1558 7588 1562 7644
rect 1562 7588 1618 7644
rect 1618 7588 1622 7644
rect 1558 7584 1622 7588
rect 1638 7644 1702 7648
rect 1638 7588 1642 7644
rect 1642 7588 1698 7644
rect 1698 7588 1702 7644
rect 1638 7584 1702 7588
rect 1718 7644 1782 7648
rect 1718 7588 1722 7644
rect 1722 7588 1778 7644
rect 1778 7588 1782 7644
rect 1718 7584 1782 7588
rect 1798 7644 1862 7648
rect 1798 7588 1802 7644
rect 1802 7588 1858 7644
rect 1858 7588 1862 7644
rect 1798 7584 1862 7588
rect 4658 7644 4722 7648
rect 4658 7588 4662 7644
rect 4662 7588 4718 7644
rect 4718 7588 4722 7644
rect 4658 7584 4722 7588
rect 4738 7644 4802 7648
rect 4738 7588 4742 7644
rect 4742 7588 4798 7644
rect 4798 7588 4802 7644
rect 4738 7584 4802 7588
rect 4818 7644 4882 7648
rect 4818 7588 4822 7644
rect 4822 7588 4878 7644
rect 4878 7588 4882 7644
rect 4818 7584 4882 7588
rect 4898 7644 4962 7648
rect 4898 7588 4902 7644
rect 4902 7588 4958 7644
rect 4958 7588 4962 7644
rect 4898 7584 4962 7588
rect 7758 7644 7822 7648
rect 7758 7588 7762 7644
rect 7762 7588 7818 7644
rect 7818 7588 7822 7644
rect 7758 7584 7822 7588
rect 7838 7644 7902 7648
rect 7838 7588 7842 7644
rect 7842 7588 7898 7644
rect 7898 7588 7902 7644
rect 7838 7584 7902 7588
rect 7918 7644 7982 7648
rect 7918 7588 7922 7644
rect 7922 7588 7978 7644
rect 7978 7588 7982 7644
rect 7918 7584 7982 7588
rect 7998 7644 8062 7648
rect 7998 7588 8002 7644
rect 8002 7588 8058 7644
rect 8058 7588 8062 7644
rect 7998 7584 8062 7588
rect 10858 7644 10922 7648
rect 10858 7588 10862 7644
rect 10862 7588 10918 7644
rect 10918 7588 10922 7644
rect 10858 7584 10922 7588
rect 10938 7644 11002 7648
rect 10938 7588 10942 7644
rect 10942 7588 10998 7644
rect 10998 7588 11002 7644
rect 10938 7584 11002 7588
rect 11018 7644 11082 7648
rect 11018 7588 11022 7644
rect 11022 7588 11078 7644
rect 11078 7588 11082 7644
rect 11018 7584 11082 7588
rect 11098 7644 11162 7648
rect 11098 7588 11102 7644
rect 11102 7588 11158 7644
rect 11158 7588 11162 7644
rect 11098 7584 11162 7588
rect 13958 7644 14022 7648
rect 13958 7588 13962 7644
rect 13962 7588 14018 7644
rect 14018 7588 14022 7644
rect 13958 7584 14022 7588
rect 14038 7644 14102 7648
rect 14038 7588 14042 7644
rect 14042 7588 14098 7644
rect 14098 7588 14102 7644
rect 14038 7584 14102 7588
rect 14118 7644 14182 7648
rect 14118 7588 14122 7644
rect 14122 7588 14178 7644
rect 14178 7588 14182 7644
rect 14118 7584 14182 7588
rect 14198 7644 14262 7648
rect 14198 7588 14202 7644
rect 14202 7588 14258 7644
rect 14258 7588 14262 7644
rect 14198 7584 14262 7588
rect 17058 7644 17122 7648
rect 17058 7588 17062 7644
rect 17062 7588 17118 7644
rect 17118 7588 17122 7644
rect 17058 7584 17122 7588
rect 17138 7644 17202 7648
rect 17138 7588 17142 7644
rect 17142 7588 17198 7644
rect 17198 7588 17202 7644
rect 17138 7584 17202 7588
rect 17218 7644 17282 7648
rect 17218 7588 17222 7644
rect 17222 7588 17278 7644
rect 17278 7588 17282 7644
rect 17218 7584 17282 7588
rect 17298 7644 17362 7648
rect 17298 7588 17302 7644
rect 17302 7588 17358 7644
rect 17358 7588 17362 7644
rect 17298 7584 17362 7588
rect 3108 7100 3172 7104
rect 3108 7044 3112 7100
rect 3112 7044 3168 7100
rect 3168 7044 3172 7100
rect 3108 7040 3172 7044
rect 3188 7100 3252 7104
rect 3188 7044 3192 7100
rect 3192 7044 3248 7100
rect 3248 7044 3252 7100
rect 3188 7040 3252 7044
rect 3268 7100 3332 7104
rect 3268 7044 3272 7100
rect 3272 7044 3328 7100
rect 3328 7044 3332 7100
rect 3268 7040 3332 7044
rect 3348 7100 3412 7104
rect 3348 7044 3352 7100
rect 3352 7044 3408 7100
rect 3408 7044 3412 7100
rect 3348 7040 3412 7044
rect 6208 7100 6272 7104
rect 6208 7044 6212 7100
rect 6212 7044 6268 7100
rect 6268 7044 6272 7100
rect 6208 7040 6272 7044
rect 6288 7100 6352 7104
rect 6288 7044 6292 7100
rect 6292 7044 6348 7100
rect 6348 7044 6352 7100
rect 6288 7040 6352 7044
rect 6368 7100 6432 7104
rect 6368 7044 6372 7100
rect 6372 7044 6428 7100
rect 6428 7044 6432 7100
rect 6368 7040 6432 7044
rect 6448 7100 6512 7104
rect 6448 7044 6452 7100
rect 6452 7044 6508 7100
rect 6508 7044 6512 7100
rect 6448 7040 6512 7044
rect 9308 7100 9372 7104
rect 9308 7044 9312 7100
rect 9312 7044 9368 7100
rect 9368 7044 9372 7100
rect 9308 7040 9372 7044
rect 9388 7100 9452 7104
rect 9388 7044 9392 7100
rect 9392 7044 9448 7100
rect 9448 7044 9452 7100
rect 9388 7040 9452 7044
rect 9468 7100 9532 7104
rect 9468 7044 9472 7100
rect 9472 7044 9528 7100
rect 9528 7044 9532 7100
rect 9468 7040 9532 7044
rect 9548 7100 9612 7104
rect 9548 7044 9552 7100
rect 9552 7044 9608 7100
rect 9608 7044 9612 7100
rect 9548 7040 9612 7044
rect 12408 7100 12472 7104
rect 12408 7044 12412 7100
rect 12412 7044 12468 7100
rect 12468 7044 12472 7100
rect 12408 7040 12472 7044
rect 12488 7100 12552 7104
rect 12488 7044 12492 7100
rect 12492 7044 12548 7100
rect 12548 7044 12552 7100
rect 12488 7040 12552 7044
rect 12568 7100 12632 7104
rect 12568 7044 12572 7100
rect 12572 7044 12628 7100
rect 12628 7044 12632 7100
rect 12568 7040 12632 7044
rect 12648 7100 12712 7104
rect 12648 7044 12652 7100
rect 12652 7044 12708 7100
rect 12708 7044 12712 7100
rect 12648 7040 12712 7044
rect 15508 7100 15572 7104
rect 15508 7044 15512 7100
rect 15512 7044 15568 7100
rect 15568 7044 15572 7100
rect 15508 7040 15572 7044
rect 15588 7100 15652 7104
rect 15588 7044 15592 7100
rect 15592 7044 15648 7100
rect 15648 7044 15652 7100
rect 15588 7040 15652 7044
rect 15668 7100 15732 7104
rect 15668 7044 15672 7100
rect 15672 7044 15728 7100
rect 15728 7044 15732 7100
rect 15668 7040 15732 7044
rect 15748 7100 15812 7104
rect 15748 7044 15752 7100
rect 15752 7044 15808 7100
rect 15808 7044 15812 7100
rect 15748 7040 15812 7044
rect 18608 7100 18672 7104
rect 18608 7044 18612 7100
rect 18612 7044 18668 7100
rect 18668 7044 18672 7100
rect 18608 7040 18672 7044
rect 18688 7100 18752 7104
rect 18688 7044 18692 7100
rect 18692 7044 18748 7100
rect 18748 7044 18752 7100
rect 18688 7040 18752 7044
rect 18768 7100 18832 7104
rect 18768 7044 18772 7100
rect 18772 7044 18828 7100
rect 18828 7044 18832 7100
rect 18768 7040 18832 7044
rect 18848 7100 18912 7104
rect 18848 7044 18852 7100
rect 18852 7044 18908 7100
rect 18908 7044 18912 7100
rect 18848 7040 18912 7044
rect 1558 6556 1622 6560
rect 1558 6500 1562 6556
rect 1562 6500 1618 6556
rect 1618 6500 1622 6556
rect 1558 6496 1622 6500
rect 1638 6556 1702 6560
rect 1638 6500 1642 6556
rect 1642 6500 1698 6556
rect 1698 6500 1702 6556
rect 1638 6496 1702 6500
rect 1718 6556 1782 6560
rect 1718 6500 1722 6556
rect 1722 6500 1778 6556
rect 1778 6500 1782 6556
rect 1718 6496 1782 6500
rect 1798 6556 1862 6560
rect 1798 6500 1802 6556
rect 1802 6500 1858 6556
rect 1858 6500 1862 6556
rect 1798 6496 1862 6500
rect 4658 6556 4722 6560
rect 4658 6500 4662 6556
rect 4662 6500 4718 6556
rect 4718 6500 4722 6556
rect 4658 6496 4722 6500
rect 4738 6556 4802 6560
rect 4738 6500 4742 6556
rect 4742 6500 4798 6556
rect 4798 6500 4802 6556
rect 4738 6496 4802 6500
rect 4818 6556 4882 6560
rect 4818 6500 4822 6556
rect 4822 6500 4878 6556
rect 4878 6500 4882 6556
rect 4818 6496 4882 6500
rect 4898 6556 4962 6560
rect 4898 6500 4902 6556
rect 4902 6500 4958 6556
rect 4958 6500 4962 6556
rect 4898 6496 4962 6500
rect 7758 6556 7822 6560
rect 7758 6500 7762 6556
rect 7762 6500 7818 6556
rect 7818 6500 7822 6556
rect 7758 6496 7822 6500
rect 7838 6556 7902 6560
rect 7838 6500 7842 6556
rect 7842 6500 7898 6556
rect 7898 6500 7902 6556
rect 7838 6496 7902 6500
rect 7918 6556 7982 6560
rect 7918 6500 7922 6556
rect 7922 6500 7978 6556
rect 7978 6500 7982 6556
rect 7918 6496 7982 6500
rect 7998 6556 8062 6560
rect 7998 6500 8002 6556
rect 8002 6500 8058 6556
rect 8058 6500 8062 6556
rect 7998 6496 8062 6500
rect 10858 6556 10922 6560
rect 10858 6500 10862 6556
rect 10862 6500 10918 6556
rect 10918 6500 10922 6556
rect 10858 6496 10922 6500
rect 10938 6556 11002 6560
rect 10938 6500 10942 6556
rect 10942 6500 10998 6556
rect 10998 6500 11002 6556
rect 10938 6496 11002 6500
rect 11018 6556 11082 6560
rect 11018 6500 11022 6556
rect 11022 6500 11078 6556
rect 11078 6500 11082 6556
rect 11018 6496 11082 6500
rect 11098 6556 11162 6560
rect 11098 6500 11102 6556
rect 11102 6500 11158 6556
rect 11158 6500 11162 6556
rect 11098 6496 11162 6500
rect 13958 6556 14022 6560
rect 13958 6500 13962 6556
rect 13962 6500 14018 6556
rect 14018 6500 14022 6556
rect 13958 6496 14022 6500
rect 14038 6556 14102 6560
rect 14038 6500 14042 6556
rect 14042 6500 14098 6556
rect 14098 6500 14102 6556
rect 14038 6496 14102 6500
rect 14118 6556 14182 6560
rect 14118 6500 14122 6556
rect 14122 6500 14178 6556
rect 14178 6500 14182 6556
rect 14118 6496 14182 6500
rect 14198 6556 14262 6560
rect 14198 6500 14202 6556
rect 14202 6500 14258 6556
rect 14258 6500 14262 6556
rect 14198 6496 14262 6500
rect 17058 6556 17122 6560
rect 17058 6500 17062 6556
rect 17062 6500 17118 6556
rect 17118 6500 17122 6556
rect 17058 6496 17122 6500
rect 17138 6556 17202 6560
rect 17138 6500 17142 6556
rect 17142 6500 17198 6556
rect 17198 6500 17202 6556
rect 17138 6496 17202 6500
rect 17218 6556 17282 6560
rect 17218 6500 17222 6556
rect 17222 6500 17278 6556
rect 17278 6500 17282 6556
rect 17218 6496 17282 6500
rect 17298 6556 17362 6560
rect 17298 6500 17302 6556
rect 17302 6500 17358 6556
rect 17358 6500 17362 6556
rect 17298 6496 17362 6500
rect 3108 6012 3172 6016
rect 3108 5956 3112 6012
rect 3112 5956 3168 6012
rect 3168 5956 3172 6012
rect 3108 5952 3172 5956
rect 3188 6012 3252 6016
rect 3188 5956 3192 6012
rect 3192 5956 3248 6012
rect 3248 5956 3252 6012
rect 3188 5952 3252 5956
rect 3268 6012 3332 6016
rect 3268 5956 3272 6012
rect 3272 5956 3328 6012
rect 3328 5956 3332 6012
rect 3268 5952 3332 5956
rect 3348 6012 3412 6016
rect 3348 5956 3352 6012
rect 3352 5956 3408 6012
rect 3408 5956 3412 6012
rect 3348 5952 3412 5956
rect 6208 6012 6272 6016
rect 6208 5956 6212 6012
rect 6212 5956 6268 6012
rect 6268 5956 6272 6012
rect 6208 5952 6272 5956
rect 6288 6012 6352 6016
rect 6288 5956 6292 6012
rect 6292 5956 6348 6012
rect 6348 5956 6352 6012
rect 6288 5952 6352 5956
rect 6368 6012 6432 6016
rect 6368 5956 6372 6012
rect 6372 5956 6428 6012
rect 6428 5956 6432 6012
rect 6368 5952 6432 5956
rect 6448 6012 6512 6016
rect 6448 5956 6452 6012
rect 6452 5956 6508 6012
rect 6508 5956 6512 6012
rect 6448 5952 6512 5956
rect 9308 6012 9372 6016
rect 9308 5956 9312 6012
rect 9312 5956 9368 6012
rect 9368 5956 9372 6012
rect 9308 5952 9372 5956
rect 9388 6012 9452 6016
rect 9388 5956 9392 6012
rect 9392 5956 9448 6012
rect 9448 5956 9452 6012
rect 9388 5952 9452 5956
rect 9468 6012 9532 6016
rect 9468 5956 9472 6012
rect 9472 5956 9528 6012
rect 9528 5956 9532 6012
rect 9468 5952 9532 5956
rect 9548 6012 9612 6016
rect 9548 5956 9552 6012
rect 9552 5956 9608 6012
rect 9608 5956 9612 6012
rect 9548 5952 9612 5956
rect 12408 6012 12472 6016
rect 12408 5956 12412 6012
rect 12412 5956 12468 6012
rect 12468 5956 12472 6012
rect 12408 5952 12472 5956
rect 12488 6012 12552 6016
rect 12488 5956 12492 6012
rect 12492 5956 12548 6012
rect 12548 5956 12552 6012
rect 12488 5952 12552 5956
rect 12568 6012 12632 6016
rect 12568 5956 12572 6012
rect 12572 5956 12628 6012
rect 12628 5956 12632 6012
rect 12568 5952 12632 5956
rect 12648 6012 12712 6016
rect 12648 5956 12652 6012
rect 12652 5956 12708 6012
rect 12708 5956 12712 6012
rect 12648 5952 12712 5956
rect 15508 6012 15572 6016
rect 15508 5956 15512 6012
rect 15512 5956 15568 6012
rect 15568 5956 15572 6012
rect 15508 5952 15572 5956
rect 15588 6012 15652 6016
rect 15588 5956 15592 6012
rect 15592 5956 15648 6012
rect 15648 5956 15652 6012
rect 15588 5952 15652 5956
rect 15668 6012 15732 6016
rect 15668 5956 15672 6012
rect 15672 5956 15728 6012
rect 15728 5956 15732 6012
rect 15668 5952 15732 5956
rect 15748 6012 15812 6016
rect 15748 5956 15752 6012
rect 15752 5956 15808 6012
rect 15808 5956 15812 6012
rect 15748 5952 15812 5956
rect 18608 6012 18672 6016
rect 18608 5956 18612 6012
rect 18612 5956 18668 6012
rect 18668 5956 18672 6012
rect 18608 5952 18672 5956
rect 18688 6012 18752 6016
rect 18688 5956 18692 6012
rect 18692 5956 18748 6012
rect 18748 5956 18752 6012
rect 18688 5952 18752 5956
rect 18768 6012 18832 6016
rect 18768 5956 18772 6012
rect 18772 5956 18828 6012
rect 18828 5956 18832 6012
rect 18768 5952 18832 5956
rect 18848 6012 18912 6016
rect 18848 5956 18852 6012
rect 18852 5956 18908 6012
rect 18908 5956 18912 6012
rect 18848 5952 18912 5956
rect 1558 5468 1622 5472
rect 1558 5412 1562 5468
rect 1562 5412 1618 5468
rect 1618 5412 1622 5468
rect 1558 5408 1622 5412
rect 1638 5468 1702 5472
rect 1638 5412 1642 5468
rect 1642 5412 1698 5468
rect 1698 5412 1702 5468
rect 1638 5408 1702 5412
rect 1718 5468 1782 5472
rect 1718 5412 1722 5468
rect 1722 5412 1778 5468
rect 1778 5412 1782 5468
rect 1718 5408 1782 5412
rect 1798 5468 1862 5472
rect 1798 5412 1802 5468
rect 1802 5412 1858 5468
rect 1858 5412 1862 5468
rect 1798 5408 1862 5412
rect 4658 5468 4722 5472
rect 4658 5412 4662 5468
rect 4662 5412 4718 5468
rect 4718 5412 4722 5468
rect 4658 5408 4722 5412
rect 4738 5468 4802 5472
rect 4738 5412 4742 5468
rect 4742 5412 4798 5468
rect 4798 5412 4802 5468
rect 4738 5408 4802 5412
rect 4818 5468 4882 5472
rect 4818 5412 4822 5468
rect 4822 5412 4878 5468
rect 4878 5412 4882 5468
rect 4818 5408 4882 5412
rect 4898 5468 4962 5472
rect 4898 5412 4902 5468
rect 4902 5412 4958 5468
rect 4958 5412 4962 5468
rect 4898 5408 4962 5412
rect 7758 5468 7822 5472
rect 7758 5412 7762 5468
rect 7762 5412 7818 5468
rect 7818 5412 7822 5468
rect 7758 5408 7822 5412
rect 7838 5468 7902 5472
rect 7838 5412 7842 5468
rect 7842 5412 7898 5468
rect 7898 5412 7902 5468
rect 7838 5408 7902 5412
rect 7918 5468 7982 5472
rect 7918 5412 7922 5468
rect 7922 5412 7978 5468
rect 7978 5412 7982 5468
rect 7918 5408 7982 5412
rect 7998 5468 8062 5472
rect 7998 5412 8002 5468
rect 8002 5412 8058 5468
rect 8058 5412 8062 5468
rect 7998 5408 8062 5412
rect 10858 5468 10922 5472
rect 10858 5412 10862 5468
rect 10862 5412 10918 5468
rect 10918 5412 10922 5468
rect 10858 5408 10922 5412
rect 10938 5468 11002 5472
rect 10938 5412 10942 5468
rect 10942 5412 10998 5468
rect 10998 5412 11002 5468
rect 10938 5408 11002 5412
rect 11018 5468 11082 5472
rect 11018 5412 11022 5468
rect 11022 5412 11078 5468
rect 11078 5412 11082 5468
rect 11018 5408 11082 5412
rect 11098 5468 11162 5472
rect 11098 5412 11102 5468
rect 11102 5412 11158 5468
rect 11158 5412 11162 5468
rect 11098 5408 11162 5412
rect 13958 5468 14022 5472
rect 13958 5412 13962 5468
rect 13962 5412 14018 5468
rect 14018 5412 14022 5468
rect 13958 5408 14022 5412
rect 14038 5468 14102 5472
rect 14038 5412 14042 5468
rect 14042 5412 14098 5468
rect 14098 5412 14102 5468
rect 14038 5408 14102 5412
rect 14118 5468 14182 5472
rect 14118 5412 14122 5468
rect 14122 5412 14178 5468
rect 14178 5412 14182 5468
rect 14118 5408 14182 5412
rect 14198 5468 14262 5472
rect 14198 5412 14202 5468
rect 14202 5412 14258 5468
rect 14258 5412 14262 5468
rect 14198 5408 14262 5412
rect 17058 5468 17122 5472
rect 17058 5412 17062 5468
rect 17062 5412 17118 5468
rect 17118 5412 17122 5468
rect 17058 5408 17122 5412
rect 17138 5468 17202 5472
rect 17138 5412 17142 5468
rect 17142 5412 17198 5468
rect 17198 5412 17202 5468
rect 17138 5408 17202 5412
rect 17218 5468 17282 5472
rect 17218 5412 17222 5468
rect 17222 5412 17278 5468
rect 17278 5412 17282 5468
rect 17218 5408 17282 5412
rect 17298 5468 17362 5472
rect 17298 5412 17302 5468
rect 17302 5412 17358 5468
rect 17358 5412 17362 5468
rect 17298 5408 17362 5412
rect 3108 4924 3172 4928
rect 3108 4868 3112 4924
rect 3112 4868 3168 4924
rect 3168 4868 3172 4924
rect 3108 4864 3172 4868
rect 3188 4924 3252 4928
rect 3188 4868 3192 4924
rect 3192 4868 3248 4924
rect 3248 4868 3252 4924
rect 3188 4864 3252 4868
rect 3268 4924 3332 4928
rect 3268 4868 3272 4924
rect 3272 4868 3328 4924
rect 3328 4868 3332 4924
rect 3268 4864 3332 4868
rect 3348 4924 3412 4928
rect 3348 4868 3352 4924
rect 3352 4868 3408 4924
rect 3408 4868 3412 4924
rect 3348 4864 3412 4868
rect 6208 4924 6272 4928
rect 6208 4868 6212 4924
rect 6212 4868 6268 4924
rect 6268 4868 6272 4924
rect 6208 4864 6272 4868
rect 6288 4924 6352 4928
rect 6288 4868 6292 4924
rect 6292 4868 6348 4924
rect 6348 4868 6352 4924
rect 6288 4864 6352 4868
rect 6368 4924 6432 4928
rect 6368 4868 6372 4924
rect 6372 4868 6428 4924
rect 6428 4868 6432 4924
rect 6368 4864 6432 4868
rect 6448 4924 6512 4928
rect 6448 4868 6452 4924
rect 6452 4868 6508 4924
rect 6508 4868 6512 4924
rect 6448 4864 6512 4868
rect 9308 4924 9372 4928
rect 9308 4868 9312 4924
rect 9312 4868 9368 4924
rect 9368 4868 9372 4924
rect 9308 4864 9372 4868
rect 9388 4924 9452 4928
rect 9388 4868 9392 4924
rect 9392 4868 9448 4924
rect 9448 4868 9452 4924
rect 9388 4864 9452 4868
rect 9468 4924 9532 4928
rect 9468 4868 9472 4924
rect 9472 4868 9528 4924
rect 9528 4868 9532 4924
rect 9468 4864 9532 4868
rect 9548 4924 9612 4928
rect 9548 4868 9552 4924
rect 9552 4868 9608 4924
rect 9608 4868 9612 4924
rect 9548 4864 9612 4868
rect 12408 4924 12472 4928
rect 12408 4868 12412 4924
rect 12412 4868 12468 4924
rect 12468 4868 12472 4924
rect 12408 4864 12472 4868
rect 12488 4924 12552 4928
rect 12488 4868 12492 4924
rect 12492 4868 12548 4924
rect 12548 4868 12552 4924
rect 12488 4864 12552 4868
rect 12568 4924 12632 4928
rect 12568 4868 12572 4924
rect 12572 4868 12628 4924
rect 12628 4868 12632 4924
rect 12568 4864 12632 4868
rect 12648 4924 12712 4928
rect 12648 4868 12652 4924
rect 12652 4868 12708 4924
rect 12708 4868 12712 4924
rect 12648 4864 12712 4868
rect 15508 4924 15572 4928
rect 15508 4868 15512 4924
rect 15512 4868 15568 4924
rect 15568 4868 15572 4924
rect 15508 4864 15572 4868
rect 15588 4924 15652 4928
rect 15588 4868 15592 4924
rect 15592 4868 15648 4924
rect 15648 4868 15652 4924
rect 15588 4864 15652 4868
rect 15668 4924 15732 4928
rect 15668 4868 15672 4924
rect 15672 4868 15728 4924
rect 15728 4868 15732 4924
rect 15668 4864 15732 4868
rect 15748 4924 15812 4928
rect 15748 4868 15752 4924
rect 15752 4868 15808 4924
rect 15808 4868 15812 4924
rect 15748 4864 15812 4868
rect 18608 4924 18672 4928
rect 18608 4868 18612 4924
rect 18612 4868 18668 4924
rect 18668 4868 18672 4924
rect 18608 4864 18672 4868
rect 18688 4924 18752 4928
rect 18688 4868 18692 4924
rect 18692 4868 18748 4924
rect 18748 4868 18752 4924
rect 18688 4864 18752 4868
rect 18768 4924 18832 4928
rect 18768 4868 18772 4924
rect 18772 4868 18828 4924
rect 18828 4868 18832 4924
rect 18768 4864 18832 4868
rect 18848 4924 18912 4928
rect 18848 4868 18852 4924
rect 18852 4868 18908 4924
rect 18908 4868 18912 4924
rect 18848 4864 18912 4868
rect 1558 4380 1622 4384
rect 1558 4324 1562 4380
rect 1562 4324 1618 4380
rect 1618 4324 1622 4380
rect 1558 4320 1622 4324
rect 1638 4380 1702 4384
rect 1638 4324 1642 4380
rect 1642 4324 1698 4380
rect 1698 4324 1702 4380
rect 1638 4320 1702 4324
rect 1718 4380 1782 4384
rect 1718 4324 1722 4380
rect 1722 4324 1778 4380
rect 1778 4324 1782 4380
rect 1718 4320 1782 4324
rect 1798 4380 1862 4384
rect 1798 4324 1802 4380
rect 1802 4324 1858 4380
rect 1858 4324 1862 4380
rect 1798 4320 1862 4324
rect 4658 4380 4722 4384
rect 4658 4324 4662 4380
rect 4662 4324 4718 4380
rect 4718 4324 4722 4380
rect 4658 4320 4722 4324
rect 4738 4380 4802 4384
rect 4738 4324 4742 4380
rect 4742 4324 4798 4380
rect 4798 4324 4802 4380
rect 4738 4320 4802 4324
rect 4818 4380 4882 4384
rect 4818 4324 4822 4380
rect 4822 4324 4878 4380
rect 4878 4324 4882 4380
rect 4818 4320 4882 4324
rect 4898 4380 4962 4384
rect 4898 4324 4902 4380
rect 4902 4324 4958 4380
rect 4958 4324 4962 4380
rect 4898 4320 4962 4324
rect 7758 4380 7822 4384
rect 7758 4324 7762 4380
rect 7762 4324 7818 4380
rect 7818 4324 7822 4380
rect 7758 4320 7822 4324
rect 7838 4380 7902 4384
rect 7838 4324 7842 4380
rect 7842 4324 7898 4380
rect 7898 4324 7902 4380
rect 7838 4320 7902 4324
rect 7918 4380 7982 4384
rect 7918 4324 7922 4380
rect 7922 4324 7978 4380
rect 7978 4324 7982 4380
rect 7918 4320 7982 4324
rect 7998 4380 8062 4384
rect 7998 4324 8002 4380
rect 8002 4324 8058 4380
rect 8058 4324 8062 4380
rect 7998 4320 8062 4324
rect 10858 4380 10922 4384
rect 10858 4324 10862 4380
rect 10862 4324 10918 4380
rect 10918 4324 10922 4380
rect 10858 4320 10922 4324
rect 10938 4380 11002 4384
rect 10938 4324 10942 4380
rect 10942 4324 10998 4380
rect 10998 4324 11002 4380
rect 10938 4320 11002 4324
rect 11018 4380 11082 4384
rect 11018 4324 11022 4380
rect 11022 4324 11078 4380
rect 11078 4324 11082 4380
rect 11018 4320 11082 4324
rect 11098 4380 11162 4384
rect 11098 4324 11102 4380
rect 11102 4324 11158 4380
rect 11158 4324 11162 4380
rect 11098 4320 11162 4324
rect 13958 4380 14022 4384
rect 13958 4324 13962 4380
rect 13962 4324 14018 4380
rect 14018 4324 14022 4380
rect 13958 4320 14022 4324
rect 14038 4380 14102 4384
rect 14038 4324 14042 4380
rect 14042 4324 14098 4380
rect 14098 4324 14102 4380
rect 14038 4320 14102 4324
rect 14118 4380 14182 4384
rect 14118 4324 14122 4380
rect 14122 4324 14178 4380
rect 14178 4324 14182 4380
rect 14118 4320 14182 4324
rect 14198 4380 14262 4384
rect 14198 4324 14202 4380
rect 14202 4324 14258 4380
rect 14258 4324 14262 4380
rect 14198 4320 14262 4324
rect 17058 4380 17122 4384
rect 17058 4324 17062 4380
rect 17062 4324 17118 4380
rect 17118 4324 17122 4380
rect 17058 4320 17122 4324
rect 17138 4380 17202 4384
rect 17138 4324 17142 4380
rect 17142 4324 17198 4380
rect 17198 4324 17202 4380
rect 17138 4320 17202 4324
rect 17218 4380 17282 4384
rect 17218 4324 17222 4380
rect 17222 4324 17278 4380
rect 17278 4324 17282 4380
rect 17218 4320 17282 4324
rect 17298 4380 17362 4384
rect 17298 4324 17302 4380
rect 17302 4324 17358 4380
rect 17358 4324 17362 4380
rect 17298 4320 17362 4324
rect 3108 3836 3172 3840
rect 3108 3780 3112 3836
rect 3112 3780 3168 3836
rect 3168 3780 3172 3836
rect 3108 3776 3172 3780
rect 3188 3836 3252 3840
rect 3188 3780 3192 3836
rect 3192 3780 3248 3836
rect 3248 3780 3252 3836
rect 3188 3776 3252 3780
rect 3268 3836 3332 3840
rect 3268 3780 3272 3836
rect 3272 3780 3328 3836
rect 3328 3780 3332 3836
rect 3268 3776 3332 3780
rect 3348 3836 3412 3840
rect 3348 3780 3352 3836
rect 3352 3780 3408 3836
rect 3408 3780 3412 3836
rect 3348 3776 3412 3780
rect 6208 3836 6272 3840
rect 6208 3780 6212 3836
rect 6212 3780 6268 3836
rect 6268 3780 6272 3836
rect 6208 3776 6272 3780
rect 6288 3836 6352 3840
rect 6288 3780 6292 3836
rect 6292 3780 6348 3836
rect 6348 3780 6352 3836
rect 6288 3776 6352 3780
rect 6368 3836 6432 3840
rect 6368 3780 6372 3836
rect 6372 3780 6428 3836
rect 6428 3780 6432 3836
rect 6368 3776 6432 3780
rect 6448 3836 6512 3840
rect 6448 3780 6452 3836
rect 6452 3780 6508 3836
rect 6508 3780 6512 3836
rect 6448 3776 6512 3780
rect 9308 3836 9372 3840
rect 9308 3780 9312 3836
rect 9312 3780 9368 3836
rect 9368 3780 9372 3836
rect 9308 3776 9372 3780
rect 9388 3836 9452 3840
rect 9388 3780 9392 3836
rect 9392 3780 9448 3836
rect 9448 3780 9452 3836
rect 9388 3776 9452 3780
rect 9468 3836 9532 3840
rect 9468 3780 9472 3836
rect 9472 3780 9528 3836
rect 9528 3780 9532 3836
rect 9468 3776 9532 3780
rect 9548 3836 9612 3840
rect 9548 3780 9552 3836
rect 9552 3780 9608 3836
rect 9608 3780 9612 3836
rect 9548 3776 9612 3780
rect 12408 3836 12472 3840
rect 12408 3780 12412 3836
rect 12412 3780 12468 3836
rect 12468 3780 12472 3836
rect 12408 3776 12472 3780
rect 12488 3836 12552 3840
rect 12488 3780 12492 3836
rect 12492 3780 12548 3836
rect 12548 3780 12552 3836
rect 12488 3776 12552 3780
rect 12568 3836 12632 3840
rect 12568 3780 12572 3836
rect 12572 3780 12628 3836
rect 12628 3780 12632 3836
rect 12568 3776 12632 3780
rect 12648 3836 12712 3840
rect 12648 3780 12652 3836
rect 12652 3780 12708 3836
rect 12708 3780 12712 3836
rect 12648 3776 12712 3780
rect 15508 3836 15572 3840
rect 15508 3780 15512 3836
rect 15512 3780 15568 3836
rect 15568 3780 15572 3836
rect 15508 3776 15572 3780
rect 15588 3836 15652 3840
rect 15588 3780 15592 3836
rect 15592 3780 15648 3836
rect 15648 3780 15652 3836
rect 15588 3776 15652 3780
rect 15668 3836 15732 3840
rect 15668 3780 15672 3836
rect 15672 3780 15728 3836
rect 15728 3780 15732 3836
rect 15668 3776 15732 3780
rect 15748 3836 15812 3840
rect 15748 3780 15752 3836
rect 15752 3780 15808 3836
rect 15808 3780 15812 3836
rect 15748 3776 15812 3780
rect 18608 3836 18672 3840
rect 18608 3780 18612 3836
rect 18612 3780 18668 3836
rect 18668 3780 18672 3836
rect 18608 3776 18672 3780
rect 18688 3836 18752 3840
rect 18688 3780 18692 3836
rect 18692 3780 18748 3836
rect 18748 3780 18752 3836
rect 18688 3776 18752 3780
rect 18768 3836 18832 3840
rect 18768 3780 18772 3836
rect 18772 3780 18828 3836
rect 18828 3780 18832 3836
rect 18768 3776 18832 3780
rect 18848 3836 18912 3840
rect 18848 3780 18852 3836
rect 18852 3780 18908 3836
rect 18908 3780 18912 3836
rect 18848 3776 18912 3780
rect 1558 3292 1622 3296
rect 1558 3236 1562 3292
rect 1562 3236 1618 3292
rect 1618 3236 1622 3292
rect 1558 3232 1622 3236
rect 1638 3292 1702 3296
rect 1638 3236 1642 3292
rect 1642 3236 1698 3292
rect 1698 3236 1702 3292
rect 1638 3232 1702 3236
rect 1718 3292 1782 3296
rect 1718 3236 1722 3292
rect 1722 3236 1778 3292
rect 1778 3236 1782 3292
rect 1718 3232 1782 3236
rect 1798 3292 1862 3296
rect 1798 3236 1802 3292
rect 1802 3236 1858 3292
rect 1858 3236 1862 3292
rect 1798 3232 1862 3236
rect 4658 3292 4722 3296
rect 4658 3236 4662 3292
rect 4662 3236 4718 3292
rect 4718 3236 4722 3292
rect 4658 3232 4722 3236
rect 4738 3292 4802 3296
rect 4738 3236 4742 3292
rect 4742 3236 4798 3292
rect 4798 3236 4802 3292
rect 4738 3232 4802 3236
rect 4818 3292 4882 3296
rect 4818 3236 4822 3292
rect 4822 3236 4878 3292
rect 4878 3236 4882 3292
rect 4818 3232 4882 3236
rect 4898 3292 4962 3296
rect 4898 3236 4902 3292
rect 4902 3236 4958 3292
rect 4958 3236 4962 3292
rect 4898 3232 4962 3236
rect 7758 3292 7822 3296
rect 7758 3236 7762 3292
rect 7762 3236 7818 3292
rect 7818 3236 7822 3292
rect 7758 3232 7822 3236
rect 7838 3292 7902 3296
rect 7838 3236 7842 3292
rect 7842 3236 7898 3292
rect 7898 3236 7902 3292
rect 7838 3232 7902 3236
rect 7918 3292 7982 3296
rect 7918 3236 7922 3292
rect 7922 3236 7978 3292
rect 7978 3236 7982 3292
rect 7918 3232 7982 3236
rect 7998 3292 8062 3296
rect 7998 3236 8002 3292
rect 8002 3236 8058 3292
rect 8058 3236 8062 3292
rect 7998 3232 8062 3236
rect 10858 3292 10922 3296
rect 10858 3236 10862 3292
rect 10862 3236 10918 3292
rect 10918 3236 10922 3292
rect 10858 3232 10922 3236
rect 10938 3292 11002 3296
rect 10938 3236 10942 3292
rect 10942 3236 10998 3292
rect 10998 3236 11002 3292
rect 10938 3232 11002 3236
rect 11018 3292 11082 3296
rect 11018 3236 11022 3292
rect 11022 3236 11078 3292
rect 11078 3236 11082 3292
rect 11018 3232 11082 3236
rect 11098 3292 11162 3296
rect 11098 3236 11102 3292
rect 11102 3236 11158 3292
rect 11158 3236 11162 3292
rect 11098 3232 11162 3236
rect 13958 3292 14022 3296
rect 13958 3236 13962 3292
rect 13962 3236 14018 3292
rect 14018 3236 14022 3292
rect 13958 3232 14022 3236
rect 14038 3292 14102 3296
rect 14038 3236 14042 3292
rect 14042 3236 14098 3292
rect 14098 3236 14102 3292
rect 14038 3232 14102 3236
rect 14118 3292 14182 3296
rect 14118 3236 14122 3292
rect 14122 3236 14178 3292
rect 14178 3236 14182 3292
rect 14118 3232 14182 3236
rect 14198 3292 14262 3296
rect 14198 3236 14202 3292
rect 14202 3236 14258 3292
rect 14258 3236 14262 3292
rect 14198 3232 14262 3236
rect 17058 3292 17122 3296
rect 17058 3236 17062 3292
rect 17062 3236 17118 3292
rect 17118 3236 17122 3292
rect 17058 3232 17122 3236
rect 17138 3292 17202 3296
rect 17138 3236 17142 3292
rect 17142 3236 17198 3292
rect 17198 3236 17202 3292
rect 17138 3232 17202 3236
rect 17218 3292 17282 3296
rect 17218 3236 17222 3292
rect 17222 3236 17278 3292
rect 17278 3236 17282 3292
rect 17218 3232 17282 3236
rect 17298 3292 17362 3296
rect 17298 3236 17302 3292
rect 17302 3236 17358 3292
rect 17358 3236 17362 3292
rect 17298 3232 17362 3236
rect 3108 2748 3172 2752
rect 3108 2692 3112 2748
rect 3112 2692 3168 2748
rect 3168 2692 3172 2748
rect 3108 2688 3172 2692
rect 3188 2748 3252 2752
rect 3188 2692 3192 2748
rect 3192 2692 3248 2748
rect 3248 2692 3252 2748
rect 3188 2688 3252 2692
rect 3268 2748 3332 2752
rect 3268 2692 3272 2748
rect 3272 2692 3328 2748
rect 3328 2692 3332 2748
rect 3268 2688 3332 2692
rect 3348 2748 3412 2752
rect 3348 2692 3352 2748
rect 3352 2692 3408 2748
rect 3408 2692 3412 2748
rect 3348 2688 3412 2692
rect 6208 2748 6272 2752
rect 6208 2692 6212 2748
rect 6212 2692 6268 2748
rect 6268 2692 6272 2748
rect 6208 2688 6272 2692
rect 6288 2748 6352 2752
rect 6288 2692 6292 2748
rect 6292 2692 6348 2748
rect 6348 2692 6352 2748
rect 6288 2688 6352 2692
rect 6368 2748 6432 2752
rect 6368 2692 6372 2748
rect 6372 2692 6428 2748
rect 6428 2692 6432 2748
rect 6368 2688 6432 2692
rect 6448 2748 6512 2752
rect 6448 2692 6452 2748
rect 6452 2692 6508 2748
rect 6508 2692 6512 2748
rect 6448 2688 6512 2692
rect 9308 2748 9372 2752
rect 9308 2692 9312 2748
rect 9312 2692 9368 2748
rect 9368 2692 9372 2748
rect 9308 2688 9372 2692
rect 9388 2748 9452 2752
rect 9388 2692 9392 2748
rect 9392 2692 9448 2748
rect 9448 2692 9452 2748
rect 9388 2688 9452 2692
rect 9468 2748 9532 2752
rect 9468 2692 9472 2748
rect 9472 2692 9528 2748
rect 9528 2692 9532 2748
rect 9468 2688 9532 2692
rect 9548 2748 9612 2752
rect 9548 2692 9552 2748
rect 9552 2692 9608 2748
rect 9608 2692 9612 2748
rect 9548 2688 9612 2692
rect 12408 2748 12472 2752
rect 12408 2692 12412 2748
rect 12412 2692 12468 2748
rect 12468 2692 12472 2748
rect 12408 2688 12472 2692
rect 12488 2748 12552 2752
rect 12488 2692 12492 2748
rect 12492 2692 12548 2748
rect 12548 2692 12552 2748
rect 12488 2688 12552 2692
rect 12568 2748 12632 2752
rect 12568 2692 12572 2748
rect 12572 2692 12628 2748
rect 12628 2692 12632 2748
rect 12568 2688 12632 2692
rect 12648 2748 12712 2752
rect 12648 2692 12652 2748
rect 12652 2692 12708 2748
rect 12708 2692 12712 2748
rect 12648 2688 12712 2692
rect 15508 2748 15572 2752
rect 15508 2692 15512 2748
rect 15512 2692 15568 2748
rect 15568 2692 15572 2748
rect 15508 2688 15572 2692
rect 15588 2748 15652 2752
rect 15588 2692 15592 2748
rect 15592 2692 15648 2748
rect 15648 2692 15652 2748
rect 15588 2688 15652 2692
rect 15668 2748 15732 2752
rect 15668 2692 15672 2748
rect 15672 2692 15728 2748
rect 15728 2692 15732 2748
rect 15668 2688 15732 2692
rect 15748 2748 15812 2752
rect 15748 2692 15752 2748
rect 15752 2692 15808 2748
rect 15808 2692 15812 2748
rect 15748 2688 15812 2692
rect 18608 2748 18672 2752
rect 18608 2692 18612 2748
rect 18612 2692 18668 2748
rect 18668 2692 18672 2748
rect 18608 2688 18672 2692
rect 18688 2748 18752 2752
rect 18688 2692 18692 2748
rect 18692 2692 18748 2748
rect 18748 2692 18752 2748
rect 18688 2688 18752 2692
rect 18768 2748 18832 2752
rect 18768 2692 18772 2748
rect 18772 2692 18828 2748
rect 18828 2692 18832 2748
rect 18768 2688 18832 2692
rect 18848 2748 18912 2752
rect 18848 2692 18852 2748
rect 18852 2692 18908 2748
rect 18908 2692 18912 2748
rect 18848 2688 18912 2692
rect 1558 2204 1622 2208
rect 1558 2148 1562 2204
rect 1562 2148 1618 2204
rect 1618 2148 1622 2204
rect 1558 2144 1622 2148
rect 1638 2204 1702 2208
rect 1638 2148 1642 2204
rect 1642 2148 1698 2204
rect 1698 2148 1702 2204
rect 1638 2144 1702 2148
rect 1718 2204 1782 2208
rect 1718 2148 1722 2204
rect 1722 2148 1778 2204
rect 1778 2148 1782 2204
rect 1718 2144 1782 2148
rect 1798 2204 1862 2208
rect 1798 2148 1802 2204
rect 1802 2148 1858 2204
rect 1858 2148 1862 2204
rect 1798 2144 1862 2148
rect 4658 2204 4722 2208
rect 4658 2148 4662 2204
rect 4662 2148 4718 2204
rect 4718 2148 4722 2204
rect 4658 2144 4722 2148
rect 4738 2204 4802 2208
rect 4738 2148 4742 2204
rect 4742 2148 4798 2204
rect 4798 2148 4802 2204
rect 4738 2144 4802 2148
rect 4818 2204 4882 2208
rect 4818 2148 4822 2204
rect 4822 2148 4878 2204
rect 4878 2148 4882 2204
rect 4818 2144 4882 2148
rect 4898 2204 4962 2208
rect 4898 2148 4902 2204
rect 4902 2148 4958 2204
rect 4958 2148 4962 2204
rect 4898 2144 4962 2148
rect 7758 2204 7822 2208
rect 7758 2148 7762 2204
rect 7762 2148 7818 2204
rect 7818 2148 7822 2204
rect 7758 2144 7822 2148
rect 7838 2204 7902 2208
rect 7838 2148 7842 2204
rect 7842 2148 7898 2204
rect 7898 2148 7902 2204
rect 7838 2144 7902 2148
rect 7918 2204 7982 2208
rect 7918 2148 7922 2204
rect 7922 2148 7978 2204
rect 7978 2148 7982 2204
rect 7918 2144 7982 2148
rect 7998 2204 8062 2208
rect 7998 2148 8002 2204
rect 8002 2148 8058 2204
rect 8058 2148 8062 2204
rect 7998 2144 8062 2148
rect 10858 2204 10922 2208
rect 10858 2148 10862 2204
rect 10862 2148 10918 2204
rect 10918 2148 10922 2204
rect 10858 2144 10922 2148
rect 10938 2204 11002 2208
rect 10938 2148 10942 2204
rect 10942 2148 10998 2204
rect 10998 2148 11002 2204
rect 10938 2144 11002 2148
rect 11018 2204 11082 2208
rect 11018 2148 11022 2204
rect 11022 2148 11078 2204
rect 11078 2148 11082 2204
rect 11018 2144 11082 2148
rect 11098 2204 11162 2208
rect 11098 2148 11102 2204
rect 11102 2148 11158 2204
rect 11158 2148 11162 2204
rect 11098 2144 11162 2148
rect 13958 2204 14022 2208
rect 13958 2148 13962 2204
rect 13962 2148 14018 2204
rect 14018 2148 14022 2204
rect 13958 2144 14022 2148
rect 14038 2204 14102 2208
rect 14038 2148 14042 2204
rect 14042 2148 14098 2204
rect 14098 2148 14102 2204
rect 14038 2144 14102 2148
rect 14118 2204 14182 2208
rect 14118 2148 14122 2204
rect 14122 2148 14178 2204
rect 14178 2148 14182 2204
rect 14118 2144 14182 2148
rect 14198 2204 14262 2208
rect 14198 2148 14202 2204
rect 14202 2148 14258 2204
rect 14258 2148 14262 2204
rect 14198 2144 14262 2148
rect 17058 2204 17122 2208
rect 17058 2148 17062 2204
rect 17062 2148 17118 2204
rect 17118 2148 17122 2204
rect 17058 2144 17122 2148
rect 17138 2204 17202 2208
rect 17138 2148 17142 2204
rect 17142 2148 17198 2204
rect 17198 2148 17202 2204
rect 17138 2144 17202 2148
rect 17218 2204 17282 2208
rect 17218 2148 17222 2204
rect 17222 2148 17278 2204
rect 17278 2148 17282 2204
rect 17218 2144 17282 2148
rect 17298 2204 17362 2208
rect 17298 2148 17302 2204
rect 17302 2148 17358 2204
rect 17358 2148 17362 2204
rect 17298 2144 17362 2148
rect 3108 1660 3172 1664
rect 3108 1604 3112 1660
rect 3112 1604 3168 1660
rect 3168 1604 3172 1660
rect 3108 1600 3172 1604
rect 3188 1660 3252 1664
rect 3188 1604 3192 1660
rect 3192 1604 3248 1660
rect 3248 1604 3252 1660
rect 3188 1600 3252 1604
rect 3268 1660 3332 1664
rect 3268 1604 3272 1660
rect 3272 1604 3328 1660
rect 3328 1604 3332 1660
rect 3268 1600 3332 1604
rect 3348 1660 3412 1664
rect 3348 1604 3352 1660
rect 3352 1604 3408 1660
rect 3408 1604 3412 1660
rect 3348 1600 3412 1604
rect 6208 1660 6272 1664
rect 6208 1604 6212 1660
rect 6212 1604 6268 1660
rect 6268 1604 6272 1660
rect 6208 1600 6272 1604
rect 6288 1660 6352 1664
rect 6288 1604 6292 1660
rect 6292 1604 6348 1660
rect 6348 1604 6352 1660
rect 6288 1600 6352 1604
rect 6368 1660 6432 1664
rect 6368 1604 6372 1660
rect 6372 1604 6428 1660
rect 6428 1604 6432 1660
rect 6368 1600 6432 1604
rect 6448 1660 6512 1664
rect 6448 1604 6452 1660
rect 6452 1604 6508 1660
rect 6508 1604 6512 1660
rect 6448 1600 6512 1604
rect 9308 1660 9372 1664
rect 9308 1604 9312 1660
rect 9312 1604 9368 1660
rect 9368 1604 9372 1660
rect 9308 1600 9372 1604
rect 9388 1660 9452 1664
rect 9388 1604 9392 1660
rect 9392 1604 9448 1660
rect 9448 1604 9452 1660
rect 9388 1600 9452 1604
rect 9468 1660 9532 1664
rect 9468 1604 9472 1660
rect 9472 1604 9528 1660
rect 9528 1604 9532 1660
rect 9468 1600 9532 1604
rect 9548 1660 9612 1664
rect 9548 1604 9552 1660
rect 9552 1604 9608 1660
rect 9608 1604 9612 1660
rect 9548 1600 9612 1604
rect 12408 1660 12472 1664
rect 12408 1604 12412 1660
rect 12412 1604 12468 1660
rect 12468 1604 12472 1660
rect 12408 1600 12472 1604
rect 12488 1660 12552 1664
rect 12488 1604 12492 1660
rect 12492 1604 12548 1660
rect 12548 1604 12552 1660
rect 12488 1600 12552 1604
rect 12568 1660 12632 1664
rect 12568 1604 12572 1660
rect 12572 1604 12628 1660
rect 12628 1604 12632 1660
rect 12568 1600 12632 1604
rect 12648 1660 12712 1664
rect 12648 1604 12652 1660
rect 12652 1604 12708 1660
rect 12708 1604 12712 1660
rect 12648 1600 12712 1604
rect 15508 1660 15572 1664
rect 15508 1604 15512 1660
rect 15512 1604 15568 1660
rect 15568 1604 15572 1660
rect 15508 1600 15572 1604
rect 15588 1660 15652 1664
rect 15588 1604 15592 1660
rect 15592 1604 15648 1660
rect 15648 1604 15652 1660
rect 15588 1600 15652 1604
rect 15668 1660 15732 1664
rect 15668 1604 15672 1660
rect 15672 1604 15728 1660
rect 15728 1604 15732 1660
rect 15668 1600 15732 1604
rect 15748 1660 15812 1664
rect 15748 1604 15752 1660
rect 15752 1604 15808 1660
rect 15808 1604 15812 1660
rect 15748 1600 15812 1604
rect 18608 1660 18672 1664
rect 18608 1604 18612 1660
rect 18612 1604 18668 1660
rect 18668 1604 18672 1660
rect 18608 1600 18672 1604
rect 18688 1660 18752 1664
rect 18688 1604 18692 1660
rect 18692 1604 18748 1660
rect 18748 1604 18752 1660
rect 18688 1600 18752 1604
rect 18768 1660 18832 1664
rect 18768 1604 18772 1660
rect 18772 1604 18828 1660
rect 18828 1604 18832 1660
rect 18768 1600 18832 1604
rect 18848 1660 18912 1664
rect 18848 1604 18852 1660
rect 18852 1604 18908 1660
rect 18908 1604 18912 1660
rect 18848 1600 18912 1604
rect 1558 1116 1622 1120
rect 1558 1060 1562 1116
rect 1562 1060 1618 1116
rect 1618 1060 1622 1116
rect 1558 1056 1622 1060
rect 1638 1116 1702 1120
rect 1638 1060 1642 1116
rect 1642 1060 1698 1116
rect 1698 1060 1702 1116
rect 1638 1056 1702 1060
rect 1718 1116 1782 1120
rect 1718 1060 1722 1116
rect 1722 1060 1778 1116
rect 1778 1060 1782 1116
rect 1718 1056 1782 1060
rect 1798 1116 1862 1120
rect 1798 1060 1802 1116
rect 1802 1060 1858 1116
rect 1858 1060 1862 1116
rect 1798 1056 1862 1060
rect 4658 1116 4722 1120
rect 4658 1060 4662 1116
rect 4662 1060 4718 1116
rect 4718 1060 4722 1116
rect 4658 1056 4722 1060
rect 4738 1116 4802 1120
rect 4738 1060 4742 1116
rect 4742 1060 4798 1116
rect 4798 1060 4802 1116
rect 4738 1056 4802 1060
rect 4818 1116 4882 1120
rect 4818 1060 4822 1116
rect 4822 1060 4878 1116
rect 4878 1060 4882 1116
rect 4818 1056 4882 1060
rect 4898 1116 4962 1120
rect 4898 1060 4902 1116
rect 4902 1060 4958 1116
rect 4958 1060 4962 1116
rect 4898 1056 4962 1060
rect 7758 1116 7822 1120
rect 7758 1060 7762 1116
rect 7762 1060 7818 1116
rect 7818 1060 7822 1116
rect 7758 1056 7822 1060
rect 7838 1116 7902 1120
rect 7838 1060 7842 1116
rect 7842 1060 7898 1116
rect 7898 1060 7902 1116
rect 7838 1056 7902 1060
rect 7918 1116 7982 1120
rect 7918 1060 7922 1116
rect 7922 1060 7978 1116
rect 7978 1060 7982 1116
rect 7918 1056 7982 1060
rect 7998 1116 8062 1120
rect 7998 1060 8002 1116
rect 8002 1060 8058 1116
rect 8058 1060 8062 1116
rect 7998 1056 8062 1060
rect 10858 1116 10922 1120
rect 10858 1060 10862 1116
rect 10862 1060 10918 1116
rect 10918 1060 10922 1116
rect 10858 1056 10922 1060
rect 10938 1116 11002 1120
rect 10938 1060 10942 1116
rect 10942 1060 10998 1116
rect 10998 1060 11002 1116
rect 10938 1056 11002 1060
rect 11018 1116 11082 1120
rect 11018 1060 11022 1116
rect 11022 1060 11078 1116
rect 11078 1060 11082 1116
rect 11018 1056 11082 1060
rect 11098 1116 11162 1120
rect 11098 1060 11102 1116
rect 11102 1060 11158 1116
rect 11158 1060 11162 1116
rect 11098 1056 11162 1060
rect 13958 1116 14022 1120
rect 13958 1060 13962 1116
rect 13962 1060 14018 1116
rect 14018 1060 14022 1116
rect 13958 1056 14022 1060
rect 14038 1116 14102 1120
rect 14038 1060 14042 1116
rect 14042 1060 14098 1116
rect 14098 1060 14102 1116
rect 14038 1056 14102 1060
rect 14118 1116 14182 1120
rect 14118 1060 14122 1116
rect 14122 1060 14178 1116
rect 14178 1060 14182 1116
rect 14118 1056 14182 1060
rect 14198 1116 14262 1120
rect 14198 1060 14202 1116
rect 14202 1060 14258 1116
rect 14258 1060 14262 1116
rect 14198 1056 14262 1060
rect 17058 1116 17122 1120
rect 17058 1060 17062 1116
rect 17062 1060 17118 1116
rect 17118 1060 17122 1116
rect 17058 1056 17122 1060
rect 17138 1116 17202 1120
rect 17138 1060 17142 1116
rect 17142 1060 17198 1116
rect 17198 1060 17202 1116
rect 17138 1056 17202 1060
rect 17218 1116 17282 1120
rect 17218 1060 17222 1116
rect 17222 1060 17278 1116
rect 17278 1060 17282 1116
rect 17218 1056 17282 1060
rect 17298 1116 17362 1120
rect 17298 1060 17302 1116
rect 17302 1060 17358 1116
rect 17358 1060 17362 1116
rect 17298 1056 17362 1060
rect 3108 572 3172 576
rect 3108 516 3112 572
rect 3112 516 3168 572
rect 3168 516 3172 572
rect 3108 512 3172 516
rect 3188 572 3252 576
rect 3188 516 3192 572
rect 3192 516 3248 572
rect 3248 516 3252 572
rect 3188 512 3252 516
rect 3268 572 3332 576
rect 3268 516 3272 572
rect 3272 516 3328 572
rect 3328 516 3332 572
rect 3268 512 3332 516
rect 3348 572 3412 576
rect 3348 516 3352 572
rect 3352 516 3408 572
rect 3408 516 3412 572
rect 3348 512 3412 516
rect 6208 572 6272 576
rect 6208 516 6212 572
rect 6212 516 6268 572
rect 6268 516 6272 572
rect 6208 512 6272 516
rect 6288 572 6352 576
rect 6288 516 6292 572
rect 6292 516 6348 572
rect 6348 516 6352 572
rect 6288 512 6352 516
rect 6368 572 6432 576
rect 6368 516 6372 572
rect 6372 516 6428 572
rect 6428 516 6432 572
rect 6368 512 6432 516
rect 6448 572 6512 576
rect 6448 516 6452 572
rect 6452 516 6508 572
rect 6508 516 6512 572
rect 6448 512 6512 516
rect 9308 572 9372 576
rect 9308 516 9312 572
rect 9312 516 9368 572
rect 9368 516 9372 572
rect 9308 512 9372 516
rect 9388 572 9452 576
rect 9388 516 9392 572
rect 9392 516 9448 572
rect 9448 516 9452 572
rect 9388 512 9452 516
rect 9468 572 9532 576
rect 9468 516 9472 572
rect 9472 516 9528 572
rect 9528 516 9532 572
rect 9468 512 9532 516
rect 9548 572 9612 576
rect 9548 516 9552 572
rect 9552 516 9608 572
rect 9608 516 9612 572
rect 9548 512 9612 516
rect 12408 572 12472 576
rect 12408 516 12412 572
rect 12412 516 12468 572
rect 12468 516 12472 572
rect 12408 512 12472 516
rect 12488 572 12552 576
rect 12488 516 12492 572
rect 12492 516 12548 572
rect 12548 516 12552 572
rect 12488 512 12552 516
rect 12568 572 12632 576
rect 12568 516 12572 572
rect 12572 516 12628 572
rect 12628 516 12632 572
rect 12568 512 12632 516
rect 12648 572 12712 576
rect 12648 516 12652 572
rect 12652 516 12708 572
rect 12708 516 12712 572
rect 12648 512 12712 516
rect 15508 572 15572 576
rect 15508 516 15512 572
rect 15512 516 15568 572
rect 15568 516 15572 572
rect 15508 512 15572 516
rect 15588 572 15652 576
rect 15588 516 15592 572
rect 15592 516 15648 572
rect 15648 516 15652 572
rect 15588 512 15652 516
rect 15668 572 15732 576
rect 15668 516 15672 572
rect 15672 516 15728 572
rect 15728 516 15732 572
rect 15668 512 15732 516
rect 15748 572 15812 576
rect 15748 516 15752 572
rect 15752 516 15808 572
rect 15808 516 15812 572
rect 15748 512 15812 516
rect 18608 572 18672 576
rect 18608 516 18612 572
rect 18612 516 18668 572
rect 18668 516 18672 572
rect 18608 512 18672 516
rect 18688 572 18752 576
rect 18688 516 18692 572
rect 18692 516 18748 572
rect 18748 516 18752 572
rect 18688 512 18752 516
rect 18768 572 18832 576
rect 18768 516 18772 572
rect 18772 516 18828 572
rect 18828 516 18832 572
rect 18768 512 18832 516
rect 18848 572 18912 576
rect 18848 516 18852 572
rect 18852 516 18908 572
rect 18908 516 18912 572
rect 18848 512 18912 516
<< metal4 >>
rect 1550 18528 1870 18544
rect 1550 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1870 18528
rect 1550 17440 1870 18464
rect 1550 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1870 17440
rect 1550 16352 1870 17376
rect 1550 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1870 16352
rect 1550 15264 1870 16288
rect 1550 15200 1558 15264
rect 1622 15200 1638 15264
rect 1702 15200 1718 15264
rect 1782 15200 1798 15264
rect 1862 15200 1870 15264
rect 1550 14176 1870 15200
rect 1550 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1870 14176
rect 1550 13088 1870 14112
rect 1550 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1870 13088
rect 1550 12000 1870 13024
rect 1550 11936 1558 12000
rect 1622 11936 1638 12000
rect 1702 11936 1718 12000
rect 1782 11936 1798 12000
rect 1862 11936 1870 12000
rect 1550 10912 1870 11936
rect 1550 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1870 10912
rect 1550 9824 1870 10848
rect 1550 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1870 9824
rect 1550 8736 1870 9760
rect 1550 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1870 8736
rect 1550 7648 1870 8672
rect 1550 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1870 7648
rect 1550 6560 1870 7584
rect 1550 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1870 6560
rect 1550 5472 1870 6496
rect 1550 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1870 5472
rect 1550 4384 1870 5408
rect 1550 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1870 4384
rect 1550 3296 1870 4320
rect 1550 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1870 3296
rect 1550 2208 1870 3232
rect 1550 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1870 2208
rect 1550 1120 1870 2144
rect 1550 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1870 1120
rect 1550 496 1870 1056
rect 3100 17984 3420 18544
rect 3100 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3420 17984
rect 3100 16896 3420 17920
rect 3100 16832 3108 16896
rect 3172 16832 3188 16896
rect 3252 16832 3268 16896
rect 3332 16832 3348 16896
rect 3412 16832 3420 16896
rect 3100 15808 3420 16832
rect 3100 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3420 15808
rect 3100 14720 3420 15744
rect 3100 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3420 14720
rect 3100 13632 3420 14656
rect 3100 13568 3108 13632
rect 3172 13568 3188 13632
rect 3252 13568 3268 13632
rect 3332 13568 3348 13632
rect 3412 13568 3420 13632
rect 3100 12544 3420 13568
rect 3100 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3420 12544
rect 3100 11456 3420 12480
rect 3100 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3420 11456
rect 3100 10368 3420 11392
rect 3100 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3420 10368
rect 3100 9280 3420 10304
rect 3100 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3420 9280
rect 3100 8192 3420 9216
rect 3100 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3420 8192
rect 3100 7104 3420 8128
rect 3100 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3420 7104
rect 3100 6016 3420 7040
rect 3100 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3420 6016
rect 3100 4928 3420 5952
rect 3100 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3420 4928
rect 3100 3840 3420 4864
rect 3100 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3420 3840
rect 3100 2752 3420 3776
rect 3100 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3420 2752
rect 3100 1664 3420 2688
rect 3100 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3420 1664
rect 3100 576 3420 1600
rect 3100 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3420 576
rect 3100 496 3420 512
rect 4650 18528 4970 18544
rect 4650 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4970 18528
rect 4650 17440 4970 18464
rect 4650 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4970 17440
rect 4650 16352 4970 17376
rect 4650 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4970 16352
rect 4650 15264 4970 16288
rect 4650 15200 4658 15264
rect 4722 15200 4738 15264
rect 4802 15200 4818 15264
rect 4882 15200 4898 15264
rect 4962 15200 4970 15264
rect 4650 14176 4970 15200
rect 4650 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4970 14176
rect 4650 13088 4970 14112
rect 4650 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4970 13088
rect 4650 12000 4970 13024
rect 4650 11936 4658 12000
rect 4722 11936 4738 12000
rect 4802 11936 4818 12000
rect 4882 11936 4898 12000
rect 4962 11936 4970 12000
rect 4650 10912 4970 11936
rect 4650 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4970 10912
rect 4650 9824 4970 10848
rect 4650 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4970 9824
rect 4650 8736 4970 9760
rect 4650 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4970 8736
rect 4650 7648 4970 8672
rect 4650 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4970 7648
rect 4650 6560 4970 7584
rect 4650 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4970 6560
rect 4650 5472 4970 6496
rect 4650 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4970 5472
rect 4650 4384 4970 5408
rect 4650 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4970 4384
rect 4650 3296 4970 4320
rect 4650 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4970 3296
rect 4650 2208 4970 3232
rect 4650 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4970 2208
rect 4650 1120 4970 2144
rect 4650 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4970 1120
rect 4650 496 4970 1056
rect 6200 17984 6520 18544
rect 6200 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6520 17984
rect 6200 16896 6520 17920
rect 6200 16832 6208 16896
rect 6272 16832 6288 16896
rect 6352 16832 6368 16896
rect 6432 16832 6448 16896
rect 6512 16832 6520 16896
rect 6200 15808 6520 16832
rect 6200 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6520 15808
rect 6200 14720 6520 15744
rect 6200 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6520 14720
rect 6200 13632 6520 14656
rect 6200 13568 6208 13632
rect 6272 13568 6288 13632
rect 6352 13568 6368 13632
rect 6432 13568 6448 13632
rect 6512 13568 6520 13632
rect 6200 12544 6520 13568
rect 6200 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6520 12544
rect 6200 11456 6520 12480
rect 6200 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6520 11456
rect 6200 10368 6520 11392
rect 6200 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6520 10368
rect 6200 9280 6520 10304
rect 6200 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6520 9280
rect 6200 8192 6520 9216
rect 6200 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6520 8192
rect 6200 7104 6520 8128
rect 6200 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6520 7104
rect 6200 6016 6520 7040
rect 6200 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6520 6016
rect 6200 4928 6520 5952
rect 6200 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6520 4928
rect 6200 3840 6520 4864
rect 6200 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6520 3840
rect 6200 2752 6520 3776
rect 6200 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6520 2752
rect 6200 1664 6520 2688
rect 6200 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6520 1664
rect 6200 576 6520 1600
rect 6200 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6520 576
rect 6200 496 6520 512
rect 7750 18528 8070 18544
rect 7750 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8070 18528
rect 7750 17440 8070 18464
rect 7750 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8070 17440
rect 7750 16352 8070 17376
rect 7750 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8070 16352
rect 7750 15264 8070 16288
rect 7750 15200 7758 15264
rect 7822 15200 7838 15264
rect 7902 15200 7918 15264
rect 7982 15200 7998 15264
rect 8062 15200 8070 15264
rect 7750 14176 8070 15200
rect 7750 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8070 14176
rect 7750 13088 8070 14112
rect 7750 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8070 13088
rect 7750 12000 8070 13024
rect 7750 11936 7758 12000
rect 7822 11936 7838 12000
rect 7902 11936 7918 12000
rect 7982 11936 7998 12000
rect 8062 11936 8070 12000
rect 7750 10912 8070 11936
rect 7750 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8070 10912
rect 7750 9824 8070 10848
rect 7750 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8070 9824
rect 7750 8736 8070 9760
rect 7750 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8070 8736
rect 7750 7648 8070 8672
rect 7750 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8070 7648
rect 7750 6560 8070 7584
rect 7750 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8070 6560
rect 7750 5472 8070 6496
rect 7750 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8070 5472
rect 7750 4384 8070 5408
rect 7750 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8070 4384
rect 7750 3296 8070 4320
rect 7750 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8070 3296
rect 7750 2208 8070 3232
rect 7750 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8070 2208
rect 7750 1120 8070 2144
rect 7750 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8070 1120
rect 7750 496 8070 1056
rect 9300 17984 9620 18544
rect 9300 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9620 17984
rect 9300 16896 9620 17920
rect 9300 16832 9308 16896
rect 9372 16832 9388 16896
rect 9452 16832 9468 16896
rect 9532 16832 9548 16896
rect 9612 16832 9620 16896
rect 9300 15808 9620 16832
rect 9300 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9620 15808
rect 9300 14720 9620 15744
rect 9300 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9620 14720
rect 9300 13632 9620 14656
rect 9300 13568 9308 13632
rect 9372 13568 9388 13632
rect 9452 13568 9468 13632
rect 9532 13568 9548 13632
rect 9612 13568 9620 13632
rect 9300 12544 9620 13568
rect 9300 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9620 12544
rect 9300 11456 9620 12480
rect 9300 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9620 11456
rect 9300 10368 9620 11392
rect 9300 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9620 10368
rect 9300 9280 9620 10304
rect 9300 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9620 9280
rect 9300 8192 9620 9216
rect 9300 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9620 8192
rect 9300 7104 9620 8128
rect 9300 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9620 7104
rect 9300 6016 9620 7040
rect 9300 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9620 6016
rect 9300 4928 9620 5952
rect 9300 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9620 4928
rect 9300 3840 9620 4864
rect 9300 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9620 3840
rect 9300 2752 9620 3776
rect 9300 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9620 2752
rect 9300 1664 9620 2688
rect 9300 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9620 1664
rect 9300 576 9620 1600
rect 9300 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9620 576
rect 9300 496 9620 512
rect 10850 18528 11170 18544
rect 10850 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11170 18528
rect 10850 17440 11170 18464
rect 10850 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11170 17440
rect 10850 16352 11170 17376
rect 10850 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11170 16352
rect 10850 15264 11170 16288
rect 10850 15200 10858 15264
rect 10922 15200 10938 15264
rect 11002 15200 11018 15264
rect 11082 15200 11098 15264
rect 11162 15200 11170 15264
rect 10850 14176 11170 15200
rect 10850 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11170 14176
rect 10850 13088 11170 14112
rect 10850 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11170 13088
rect 10850 12000 11170 13024
rect 10850 11936 10858 12000
rect 10922 11936 10938 12000
rect 11002 11936 11018 12000
rect 11082 11936 11098 12000
rect 11162 11936 11170 12000
rect 10850 10912 11170 11936
rect 10850 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11170 10912
rect 10850 9824 11170 10848
rect 10850 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11170 9824
rect 10850 8736 11170 9760
rect 10850 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11170 8736
rect 10850 7648 11170 8672
rect 10850 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11170 7648
rect 10850 6560 11170 7584
rect 10850 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11170 6560
rect 10850 5472 11170 6496
rect 10850 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11170 5472
rect 10850 4384 11170 5408
rect 10850 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11170 4384
rect 10850 3296 11170 4320
rect 10850 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11170 3296
rect 10850 2208 11170 3232
rect 10850 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11170 2208
rect 10850 1120 11170 2144
rect 10850 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11170 1120
rect 10850 496 11170 1056
rect 12400 17984 12720 18544
rect 12400 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12720 17984
rect 12400 16896 12720 17920
rect 12400 16832 12408 16896
rect 12472 16832 12488 16896
rect 12552 16832 12568 16896
rect 12632 16832 12648 16896
rect 12712 16832 12720 16896
rect 12400 15808 12720 16832
rect 12400 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12720 15808
rect 12400 14720 12720 15744
rect 12400 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12720 14720
rect 12400 13632 12720 14656
rect 12400 13568 12408 13632
rect 12472 13568 12488 13632
rect 12552 13568 12568 13632
rect 12632 13568 12648 13632
rect 12712 13568 12720 13632
rect 12400 12544 12720 13568
rect 12400 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12720 12544
rect 12400 11456 12720 12480
rect 12400 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12720 11456
rect 12400 10368 12720 11392
rect 12400 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12720 10368
rect 12400 9280 12720 10304
rect 12400 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12720 9280
rect 12400 8192 12720 9216
rect 12400 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12720 8192
rect 12400 7104 12720 8128
rect 12400 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12720 7104
rect 12400 6016 12720 7040
rect 12400 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12720 6016
rect 12400 4928 12720 5952
rect 12400 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12720 4928
rect 12400 3840 12720 4864
rect 12400 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12720 3840
rect 12400 2752 12720 3776
rect 12400 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12720 2752
rect 12400 1664 12720 2688
rect 12400 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12720 1664
rect 12400 576 12720 1600
rect 12400 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12720 576
rect 12400 496 12720 512
rect 13950 18528 14270 18544
rect 13950 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14270 18528
rect 13950 17440 14270 18464
rect 13950 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14270 17440
rect 13950 16352 14270 17376
rect 13950 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14270 16352
rect 13950 15264 14270 16288
rect 13950 15200 13958 15264
rect 14022 15200 14038 15264
rect 14102 15200 14118 15264
rect 14182 15200 14198 15264
rect 14262 15200 14270 15264
rect 13950 14176 14270 15200
rect 13950 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14270 14176
rect 13950 13088 14270 14112
rect 13950 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14270 13088
rect 13950 12000 14270 13024
rect 13950 11936 13958 12000
rect 14022 11936 14038 12000
rect 14102 11936 14118 12000
rect 14182 11936 14198 12000
rect 14262 11936 14270 12000
rect 13950 10912 14270 11936
rect 13950 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14270 10912
rect 13950 9824 14270 10848
rect 13950 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14270 9824
rect 13950 8736 14270 9760
rect 13950 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14270 8736
rect 13950 7648 14270 8672
rect 13950 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14270 7648
rect 13950 6560 14270 7584
rect 13950 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14270 6560
rect 13950 5472 14270 6496
rect 13950 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14270 5472
rect 13950 4384 14270 5408
rect 13950 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14270 4384
rect 13950 3296 14270 4320
rect 13950 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14270 3296
rect 13950 2208 14270 3232
rect 13950 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14270 2208
rect 13950 1120 14270 2144
rect 13950 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14270 1120
rect 13950 496 14270 1056
rect 15500 17984 15820 18544
rect 15500 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15820 17984
rect 15500 16896 15820 17920
rect 15500 16832 15508 16896
rect 15572 16832 15588 16896
rect 15652 16832 15668 16896
rect 15732 16832 15748 16896
rect 15812 16832 15820 16896
rect 15500 15808 15820 16832
rect 15500 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15820 15808
rect 15500 14720 15820 15744
rect 15500 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15820 14720
rect 15500 13632 15820 14656
rect 15500 13568 15508 13632
rect 15572 13568 15588 13632
rect 15652 13568 15668 13632
rect 15732 13568 15748 13632
rect 15812 13568 15820 13632
rect 15500 12544 15820 13568
rect 15500 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15820 12544
rect 15500 11456 15820 12480
rect 15500 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15820 11456
rect 15500 10368 15820 11392
rect 15500 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15820 10368
rect 15500 9280 15820 10304
rect 15500 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15820 9280
rect 15500 8192 15820 9216
rect 15500 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15820 8192
rect 15500 7104 15820 8128
rect 15500 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15820 7104
rect 15500 6016 15820 7040
rect 15500 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15820 6016
rect 15500 4928 15820 5952
rect 15500 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15820 4928
rect 15500 3840 15820 4864
rect 15500 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15820 3840
rect 15500 2752 15820 3776
rect 15500 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15820 2752
rect 15500 1664 15820 2688
rect 15500 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15820 1664
rect 15500 576 15820 1600
rect 15500 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15820 576
rect 15500 496 15820 512
rect 17050 18528 17370 18544
rect 17050 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17370 18528
rect 17050 17440 17370 18464
rect 17050 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17370 17440
rect 17050 16352 17370 17376
rect 17050 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17370 16352
rect 17050 15264 17370 16288
rect 17050 15200 17058 15264
rect 17122 15200 17138 15264
rect 17202 15200 17218 15264
rect 17282 15200 17298 15264
rect 17362 15200 17370 15264
rect 17050 14176 17370 15200
rect 17050 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17370 14176
rect 17050 13088 17370 14112
rect 17050 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17370 13088
rect 17050 12000 17370 13024
rect 17050 11936 17058 12000
rect 17122 11936 17138 12000
rect 17202 11936 17218 12000
rect 17282 11936 17298 12000
rect 17362 11936 17370 12000
rect 17050 10912 17370 11936
rect 17050 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17370 10912
rect 17050 9824 17370 10848
rect 17050 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17370 9824
rect 17050 8736 17370 9760
rect 17050 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17370 8736
rect 17050 7648 17370 8672
rect 17050 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17370 7648
rect 17050 6560 17370 7584
rect 17050 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17370 6560
rect 17050 5472 17370 6496
rect 17050 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17370 5472
rect 17050 4384 17370 5408
rect 17050 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17370 4384
rect 17050 3296 17370 4320
rect 17050 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17370 3296
rect 17050 2208 17370 3232
rect 17050 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17370 2208
rect 17050 1120 17370 2144
rect 17050 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17370 1120
rect 17050 496 17370 1056
rect 18600 17984 18920 18544
rect 18600 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18920 17984
rect 18600 16896 18920 17920
rect 18600 16832 18608 16896
rect 18672 16832 18688 16896
rect 18752 16832 18768 16896
rect 18832 16832 18848 16896
rect 18912 16832 18920 16896
rect 18600 15808 18920 16832
rect 18600 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18920 15808
rect 18600 14720 18920 15744
rect 18600 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18920 14720
rect 18600 13632 18920 14656
rect 18600 13568 18608 13632
rect 18672 13568 18688 13632
rect 18752 13568 18768 13632
rect 18832 13568 18848 13632
rect 18912 13568 18920 13632
rect 18600 12544 18920 13568
rect 18600 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18920 12544
rect 18600 11456 18920 12480
rect 18600 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18920 11456
rect 18600 10368 18920 11392
rect 18600 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18920 10368
rect 18600 9280 18920 10304
rect 18600 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18920 9280
rect 18600 8192 18920 9216
rect 18600 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18920 8192
rect 18600 7104 18920 8128
rect 18600 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18920 7104
rect 18600 6016 18920 7040
rect 18600 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18920 6016
rect 18600 4928 18920 5952
rect 18600 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18920 4928
rect 18600 3840 18920 4864
rect 18600 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18920 3840
rect 18600 2752 18920 3776
rect 18600 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18920 2752
rect 18600 1664 18920 2688
rect 18600 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18920 1664
rect 18600 576 18920 1600
rect 18600 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18920 576
rect 18600 496 18920 512
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6348 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A1
timestamp 1673029049
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1673029049
transform -1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A1
timestamp 1673029049
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1673029049
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1
timestamp 1673029049
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1673029049
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1673029049
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A1
timestamp 1673029049
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1673029049
transform 1 0 14168 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A1
timestamp 1673029049
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1673029049
transform -1 0 18492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A1
timestamp 1673029049
transform -1 0 16100 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1673029049
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B
timestamp 1673029049
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A1
timestamp 1673029049
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2
timestamp 1673029049
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1673029049
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 1673029049
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__B
timestamp 1673029049
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A2
timestamp 1673029049
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1673029049
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1673029049
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A2
timestamp 1673029049
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1673029049
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1673029049
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__B
timestamp 1673029049
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1673029049
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__B
timestamp 1673029049
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__C
timestamp 1673029049
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__B1
timestamp 1673029049
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1673029049
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A2
timestamp 1673029049
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__B1
timestamp 1673029049
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1673029049
transform -1 0 18492 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A_N
timestamp 1673029049
transform -1 0 18492 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__B
timestamp 1673029049
transform -1 0 18492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1673029049
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1673029049
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A2
timestamp 1673029049
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__S
timestamp 1673029049
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__S
timestamp 1673029049
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1673029049
transform 1 0 15548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A1
timestamp 1673029049
transform -1 0 15640 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__SET_B
timestamp 1673029049
transform -1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__D
timestamp 1673029049
transform -1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__RESET_B
timestamp 1673029049
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__SET_B
timestamp 1673029049
transform -1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__RESET_B
timestamp 1673029049
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__SET_B
timestamp 1673029049
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1673029049
transform -1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1673029049
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1673029049
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__SET_B
timestamp 1673029049
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__RESET_B
timestamp 1673029049
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__D
timestamp 1673029049
transform -1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__D
timestamp 1673029049
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__D
timestamp 1673029049
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1673029049
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1673029049
transform -1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1673029049
transform -1 0 18492 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1673029049
transform -1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1673029049
transform -1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1673029049
transform -1 0 18492 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1673029049
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1673029049
transform -1 0 1196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1673029049
transform -1 0 2208 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1673029049
transform -1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1673029049
transform -1 0 18492 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1673029049
transform -1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1673029049
transform -1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1673029049
transform -1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1673029049
transform -1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 460 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1196 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1472 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27
timestamp 1673029049
transform 1 0 2668 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 1673029049
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53
timestamp 1673029049
transform 1 0 5060 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66
timestamp 1673029049
transform 1 0 6256 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79
timestamp 1673029049
transform 1 0 7452 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92
timestamp 1673029049
transform 1 0 8648 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105
timestamp 1673029049
transform 1 0 9844 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118
timestamp 1673029049
transform 1 0 11040 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131
timestamp 1673029049
transform 1 0 12236 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144
timestamp 1673029049
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_157
timestamp 1673029049
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_170
timestamp 1673029049
transform 1 0 15824 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_183
timestamp 1673029049
transform 1 0 17020 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 18216 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1673029049
transform 1 0 460 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1673029049
transform 1 0 1564 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1673029049
transform 1 0 2668 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3036 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1673029049
transform 1 0 3588 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_43
timestamp 1673029049
transform 1 0 4140 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_49
timestamp 1673029049
transform 1 0 4692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1673029049
transform 1 0 5060 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_63
timestamp 1673029049
transform 1 0 5980 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp 1673029049
transform 1 0 7084 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7452 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_94
timestamp 1673029049
transform 1 0 8832 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1673029049
transform 1 0 9568 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1673029049
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_111
timestamp 1673029049
transform 1 0 10396 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_123
timestamp 1673029049
transform 1 0 11500 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 1673029049
transform 1 0 12052 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_131
timestamp 1673029049
transform 1 0 12236 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139
timestamp 1673029049
transform 1 0 12972 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_145
timestamp 1673029049
transform 1 0 13524 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_153
timestamp 1673029049
transform 1 0 14260 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp 1673029049
transform 1 0 14628 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_163
timestamp 1673029049
transform 1 0 15180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_168
timestamp 1673029049
transform 1 0 15640 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1673029049
transform 1 0 16100 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 1673029049
transform 1 0 16836 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1673029049
transform 1 0 17020 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_191
timestamp 1673029049
transform 1 0 17756 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1673029049
transform 1 0 18492 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1673029049
transform 1 0 460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1673029049
transform 1 0 1196 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1673029049
transform 1 0 1472 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1673029049
transform 1 0 2116 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1673029049
transform 1 0 3680 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1673029049
transform 1 0 3864 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1673029049
transform 1 0 4876 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1673029049
transform 1 0 6072 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_66
timestamp 1673029049
transform 1 0 6256 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1673029049
transform 1 0 6532 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_82
timestamp 1673029049
transform 1 0 7728 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_90
timestamp 1673029049
transform 1 0 8464 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_92
timestamp 1673029049
transform 1 0 8648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_102
timestamp 1673029049
transform 1 0 9568 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_108
timestamp 1673029049
transform 1 0 10120 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_116
timestamp 1673029049
transform 1 0 10856 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_118
timestamp 1673029049
transform 1 0 11040 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_131
timestamp 1673029049
transform 1 0 12236 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1673029049
transform 1 0 13156 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1673029049
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_149
timestamp 1673029049
transform 1 0 13892 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_154
timestamp 1673029049
transform 1 0 14352 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp 1673029049
transform 1 0 15456 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_170
timestamp 1673029049
transform 1 0 15824 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1673029049
transform 1 0 16928 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_194
timestamp 1673029049
transform 1 0 18032 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196
timestamp 1673029049
transform 1 0 18216 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1673029049
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1673029049
transform 1 0 460 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1673029049
transform 1 0 1564 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_25
timestamp 1673029049
transform 1 0 2484 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1673029049
transform 1 0 2668 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1673029049
transform 1 0 3772 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_51
timestamp 1673029049
transform 1 0 4876 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_53
timestamp 1673029049
transform 1 0 5060 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1673029049
transform 1 0 5428 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp 1673029049
transform 1 0 6164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1673029049
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_79
timestamp 1673029049
transform 1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1673029049
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1673029049
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_105
timestamp 1673029049
transform 1 0 9844 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1673029049
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_116
timestamp 1673029049
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1673029049
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_131
timestamp 1673029049
transform 1 0 12236 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1673029049
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 1673029049
transform 1 0 14628 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1673029049
transform 1 0 15364 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1673029049
transform 1 0 15732 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp 1673029049
transform 1 0 16836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1673029049
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_189
timestamp 1673029049
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1673029049
transform 1 0 18124 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1673029049
transform 1 0 18492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1673029049
transform 1 0 460 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_10
timestamp 1673029049
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_14
timestamp 1673029049
transform 1 0 1472 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_24
timestamp 1673029049
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_36
timestamp 1673029049
transform 1 0 3496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1673029049
transform 1 0 3864 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1673029049
transform 1 0 4232 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_52
timestamp 1673029049
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1673029049
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_66
timestamp 1673029049
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1673029049
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1673029049
transform 1 0 7636 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_89
timestamp 1673029049
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_92
timestamp 1673029049
transform 1 0 8648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1673029049
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp 1673029049
transform 1 0 10580 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_118
timestamp 1673029049
transform 1 0 11040 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1673029049
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1673029049
transform 1 0 12604 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1673029049
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_144
timestamp 1673029049
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1673029049
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_157
timestamp 1673029049
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_170
timestamp 1673029049
transform 1 0 15824 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1673029049
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_184
timestamp 1673029049
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1673029049
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_194
timestamp 1673029049
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_196
timestamp 1673029049
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1673029049
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1673029049
transform 1 0 460 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1673029049
transform 1 0 1564 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1673029049
transform 1 0 2300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1673029049
transform 1 0 2668 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1673029049
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 1673029049
transform 1 0 3956 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1673029049
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_53
timestamp 1673029049
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_61
timestamp 1673029049
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1673029049
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1673029049
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_79
timestamp 1673029049
transform 1 0 7452 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_91
timestamp 1673029049
transform 1 0 8556 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1673029049
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_105
timestamp 1673029049
transform 1 0 9844 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_117
timestamp 1673029049
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1673029049
transform 1 0 12052 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1673029049
transform 1 0 12236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1673029049
transform 1 0 13156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1673029049
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1673029049
transform 1 0 14628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1673029049
transform 1 0 16560 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1673029049
transform 1 0 17020 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1673029049
transform 1 0 17940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1673029049
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1673029049
transform 1 0 460 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1673029049
transform 1 0 1196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_14
timestamp 1673029049
transform 1 0 1472 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_24
timestamp 1673029049
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1673029049
transform 1 0 3128 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1673029049
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_40
timestamp 1673029049
transform 1 0 3864 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_52
timestamp 1673029049
transform 1 0 4968 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1673029049
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1673029049
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1673029049
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1673029049
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1673029049
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp 1673029049
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1673029049
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_107
timestamp 1673029049
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1673029049
transform 1 0 10396 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_118
timestamp 1673029049
transform 1 0 11040 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1673029049
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1673029049
transform 1 0 12328 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1673029049
transform 1 0 13248 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1673029049
transform 1 0 13432 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1673029049
transform 1 0 15640 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1673029049
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp 1673029049
transform 1 0 17020 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_194
timestamp 1673029049
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1673029049
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1673029049
transform 1 0 460 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1673029049
transform 1 0 1012 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_13
timestamp 1673029049
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_18
timestamp 1673029049
transform 1 0 1840 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1673029049
transform 1 0 2668 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1673029049
transform 1 0 3772 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1673029049
transform 1 0 4140 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1673029049
transform 1 0 4876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1673029049
transform 1 0 5060 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_56
timestamp 1673029049
transform 1 0 5336 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1673029049
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp 1673029049
transform 1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_79
timestamp 1673029049
transform 1 0 7452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1673029049
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_95
timestamp 1673029049
transform 1 0 8924 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1673029049
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1673029049
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_112
timestamp 1673029049
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_116
timestamp 1673029049
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1673029049
transform 1 0 11776 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_131
timestamp 1673029049
transform 1 0 12236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1673029049
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_150
timestamp 1673029049
transform 1 0 13984 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_157
timestamp 1673029049
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1673029049
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_183
timestamp 1673029049
transform 1 0 17020 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1673029049
transform 1 0 17296 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_196
timestamp 1673029049
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1673029049
transform 1 0 460 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1673029049
transform 1 0 1196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_14
timestamp 1673029049
transform 1 0 1472 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_19
timestamp 1673029049
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1673029049
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1673029049
transform 1 0 3680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1673029049
transform 1 0 3864 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1673029049
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_54
timestamp 1673029049
transform 1 0 5152 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1673029049
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1673029049
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1673029049
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_74
timestamp 1673029049
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1673029049
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1673029049
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp 1673029049
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_92
timestamp 1673029049
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1673029049
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1673029049
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp 1673029049
transform 1 0 11040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1673029049
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1673029049
transform 1 0 12328 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_140
timestamp 1673029049
transform 1 0 13064 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1673029049
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1673029049
transform 1 0 15364 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_170
timestamp 1673029049
transform 1 0 15824 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_182
timestamp 1673029049
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_194
timestamp 1673029049
transform 1 0 18032 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1673029049
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1673029049
transform 1 0 460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1673029049
transform 1 0 1564 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1673029049
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_24
timestamp 1673029049
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 1673029049
transform 1 0 2668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1673029049
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1673029049
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_53
timestamp 1673029049
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp 1673029049
transform 1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1673029049
transform 1 0 7452 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1673029049
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp 1673029049
transform 1 0 9844 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_108
timestamp 1673029049
transform 1 0 10120 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1673029049
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1673029049
transform 1 0 12052 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1673029049
transform 1 0 12236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp 1673029049
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_157
timestamp 1673029049
transform 1 0 14628 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1673029049
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_183
timestamp 1673029049
transform 1 0 17020 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_191
timestamp 1673029049
transform 1 0 17756 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_194
timestamp 1673029049
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp 1673029049
transform 1 0 18492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1673029049
transform 1 0 460 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1673029049
transform 1 0 1196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_14
timestamp 1673029049
transform 1 0 1472 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1673029049
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_26
timestamp 1673029049
transform 1 0 2576 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1673029049
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 1673029049
transform 1 0 3864 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp 1673029049
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1673029049
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1673029049
transform 1 0 6072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1673029049
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1673029049
transform 1 0 8280 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_92
timestamp 1673029049
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1673029049
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_105
timestamp 1673029049
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1673029049
transform 1 0 11040 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_139
timestamp 1673029049
transform 1 0 12972 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_144
timestamp 1673029049
transform 1 0 13432 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1673029049
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_166
timestamp 1673029049
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_170
timestamp 1673029049
transform 1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1673029049
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_196
timestamp 1673029049
transform 1 0 18216 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_199
timestamp 1673029049
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1673029049
transform 1 0 460 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1673029049
transform 1 0 1012 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_19
timestamp 1673029049
transform 1 0 1932 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1673029049
transform 1 0 2484 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1673029049
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_49
timestamp 1673029049
transform 1 0 4692 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1673029049
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_75
timestamp 1673029049
transform 1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_79
timestamp 1673029049
transform 1 0 7452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1673029049
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_105
timestamp 1673029049
transform 1 0 9844 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_117
timestamp 1673029049
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_124
timestamp 1673029049
transform 1 0 11592 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_131
timestamp 1673029049
transform 1 0 12236 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1673029049
transform 1 0 12788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_145
timestamp 1673029049
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_153
timestamp 1673029049
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_157
timestamp 1673029049
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1673029049
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1673029049
transform 1 0 15456 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1673029049
transform 1 0 15824 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1673029049
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1673029049
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1673029049
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1673029049
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_187
timestamp 1673029049
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1673029049
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1673029049
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1673029049
transform 1 0 460 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1673029049
transform 1 0 1196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1673029049
transform 1 0 1472 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1673029049
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1673029049
transform 1 0 3864 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_43
timestamp 1673029049
transform 1 0 4140 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1673029049
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1673029049
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1673029049
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_66
timestamp 1673029049
transform 1 0 6256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_78
timestamp 1673029049
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_82
timestamp 1673029049
transform 1 0 7728 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp 1673029049
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1673029049
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1673029049
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_103
timestamp 1673029049
transform 1 0 9660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1673029049
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1673029049
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_123
timestamp 1673029049
transform 1 0 11500 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1673029049
transform 1 0 12604 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_144
timestamp 1673029049
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1673029049
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_170
timestamp 1673029049
transform 1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1673029049
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_194
timestamp 1673029049
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_196
timestamp 1673029049
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1673029049
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1673029049
transform 1 0 460 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_13
timestamp 1673029049
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1673029049
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1673029049
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1673029049
transform 1 0 3772 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_51
timestamp 1673029049
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1673029049
transform 1 0 5060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_75
timestamp 1673029049
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1673029049
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1673029049
transform 1 0 7728 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1673029049
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_95
timestamp 1673029049
transform 1 0 8924 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1673029049
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_105
timestamp 1673029049
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1673029049
transform 1 0 12052 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1673029049
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1673029049
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1673029049
transform 1 0 13892 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1673029049
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1673029049
transform 1 0 14628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1673029049
transform 1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_183
timestamp 1673029049
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1673029049
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_197
timestamp 1673029049
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1673029049
transform 1 0 460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1673029049
transform 1 0 1012 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_14
timestamp 1673029049
transform 1 0 1472 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_24
timestamp 1673029049
transform 1 0 2392 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_36
timestamp 1673029049
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1673029049
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 1673029049
transform 1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 1673029049
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1673029049
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1673029049
transform 1 0 6256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1673029049
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1673029049
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_89
timestamp 1673029049
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_92
timestamp 1673029049
transform 1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1673029049
transform 1 0 10856 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1673029049
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_125
timestamp 1673029049
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1673029049
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1673029049
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1673029049
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1673029049
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1673029049
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1673029049
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_173
timestamp 1673029049
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_192
timestamp 1673029049
transform 1 0 17848 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_196
timestamp 1673029049
transform 1 0 18216 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_199
timestamp 1673029049
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1673029049
transform 1 0 460 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1673029049
transform 1 0 1564 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1673029049
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_25
timestamp 1673029049
transform 1 0 2484 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 1673029049
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_34
timestamp 1673029049
transform 1 0 3312 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1673029049
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1673029049
transform 1 0 5060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1673029049
transform 1 0 5428 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1673029049
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_65
timestamp 1673029049
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1673029049
transform 1 0 6900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1673029049
transform 1 0 7268 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 1673029049
transform 1 0 7452 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1673029049
transform 1 0 8096 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1673029049
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_96
timestamp 1673029049
transform 1 0 9016 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_105
timestamp 1673029049
transform 1 0 9844 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1673029049
transform 1 0 11776 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_131
timestamp 1673029049
transform 1 0 12236 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1673029049
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1673029049
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1673029049
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_153
timestamp 1673029049
transform 1 0 14260 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_157
timestamp 1673029049
transform 1 0 14628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1673029049
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1673029049
transform 1 0 17020 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_190
timestamp 1673029049
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1673029049
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1673029049
transform 1 0 460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_12
timestamp 1673029049
transform 1 0 1288 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_14
timestamp 1673029049
transform 1 0 1472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_25
timestamp 1673029049
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_30
timestamp 1673029049
transform 1 0 2944 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1673029049
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1673029049
transform 1 0 3864 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1673029049
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1673029049
transform 1 0 5152 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_62
timestamp 1673029049
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_66
timestamp 1673029049
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_90
timestamp 1673029049
transform 1 0 8464 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1673029049
transform 1 0 8648 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_116
timestamp 1673029049
transform 1 0 10856 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1673029049
transform 1 0 11040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1673029049
transform 1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp 1673029049
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1673029049
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_155
timestamp 1673029049
transform 1 0 14444 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_163
timestamp 1673029049
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_168
timestamp 1673029049
transform 1 0 15640 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1673029049
transform 1 0 15824 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1673029049
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1673029049
transform 1 0 17940 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_196
timestamp 1673029049
transform 1 0 18216 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_199
timestamp 1673029049
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1673029049
transform 1 0 460 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1673029049
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1673029049
transform 1 0 1196 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1673029049
transform 1 0 1564 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_25
timestamp 1673029049
transform 1 0 2484 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1673029049
transform 1 0 2668 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 1673029049
transform 1 0 4600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_53
timestamp 1673029049
transform 1 0 5060 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_61
timestamp 1673029049
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 1673029049
transform 1 0 6348 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1673029049
transform 1 0 7268 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_79
timestamp 1673029049
transform 1 0 7452 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_91
timestamp 1673029049
transform 1 0 8556 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1673029049
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_103
timestamp 1673029049
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_105
timestamp 1673029049
transform 1 0 9844 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_117
timestamp 1673029049
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1673029049
transform 1 0 12052 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_131
timestamp 1673029049
transform 1 0 12236 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1673029049
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_150
timestamp 1673029049
transform 1 0 13984 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_157
timestamp 1673029049
transform 1 0 14628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_179
timestamp 1673029049
transform 1 0 16652 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_183
timestamp 1673029049
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_192
timestamp 1673029049
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1673029049
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1673029049
transform 1 0 460 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1673029049
transform 1 0 1196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1673029049
transform 1 0 1472 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1673029049
transform 1 0 3680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1673029049
transform 1 0 3864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_57
timestamp 1673029049
transform 1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_66
timestamp 1673029049
transform 1 0 6256 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1673029049
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_90
timestamp 1673029049
transform 1 0 8464 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_92
timestamp 1673029049
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1673029049
transform 1 0 9752 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1673029049
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_116
timestamp 1673029049
transform 1 0 10856 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1673029049
transform 1 0 11040 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1673029049
transform 1 0 13248 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_144
timestamp 1673029049
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1673029049
transform 1 0 15364 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1673029049
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1673029049
transform 1 0 16652 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1673029049
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_192
timestamp 1673029049
transform 1 0 17848 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_196
timestamp 1673029049
transform 1 0 18216 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1673029049
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1673029049
transform 1 0 460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1673029049
transform 1 0 1196 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1673029049
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1673029049
transform 1 0 2484 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 1673029049
transform 1 0 2668 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_48
timestamp 1673029049
transform 1 0 4600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_53
timestamp 1673029049
transform 1 0 5060 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1673029049
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_79
timestamp 1673029049
transform 1 0 7452 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1673029049
transform 1 0 8004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1673029049
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1673029049
transform 1 0 9292 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1673029049
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1673029049
transform 1 0 9844 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_127
timestamp 1673029049
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1673029049
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1673029049
transform 1 0 13340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1673029049
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1673029049
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_162
timestamp 1673029049
transform 1 0 15088 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_166
timestamp 1673029049
transform 1 0 15456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1673029049
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_181
timestamp 1673029049
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_183
timestamp 1673029049
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_186
timestamp 1673029049
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1673029049
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_194
timestamp 1673029049
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1673029049
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1673029049
transform 1 0 460 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1673029049
transform 1 0 1196 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_14
timestamp 1673029049
transform 1 0 1472 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_24
timestamp 1673029049
transform 1 0 2392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1673029049
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_40
timestamp 1673029049
transform 1 0 3864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_52
timestamp 1673029049
transform 1 0 4968 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1673029049
transform 1 0 5704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1673029049
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1673029049
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1673029049
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_92
timestamp 1673029049
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1673029049
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_116
timestamp 1673029049
transform 1 0 10856 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_118
timestamp 1673029049
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1673029049
transform 1 0 11408 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_134
timestamp 1673029049
transform 1 0 12512 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1673029049
transform 1 0 13248 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_144
timestamp 1673029049
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1673029049
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_170
timestamp 1673029049
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1673029049
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1673029049
transform 1 0 18216 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1673029049
transform 1 0 460 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_11
timestamp 1673029049
transform 1 0 1196 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_22
timestamp 1673029049
transform 1 0 2208 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1673029049
transform 1 0 2668 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1673029049
transform 1 0 3772 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_51
timestamp 1673029049
transform 1 0 4876 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_53
timestamp 1673029049
transform 1 0 5060 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_59
timestamp 1673029049
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1673029049
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_71
timestamp 1673029049
transform 1 0 6716 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1673029049
transform 1 0 7268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_79
timestamp 1673029049
transform 1 0 7452 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1673029049
transform 1 0 9384 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1673029049
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1673029049
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1673029049
transform 1 0 11500 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1673029049
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1673029049
transform 1 0 12236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1673029049
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_153
timestamp 1673029049
transform 1 0 14260 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1673029049
transform 1 0 14628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1673029049
transform 1 0 14904 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1673029049
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1673029049
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1673029049
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_183
timestamp 1673029049
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_187
timestamp 1673029049
transform 1 0 17388 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_199
timestamp 1673029049
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1673029049
transform 1 0 460 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1673029049
transform 1 0 1196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_14
timestamp 1673029049
transform 1 0 1472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1673029049
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1673029049
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1673029049
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_62
timestamp 1673029049
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_66
timestamp 1673029049
transform 1 0 6256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1673029049
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1673029049
transform 1 0 8188 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_92
timestamp 1673029049
transform 1 0 8648 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1673029049
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1673029049
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1673029049
transform 1 0 11040 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1673029049
transform 1 0 13248 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1673029049
transform 1 0 13432 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_168
timestamp 1673029049
transform 1 0 15640 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_170
timestamp 1673029049
transform 1 0 15824 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1673029049
transform 1 0 16836 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_190
timestamp 1673029049
transform 1 0 17664 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1673029049
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_196
timestamp 1673029049
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1673029049
transform 1 0 460 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1673029049
transform 1 0 1012 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_19
timestamp 1673029049
transform 1 0 1932 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1673029049
transform 1 0 2484 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_27
timestamp 1673029049
transform 1 0 2668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_33
timestamp 1673029049
transform 1 0 3220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_38
timestamp 1673029049
transform 1 0 3680 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_50
timestamp 1673029049
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1673029049
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_71
timestamp 1673029049
transform 1 0 6716 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1673029049
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1673029049
transform 1 0 7452 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_103
timestamp 1673029049
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_105
timestamp 1673029049
transform 1 0 9844 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_112
timestamp 1673029049
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_120
timestamp 1673029049
transform 1 0 11224 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1673029049
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1673029049
transform 1 0 12236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_141
timestamp 1673029049
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1673029049
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1673029049
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1673029049
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1673029049
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1673029049
transform 1 0 17020 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1673029049
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1673029049
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1673029049
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1673029049
transform 1 0 460 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1673029049
transform 1 0 1196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_14
timestamp 1673029049
transform 1 0 1472 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1673029049
transform 1 0 3680 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_40
timestamp 1673029049
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1673029049
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_66
timestamp 1673029049
transform 1 0 6256 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_74
timestamp 1673029049
transform 1 0 6992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1673029049
transform 1 0 7820 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 1673029049
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1673029049
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1673029049
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1673029049
transform 1 0 10488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_116
timestamp 1673029049
transform 1 0 10856 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1673029049
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_140
timestamp 1673029049
transform 1 0 13064 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1673029049
transform 1 0 13432 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_152
timestamp 1673029049
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1673029049
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_166
timestamp 1673029049
transform 1 0 15456 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1673029049
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_194
timestamp 1673029049
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1673029049
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1673029049
transform 1 0 460 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_16
timestamp 1673029049
transform 1 0 1656 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_24
timestamp 1673029049
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1673029049
transform 1 0 2668 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_40
timestamp 1673029049
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1673029049
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_75
timestamp 1673029049
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_79
timestamp 1673029049
transform 1 0 7452 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1673029049
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_103
timestamp 1673029049
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_105
timestamp 1673029049
transform 1 0 9844 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_108
timestamp 1673029049
transform 1 0 10120 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1673029049
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1673029049
transform 1 0 12052 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1673029049
transform 1 0 12236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1673029049
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1673029049
transform 1 0 13432 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_148
timestamp 1673029049
transform 1 0 13800 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp 1673029049
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_157
timestamp 1673029049
transform 1 0 14628 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1673029049
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_183
timestamp 1673029049
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1673029049
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_197
timestamp 1673029049
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1673029049
transform 1 0 460 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1673029049
transform 1 0 1196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_14
timestamp 1673029049
transform 1 0 1472 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1673029049
transform 1 0 3680 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1673029049
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_44
timestamp 1673029049
transform 1 0 4232 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1673029049
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_64
timestamp 1673029049
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1673029049
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1673029049
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_92
timestamp 1673029049
transform 1 0 8648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1673029049
transform 1 0 9568 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_111
timestamp 1673029049
transform 1 0 10396 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1673029049
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1673029049
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_136
timestamp 1673029049
transform 1 0 12696 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1673029049
transform 1 0 13248 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_144
timestamp 1673029049
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1673029049
transform 1 0 14536 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1673029049
transform 1 0 14904 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_168
timestamp 1673029049
transform 1 0 15640 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_170
timestamp 1673029049
transform 1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_194
timestamp 1673029049
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_196
timestamp 1673029049
transform 1 0 18216 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_199
timestamp 1673029049
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1673029049
transform 1 0 460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1673029049
transform 1 0 1012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_20
timestamp 1673029049
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1673029049
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1673029049
transform 1 0 3772 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_51
timestamp 1673029049
transform 1 0 4876 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1673029049
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_75
timestamp 1673029049
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1673029049
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_103
timestamp 1673029049
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_105
timestamp 1673029049
transform 1 0 9844 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1673029049
transform 1 0 10580 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1673029049
transform 1 0 11132 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_129
timestamp 1673029049
transform 1 0 12052 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1673029049
transform 1 0 12236 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1673029049
transform 1 0 13156 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1673029049
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_155
timestamp 1673029049
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1673029049
transform 1 0 14628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1673029049
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_183
timestamp 1673029049
transform 1 0 17020 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1673029049
transform 1 0 17848 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1673029049
transform 1 0 18492 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1673029049
transform 1 0 460 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1673029049
transform 1 0 1196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_14
timestamp 1673029049
transform 1 0 1472 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_24
timestamp 1673029049
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1673029049
transform 1 0 2852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1673029049
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_40
timestamp 1673029049
transform 1 0 3864 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_62
timestamp 1673029049
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp 1673029049
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_77
timestamp 1673029049
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_84
timestamp 1673029049
transform 1 0 7912 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_90
timestamp 1673029049
transform 1 0 8464 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_92
timestamp 1673029049
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1673029049
transform 1 0 9476 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_105
timestamp 1673029049
transform 1 0 9844 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_111
timestamp 1673029049
transform 1 0 10396 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1673029049
transform 1 0 11040 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1673029049
transform 1 0 12972 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_144
timestamp 1673029049
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1673029049
transform 1 0 15364 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1673029049
transform 1 0 15824 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_192
timestamp 1673029049
transform 1 0 17848 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1673029049
transform 1 0 18216 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1673029049
transform 1 0 460 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_15
timestamp 1673029049
transform 1 0 1564 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_23
timestamp 1673029049
transform 1 0 2300 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_27
timestamp 1673029049
transform 1 0 2668 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_48
timestamp 1673029049
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1673029049
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1673029049
transform 1 0 7084 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1673029049
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1673029049
transform 1 0 9568 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1673029049
transform 1 0 9844 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1673029049
transform 1 0 11776 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1673029049
transform 1 0 12236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1673029049
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1673029049
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1673029049
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1673029049
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1673029049
transform 1 0 14628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_167
timestamp 1673029049
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1673029049
transform 1 0 16008 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_180
timestamp 1673029049
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_183
timestamp 1673029049
transform 1 0 17020 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_191
timestamp 1673029049
transform 1 0 17756 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_194
timestamp 1673029049
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1673029049
transform 1 0 18492 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1673029049
transform 1 0 460 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1673029049
transform 1 0 1196 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_14
timestamp 1673029049
transform 1 0 1472 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_21
timestamp 1673029049
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_28
timestamp 1673029049
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_33
timestamp 1673029049
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1673029049
transform 1 0 3680 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1673029049
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1673029049
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1673029049
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_66
timestamp 1673029049
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_88
timestamp 1673029049
transform 1 0 8280 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_92
timestamp 1673029049
transform 1 0 8648 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_116
timestamp 1673029049
transform 1 0 10856 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 1673029049
transform 1 0 11040 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_126
timestamp 1673029049
transform 1 0 11776 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1673029049
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_140
timestamp 1673029049
transform 1 0 13064 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_144
timestamp 1673029049
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_160
timestamp 1673029049
transform 1 0 14904 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1673029049
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1673029049
transform 1 0 15824 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_192
timestamp 1673029049
transform 1 0 17848 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1673029049
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1673029049
transform 1 0 460 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_15
timestamp 1673029049
transform 1 0 1564 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_23
timestamp 1673029049
transform 1 0 2300 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1673029049
transform 1 0 2668 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_48
timestamp 1673029049
transform 1 0 4600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_53
timestamp 1673029049
transform 1 0 5060 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_77
timestamp 1673029049
transform 1 0 7268 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_79
timestamp 1673029049
transform 1 0 7452 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1673029049
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1673029049
transform 1 0 9844 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1673029049
transform 1 0 11776 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_131
timestamp 1673029049
transform 1 0 12236 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_137
timestamp 1673029049
transform 1 0 12788 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1673029049
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1673029049
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp 1673029049
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_183
timestamp 1673029049
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1673029049
transform 1 0 17940 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1673029049
transform 1 0 18492 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1673029049
transform 1 0 460 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1673029049
transform 1 0 1196 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_14
timestamp 1673029049
transform 1 0 1472 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1673029049
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_22
timestamp 1673029049
transform 1 0 2208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_27
timestamp 1673029049
transform 1 0 2668 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1673029049
transform 1 0 3404 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1673029049
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_40
timestamp 1673029049
transform 1 0 3864 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_51
timestamp 1673029049
transform 1 0 4876 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1673029049
transform 1 0 5060 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_56
timestamp 1673029049
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1673029049
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_66
timestamp 1673029049
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1673029049
transform 1 0 6900 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_77
timestamp 1673029049
transform 1 0 7268 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1673029049
transform 1 0 7452 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_88
timestamp 1673029049
transform 1 0 8280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_92
timestamp 1673029049
transform 1 0 8648 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_101
timestamp 1673029049
transform 1 0 9476 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_105
timestamp 1673029049
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1673029049
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_118
timestamp 1673029049
transform 1 0 11040 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_126
timestamp 1673029049
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_131
timestamp 1673029049
transform 1 0 12236 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_144
timestamp 1673029049
transform 1 0 13432 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_155
timestamp 1673029049
transform 1 0 14444 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1673029049
transform 1 0 14628 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1673029049
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1673029049
transform 1 0 15824 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_175
timestamp 1673029049
transform 1 0 16284 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_181
timestamp 1673029049
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_183
timestamp 1673029049
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_194
timestamp 1673029049
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_196
timestamp 1673029049
transform 1 0 18216 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1673029049
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 184 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 18860 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 184 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1673029049
transform 1 0 184 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1673029049
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1673029049
transform 1 0 184 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1673029049
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1673029049
transform 1 0 184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1673029049
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1673029049
transform 1 0 184 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1673029049
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1673029049
transform 1 0 184 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1673029049
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1673029049
transform 1 0 184 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1673029049
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1673029049
transform 1 0 184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1673029049
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1673029049
transform 1 0 184 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1673029049
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1673029049
transform 1 0 184 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1673029049
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1673029049
transform 1 0 184 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1673029049
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1673029049
transform 1 0 184 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1673029049
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1673029049
transform 1 0 184 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1673029049
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1673029049
transform 1 0 184 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1673029049
transform -1 0 18860 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1673029049
transform 1 0 184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1673029049
transform -1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1673029049
transform 1 0 184 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1673029049
transform -1 0 18860 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1673029049
transform 1 0 184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1673029049
transform -1 0 18860 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1673029049
transform 1 0 184 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1673029049
transform -1 0 18860 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1673029049
transform 1 0 184 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1673029049
transform -1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1673029049
transform 1 0 184 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1673029049
transform -1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1673029049
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1673029049
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1673029049
transform 1 0 4968 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1673029049
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1673029049
transform 1 0 7360 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1673029049
transform 1 0 8556 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1673029049
transform 1 0 9752 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1673029049
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1673029049
transform 1 0 12144 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1673029049
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1673029049
transform 1 0 14536 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1673029049
transform 1 0 15732 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1673029049
transform 1 0 16928 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1673029049
transform 1 0 18124 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1673029049
transform 1 0 2576 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1673029049
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1673029049
transform 1 0 7360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1673029049
transform 1 0 9752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1673029049
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1673029049
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1673029049
transform 1 0 16928 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1673029049
transform 1 0 1380 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1673029049
transform 1 0 3772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1673029049
transform 1 0 6164 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1673029049
transform 1 0 8556 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1673029049
transform 1 0 10948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1673029049
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1673029049
transform 1 0 15732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1673029049
transform 1 0 18124 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1673029049
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1673029049
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1673029049
transform 1 0 7360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1673029049
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1673029049
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1673029049
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1673029049
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1673029049
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1673029049
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1673029049
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1673029049
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1673029049
transform 1 0 10948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1673029049
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1673029049
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1673029049
transform 1 0 18124 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1673029049
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1673029049
transform 1 0 4968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1673029049
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1673029049
transform 1 0 9752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1673029049
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1673029049
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1673029049
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1673029049
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1673029049
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1673029049
transform 1 0 6164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1673029049
transform 1 0 8556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1673029049
transform 1 0 10948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1673029049
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1673029049
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1673029049
transform 1 0 18124 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1673029049
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1673029049
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1673029049
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1673029049
transform 1 0 9752 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1673029049
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1673029049
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1673029049
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1673029049
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1673029049
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1673029049
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1673029049
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1673029049
transform 1 0 10948 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1673029049
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1673029049
transform 1 0 15732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1673029049
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1673029049
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1673029049
transform 1 0 4968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1673029049
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1673029049
transform 1 0 9752 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1673029049
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1673029049
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1673029049
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1673029049
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1673029049
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1673029049
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1673029049
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1673029049
transform 1 0 10948 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1673029049
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1673029049
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1673029049
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1673029049
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1673029049
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1673029049
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1673029049
transform 1 0 9752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1673029049
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1673029049
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1673029049
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1673029049
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1673029049
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1673029049
transform 1 0 6164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1673029049
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1673029049
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1673029049
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1673029049
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1673029049
transform 1 0 18124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1673029049
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1673029049
transform 1 0 4968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1673029049
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1673029049
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1673029049
transform 1 0 12144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1673029049
transform 1 0 14536 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1673029049
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1673029049
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1673029049
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1673029049
transform 1 0 6164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1673029049
transform 1 0 8556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1673029049
transform 1 0 10948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1673029049
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1673029049
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1673029049
transform 1 0 18124 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1673029049
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1673029049
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1673029049
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1673029049
transform 1 0 9752 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1673029049
transform 1 0 12144 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1673029049
transform 1 0 14536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1673029049
transform 1 0 16928 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1673029049
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1673029049
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1673029049
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1673029049
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1673029049
transform 1 0 10948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1673029049
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1673029049
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1673029049
transform 1 0 18124 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1673029049
transform 1 0 2576 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1673029049
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1673029049
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1673029049
transform 1 0 9752 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1673029049
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1673029049
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1673029049
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1673029049
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1673029049
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1673029049
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1673029049
transform 1 0 8556 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1673029049
transform 1 0 10948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1673029049
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1673029049
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1673029049
transform 1 0 18124 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1673029049
transform 1 0 2576 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1673029049
transform 1 0 4968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1673029049
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1673029049
transform 1 0 9752 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1673029049
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1673029049
transform 1 0 14536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1673029049
transform 1 0 16928 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1673029049
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1673029049
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1673029049
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1673029049
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1673029049
transform 1 0 10948 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1673029049
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1673029049
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1673029049
transform 1 0 18124 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1673029049
transform 1 0 2576 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1673029049
transform 1 0 4968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1673029049
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1673029049
transform 1 0 9752 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1673029049
transform 1 0 12144 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1673029049
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1673029049
transform 1 0 16928 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1673029049
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1673029049
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1673029049
transform 1 0 6164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1673029049
transform 1 0 8556 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1673029049
transform 1 0 10948 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1673029049
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1673029049
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1673029049
transform 1 0 18124 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1673029049
transform 1 0 2576 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1673029049
transform 1 0 4968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1673029049
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1673029049
transform 1 0 9752 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1673029049
transform 1 0 12144 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1673029049
transform 1 0 14536 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1673029049
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1673029049
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1673029049
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1673029049
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1673029049
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1673029049
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1673029049
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1673029049
transform 1 0 15732 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1673029049
transform 1 0 18124 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1673029049
transform 1 0 2576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1673029049
transform 1 0 4968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1673029049
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1673029049
transform 1 0 9752 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1673029049
transform 1 0 12144 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1673029049
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1673029049
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1673029049
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1673029049
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1673029049
transform 1 0 6164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1673029049
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1673029049
transform 1 0 10948 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1673029049
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1673029049
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1673029049
transform 1 0 18124 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1673029049
transform 1 0 2576 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1673029049
transform 1 0 4968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1673029049
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1673029049
transform 1 0 9752 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1673029049
transform 1 0 12144 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1673029049
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1673029049
transform 1 0 16928 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1673029049
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1673029049
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1673029049
transform 1 0 6164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1673029049
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1673029049
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1673029049
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1673029049
transform 1 0 15732 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1673029049
transform 1 0 18124 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1673029049
transform 1 0 2576 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1673029049
transform 1 0 4968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1673029049
transform 1 0 7360 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1673029049
transform 1 0 9752 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1673029049
transform 1 0 12144 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1673029049
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1673029049
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1673029049
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1673029049
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1673029049
transform 1 0 6164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1673029049
transform 1 0 8556 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1673029049
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1673029049
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1673029049
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1673029049
transform 1 0 18124 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1673029049
transform 1 0 2576 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1673029049
transform 1 0 4968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1673029049
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1673029049
transform 1 0 9752 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1673029049
transform 1 0 12144 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1673029049
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1673029049
transform 1 0 16928 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1673029049
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1673029049
transform 1 0 2576 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1673029049
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1673029049
transform 1 0 4968 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1673029049
transform 1 0 6164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1673029049
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1673029049
transform 1 0 8556 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1673029049
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1673029049
transform 1 0 10948 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1673029049
transform 1 0 12144 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1673029049
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1673029049
transform 1 0 14536 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1673029049
transform 1 0 15732 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1673029049
transform 1 0 16928 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1673029049
transform 1 0 18124 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3956 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1673029049
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1673029049
transform -1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1673029049
transform -1 0 7268 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1673029049
transform -1 0 9568 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1673029049
transform 1 0 16008 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1673029049
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1673029049
transform -1 0 1932 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1673029049
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1673029049
transform -1 0 2392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1673029049
transform -1 0 2392 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1673029049
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1673029049
transform 1 0 5244 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1673029049
transform 1 0 5244 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1673029049
transform 1 0 2852 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1673029049
transform 1 0 1656 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1673029049
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1673029049
transform 1 0 6440 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1673029049
transform 1 0 9384 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1673029049
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1673029049
transform 1 0 8004 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1673029049
transform 1 0 6900 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1673029049
transform 1 0 1104 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1673029049
transform -1 0 2024 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1673029049
transform -1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1673029049
transform -1 0 9292 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1673029049
transform -1 0 10856 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1673029049
transform -1 0 15548 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1673029049
transform -1 0 15548 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1673029049
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1673029049
transform 1 0 11132 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1673029049
transform -1 0 14444 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1673029049
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1673029049
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1673029049
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1673029049
transform 1 0 12328 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1673029049
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1673029049
transform -1 0 14168 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1673029049
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1673029049
transform 1 0 17112 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1673029049
transform 1 0 16100 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 17480 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _246_
timestamp 1673029049
transform -1 0 6992 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1012 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1673029049
transform -1 0 1012 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2116 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _250_
timestamp 1673029049
transform -1 0 9568 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1673029049
transform 1 0 17848 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1673029049
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _253_
timestamp 1673029049
transform 1 0 14168 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _254_
timestamp 1673029049
transform -1 0 12604 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _255_
timestamp 1673029049
transform -1 0 13524 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _256_
timestamp 1673029049
transform 1 0 11132 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _257__7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 8280 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1673029049
transform -1 0 1012 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _259__4
timestamp 1673029049
transform -1 0 5704 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1673029049
transform -1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1673029049
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _262__1
timestamp 1673029049
transform -1 0 11684 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1673029049
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1673029049
transform -1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13524 0 1 16864
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 11224 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15088 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14260 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1673029049
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15640 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15456 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13340 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 10396 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _277_
timestamp 1673029049
transform -1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 9936 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1673029049
transform -1 0 2116 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _280_
timestamp 1673029049
transform 1 0 5152 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 4876 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _282_
timestamp 1673029049
transform -1 0 2116 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _283_
timestamp 1673029049
transform -1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5060 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5428 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _286_
timestamp 1673029049
transform -1 0 4508 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1673029049
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 4784 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _289_
timestamp 1673029049
transform 1 0 2024 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _290_
timestamp 1673029049
transform 1 0 3496 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _291_
timestamp 1673029049
transform 1 0 5152 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _292_
timestamp 1673029049
transform 1 0 4232 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 1673029049
transform -1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _294_
timestamp 1673029049
transform -1 0 4784 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 1673029049
transform 1 0 2944 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1673029049
transform -1 0 2852 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp 1673029049
transform 1 0 6624 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _298_
timestamp 1673029049
transform 1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 9660 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16836 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _301_
timestamp 1673029049
transform -1 0 13984 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1673029049
transform -1 0 13248 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _303_
timestamp 1673029049
transform -1 0 14260 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7820 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7452 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1673029049
transform -1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7544 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _308_
timestamp 1673029049
transform 1 0 15824 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _309_
timestamp 1673029049
transform -1 0 17664 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _310_
timestamp 1673029049
transform 1 0 17112 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16836 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2208 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _313_
timestamp 1673029049
transform 1 0 552 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _314_
timestamp 1673029049
transform 1 0 2944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _315_
timestamp 1673029049
transform 1 0 2944 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _316_
timestamp 1673029049
transform 1 0 2668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1673029049
transform -1 0 1288 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 828 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _319_
timestamp 1673029049
transform 1 0 5336 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _320_
timestamp 1673029049
transform 1 0 4324 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _321_
timestamp 1673029049
transform -1 0 4140 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _322_
timestamp 1673029049
transform -1 0 3588 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _323_
timestamp 1673029049
transform -1 0 10856 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _324_
timestamp 1673029049
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _325_
timestamp 1673029049
transform -1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _326_
timestamp 1673029049
transform -1 0 10396 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _327_
timestamp 1673029049
transform 1 0 552 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _328_
timestamp 1673029049
transform 1 0 8004 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _329_
timestamp 1673029049
transform 1 0 7544 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _330_
timestamp 1673029049
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _331_
timestamp 1673029049
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _332_
timestamp 1673029049
transform 1 0 10580 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _333_
timestamp 1673029049
transform -1 0 9752 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _334_
timestamp 1673029049
transform -1 0 10488 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _335_
timestamp 1673029049
transform 1 0 11132 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _336_
timestamp 1673029049
transform -1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _337_
timestamp 1673029049
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _338_
timestamp 1673029049
transform 1 0 12604 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _339_
timestamp 1673029049
transform 1 0 11592 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _340_
timestamp 1673029049
transform -1 0 13156 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _341_
timestamp 1673029049
transform -1 0 13892 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _342_
timestamp 1673029049
transform 1 0 13064 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _343_
timestamp 1673029049
transform -1 0 17756 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4232 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _346_
timestamp 1673029049
transform 1 0 15272 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _347_
timestamp 1673029049
transform -1 0 15548 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand4bb_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 3864 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _349_
timestamp 1673029049
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _350_
timestamp 1673029049
transform 1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _351_
timestamp 1673029049
transform 1 0 5244 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _352_
timestamp 1673029049
transform 1 0 5704 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6716 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1673029049
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1673029049
transform 1 0 4232 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _356_
timestamp 1673029049
transform -1 0 4784 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5796 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 3312 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _359_
timestamp 1673029049
transform 1 0 1564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _360_
timestamp 1673029049
transform -1 0 3128 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1673029049
transform 1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1673029049
transform -1 0 2484 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1673029049
transform -1 0 2484 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _364_
timestamp 1673029049
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _365_
timestamp 1673029049
transform -1 0 7728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _366_
timestamp 1673029049
transform -1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 8464 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _368_
timestamp 1673029049
transform -1 0 8188 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _369_
timestamp 1673029049
transform 1 0 6440 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1673029049
transform -1 0 1656 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1673029049
transform -1 0 2392 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2300 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _373_
timestamp 1673029049
transform 1 0 1564 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _374_
timestamp 1673029049
transform -1 0 2300 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6072 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _376_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 4968 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _377_
timestamp 1673029049
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _378_
timestamp 1673029049
transform 1 0 17664 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _379_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 17296 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _380_
timestamp 1673029049
transform -1 0 18400 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _381_
timestamp 1673029049
transform -1 0 18492 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _382_
timestamp 1673029049
transform 1 0 17388 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _383_
timestamp 1673029049
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _384_
timestamp 1673029049
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _385_
timestamp 1673029049
transform 1 0 17572 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _386_
timestamp 1673029049
transform -1 0 18308 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _387_
timestamp 1673029049
transform 1 0 17112 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _388_
timestamp 1673029049
transform 1 0 12604 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _389_
timestamp 1673029049
transform -1 0 13708 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _390_
timestamp 1673029049
transform 1 0 12144 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _391_
timestamp 1673029049
transform 1 0 13064 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1673029049
transform -1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1673029049
transform -1 0 11500 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _394_
timestamp 1673029049
transform -1 0 11592 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _395_
timestamp 1673029049
transform -1 0 12788 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 10672 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 12052 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _398_
timestamp 1673029049
transform -1 0 13156 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _399_
timestamp 1673029049
transform -1 0 13984 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _400_
timestamp 1673029049
transform -1 0 9844 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _401_
timestamp 1673029049
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _402_
timestamp 1673029049
transform 1 0 8740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1673029049
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1673029049
transform -1 0 16744 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _405_
timestamp 1673029049
transform 1 0 14904 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _406_
timestamp 1673029049
transform -1 0 15456 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _407_
timestamp 1673029049
transform -1 0 15180 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _408__8
timestamp 1673029049
transform -1 0 10396 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _409__9
timestamp 1673029049
transform -1 0 7912 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _410__5
timestamp 1673029049
transform -1 0 5704 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _411__6
timestamp 1673029049
transform -1 0 2208 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _412__2
timestamp 1673029049
transform -1 0 16652 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _413__3
timestamp 1673029049
transform -1 0 10488 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7728 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _415_
timestamp 1673029049
transform -1 0 9568 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _416_
timestamp 1673029049
transform 1 0 6348 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _416__32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 9384 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _418_
timestamp 1673029049
transform 1 0 6348 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _419_
timestamp 1673029049
transform 1 0 14720 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp 1673029049
transform 1 0 5244 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5244 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1673029049
transform 1 0 4048 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1673029049
transform 1 0 3956 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _424_
timestamp 1673029049
transform 1 0 4140 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1673029049
transform 1 0 5152 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1840 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5152 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _428_
timestamp 1673029049
transform 1 0 2852 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _429_
timestamp 1673029049
transform 1 0 5152 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _430_
timestamp 1673029049
transform -1 0 3680 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _431_
timestamp 1673029049
transform 1 0 1656 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _432_
timestamp 1673029049
transform -1 0 4600 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _433_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7544 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _434_
timestamp 1673029049
transform 1 0 7728 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6348 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _436_
timestamp 1673029049
transform 1 0 1748 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _437_
timestamp 1673029049
transform 1 0 1748 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _438_
timestamp 1673029049
transform -1 0 4600 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp 1673029049
transform -1 0 12972 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _440_
timestamp 1673029049
transform -1 0 12052 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1673029049
transform -1 0 12972 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _442_
timestamp 1673029049
transform -1 0 11776 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _443_
timestamp 1673029049
transform -1 0 10856 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _444_
timestamp 1673029049
transform -1 0 10856 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1673029049
transform 1 0 4416 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1673029049
transform 1 0 16376 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1673029049
transform 1 0 15916 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1673029049
transform 1 0 16100 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1673029049
transform 1 0 16100 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _450_
timestamp 1673029049
transform -1 0 16560 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _451_
timestamp 1673029049
transform -1 0 15640 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _452_
timestamp 1673029049
transform 1 0 11132 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _453_
timestamp 1673029049
transform 1 0 13524 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1673029049
transform 1 0 16100 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _455_
timestamp 1673029049
transform -1 0 13248 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _456_
timestamp 1673029049
transform 1 0 9936 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _457_
timestamp 1673029049
transform -1 0 13248 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _458_
timestamp 1673029049
transform 1 0 13524 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _459_
timestamp 1673029049
transform -1 0 14260 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1673029049
transform -1 0 15640 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1673029049
transform 1 0 6532 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _462_
timestamp 1673029049
transform -1 0 16836 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1673029049
transform -1 0 16836 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 1673029049
transform 1 0 14720 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1673029049
transform 1 0 16192 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1673029049
transform 1 0 16100 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1673029049
transform 1 0 14996 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1673029049
transform -1 0 16836 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _469_
timestamp 1673029049
transform 1 0 15916 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1673029049
transform -1 0 17848 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 9016 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_0_divider.out $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider2.out
timestamp 1673029049
transform -1 0 16560 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1673029049
transform 1 0 5428 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net11
timestamp 1673029049
transform 1 0 9936 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk
timestamp 1673029049
transform -1 0 8188 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1673029049
transform -1 0 16560 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__037_
timestamp 1673029049
transform -1 0 9660 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0__f_divider.out $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider2.out
timestamp 1673029049
transform -1 0 15364 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_ext_clk
timestamp 1673029049
transform -1 0 4600 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net11
timestamp 1673029049
transform -1 0 7084 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk
timestamp 1673029049
transform -1 0 7084 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk90
timestamp 1673029049
transform -1 0 15364 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__037_
timestamp 1673029049
transform 1 0 11132 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1__f_divider.out
timestamp 1673029049
transform 1 0 9384 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider2.out
timestamp 1673029049
transform 1 0 14996 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_ext_clk
timestamp 1673029049
transform 1 0 5244 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net11
timestamp 1673029049
transform -1 0 9660 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk90
timestamp 1673029049
transform -1 0 15364 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk
timestamp 1673029049
transform -1 0 4600 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14444 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 17296 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout16
timestamp 1673029049
transform 1 0 17848 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16284 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1673029049
transform -1 0 6900 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout19
timestamp 1673029049
transform -1 0 10580 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout20
timestamp 1673029049
transform -1 0 10488 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1673029049
transform -1 0 7268 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1673029049
transform -1 0 14444 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1673029049
transform 1 0 17112 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1673029049
transform 1 0 8924 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1673029049
transform -1 0 7544 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1673029049
transform -1 0 6348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1673029049
transform -1 0 6072 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout28
timestamp 1673029049
transform -1 0 6900 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout29
timestamp 1673029049
transform -1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout30
timestamp 1673029049
transform 1 0 12328 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1673029049
transform 1 0 4784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 17204 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1673029049
transform -1 0 17848 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1673029049
transform -1 0 17848 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1673029049
transform -1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1673029049
transform -1 0 6072 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1673029049
transform -1 0 7820 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1673029049
transform 1 0 8740 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 18032 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1673029049
transform 1 0 17756 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1673029049
transform -1 0 828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1673029049
transform -1 0 1840 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1673029049
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1673029049
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1673029049
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1673029049
transform 1 0 17756 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1673029049
transform 1 0 18216 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1673029049
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12880 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  user_clk_out_buffer
timestamp 1673029049
transform 1 0 9936 0 -1 16864
box -38 -48 1878 592
<< labels >>
flabel metal4 s 3100 496 3420 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6200 496 6520 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9300 496 9620 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12400 496 12720 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15500 496 15820 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 18600 496 18920 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1550 496 1870 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4650 496 4970 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7750 496 8070 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10850 496 11170 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13950 496 14270 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17050 496 17370 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7102 19200 7158 20000 0 FreeSans 224 90 0 0 core_clk
port 2 nsew signal tristate
flabel metal2 s 4250 19200 4306 20000 0 FreeSans 224 90 0 0 ext_clk
port 3 nsew signal input
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 ext_clk_sel
port 4 nsew signal input
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 ext_reset
port 5 nsew signal input
flabel metal2 s 15658 19200 15714 20000 0 FreeSans 224 90 0 0 pll_clk
port 6 nsew signal input
flabel metal2 s 18510 19200 18566 20000 0 FreeSans 224 90 0 0 pll_clk90
port 7 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 porb
port 8 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 resetb
port 9 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 resetb_sync
port 10 nsew signal tristate
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 sel2[0]
port 11 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 sel2[1]
port 12 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 sel2[2]
port 13 nsew signal input
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 sel[0]
port 14 nsew signal input
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 sel[1]
port 15 nsew signal input
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 sel[2]
port 16 nsew signal input
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 user_clk
port 17 nsew signal tristate
rlabel metal1 9552 17952 9552 17952 0 VGND
rlabel metal1 9522 18496 9522 18496 0 VPWR
rlabel metal1 13018 13362 13018 13362 0 _000_
rlabel metal1 5658 6120 5658 6120 0 _001_
rlabel metal1 9568 11730 9568 11730 0 _002_
rlabel metal1 3128 6426 3128 6426 0 _003_
rlabel metal1 1196 13498 1196 13498 0 _004_
rlabel metal2 1978 15776 1978 15776 0 _005_
rlabel metal1 1288 3910 1288 3910 0 _006_
rlabel metal2 5290 3366 5290 3366 0 _007_
rlabel metal1 1380 2618 1380 2618 0 _008_
rlabel metal1 6256 2618 6256 2618 0 _009_
rlabel metal2 8786 4386 8786 4386 0 _010_
rlabel metal1 6992 2074 6992 2074 0 _011_
rlabel metal1 1932 6698 1932 6698 0 _012_
rlabel metal2 1610 11424 1610 11424 0 _013_
rlabel metal2 2346 9316 2346 9316 0 _014_
rlabel metal1 16882 3706 16882 3706 0 _015_
rlabel metal1 16238 2074 16238 2074 0 _016_
rlabel metal1 15594 16626 15594 16626 0 _017_
rlabel metal1 11270 15130 11270 15130 0 _018_
rlabel metal1 13478 14926 13478 14926 0 _019_
rlabel metal1 11178 4794 11178 4794 0 _020_
rlabel metal1 11224 5338 11224 5338 0 _021_
rlabel metal1 13340 3706 13340 3706 0 _022_
rlabel metal1 10212 12818 10212 12818 0 _023_
rlabel metal1 9200 11322 9200 11322 0 _024_
rlabel metal1 10764 11866 10764 11866 0 _025_
rlabel metal2 7222 9894 7222 9894 0 _026_
rlabel metal1 16606 11084 16606 11084 0 _027_
rlabel metal2 1426 14382 1426 14382 0 _028_
rlabel metal1 3864 5338 3864 5338 0 _029_
rlabel metal2 4554 3366 4554 3366 0 _030_
rlabel metal1 9292 2618 9292 2618 0 _031_
rlabel metal1 16836 1938 16836 1938 0 _032_
rlabel metal1 12926 13260 12926 13260 0 _033_
rlabel metal1 14812 16558 14812 16558 0 _034_
rlabel metal1 11914 3536 11914 3536 0 _035_
rlabel metal1 8234 10676 8234 10676 0 _036_
rlabel metal1 8142 16218 8142 16218 0 _037_
rlabel metal2 16054 11764 16054 11764 0 _038_
rlabel metal2 1242 8160 1242 8160 0 _039_
rlabel metal1 1564 6426 1564 6426 0 _040_
rlabel metal1 1518 11662 1518 11662 0 _041_
rlabel metal1 2438 9554 2438 9554 0 _042_
rlabel metal1 1012 7990 1012 7990 0 _043_
rlabel metal1 2438 8466 2438 8466 0 _044_
rlabel via1 1955 2074 1955 2074 0 _045_
rlabel metal1 2162 3162 2162 3162 0 _046_
rlabel metal1 5796 1530 5796 1530 0 _047_
rlabel metal1 5474 2074 5474 2074 0 _048_
rlabel metal1 3082 1530 3082 1530 0 _049_
rlabel metal2 2898 2278 2898 2278 0 _050_
rlabel metal1 7912 2550 7912 2550 0 _051_
rlabel metal1 7314 2618 7314 2618 0 _052_
rlabel metal1 10028 2006 10028 2006 0 _053_
rlabel metal1 9292 3162 9292 3162 0 _054_
rlabel metal1 9660 1326 9660 1326 0 _055_
rlabel metal1 7682 1530 7682 1530 0 _056_
rlabel metal1 1472 13498 1472 13498 0 _057_
rlabel metal1 1334 15674 1334 15674 0 _058_
rlabel metal1 9476 13838 9476 13838 0 _059_
rlabel metal1 8878 14586 8878 14586 0 _060_
rlabel metal1 8510 12614 8510 12614 0 _061_
rlabel metal2 10626 10948 10626 10948 0 _062_
rlabel metal2 10442 12410 10442 12410 0 _063_
rlabel metal1 10672 10574 10672 10574 0 _064_
rlabel metal1 14996 16762 14996 16762 0 _065_
rlabel metal1 15364 16762 15364 16762 0 _066_
rlabel metal1 11684 15674 11684 15674 0 _067_
rlabel metal1 11408 14926 11408 14926 0 _068_
rlabel metal1 14168 15674 14168 15674 0 _069_
rlabel metal1 14260 14926 14260 14926 0 _070_
rlabel metal1 12650 3672 12650 3672 0 _071_
rlabel metal1 11316 3706 11316 3706 0 _072_
rlabel metal1 12512 2006 12512 2006 0 _073_
rlabel metal1 11960 3706 11960 3706 0 _074_
rlabel metal1 13616 1530 13616 1530 0 _075_
rlabel metal1 13984 2618 13984 2618 0 _076_
rlabel metal1 17388 2346 17388 2346 0 _077_
rlabel metal1 16606 1360 16606 1360 0 _078_
rlabel metal1 15364 8602 15364 8602 0 _088_
rlabel metal2 4554 14314 4554 14314 0 _089_
rlabel metal1 5612 10234 5612 10234 0 _090_
rlabel metal1 1978 5270 1978 5270 0 _091_
rlabel metal2 4370 4590 4370 4590 0 _092_
rlabel metal1 2346 4794 2346 4794 0 _093_
rlabel metal1 4784 4794 4784 4794 0 _094_
rlabel metal1 2668 9622 2668 9622 0 _095_
rlabel metal1 2024 11322 2024 11322 0 _096_
rlabel metal1 2438 10200 2438 10200 0 _097_
rlabel metal2 7406 4896 7406 4896 0 _098_
rlabel metal2 8418 5780 8418 5780 0 _099_
rlabel metal1 6578 3910 6578 3910 0 _100_
rlabel metal2 2162 14076 2162 14076 0 _101_
rlabel metal1 2208 14858 2208 14858 0 _102_
rlabel metal2 2898 17034 2898 17034 0 _103_
rlabel metal1 4636 16014 4636 16014 0 _104_
rlabel metal1 18124 3706 18124 3706 0 _105_
rlabel metal1 16698 7854 16698 7854 0 _106_
rlabel metal1 15272 12682 15272 12682 0 _107_
rlabel metal2 11546 14654 11546 14654 0 _108_
rlabel metal1 13570 14246 13570 14246 0 _109_
rlabel metal1 17342 11730 17342 11730 0 _110_
rlabel metal1 10718 12852 10718 12852 0 _111_
rlabel metal1 10304 11186 10304 11186 0 _112_
rlabel metal2 12926 11356 12926 11356 0 _113_
rlabel metal1 13192 7514 13192 7514 0 _114_
rlabel metal1 12926 5678 12926 5678 0 _115_
rlabel metal1 15140 4250 15140 4250 0 _116_
rlabel metal2 8970 8534 8970 8534 0 _117_
rlabel metal2 16238 4794 16238 4794 0 _118_
rlabel metal2 16698 3808 16698 3808 0 _119_
rlabel metal1 14766 3468 14766 3468 0 _120_
rlabel metal1 15226 13838 15226 13838 0 _121_
rlabel metal2 4830 4862 4830 4862 0 _122_
rlabel metal2 874 4964 874 4964 0 _123_
rlabel metal1 1012 3162 1012 3162 0 _124_
rlabel metal1 13938 16626 13938 16626 0 _125_
rlabel metal2 13110 14620 13110 14620 0 _126_
rlabel metal1 15042 13940 15042 13940 0 _127_
rlabel metal2 11638 6256 11638 6256 0 _128_
rlabel metal1 15410 12614 15410 12614 0 _129_
rlabel metal2 11822 12784 11822 12784 0 _130_
rlabel metal2 18078 14620 18078 14620 0 _131_
rlabel metal1 16146 13702 16146 13702 0 _132_
rlabel metal1 13386 14450 13386 14450 0 _133_
rlabel metal1 10120 15130 10120 15130 0 _134_
rlabel metal2 12098 16116 12098 16116 0 _135_
rlabel metal1 5428 2618 5428 2618 0 _136_
rlabel metal1 3358 5780 3358 5780 0 _137_
rlabel metal1 5474 4250 5474 4250 0 _138_
rlabel metal1 5980 6358 5980 6358 0 _139_
rlabel metal2 2990 3264 2990 3264 0 _140_
rlabel metal2 4738 4828 4738 4828 0 _141_
rlabel metal1 1886 5338 1886 5338 0 _142_
rlabel via1 4278 3706 4278 3706 0 _143_
rlabel metal2 5198 4216 5198 4216 0 _144_
rlabel metal2 4186 3366 4186 3366 0 _145_
rlabel metal2 2806 15266 2806 15266 0 _146_
rlabel metal2 9798 4692 9798 4692 0 _147_
rlabel metal2 13202 4692 13202 4692 0 _148_
rlabel metal1 8096 9010 8096 9010 0 _149_
rlabel metal1 8004 8602 8004 8602 0 _150_
rlabel metal2 8326 8772 8326 8772 0 _151_
rlabel metal1 16054 12750 16054 12750 0 _152_
rlabel metal1 16330 12716 16330 12716 0 _153_
rlabel metal1 17020 12410 17020 12410 0 _154_
rlabel metal2 2898 9316 2898 9316 0 _155_
rlabel metal2 1058 8636 1058 8636 0 _156_
rlabel metal1 3542 1326 3542 1326 0 _157_
rlabel viali 3449 1394 3449 1394 0 _158_
rlabel metal2 10350 1836 10350 1836 0 _159_
rlabel metal1 10135 1394 10135 1394 0 _160_
rlabel metal1 11132 10574 11132 10574 0 _161_
rlabel metal2 9706 13124 9706 13124 0 _162_
rlabel metal1 12650 17204 12650 17204 0 _163_
rlabel metal1 12742 16762 12742 16762 0 _164_
rlabel metal2 13110 1564 13110 1564 0 _165_
rlabel metal1 13417 1394 13417 1394 0 _166_
rlabel metal1 15226 8398 15226 8398 0 _167_
rlabel metal2 15226 9044 15226 9044 0 _168_
rlabel metal1 3772 14586 3772 14586 0 _169_
rlabel metal1 3818 13498 3818 13498 0 _170_
rlabel metal1 6026 11798 6026 11798 0 _171_
rlabel metal1 6302 12342 6302 12342 0 _172_
rlabel metal2 5566 11084 5566 11084 0 _173_
rlabel metal2 4738 9180 4738 9180 0 _174_
rlabel metal2 4646 9180 4646 9180 0 _175_
rlabel metal1 4968 9146 4968 9146 0 _176_
rlabel metal2 2806 4454 2806 4454 0 _177_
rlabel metal2 2622 4420 2622 4420 0 _178_
rlabel metal1 6578 4046 6578 4046 0 _179_
rlabel viali 8142 4658 8142 4658 0 _180_
rlabel metal1 7498 4080 7498 4080 0 _181_
rlabel metal2 2438 17340 2438 17340 0 _182_
rlabel metal2 1978 17510 1978 17510 0 _183_
rlabel metal1 5520 17034 5520 17034 0 _184_
rlabel metal1 17526 2618 17526 2618 0 _185_
rlabel metal2 18170 4012 18170 4012 0 _186_
rlabel metal2 18354 3740 18354 3740 0 _187_
rlabel metal2 17894 9724 17894 9724 0 _188_
rlabel metal2 17802 9962 17802 9962 0 _189_
rlabel metal2 17342 8211 17342 8211 0 _190_
rlabel metal1 18308 6970 18308 6970 0 _191_
rlabel metal1 18078 6970 18078 6970 0 _192_
rlabel metal1 17434 7956 17434 7956 0 _193_
rlabel metal1 13248 15674 13248 15674 0 _194_
rlabel metal1 13156 14382 13156 14382 0 _195_
rlabel metal2 12834 7276 12834 7276 0 _196_
rlabel metal1 11546 5780 11546 5780 0 _197_
rlabel metal1 13202 4658 13202 4658 0 _198_
rlabel metal1 8970 5270 8970 5270 0 _199_
rlabel metal1 9200 7378 9200 7378 0 _200_
rlabel metal1 15134 1428 15134 1428 0 _201_
rlabel via1 15041 1394 15041 1394 0 _202_
rlabel metal1 11178 15912 11178 15912 0 clknet_0__037_
rlabel metal1 11316 11526 11316 11526 0 clknet_0_divider.out
rlabel metal1 15134 15334 15134 15334 0 clknet_0_divider2.out
rlabel metal1 5658 17714 5658 17714 0 clknet_0_ext_clk
rlabel metal1 9660 15606 9660 15606 0 clknet_0_net11
rlabel metal2 7038 10846 7038 10846 0 clknet_0_pll_clk
rlabel metal1 15272 8806 15272 8806 0 clknet_0_pll_clk90
rlabel metal2 9154 14144 9154 14144 0 clknet_1_0__leaf__037_
rlabel metal1 11822 9010 11822 9010 0 clknet_1_0__leaf_divider.out
rlabel metal1 14996 17714 14996 17714 0 clknet_1_0__leaf_divider2.out
rlabel metal2 5290 17306 5290 17306 0 clknet_1_0__leaf_ext_clk
rlabel metal1 4324 6630 4324 6630 0 clknet_1_0__leaf_pll_clk
rlabel metal1 16192 8466 16192 8466 0 clknet_1_0__leaf_pll_clk90
rlabel metal2 10350 17136 10350 17136 0 clknet_1_1__leaf__037_
rlabel metal1 9246 10234 9246 10234 0 clknet_1_1__leaf_divider.out
rlabel metal1 17296 14450 17296 14450 0 clknet_1_1__leaf_divider2.out
rlabel metal2 6854 16218 6854 16218 0 clknet_1_1__leaf_ext_clk
rlabel metal1 8280 15674 8280 15674 0 clknet_1_1__leaf_net11
rlabel metal2 3634 10404 3634 10404 0 clknet_1_1__leaf_pll_clk
rlabel metal1 10442 12308 10442 12308 0 clknet_1_1__leaf_pll_clk90
rlabel metal1 7406 16014 7406 16014 0 core_clk
rlabel metal1 10212 4658 10212 4658 0 divider.even_0.N\[0\]
rlabel via1 5842 12274 5842 12274 0 divider.even_0.N\[1\]
rlabel metal1 3036 9078 3036 9078 0 divider.even_0.N\[2\]
rlabel metal1 1380 17170 1380 17170 0 divider.even_0.counter\[0\]
rlabel metal1 1265 17238 1265 17238 0 divider.even_0.counter\[1\]
rlabel metal1 2208 17102 2208 17102 0 divider.even_0.counter\[2\]
rlabel metal1 7176 10438 7176 10438 0 divider.even_0.out_counter
rlabel metal1 4922 14926 4922 14926 0 divider.even_0.resetb
rlabel metal1 3082 3604 3082 3604 0 divider.odd_0.counter2\[0\]
rlabel metal1 5474 1394 5474 1394 0 divider.odd_0.counter2\[1\]
rlabel metal1 2898 3967 2898 3967 0 divider.odd_0.counter2\[2\]
rlabel metal2 9614 5406 9614 5406 0 divider.odd_0.counter\[0\]
rlabel metal1 8924 4658 8924 4658 0 divider.odd_0.counter\[1\]
rlabel metal1 8096 4046 8096 4046 0 divider.odd_0.counter\[2\]
rlabel metal1 1656 10778 1656 10778 0 divider.odd_0.initial_begin\[0\]
rlabel metal1 1150 12274 1150 12274 0 divider.odd_0.initial_begin\[1\]
rlabel metal1 2116 10234 2116 10234 0 divider.odd_0.initial_begin\[2\]
rlabel metal2 6670 12750 6670 12750 0 divider.odd_0.old_N\[0\]
rlabel metal1 5612 12274 5612 12274 0 divider.odd_0.old_N\[1\]
rlabel metal1 4968 9486 4968 9486 0 divider.odd_0.old_N\[2\]
rlabel metal1 8786 7276 8786 7276 0 divider.odd_0.out_counter
rlabel metal1 6900 5134 6900 5134 0 divider.odd_0.out_counter2
rlabel metal2 6946 10540 6946 10540 0 divider.odd_0.rst_pulse
rlabel metal1 9706 9146 9706 9146 0 divider.out
rlabel metal1 11270 6426 11270 6426 0 divider.syncNp\[0\]
rlabel metal1 10327 8058 10327 8058 0 divider.syncNp\[1\]
rlabel metal1 10534 9384 10534 9384 0 divider.syncNp\[2\]
rlabel metal1 16376 14246 16376 14246 0 divider2.even_0.N\[0\]
rlabel via1 17733 15878 17733 15878 0 divider2.even_0.N\[1\]
rlabel metal2 14214 14705 14214 14705 0 divider2.even_0.N\[2\]
rlabel metal2 17894 1904 17894 1904 0 divider2.even_0.counter\[0\]
rlabel metal1 17480 1394 17480 1394 0 divider2.even_0.counter\[1\]
rlabel metal1 16468 1326 16468 1326 0 divider2.even_0.counter\[2\]
rlabel metal1 17457 6086 17457 6086 0 divider2.even_0.out_counter
rlabel metal1 12650 16422 12650 16422 0 divider2.odd_0.counter2\[0\]
rlabel metal2 13110 16439 13110 16439 0 divider2.odd_0.counter2\[1\]
rlabel metal1 12558 17102 12558 17102 0 divider2.odd_0.counter2\[2\]
rlabel metal1 14168 2074 14168 2074 0 divider2.odd_0.counter\[0\]
rlabel metal1 11730 5644 11730 5644 0 divider2.odd_0.counter\[1\]
rlabel metal1 13616 1938 13616 1938 0 divider2.odd_0.counter\[2\]
rlabel metal1 10902 12614 10902 12614 0 divider2.odd_0.initial_begin\[0\]
rlabel metal1 11661 11322 11661 11322 0 divider2.odd_0.initial_begin\[1\]
rlabel metal1 11270 12274 11270 12274 0 divider2.odd_0.initial_begin\[2\]
rlabel metal1 17710 8602 17710 8602 0 divider2.odd_0.old_N\[0\]
rlabel metal2 17434 10132 17434 10132 0 divider2.odd_0.old_N\[1\]
rlabel metal1 17664 6834 17664 6834 0 divider2.odd_0.old_N\[2\]
rlabel metal1 17296 12750 17296 12750 0 divider2.odd_0.out_counter
rlabel metal2 17618 13090 17618 13090 0 divider2.odd_0.out_counter2
rlabel metal1 14766 18258 14766 18258 0 divider2.odd_0.rst_pulse
rlabel metal2 16330 14212 16330 14212 0 divider2.out
rlabel metal2 17986 14212 17986 14212 0 divider2.syncNp\[0\]
rlabel via1 17917 15130 17917 15130 0 divider2.syncNp\[1\]
rlabel metal1 17020 17646 17020 17646 0 divider2.syncNp\[2\]
rlabel metal1 3956 18394 3956 18394 0 ext_clk
rlabel metal2 18446 1581 18446 1581 0 ext_clk_sel
rlabel metal2 7038 15232 7038 15232 0 ext_clk_syncd
rlabel metal1 5796 16218 5796 16218 0 ext_clk_syncd_pre
rlabel metal2 18446 18479 18446 18479 0 ext_reset
rlabel metal1 17342 1938 17342 1938 0 net1
rlabel metal1 17342 7514 17342 7514 0 net10
rlabel metal1 9384 15130 9384 15130 0 net11
rlabel metal2 12926 17952 12926 17952 0 net12
rlabel metal2 17526 17340 17526 17340 0 net13
rlabel metal1 13800 2550 13800 2550 0 net14
rlabel metal1 11960 4998 11960 4998 0 net15
rlabel metal1 17940 2414 17940 2414 0 net16
rlabel metal1 14996 16558 14996 16558 0 net17
rlabel metal2 3358 2176 3358 2176 0 net18
rlabel metal1 2208 6222 2208 6222 0 net19
rlabel metal2 6026 17714 6026 17714 0 net2
rlabel metal2 2070 3434 2070 3434 0 net20
rlabel metal1 2162 17034 2162 17034 0 net21
rlabel metal1 8694 11152 8694 11152 0 net22
rlabel metal1 11638 4624 11638 4624 0 net23
rlabel metal2 9246 6800 9246 6800 0 net24
rlabel metal2 6854 3485 6854 3485 0 net25
rlabel metal1 1242 6800 1242 6800 0 net26
rlabel metal1 3029 11254 3029 11254 0 net27
rlabel metal1 5842 5848 5842 5848 0 net28
rlabel metal2 12190 5984 12190 5984 0 net29
rlabel metal1 2576 9894 2576 9894 0 net3
rlabel metal1 12006 8398 12006 8398 0 net30
rlabel metal2 16514 16082 16514 16082 0 net31
rlabel metal1 6532 17102 6532 17102 0 net32
rlabel metal1 11270 13906 11270 13906 0 net33
rlabel metal2 16146 11220 16146 11220 0 net34
rlabel metal2 9982 11628 9982 11628 0 net35
rlabel metal2 5198 5508 5198 5508 0 net36
rlabel metal1 5244 7922 5244 7922 0 net37
rlabel metal2 1702 12546 1702 12546 0 net38
rlabel metal1 7820 17714 7820 17714 0 net39
rlabel metal2 5474 17544 5474 17544 0 net4
rlabel metal1 9798 16626 9798 16626 0 net40
rlabel metal1 6946 17170 6946 17170 0 net41
rlabel metal1 16744 15674 16744 15674 0 net42
rlabel metal1 16836 14382 16836 14382 0 net43
rlabel metal1 8234 17646 8234 17646 0 net44
rlabel metal2 5566 14654 5566 14654 0 net45
rlabel metal1 7038 14042 7038 14042 0 net46
rlabel metal1 9292 16218 9292 16218 0 net47
rlabel metal1 18032 13974 18032 13974 0 net5
rlabel metal1 16560 14926 16560 14926 0 net6
rlabel metal1 17480 16762 17480 16762 0 net7
rlabel metal1 17710 3162 17710 3162 0 net8
rlabel metal1 12006 7854 12006 7854 0 net9
rlabel metal2 8234 11458 8234 11458 0 pll_clk
rlabel metal1 18492 8602 18492 8602 0 pll_clk90
rlabel metal1 10626 12172 10626 12172 0 pll_clk_sel
rlabel metal1 782 10098 782 10098 0 porb
rlabel metal1 9637 17850 9637 17850 0 reset_delay\[0\]
rlabel metal1 8073 16762 8073 16762 0 reset_delay\[1\]
rlabel metal2 8786 16524 8786 16524 0 reset_delay\[2\]
rlabel metal1 1518 18190 1518 18190 0 resetb
rlabel metal1 13110 17646 13110 17646 0 resetb_sync
rlabel via2 18446 11203 18446 11203 0 sel2[0]
rlabel metal1 18768 14790 18768 14790 0 sel2[1]
rlabel metal2 18446 16371 18446 16371 0 sel2[2]
rlabel metal1 18538 2958 18538 2958 0 sel[0]
rlabel metal2 18446 6035 18446 6035 0 sel[1]
rlabel metal2 17986 8041 17986 8041 0 sel[2]
rlabel metal1 7636 12138 7636 12138 0 use_pll_first
rlabel metal1 9752 14994 9752 14994 0 use_pll_second
rlabel metal1 10580 16490 10580 16490 0 user_clk
rlabel metal2 9982 17374 9982 17374 0 user_clk_buffered
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
