magic
tech sky130A
timestamp 1605994897
<< pwell >>
rect -154 -229 154 229
<< mvnmos >>
rect -40 -100 40 100
<< mvndiff >>
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
<< mvndiffc >>
rect -63 -94 -46 94
rect 46 -94 63 94
<< mvpsubdiff >>
rect -136 205 136 211
rect -136 188 -82 205
rect 82 188 136 205
rect -136 182 136 188
rect -136 -182 -107 182
rect 107 157 136 182
rect 107 -157 113 157
rect 130 -157 136 157
rect 107 -182 136 -157
rect -136 -188 136 -182
rect -136 -205 -82 -188
rect 82 -205 136 -188
rect -136 -211 136 -205
<< mvpsubdiffcont >>
rect -82 188 82 205
rect 113 -157 130 157
rect -82 -205 82 -188
<< poly >>
rect -40 136 40 144
rect -40 119 -32 136
rect 32 119 40 136
rect -40 100 40 119
rect -40 -119 40 -100
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect -40 -144 40 -136
<< polycont >>
rect -32 119 32 136
rect -32 -136 32 -119
<< locali >>
rect -130 188 -82 205
rect 82 188 130 205
rect -130 -188 -113 188
rect 113 157 130 188
rect -40 119 -32 136
rect 32 119 40 136
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect -40 -136 -32 -119
rect 32 -136 40 -119
rect 113 -188 130 -157
rect -130 -205 -82 -188
rect 82 -205 130 -188
<< viali >>
rect -32 119 32 136
rect -63 -94 -46 94
rect 46 -94 63 94
rect -32 -136 32 -119
<< metal1 >>
rect -38 136 38 139
rect -38 119 -32 136
rect 32 119 38 136
rect -38 116 38 119
rect -66 94 -43 100
rect -66 -94 -63 94
rect -46 -94 -43 94
rect -66 -100 -43 -94
rect 43 94 66 100
rect 43 -94 46 94
rect 63 -94 66 94
rect 43 -100 66 -94
rect -38 -119 38 -116
rect -38 -136 -32 -119
rect 32 -136 38 -119
rect -38 -139 38 -136
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -121 -196 121 196
string parameters w 2.00 l 0.80 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
