magic
tech sky130A
timestamp 1637147503
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4365 -480 4421 240
rect 4963 -480 5019 240
rect 5561 -480 5617 240
rect 6159 -480 6215 240
rect 6757 -480 6813 240
rect 7355 -480 7411 240
rect 7953 -480 8009 240
rect 8505 -480 8561 240
rect 9103 -480 9159 240
rect 9701 -480 9757 240
rect 10299 -480 10355 240
rect 10897 -480 10953 240
rect 11495 -480 11551 240
rect 12093 -480 12149 240
rect 12645 -480 12701 240
rect 13243 -480 13299 240
rect 13841 -480 13897 240
rect 14439 -480 14495 240
rect 15037 -480 15093 240
rect 15635 -480 15691 240
rect 16187 -480 16243 240
rect 16785 -480 16841 240
rect 17383 -480 17439 240
rect 17981 -480 18037 240
rect 18579 -480 18635 240
rect 19177 -480 19233 240
rect 19775 -480 19831 240
rect 20327 -480 20383 240
rect 20925 -480 20981 240
rect 21523 -480 21579 240
rect 22121 -480 22177 240
rect 22719 -480 22775 240
rect 23317 -480 23373 240
rect 23915 -480 23971 240
rect 24467 -480 24523 240
rect 25065 -480 25121 240
rect 25663 -480 25719 240
rect 26261 -480 26317 240
rect 26859 -480 26915 240
rect 27457 -480 27513 240
rect 28009 -480 28065 240
rect 28607 -480 28663 240
rect 29205 -480 29261 240
rect 29803 -480 29859 240
rect 30401 -480 30457 240
rect 30999 -480 31055 240
rect 31597 -480 31653 240
rect 32149 -480 32205 240
rect 32747 -480 32803 240
rect 33345 -480 33401 240
rect 33943 -480 33999 240
rect 34541 -480 34597 240
rect 35139 -480 35195 240
rect 35737 -480 35793 240
rect 36289 -480 36345 240
rect 36887 -480 36943 240
rect 37485 -480 37541 240
rect 38083 -480 38139 240
rect 38681 -480 38737 240
rect 39279 -480 39335 240
rect 39831 -480 39887 240
rect 40429 -480 40485 240
rect 41027 -480 41083 240
rect 41625 -480 41681 240
rect 42223 -480 42279 240
rect 42821 -480 42877 240
rect 43419 -480 43475 240
rect 43971 -480 44027 240
rect 44569 -480 44625 240
rect 45167 -480 45223 240
rect 45765 -480 45821 240
rect 46363 -480 46419 240
rect 46961 -480 47017 240
rect 47559 -480 47615 240
rect 48111 -480 48167 240
rect 48709 -480 48765 240
rect 49307 -480 49363 240
rect 49905 -480 49961 240
rect 50503 -480 50559 240
rect 51101 -480 51157 240
rect 51653 -480 51709 240
rect 52251 -480 52307 240
rect 52849 -480 52905 240
rect 53447 -480 53503 240
rect 54045 -480 54101 240
rect 54643 -480 54699 240
rect 55241 -480 55297 240
rect 55793 -480 55849 240
rect 56391 -480 56447 240
rect 56989 -480 57045 240
rect 57587 -480 57643 240
rect 58185 -480 58241 240
rect 58783 -480 58839 240
rect 59381 -480 59437 240
rect 59933 -480 59989 240
rect 60531 -480 60587 240
rect 61129 -480 61185 240
rect 61727 -480 61783 240
rect 62325 -480 62381 240
rect 62923 -480 62979 240
rect 63475 -480 63531 240
rect 64073 -480 64129 240
rect 64671 -480 64727 240
rect 65269 -480 65325 240
rect 65867 -480 65923 240
rect 66465 -480 66521 240
rect 67063 -480 67119 240
rect 67615 -480 67671 240
rect 68213 -480 68269 240
rect 68811 -480 68867 240
rect 69409 -480 69465 240
rect 70007 -480 70063 240
rect 70605 -480 70661 240
rect 71203 -480 71259 240
rect 71755 -480 71811 240
rect 72353 -480 72409 240
rect 72951 -480 73007 240
rect 73549 -480 73605 240
rect 74147 -480 74203 240
rect 74745 -480 74801 240
rect 75297 -480 75353 240
rect 75895 -480 75951 240
rect 76493 -480 76549 240
rect 77091 -480 77147 240
rect 77689 -480 77745 240
rect 78287 -480 78343 240
rect 78885 -480 78941 240
rect 79437 -480 79493 240
rect 80035 -480 80091 240
rect 80633 -480 80689 240
rect 81231 -480 81287 240
rect 81829 -480 81885 240
rect 82427 -480 82483 240
rect 83025 -480 83081 240
rect 83577 -480 83633 240
rect 84175 -480 84231 240
rect 84773 -480 84829 240
rect 85371 -480 85427 240
rect 85969 -480 86025 240
rect 86567 -480 86623 240
rect 87119 -480 87175 240
rect 87717 -480 87773 240
rect 88315 -480 88371 240
rect 88913 -480 88969 240
rect 89511 -480 89567 240
rect 90109 -480 90165 240
rect 90707 -480 90763 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92455 -480 92511 240
rect 93053 -480 93109 240
rect 93651 -480 93707 240
rect 94249 -480 94305 240
rect 94847 -480 94903 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98941 -480 98997 240
rect 99539 -480 99595 240
rect 100137 -480 100193 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103081 -480 103137 240
rect 103679 -480 103735 240
rect 104277 -480 104333 240
rect 104875 -480 104931 240
rect 105473 -480 105529 240
rect 106071 -480 106127 240
rect 106669 -480 106725 240
rect 107221 -480 107277 240
rect 107819 -480 107875 240
rect 108417 -480 108473 240
rect 109015 -480 109071 240
rect 109613 -480 109669 240
rect 110211 -480 110267 240
rect 110763 -480 110819 240
rect 111361 -480 111417 240
rect 111959 -480 112015 240
rect 112557 -480 112613 240
rect 113155 -480 113211 240
rect 113753 -480 113809 240
rect 114351 -480 114407 240
rect 114903 -480 114959 240
rect 115501 -480 115557 240
rect 116099 -480 116155 240
rect 116697 -480 116753 240
rect 117295 -480 117351 240
rect 117893 -480 117949 240
rect 118491 -480 118547 240
rect 119043 -480 119099 240
rect 119641 -480 119697 240
rect 120239 -480 120295 240
rect 120837 -480 120893 240
rect 121435 -480 121491 240
rect 122033 -480 122089 240
rect 122585 -480 122641 240
rect 123183 -480 123239 240
rect 123781 -480 123837 240
rect 124379 -480 124435 240
rect 124977 -480 125033 240
rect 125575 -480 125631 240
rect 126173 -480 126229 240
rect 126725 -480 126781 240
rect 127323 -480 127379 240
rect 127921 -480 127977 240
rect 128519 -480 128575 240
rect 129117 -480 129173 240
rect 129715 -480 129771 240
rect 130313 -480 130369 240
rect 130865 -480 130921 240
rect 131463 -480 131519 240
rect 132061 -480 132117 240
rect 132659 -480 132715 240
rect 133257 -480 133313 240
rect 133855 -480 133911 240
rect 134407 -480 134463 240
rect 135005 -480 135061 240
rect 135603 -480 135659 240
rect 136201 -480 136257 240
rect 136799 -480 136855 240
rect 137397 -480 137453 240
rect 137995 -480 138051 240
rect 138547 -480 138603 240
rect 139145 -480 139201 240
rect 139743 -480 139799 240
rect 140341 -480 140397 240
rect 140939 -480 140995 240
rect 141537 -480 141593 240
rect 142135 -480 142191 240
rect 142687 -480 142743 240
rect 143285 -480 143341 240
rect 143883 -480 143939 240
rect 144481 -480 144537 240
rect 145079 -480 145135 240
rect 145677 -480 145733 240
rect 146275 -480 146331 240
rect 146827 -480 146883 240
rect 147425 -480 147481 240
rect 148023 -480 148079 240
rect 148621 -480 148677 240
rect 149219 -480 149275 240
rect 149817 -480 149873 240
rect 150369 -480 150425 240
rect 150967 -480 151023 240
rect 151565 -480 151621 240
rect 152163 -480 152219 240
rect 152761 -480 152817 240
rect 153359 -480 153415 240
rect 153957 -480 154013 240
rect 154509 -480 154565 240
rect 155107 -480 155163 240
rect 155705 -480 155761 240
rect 156303 -480 156359 240
rect 156901 -480 156957 240
rect 157499 -480 157555 240
rect 158097 -480 158153 240
rect 158649 -480 158705 240
rect 159247 -480 159303 240
rect 159845 -480 159901 240
rect 160443 -480 160499 240
rect 161041 -480 161097 240
rect 161639 -480 161695 240
rect 162191 -480 162247 240
rect 162789 -480 162845 240
rect 163387 -480 163443 240
rect 163985 -480 164041 240
rect 164583 -480 164639 240
rect 165181 -480 165237 240
rect 165779 -480 165835 240
rect 166331 -480 166387 240
rect 166929 -480 166985 240
rect 167527 -480 167583 240
rect 168125 -480 168181 240
rect 168723 -480 168779 240
rect 169321 -480 169377 240
rect 169919 -480 169975 240
rect 170471 -480 170527 240
rect 171069 -480 171125 240
rect 171667 -480 171723 240
rect 172265 -480 172321 240
rect 172863 -480 172919 240
rect 173461 -480 173517 240
rect 174013 -480 174069 240
rect 174611 -480 174667 240
rect 175209 -480 175265 240
rect 175807 -480 175863 240
rect 176405 -480 176461 240
rect 177003 -480 177059 240
rect 177601 -480 177657 240
rect 178153 -480 178209 240
rect 178751 -480 178807 240
rect 179349 -480 179405 240
rect 179947 -480 180003 240
rect 180545 -480 180601 240
rect 181143 -480 181199 240
rect 181741 -480 181797 240
rect 182293 -480 182349 240
rect 182891 -480 182947 240
rect 183489 -480 183545 240
rect 184087 -480 184143 240
rect 184685 -480 184741 240
rect 185283 -480 185339 240
rect 185835 -480 185891 240
rect 186433 -480 186489 240
rect 187031 -480 187087 240
rect 187629 -480 187685 240
rect 188227 -480 188283 240
rect 188825 -480 188881 240
rect 189423 -480 189479 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192367 -480 192423 240
rect 192965 -480 193021 240
rect 193563 -480 193619 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197657 -480 197713 240
rect 198255 -480 198311 240
rect 198853 -480 198909 240
rect 199451 -480 199507 240
rect 200049 -480 200105 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201797 -480 201853 240
rect 202395 -480 202451 240
rect 202993 -480 203049 240
rect 203591 -480 203647 240
rect 204189 -480 204245 240
rect 204787 -480 204843 240
rect 205385 -480 205441 240
rect 205937 -480 205993 240
rect 206535 -480 206591 240
rect 207133 -480 207189 240
rect 207731 -480 207787 240
rect 208329 -480 208385 240
rect 208927 -480 208983 240
rect 209479 -480 209535 240
rect 210077 -480 210133 240
rect 210675 -480 210731 240
rect 211273 -480 211329 240
rect 211871 -480 211927 240
rect 212469 -480 212525 240
rect 213067 -480 213123 240
rect 213619 -480 213675 240
rect 214217 -480 214273 240
rect 214815 -480 214871 240
rect 215413 -480 215469 240
rect 216011 -480 216067 240
rect 216609 -480 216665 240
rect 217207 -480 217263 240
rect 217759 -480 217815 240
rect 218357 -480 218413 240
rect 218955 -480 219011 240
rect 219553 -480 219609 240
rect 220151 -480 220207 240
rect 220749 -480 220805 240
rect 221301 -480 221357 240
rect 221899 -480 221955 240
rect 222497 -480 222553 240
rect 223095 -480 223151 240
rect 223693 -480 223749 240
rect 224291 -480 224347 240
rect 224889 -480 224945 240
rect 225441 -480 225497 240
rect 226039 -480 226095 240
rect 226637 -480 226693 240
rect 227235 -480 227291 240
rect 227833 -480 227889 240
rect 228431 -480 228487 240
rect 229029 -480 229085 240
rect 229581 -480 229637 240
rect 230179 -480 230235 240
rect 230777 -480 230833 240
rect 231375 -480 231431 240
rect 231973 -480 232029 240
rect 232571 -480 232627 240
rect 233123 -480 233179 240
rect 233721 -480 233777 240
rect 234319 -480 234375 240
rect 234917 -480 234973 240
rect 235515 -480 235571 240
rect 236113 -480 236169 240
rect 236711 -480 236767 240
rect 237263 -480 237319 240
rect 237861 -480 237917 240
rect 238459 -480 238515 240
rect 239057 -480 239113 240
rect 239655 -480 239711 240
rect 240253 -480 240309 240
rect 240851 -480 240907 240
rect 241403 -480 241459 240
rect 242001 -480 242057 240
rect 242599 -480 242655 240
rect 243197 -480 243253 240
rect 243795 -480 243851 240
rect 244393 -480 244449 240
rect 244945 -480 245001 240
rect 245543 -480 245599 240
rect 246141 -480 246197 240
rect 246739 -480 246795 240
rect 247337 -480 247393 240
rect 247935 -480 247991 240
rect 248533 -480 248589 240
rect 249085 -480 249141 240
rect 249683 -480 249739 240
rect 250281 -480 250337 240
rect 250879 -480 250935 240
rect 251477 -480 251533 240
rect 252075 -480 252131 240
rect 252673 -480 252729 240
rect 253225 -480 253281 240
rect 253823 -480 253879 240
rect 254421 -480 254477 240
rect 255019 -480 255075 240
rect 255617 -480 255673 240
rect 256215 -480 256271 240
rect 256767 -480 256823 240
rect 257365 -480 257421 240
rect 257963 -480 258019 240
rect 258561 -480 258617 240
rect 259159 -480 259215 240
rect 259757 -480 259813 240
rect 260355 -480 260411 240
rect 260907 -480 260963 240
rect 261505 -480 261561 240
rect 262103 -480 262159 240
rect 262701 -480 262757 240
rect 263299 -480 263355 240
rect 263897 -480 263953 240
rect 264495 -480 264551 240
rect 265047 -480 265103 240
rect 265645 -480 265701 240
rect 266243 -480 266299 240
rect 266841 -480 266897 240
rect 267439 -480 267495 240
rect 268037 -480 268093 240
rect 268589 -480 268645 240
rect 269187 -480 269243 240
rect 269785 -480 269841 240
rect 270383 -480 270439 240
rect 270981 -480 271037 240
rect 271579 -480 271635 240
rect 272177 -480 272233 240
rect 272729 -480 272785 240
rect 273327 -480 273383 240
rect 273925 -480 273981 240
rect 274523 -480 274579 240
rect 275121 -480 275177 240
rect 275719 -480 275775 240
rect 276317 -480 276373 240
rect 276869 -480 276925 240
rect 277467 -480 277523 240
rect 278065 -480 278121 240
rect 278663 -480 278719 240
rect 279261 -480 279317 240
rect 279859 -480 279915 240
rect 280411 -480 280467 240
rect 281009 -480 281065 240
rect 281607 -480 281663 240
rect 282205 -480 282261 240
rect 282803 -480 282859 240
rect 283401 -480 283457 240
rect 283999 -480 284055 240
rect 284551 -480 284607 240
rect 285149 -480 285205 240
rect 285747 -480 285803 240
rect 286345 -480 286401 240
rect 286943 -480 286999 240
rect 287541 -480 287597 240
rect 288139 -480 288195 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect -480 348610 240 348730
rect 291760 348542 292480 348662
rect -480 342082 240 342202
rect 291760 341878 292480 341998
rect -480 335554 240 335674
rect 291760 335282 292480 335402
rect -480 329026 240 329146
rect 291760 328618 292480 328738
rect -480 322498 240 322618
rect 291760 321954 292480 322074
rect -480 315970 240 316090
rect 291760 315358 292480 315478
rect -480 309510 240 309630
rect 291760 308694 292480 308814
rect -480 302982 240 303102
rect 291760 302030 292480 302150
rect -480 296454 240 296574
rect 291760 295434 292480 295554
rect -480 289926 240 290046
rect 291760 288770 292480 288890
rect -480 283398 240 283518
rect 291760 282106 292480 282226
rect -480 276870 240 276990
rect 291760 275510 292480 275630
rect -480 270342 240 270462
rect 291760 268846 292480 268966
rect -480 263882 240 264002
rect 291760 262182 292480 262302
rect -480 257354 240 257474
rect 291760 255586 292480 255706
rect -480 250826 240 250946
rect 291760 248922 292480 249042
rect -480 244298 240 244418
rect 291760 242258 292480 242378
rect -480 237770 240 237890
rect 291760 235662 292480 235782
rect -480 231242 240 231362
rect 291760 228998 292480 229118
rect -480 224714 240 224834
rect 291760 222334 292480 222454
rect -480 218254 240 218374
rect 291760 215738 292480 215858
rect -480 211726 240 211846
rect 291760 209074 292480 209194
rect -480 205198 240 205318
rect 291760 202410 292480 202530
rect -480 198670 240 198790
rect 291760 195814 292480 195934
rect -480 192142 240 192262
rect 291760 189150 292480 189270
rect -480 185614 240 185734
rect 291760 182486 292480 182606
rect -480 179154 240 179274
rect 291760 175890 292480 176010
rect -480 172626 240 172746
rect 291760 169226 292480 169346
rect -480 166098 240 166218
rect 291760 162562 292480 162682
rect -480 159570 240 159690
rect 291760 155966 292480 156086
rect -480 153042 240 153162
rect 291760 149302 292480 149422
rect -480 146514 240 146634
rect 291760 142638 292480 142758
rect -480 139986 240 140106
rect 291760 136042 292480 136162
rect -480 133526 240 133646
rect 291760 129378 292480 129498
rect -480 126998 240 127118
rect 291760 122714 292480 122834
rect -480 120470 240 120590
rect 291760 116118 292480 116238
rect -480 113942 240 114062
rect 291760 109454 292480 109574
rect -480 107414 240 107534
rect 291760 102790 292480 102910
rect -480 100886 240 101006
rect 291760 96194 292480 96314
rect -480 94358 240 94478
rect 291760 89530 292480 89650
rect -480 87898 240 88018
rect 291760 82866 292480 82986
rect -480 81370 240 81490
rect 291760 76270 292480 76390
rect -480 74842 240 74962
rect 291760 69606 292480 69726
rect -480 68314 240 68434
rect 291760 62942 292480 63062
rect -480 61786 240 61906
rect 291760 56346 292480 56466
rect -480 55258 240 55378
rect 291760 49682 292480 49802
rect -480 48730 240 48850
rect 291760 43018 292480 43138
rect -480 42270 240 42390
rect 291760 36422 292480 36542
rect -480 35742 240 35862
rect 291760 29758 292480 29878
rect -480 29214 240 29334
rect 291760 23094 292480 23214
rect -480 22686 240 22806
rect 291760 16498 292480 16618
rect -480 16158 240 16278
rect 291760 9834 292480 9954
rect -480 9630 240 9750
rect -480 3170 240 3290
rect 291760 3238 292480 3358
<< metal4 >>
rect -4363 355779 -4053 355795
rect -4363 355661 -4347 355779
rect -4229 355661 -4187 355779
rect -4069 355661 -4053 355779
rect -4363 355619 -4053 355661
rect -4363 355501 -4347 355619
rect -4229 355501 -4187 355619
rect -4069 355501 -4053 355619
rect -4363 340307 -4053 355501
rect -4363 340189 -4347 340307
rect -4229 340189 -4187 340307
rect -4069 340189 -4053 340307
rect -4363 340147 -4053 340189
rect -4363 340029 -4347 340147
rect -4229 340029 -4187 340147
rect -4069 340029 -4053 340147
rect -4363 322307 -4053 340029
rect -4363 322189 -4347 322307
rect -4229 322189 -4187 322307
rect -4069 322189 -4053 322307
rect -4363 322147 -4053 322189
rect -4363 322029 -4347 322147
rect -4229 322029 -4187 322147
rect -4069 322029 -4053 322147
rect -4363 304307 -4053 322029
rect -4363 304189 -4347 304307
rect -4229 304189 -4187 304307
rect -4069 304189 -4053 304307
rect -4363 304147 -4053 304189
rect -4363 304029 -4347 304147
rect -4229 304029 -4187 304147
rect -4069 304029 -4053 304147
rect -4363 286307 -4053 304029
rect -4363 286189 -4347 286307
rect -4229 286189 -4187 286307
rect -4069 286189 -4053 286307
rect -4363 286147 -4053 286189
rect -4363 286029 -4347 286147
rect -4229 286029 -4187 286147
rect -4069 286029 -4053 286147
rect -4363 268307 -4053 286029
rect -4363 268189 -4347 268307
rect -4229 268189 -4187 268307
rect -4069 268189 -4053 268307
rect -4363 268147 -4053 268189
rect -4363 268029 -4347 268147
rect -4229 268029 -4187 268147
rect -4069 268029 -4053 268147
rect -4363 250307 -4053 268029
rect -4363 250189 -4347 250307
rect -4229 250189 -4187 250307
rect -4069 250189 -4053 250307
rect -4363 250147 -4053 250189
rect -4363 250029 -4347 250147
rect -4229 250029 -4187 250147
rect -4069 250029 -4053 250147
rect -4363 232307 -4053 250029
rect -4363 232189 -4347 232307
rect -4229 232189 -4187 232307
rect -4069 232189 -4053 232307
rect -4363 232147 -4053 232189
rect -4363 232029 -4347 232147
rect -4229 232029 -4187 232147
rect -4069 232029 -4053 232147
rect -4363 214307 -4053 232029
rect -4363 214189 -4347 214307
rect -4229 214189 -4187 214307
rect -4069 214189 -4053 214307
rect -4363 214147 -4053 214189
rect -4363 214029 -4347 214147
rect -4229 214029 -4187 214147
rect -4069 214029 -4053 214147
rect -4363 196307 -4053 214029
rect -4363 196189 -4347 196307
rect -4229 196189 -4187 196307
rect -4069 196189 -4053 196307
rect -4363 196147 -4053 196189
rect -4363 196029 -4347 196147
rect -4229 196029 -4187 196147
rect -4069 196029 -4053 196147
rect -4363 178307 -4053 196029
rect -4363 178189 -4347 178307
rect -4229 178189 -4187 178307
rect -4069 178189 -4053 178307
rect -4363 178147 -4053 178189
rect -4363 178029 -4347 178147
rect -4229 178029 -4187 178147
rect -4069 178029 -4053 178147
rect -4363 160307 -4053 178029
rect -4363 160189 -4347 160307
rect -4229 160189 -4187 160307
rect -4069 160189 -4053 160307
rect -4363 160147 -4053 160189
rect -4363 160029 -4347 160147
rect -4229 160029 -4187 160147
rect -4069 160029 -4053 160147
rect -4363 142307 -4053 160029
rect -4363 142189 -4347 142307
rect -4229 142189 -4187 142307
rect -4069 142189 -4053 142307
rect -4363 142147 -4053 142189
rect -4363 142029 -4347 142147
rect -4229 142029 -4187 142147
rect -4069 142029 -4053 142147
rect -4363 124307 -4053 142029
rect -4363 124189 -4347 124307
rect -4229 124189 -4187 124307
rect -4069 124189 -4053 124307
rect -4363 124147 -4053 124189
rect -4363 124029 -4347 124147
rect -4229 124029 -4187 124147
rect -4069 124029 -4053 124147
rect -4363 106307 -4053 124029
rect -4363 106189 -4347 106307
rect -4229 106189 -4187 106307
rect -4069 106189 -4053 106307
rect -4363 106147 -4053 106189
rect -4363 106029 -4347 106147
rect -4229 106029 -4187 106147
rect -4069 106029 -4053 106147
rect -4363 88307 -4053 106029
rect -4363 88189 -4347 88307
rect -4229 88189 -4187 88307
rect -4069 88189 -4053 88307
rect -4363 88147 -4053 88189
rect -4363 88029 -4347 88147
rect -4229 88029 -4187 88147
rect -4069 88029 -4053 88147
rect -4363 70307 -4053 88029
rect -4363 70189 -4347 70307
rect -4229 70189 -4187 70307
rect -4069 70189 -4053 70307
rect -4363 70147 -4053 70189
rect -4363 70029 -4347 70147
rect -4229 70029 -4187 70147
rect -4069 70029 -4053 70147
rect -4363 52307 -4053 70029
rect -4363 52189 -4347 52307
rect -4229 52189 -4187 52307
rect -4069 52189 -4053 52307
rect -4363 52147 -4053 52189
rect -4363 52029 -4347 52147
rect -4229 52029 -4187 52147
rect -4069 52029 -4053 52147
rect -4363 34307 -4053 52029
rect -4363 34189 -4347 34307
rect -4229 34189 -4187 34307
rect -4069 34189 -4053 34307
rect -4363 34147 -4053 34189
rect -4363 34029 -4347 34147
rect -4229 34029 -4187 34147
rect -4069 34029 -4053 34147
rect -4363 16307 -4053 34029
rect -4363 16189 -4347 16307
rect -4229 16189 -4187 16307
rect -4069 16189 -4053 16307
rect -4363 16147 -4053 16189
rect -4363 16029 -4347 16147
rect -4229 16029 -4187 16147
rect -4069 16029 -4053 16147
rect -4363 -3533 -4053 16029
rect -3883 355299 -3573 355315
rect -3883 355181 -3867 355299
rect -3749 355181 -3707 355299
rect -3589 355181 -3573 355299
rect -3883 355139 -3573 355181
rect -3883 355021 -3867 355139
rect -3749 355021 -3707 355139
rect -3589 355021 -3573 355139
rect -3883 349307 -3573 355021
rect 6477 355299 6787 355795
rect 6477 355181 6493 355299
rect 6611 355181 6653 355299
rect 6771 355181 6787 355299
rect 6477 355139 6787 355181
rect 6477 355021 6493 355139
rect 6611 355021 6653 355139
rect 6771 355021 6787 355139
rect -3883 349189 -3867 349307
rect -3749 349189 -3707 349307
rect -3589 349189 -3573 349307
rect -3883 349147 -3573 349189
rect -3883 349029 -3867 349147
rect -3749 349029 -3707 349147
rect -3589 349029 -3573 349147
rect -3883 331307 -3573 349029
rect -3883 331189 -3867 331307
rect -3749 331189 -3707 331307
rect -3589 331189 -3573 331307
rect -3883 331147 -3573 331189
rect -3883 331029 -3867 331147
rect -3749 331029 -3707 331147
rect -3589 331029 -3573 331147
rect -3883 313307 -3573 331029
rect -3883 313189 -3867 313307
rect -3749 313189 -3707 313307
rect -3589 313189 -3573 313307
rect -3883 313147 -3573 313189
rect -3883 313029 -3867 313147
rect -3749 313029 -3707 313147
rect -3589 313029 -3573 313147
rect -3883 295307 -3573 313029
rect -3883 295189 -3867 295307
rect -3749 295189 -3707 295307
rect -3589 295189 -3573 295307
rect -3883 295147 -3573 295189
rect -3883 295029 -3867 295147
rect -3749 295029 -3707 295147
rect -3589 295029 -3573 295147
rect -3883 277307 -3573 295029
rect -3883 277189 -3867 277307
rect -3749 277189 -3707 277307
rect -3589 277189 -3573 277307
rect -3883 277147 -3573 277189
rect -3883 277029 -3867 277147
rect -3749 277029 -3707 277147
rect -3589 277029 -3573 277147
rect -3883 259307 -3573 277029
rect -3883 259189 -3867 259307
rect -3749 259189 -3707 259307
rect -3589 259189 -3573 259307
rect -3883 259147 -3573 259189
rect -3883 259029 -3867 259147
rect -3749 259029 -3707 259147
rect -3589 259029 -3573 259147
rect -3883 241307 -3573 259029
rect -3883 241189 -3867 241307
rect -3749 241189 -3707 241307
rect -3589 241189 -3573 241307
rect -3883 241147 -3573 241189
rect -3883 241029 -3867 241147
rect -3749 241029 -3707 241147
rect -3589 241029 -3573 241147
rect -3883 223307 -3573 241029
rect -3883 223189 -3867 223307
rect -3749 223189 -3707 223307
rect -3589 223189 -3573 223307
rect -3883 223147 -3573 223189
rect -3883 223029 -3867 223147
rect -3749 223029 -3707 223147
rect -3589 223029 -3573 223147
rect -3883 205307 -3573 223029
rect -3883 205189 -3867 205307
rect -3749 205189 -3707 205307
rect -3589 205189 -3573 205307
rect -3883 205147 -3573 205189
rect -3883 205029 -3867 205147
rect -3749 205029 -3707 205147
rect -3589 205029 -3573 205147
rect -3883 187307 -3573 205029
rect -3883 187189 -3867 187307
rect -3749 187189 -3707 187307
rect -3589 187189 -3573 187307
rect -3883 187147 -3573 187189
rect -3883 187029 -3867 187147
rect -3749 187029 -3707 187147
rect -3589 187029 -3573 187147
rect -3883 169307 -3573 187029
rect -3883 169189 -3867 169307
rect -3749 169189 -3707 169307
rect -3589 169189 -3573 169307
rect -3883 169147 -3573 169189
rect -3883 169029 -3867 169147
rect -3749 169029 -3707 169147
rect -3589 169029 -3573 169147
rect -3883 151307 -3573 169029
rect -3883 151189 -3867 151307
rect -3749 151189 -3707 151307
rect -3589 151189 -3573 151307
rect -3883 151147 -3573 151189
rect -3883 151029 -3867 151147
rect -3749 151029 -3707 151147
rect -3589 151029 -3573 151147
rect -3883 133307 -3573 151029
rect -3883 133189 -3867 133307
rect -3749 133189 -3707 133307
rect -3589 133189 -3573 133307
rect -3883 133147 -3573 133189
rect -3883 133029 -3867 133147
rect -3749 133029 -3707 133147
rect -3589 133029 -3573 133147
rect -3883 115307 -3573 133029
rect -3883 115189 -3867 115307
rect -3749 115189 -3707 115307
rect -3589 115189 -3573 115307
rect -3883 115147 -3573 115189
rect -3883 115029 -3867 115147
rect -3749 115029 -3707 115147
rect -3589 115029 -3573 115147
rect -3883 97307 -3573 115029
rect -3883 97189 -3867 97307
rect -3749 97189 -3707 97307
rect -3589 97189 -3573 97307
rect -3883 97147 -3573 97189
rect -3883 97029 -3867 97147
rect -3749 97029 -3707 97147
rect -3589 97029 -3573 97147
rect -3883 79307 -3573 97029
rect -3883 79189 -3867 79307
rect -3749 79189 -3707 79307
rect -3589 79189 -3573 79307
rect -3883 79147 -3573 79189
rect -3883 79029 -3867 79147
rect -3749 79029 -3707 79147
rect -3589 79029 -3573 79147
rect -3883 61307 -3573 79029
rect -3883 61189 -3867 61307
rect -3749 61189 -3707 61307
rect -3589 61189 -3573 61307
rect -3883 61147 -3573 61189
rect -3883 61029 -3867 61147
rect -3749 61029 -3707 61147
rect -3589 61029 -3573 61147
rect -3883 43307 -3573 61029
rect -3883 43189 -3867 43307
rect -3749 43189 -3707 43307
rect -3589 43189 -3573 43307
rect -3883 43147 -3573 43189
rect -3883 43029 -3867 43147
rect -3749 43029 -3707 43147
rect -3589 43029 -3573 43147
rect -3883 25307 -3573 43029
rect -3883 25189 -3867 25307
rect -3749 25189 -3707 25307
rect -3589 25189 -3573 25307
rect -3883 25147 -3573 25189
rect -3883 25029 -3867 25147
rect -3749 25029 -3707 25147
rect -3589 25029 -3573 25147
rect -3883 7307 -3573 25029
rect -3883 7189 -3867 7307
rect -3749 7189 -3707 7307
rect -3589 7189 -3573 7307
rect -3883 7147 -3573 7189
rect -3883 7029 -3867 7147
rect -3749 7029 -3707 7147
rect -3589 7029 -3573 7147
rect -3883 -3053 -3573 7029
rect -3403 354819 -3093 354835
rect -3403 354701 -3387 354819
rect -3269 354701 -3227 354819
rect -3109 354701 -3093 354819
rect -3403 354659 -3093 354701
rect -3403 354541 -3387 354659
rect -3269 354541 -3227 354659
rect -3109 354541 -3093 354659
rect -3403 338447 -3093 354541
rect -3403 338329 -3387 338447
rect -3269 338329 -3227 338447
rect -3109 338329 -3093 338447
rect -3403 338287 -3093 338329
rect -3403 338169 -3387 338287
rect -3269 338169 -3227 338287
rect -3109 338169 -3093 338287
rect -3403 320447 -3093 338169
rect -3403 320329 -3387 320447
rect -3269 320329 -3227 320447
rect -3109 320329 -3093 320447
rect -3403 320287 -3093 320329
rect -3403 320169 -3387 320287
rect -3269 320169 -3227 320287
rect -3109 320169 -3093 320287
rect -3403 302447 -3093 320169
rect -3403 302329 -3387 302447
rect -3269 302329 -3227 302447
rect -3109 302329 -3093 302447
rect -3403 302287 -3093 302329
rect -3403 302169 -3387 302287
rect -3269 302169 -3227 302287
rect -3109 302169 -3093 302287
rect -3403 284447 -3093 302169
rect -3403 284329 -3387 284447
rect -3269 284329 -3227 284447
rect -3109 284329 -3093 284447
rect -3403 284287 -3093 284329
rect -3403 284169 -3387 284287
rect -3269 284169 -3227 284287
rect -3109 284169 -3093 284287
rect -3403 266447 -3093 284169
rect -3403 266329 -3387 266447
rect -3269 266329 -3227 266447
rect -3109 266329 -3093 266447
rect -3403 266287 -3093 266329
rect -3403 266169 -3387 266287
rect -3269 266169 -3227 266287
rect -3109 266169 -3093 266287
rect -3403 248447 -3093 266169
rect -3403 248329 -3387 248447
rect -3269 248329 -3227 248447
rect -3109 248329 -3093 248447
rect -3403 248287 -3093 248329
rect -3403 248169 -3387 248287
rect -3269 248169 -3227 248287
rect -3109 248169 -3093 248287
rect -3403 230447 -3093 248169
rect -3403 230329 -3387 230447
rect -3269 230329 -3227 230447
rect -3109 230329 -3093 230447
rect -3403 230287 -3093 230329
rect -3403 230169 -3387 230287
rect -3269 230169 -3227 230287
rect -3109 230169 -3093 230287
rect -3403 212447 -3093 230169
rect -3403 212329 -3387 212447
rect -3269 212329 -3227 212447
rect -3109 212329 -3093 212447
rect -3403 212287 -3093 212329
rect -3403 212169 -3387 212287
rect -3269 212169 -3227 212287
rect -3109 212169 -3093 212287
rect -3403 194447 -3093 212169
rect -3403 194329 -3387 194447
rect -3269 194329 -3227 194447
rect -3109 194329 -3093 194447
rect -3403 194287 -3093 194329
rect -3403 194169 -3387 194287
rect -3269 194169 -3227 194287
rect -3109 194169 -3093 194287
rect -3403 176447 -3093 194169
rect -3403 176329 -3387 176447
rect -3269 176329 -3227 176447
rect -3109 176329 -3093 176447
rect -3403 176287 -3093 176329
rect -3403 176169 -3387 176287
rect -3269 176169 -3227 176287
rect -3109 176169 -3093 176287
rect -3403 158447 -3093 176169
rect -3403 158329 -3387 158447
rect -3269 158329 -3227 158447
rect -3109 158329 -3093 158447
rect -3403 158287 -3093 158329
rect -3403 158169 -3387 158287
rect -3269 158169 -3227 158287
rect -3109 158169 -3093 158287
rect -3403 140447 -3093 158169
rect -3403 140329 -3387 140447
rect -3269 140329 -3227 140447
rect -3109 140329 -3093 140447
rect -3403 140287 -3093 140329
rect -3403 140169 -3387 140287
rect -3269 140169 -3227 140287
rect -3109 140169 -3093 140287
rect -3403 122447 -3093 140169
rect -3403 122329 -3387 122447
rect -3269 122329 -3227 122447
rect -3109 122329 -3093 122447
rect -3403 122287 -3093 122329
rect -3403 122169 -3387 122287
rect -3269 122169 -3227 122287
rect -3109 122169 -3093 122287
rect -3403 104447 -3093 122169
rect -3403 104329 -3387 104447
rect -3269 104329 -3227 104447
rect -3109 104329 -3093 104447
rect -3403 104287 -3093 104329
rect -3403 104169 -3387 104287
rect -3269 104169 -3227 104287
rect -3109 104169 -3093 104287
rect -3403 86447 -3093 104169
rect -3403 86329 -3387 86447
rect -3269 86329 -3227 86447
rect -3109 86329 -3093 86447
rect -3403 86287 -3093 86329
rect -3403 86169 -3387 86287
rect -3269 86169 -3227 86287
rect -3109 86169 -3093 86287
rect -3403 68447 -3093 86169
rect -3403 68329 -3387 68447
rect -3269 68329 -3227 68447
rect -3109 68329 -3093 68447
rect -3403 68287 -3093 68329
rect -3403 68169 -3387 68287
rect -3269 68169 -3227 68287
rect -3109 68169 -3093 68287
rect -3403 50447 -3093 68169
rect -3403 50329 -3387 50447
rect -3269 50329 -3227 50447
rect -3109 50329 -3093 50447
rect -3403 50287 -3093 50329
rect -3403 50169 -3387 50287
rect -3269 50169 -3227 50287
rect -3109 50169 -3093 50287
rect -3403 32447 -3093 50169
rect -3403 32329 -3387 32447
rect -3269 32329 -3227 32447
rect -3109 32329 -3093 32447
rect -3403 32287 -3093 32329
rect -3403 32169 -3387 32287
rect -3269 32169 -3227 32287
rect -3109 32169 -3093 32287
rect -3403 14447 -3093 32169
rect -3403 14329 -3387 14447
rect -3269 14329 -3227 14447
rect -3109 14329 -3093 14447
rect -3403 14287 -3093 14329
rect -3403 14169 -3387 14287
rect -3269 14169 -3227 14287
rect -3109 14169 -3093 14287
rect -3403 -2573 -3093 14169
rect -2923 354339 -2613 354355
rect -2923 354221 -2907 354339
rect -2789 354221 -2747 354339
rect -2629 354221 -2613 354339
rect -2923 354179 -2613 354221
rect -2923 354061 -2907 354179
rect -2789 354061 -2747 354179
rect -2629 354061 -2613 354179
rect -2923 347447 -2613 354061
rect 4617 354339 4927 354835
rect 4617 354221 4633 354339
rect 4751 354221 4793 354339
rect 4911 354221 4927 354339
rect 4617 354179 4927 354221
rect 4617 354061 4633 354179
rect 4751 354061 4793 354179
rect 4911 354061 4927 354179
rect -2923 347329 -2907 347447
rect -2789 347329 -2747 347447
rect -2629 347329 -2613 347447
rect -2923 347287 -2613 347329
rect -2923 347169 -2907 347287
rect -2789 347169 -2747 347287
rect -2629 347169 -2613 347287
rect -2923 329447 -2613 347169
rect -2923 329329 -2907 329447
rect -2789 329329 -2747 329447
rect -2629 329329 -2613 329447
rect -2923 329287 -2613 329329
rect -2923 329169 -2907 329287
rect -2789 329169 -2747 329287
rect -2629 329169 -2613 329287
rect -2923 311447 -2613 329169
rect -2923 311329 -2907 311447
rect -2789 311329 -2747 311447
rect -2629 311329 -2613 311447
rect -2923 311287 -2613 311329
rect -2923 311169 -2907 311287
rect -2789 311169 -2747 311287
rect -2629 311169 -2613 311287
rect -2923 293447 -2613 311169
rect -2923 293329 -2907 293447
rect -2789 293329 -2747 293447
rect -2629 293329 -2613 293447
rect -2923 293287 -2613 293329
rect -2923 293169 -2907 293287
rect -2789 293169 -2747 293287
rect -2629 293169 -2613 293287
rect -2923 275447 -2613 293169
rect -2923 275329 -2907 275447
rect -2789 275329 -2747 275447
rect -2629 275329 -2613 275447
rect -2923 275287 -2613 275329
rect -2923 275169 -2907 275287
rect -2789 275169 -2747 275287
rect -2629 275169 -2613 275287
rect -2923 257447 -2613 275169
rect -2923 257329 -2907 257447
rect -2789 257329 -2747 257447
rect -2629 257329 -2613 257447
rect -2923 257287 -2613 257329
rect -2923 257169 -2907 257287
rect -2789 257169 -2747 257287
rect -2629 257169 -2613 257287
rect -2923 239447 -2613 257169
rect -2923 239329 -2907 239447
rect -2789 239329 -2747 239447
rect -2629 239329 -2613 239447
rect -2923 239287 -2613 239329
rect -2923 239169 -2907 239287
rect -2789 239169 -2747 239287
rect -2629 239169 -2613 239287
rect -2923 221447 -2613 239169
rect -2923 221329 -2907 221447
rect -2789 221329 -2747 221447
rect -2629 221329 -2613 221447
rect -2923 221287 -2613 221329
rect -2923 221169 -2907 221287
rect -2789 221169 -2747 221287
rect -2629 221169 -2613 221287
rect -2923 203447 -2613 221169
rect -2923 203329 -2907 203447
rect -2789 203329 -2747 203447
rect -2629 203329 -2613 203447
rect -2923 203287 -2613 203329
rect -2923 203169 -2907 203287
rect -2789 203169 -2747 203287
rect -2629 203169 -2613 203287
rect -2923 185447 -2613 203169
rect -2923 185329 -2907 185447
rect -2789 185329 -2747 185447
rect -2629 185329 -2613 185447
rect -2923 185287 -2613 185329
rect -2923 185169 -2907 185287
rect -2789 185169 -2747 185287
rect -2629 185169 -2613 185287
rect -2923 167447 -2613 185169
rect -2923 167329 -2907 167447
rect -2789 167329 -2747 167447
rect -2629 167329 -2613 167447
rect -2923 167287 -2613 167329
rect -2923 167169 -2907 167287
rect -2789 167169 -2747 167287
rect -2629 167169 -2613 167287
rect -2923 149447 -2613 167169
rect -2923 149329 -2907 149447
rect -2789 149329 -2747 149447
rect -2629 149329 -2613 149447
rect -2923 149287 -2613 149329
rect -2923 149169 -2907 149287
rect -2789 149169 -2747 149287
rect -2629 149169 -2613 149287
rect -2923 131447 -2613 149169
rect -2923 131329 -2907 131447
rect -2789 131329 -2747 131447
rect -2629 131329 -2613 131447
rect -2923 131287 -2613 131329
rect -2923 131169 -2907 131287
rect -2789 131169 -2747 131287
rect -2629 131169 -2613 131287
rect -2923 113447 -2613 131169
rect -2923 113329 -2907 113447
rect -2789 113329 -2747 113447
rect -2629 113329 -2613 113447
rect -2923 113287 -2613 113329
rect -2923 113169 -2907 113287
rect -2789 113169 -2747 113287
rect -2629 113169 -2613 113287
rect -2923 95447 -2613 113169
rect -2923 95329 -2907 95447
rect -2789 95329 -2747 95447
rect -2629 95329 -2613 95447
rect -2923 95287 -2613 95329
rect -2923 95169 -2907 95287
rect -2789 95169 -2747 95287
rect -2629 95169 -2613 95287
rect -2923 77447 -2613 95169
rect -2923 77329 -2907 77447
rect -2789 77329 -2747 77447
rect -2629 77329 -2613 77447
rect -2923 77287 -2613 77329
rect -2923 77169 -2907 77287
rect -2789 77169 -2747 77287
rect -2629 77169 -2613 77287
rect -2923 59447 -2613 77169
rect -2923 59329 -2907 59447
rect -2789 59329 -2747 59447
rect -2629 59329 -2613 59447
rect -2923 59287 -2613 59329
rect -2923 59169 -2907 59287
rect -2789 59169 -2747 59287
rect -2629 59169 -2613 59287
rect -2923 41447 -2613 59169
rect -2923 41329 -2907 41447
rect -2789 41329 -2747 41447
rect -2629 41329 -2613 41447
rect -2923 41287 -2613 41329
rect -2923 41169 -2907 41287
rect -2789 41169 -2747 41287
rect -2629 41169 -2613 41287
rect -2923 23447 -2613 41169
rect -2923 23329 -2907 23447
rect -2789 23329 -2747 23447
rect -2629 23329 -2613 23447
rect -2923 23287 -2613 23329
rect -2923 23169 -2907 23287
rect -2789 23169 -2747 23287
rect -2629 23169 -2613 23287
rect -2923 5447 -2613 23169
rect -2923 5329 -2907 5447
rect -2789 5329 -2747 5447
rect -2629 5329 -2613 5447
rect -2923 5287 -2613 5329
rect -2923 5169 -2907 5287
rect -2789 5169 -2747 5287
rect -2629 5169 -2613 5287
rect -2923 -2093 -2613 5169
rect -2443 353859 -2133 353875
rect -2443 353741 -2427 353859
rect -2309 353741 -2267 353859
rect -2149 353741 -2133 353859
rect -2443 353699 -2133 353741
rect -2443 353581 -2427 353699
rect -2309 353581 -2267 353699
rect -2149 353581 -2133 353699
rect -2443 336587 -2133 353581
rect -2443 336469 -2427 336587
rect -2309 336469 -2267 336587
rect -2149 336469 -2133 336587
rect -2443 336427 -2133 336469
rect -2443 336309 -2427 336427
rect -2309 336309 -2267 336427
rect -2149 336309 -2133 336427
rect -2443 318587 -2133 336309
rect -2443 318469 -2427 318587
rect -2309 318469 -2267 318587
rect -2149 318469 -2133 318587
rect -2443 318427 -2133 318469
rect -2443 318309 -2427 318427
rect -2309 318309 -2267 318427
rect -2149 318309 -2133 318427
rect -2443 300587 -2133 318309
rect -2443 300469 -2427 300587
rect -2309 300469 -2267 300587
rect -2149 300469 -2133 300587
rect -2443 300427 -2133 300469
rect -2443 300309 -2427 300427
rect -2309 300309 -2267 300427
rect -2149 300309 -2133 300427
rect -2443 282587 -2133 300309
rect -2443 282469 -2427 282587
rect -2309 282469 -2267 282587
rect -2149 282469 -2133 282587
rect -2443 282427 -2133 282469
rect -2443 282309 -2427 282427
rect -2309 282309 -2267 282427
rect -2149 282309 -2133 282427
rect -2443 264587 -2133 282309
rect -2443 264469 -2427 264587
rect -2309 264469 -2267 264587
rect -2149 264469 -2133 264587
rect -2443 264427 -2133 264469
rect -2443 264309 -2427 264427
rect -2309 264309 -2267 264427
rect -2149 264309 -2133 264427
rect -2443 246587 -2133 264309
rect -2443 246469 -2427 246587
rect -2309 246469 -2267 246587
rect -2149 246469 -2133 246587
rect -2443 246427 -2133 246469
rect -2443 246309 -2427 246427
rect -2309 246309 -2267 246427
rect -2149 246309 -2133 246427
rect -2443 228587 -2133 246309
rect -2443 228469 -2427 228587
rect -2309 228469 -2267 228587
rect -2149 228469 -2133 228587
rect -2443 228427 -2133 228469
rect -2443 228309 -2427 228427
rect -2309 228309 -2267 228427
rect -2149 228309 -2133 228427
rect -2443 210587 -2133 228309
rect -2443 210469 -2427 210587
rect -2309 210469 -2267 210587
rect -2149 210469 -2133 210587
rect -2443 210427 -2133 210469
rect -2443 210309 -2427 210427
rect -2309 210309 -2267 210427
rect -2149 210309 -2133 210427
rect -2443 192587 -2133 210309
rect -2443 192469 -2427 192587
rect -2309 192469 -2267 192587
rect -2149 192469 -2133 192587
rect -2443 192427 -2133 192469
rect -2443 192309 -2427 192427
rect -2309 192309 -2267 192427
rect -2149 192309 -2133 192427
rect -2443 174587 -2133 192309
rect -2443 174469 -2427 174587
rect -2309 174469 -2267 174587
rect -2149 174469 -2133 174587
rect -2443 174427 -2133 174469
rect -2443 174309 -2427 174427
rect -2309 174309 -2267 174427
rect -2149 174309 -2133 174427
rect -2443 156587 -2133 174309
rect -2443 156469 -2427 156587
rect -2309 156469 -2267 156587
rect -2149 156469 -2133 156587
rect -2443 156427 -2133 156469
rect -2443 156309 -2427 156427
rect -2309 156309 -2267 156427
rect -2149 156309 -2133 156427
rect -2443 138587 -2133 156309
rect -2443 138469 -2427 138587
rect -2309 138469 -2267 138587
rect -2149 138469 -2133 138587
rect -2443 138427 -2133 138469
rect -2443 138309 -2427 138427
rect -2309 138309 -2267 138427
rect -2149 138309 -2133 138427
rect -2443 120587 -2133 138309
rect -2443 120469 -2427 120587
rect -2309 120469 -2267 120587
rect -2149 120469 -2133 120587
rect -2443 120427 -2133 120469
rect -2443 120309 -2427 120427
rect -2309 120309 -2267 120427
rect -2149 120309 -2133 120427
rect -2443 102587 -2133 120309
rect -2443 102469 -2427 102587
rect -2309 102469 -2267 102587
rect -2149 102469 -2133 102587
rect -2443 102427 -2133 102469
rect -2443 102309 -2427 102427
rect -2309 102309 -2267 102427
rect -2149 102309 -2133 102427
rect -2443 84587 -2133 102309
rect -2443 84469 -2427 84587
rect -2309 84469 -2267 84587
rect -2149 84469 -2133 84587
rect -2443 84427 -2133 84469
rect -2443 84309 -2427 84427
rect -2309 84309 -2267 84427
rect -2149 84309 -2133 84427
rect -2443 66587 -2133 84309
rect -2443 66469 -2427 66587
rect -2309 66469 -2267 66587
rect -2149 66469 -2133 66587
rect -2443 66427 -2133 66469
rect -2443 66309 -2427 66427
rect -2309 66309 -2267 66427
rect -2149 66309 -2133 66427
rect -2443 48587 -2133 66309
rect -2443 48469 -2427 48587
rect -2309 48469 -2267 48587
rect -2149 48469 -2133 48587
rect -2443 48427 -2133 48469
rect -2443 48309 -2427 48427
rect -2309 48309 -2267 48427
rect -2149 48309 -2133 48427
rect -2443 30587 -2133 48309
rect -2443 30469 -2427 30587
rect -2309 30469 -2267 30587
rect -2149 30469 -2133 30587
rect -2443 30427 -2133 30469
rect -2443 30309 -2427 30427
rect -2309 30309 -2267 30427
rect -2149 30309 -2133 30427
rect -2443 12587 -2133 30309
rect -2443 12469 -2427 12587
rect -2309 12469 -2267 12587
rect -2149 12469 -2133 12587
rect -2443 12427 -2133 12469
rect -2443 12309 -2427 12427
rect -2309 12309 -2267 12427
rect -2149 12309 -2133 12427
rect -2443 -1613 -2133 12309
rect -1963 353379 -1653 353395
rect -1963 353261 -1947 353379
rect -1829 353261 -1787 353379
rect -1669 353261 -1653 353379
rect -1963 353219 -1653 353261
rect -1963 353101 -1947 353219
rect -1829 353101 -1787 353219
rect -1669 353101 -1653 353219
rect -1963 345587 -1653 353101
rect 2757 353379 3067 353875
rect 2757 353261 2773 353379
rect 2891 353261 2933 353379
rect 3051 353261 3067 353379
rect 2757 353219 3067 353261
rect 2757 353101 2773 353219
rect 2891 353101 2933 353219
rect 3051 353101 3067 353219
rect -1963 345469 -1947 345587
rect -1829 345469 -1787 345587
rect -1669 345469 -1653 345587
rect -1963 345427 -1653 345469
rect -1963 345309 -1947 345427
rect -1829 345309 -1787 345427
rect -1669 345309 -1653 345427
rect -1963 327587 -1653 345309
rect -1963 327469 -1947 327587
rect -1829 327469 -1787 327587
rect -1669 327469 -1653 327587
rect -1963 327427 -1653 327469
rect -1963 327309 -1947 327427
rect -1829 327309 -1787 327427
rect -1669 327309 -1653 327427
rect -1963 309587 -1653 327309
rect -1963 309469 -1947 309587
rect -1829 309469 -1787 309587
rect -1669 309469 -1653 309587
rect -1963 309427 -1653 309469
rect -1963 309309 -1947 309427
rect -1829 309309 -1787 309427
rect -1669 309309 -1653 309427
rect -1963 291587 -1653 309309
rect -1963 291469 -1947 291587
rect -1829 291469 -1787 291587
rect -1669 291469 -1653 291587
rect -1963 291427 -1653 291469
rect -1963 291309 -1947 291427
rect -1829 291309 -1787 291427
rect -1669 291309 -1653 291427
rect -1963 273587 -1653 291309
rect -1963 273469 -1947 273587
rect -1829 273469 -1787 273587
rect -1669 273469 -1653 273587
rect -1963 273427 -1653 273469
rect -1963 273309 -1947 273427
rect -1829 273309 -1787 273427
rect -1669 273309 -1653 273427
rect -1963 255587 -1653 273309
rect -1963 255469 -1947 255587
rect -1829 255469 -1787 255587
rect -1669 255469 -1653 255587
rect -1963 255427 -1653 255469
rect -1963 255309 -1947 255427
rect -1829 255309 -1787 255427
rect -1669 255309 -1653 255427
rect -1963 237587 -1653 255309
rect -1963 237469 -1947 237587
rect -1829 237469 -1787 237587
rect -1669 237469 -1653 237587
rect -1963 237427 -1653 237469
rect -1963 237309 -1947 237427
rect -1829 237309 -1787 237427
rect -1669 237309 -1653 237427
rect -1963 219587 -1653 237309
rect -1963 219469 -1947 219587
rect -1829 219469 -1787 219587
rect -1669 219469 -1653 219587
rect -1963 219427 -1653 219469
rect -1963 219309 -1947 219427
rect -1829 219309 -1787 219427
rect -1669 219309 -1653 219427
rect -1963 201587 -1653 219309
rect -1963 201469 -1947 201587
rect -1829 201469 -1787 201587
rect -1669 201469 -1653 201587
rect -1963 201427 -1653 201469
rect -1963 201309 -1947 201427
rect -1829 201309 -1787 201427
rect -1669 201309 -1653 201427
rect -1963 183587 -1653 201309
rect -1963 183469 -1947 183587
rect -1829 183469 -1787 183587
rect -1669 183469 -1653 183587
rect -1963 183427 -1653 183469
rect -1963 183309 -1947 183427
rect -1829 183309 -1787 183427
rect -1669 183309 -1653 183427
rect -1963 165587 -1653 183309
rect -1963 165469 -1947 165587
rect -1829 165469 -1787 165587
rect -1669 165469 -1653 165587
rect -1963 165427 -1653 165469
rect -1963 165309 -1947 165427
rect -1829 165309 -1787 165427
rect -1669 165309 -1653 165427
rect -1963 147587 -1653 165309
rect -1963 147469 -1947 147587
rect -1829 147469 -1787 147587
rect -1669 147469 -1653 147587
rect -1963 147427 -1653 147469
rect -1963 147309 -1947 147427
rect -1829 147309 -1787 147427
rect -1669 147309 -1653 147427
rect -1963 129587 -1653 147309
rect -1963 129469 -1947 129587
rect -1829 129469 -1787 129587
rect -1669 129469 -1653 129587
rect -1963 129427 -1653 129469
rect -1963 129309 -1947 129427
rect -1829 129309 -1787 129427
rect -1669 129309 -1653 129427
rect -1963 111587 -1653 129309
rect -1963 111469 -1947 111587
rect -1829 111469 -1787 111587
rect -1669 111469 -1653 111587
rect -1963 111427 -1653 111469
rect -1963 111309 -1947 111427
rect -1829 111309 -1787 111427
rect -1669 111309 -1653 111427
rect -1963 93587 -1653 111309
rect -1963 93469 -1947 93587
rect -1829 93469 -1787 93587
rect -1669 93469 -1653 93587
rect -1963 93427 -1653 93469
rect -1963 93309 -1947 93427
rect -1829 93309 -1787 93427
rect -1669 93309 -1653 93427
rect -1963 75587 -1653 93309
rect -1963 75469 -1947 75587
rect -1829 75469 -1787 75587
rect -1669 75469 -1653 75587
rect -1963 75427 -1653 75469
rect -1963 75309 -1947 75427
rect -1829 75309 -1787 75427
rect -1669 75309 -1653 75427
rect -1963 57587 -1653 75309
rect -1963 57469 -1947 57587
rect -1829 57469 -1787 57587
rect -1669 57469 -1653 57587
rect -1963 57427 -1653 57469
rect -1963 57309 -1947 57427
rect -1829 57309 -1787 57427
rect -1669 57309 -1653 57427
rect -1963 39587 -1653 57309
rect -1963 39469 -1947 39587
rect -1829 39469 -1787 39587
rect -1669 39469 -1653 39587
rect -1963 39427 -1653 39469
rect -1963 39309 -1947 39427
rect -1829 39309 -1787 39427
rect -1669 39309 -1653 39427
rect -1963 21587 -1653 39309
rect -1963 21469 -1947 21587
rect -1829 21469 -1787 21587
rect -1669 21469 -1653 21587
rect -1963 21427 -1653 21469
rect -1963 21309 -1947 21427
rect -1829 21309 -1787 21427
rect -1669 21309 -1653 21427
rect -1963 3587 -1653 21309
rect -1963 3469 -1947 3587
rect -1829 3469 -1787 3587
rect -1669 3469 -1653 3587
rect -1963 3427 -1653 3469
rect -1963 3309 -1947 3427
rect -1829 3309 -1787 3427
rect -1669 3309 -1653 3427
rect -1963 -1133 -1653 3309
rect -1483 352899 -1173 352915
rect -1483 352781 -1467 352899
rect -1349 352781 -1307 352899
rect -1189 352781 -1173 352899
rect -1483 352739 -1173 352781
rect -1483 352621 -1467 352739
rect -1349 352621 -1307 352739
rect -1189 352621 -1173 352739
rect -1483 334727 -1173 352621
rect -1483 334609 -1467 334727
rect -1349 334609 -1307 334727
rect -1189 334609 -1173 334727
rect -1483 334567 -1173 334609
rect -1483 334449 -1467 334567
rect -1349 334449 -1307 334567
rect -1189 334449 -1173 334567
rect -1483 316727 -1173 334449
rect -1483 316609 -1467 316727
rect -1349 316609 -1307 316727
rect -1189 316609 -1173 316727
rect -1483 316567 -1173 316609
rect -1483 316449 -1467 316567
rect -1349 316449 -1307 316567
rect -1189 316449 -1173 316567
rect -1483 298727 -1173 316449
rect -1483 298609 -1467 298727
rect -1349 298609 -1307 298727
rect -1189 298609 -1173 298727
rect -1483 298567 -1173 298609
rect -1483 298449 -1467 298567
rect -1349 298449 -1307 298567
rect -1189 298449 -1173 298567
rect -1483 280727 -1173 298449
rect -1483 280609 -1467 280727
rect -1349 280609 -1307 280727
rect -1189 280609 -1173 280727
rect -1483 280567 -1173 280609
rect -1483 280449 -1467 280567
rect -1349 280449 -1307 280567
rect -1189 280449 -1173 280567
rect -1483 262727 -1173 280449
rect -1483 262609 -1467 262727
rect -1349 262609 -1307 262727
rect -1189 262609 -1173 262727
rect -1483 262567 -1173 262609
rect -1483 262449 -1467 262567
rect -1349 262449 -1307 262567
rect -1189 262449 -1173 262567
rect -1483 244727 -1173 262449
rect -1483 244609 -1467 244727
rect -1349 244609 -1307 244727
rect -1189 244609 -1173 244727
rect -1483 244567 -1173 244609
rect -1483 244449 -1467 244567
rect -1349 244449 -1307 244567
rect -1189 244449 -1173 244567
rect -1483 226727 -1173 244449
rect -1483 226609 -1467 226727
rect -1349 226609 -1307 226727
rect -1189 226609 -1173 226727
rect -1483 226567 -1173 226609
rect -1483 226449 -1467 226567
rect -1349 226449 -1307 226567
rect -1189 226449 -1173 226567
rect -1483 208727 -1173 226449
rect -1483 208609 -1467 208727
rect -1349 208609 -1307 208727
rect -1189 208609 -1173 208727
rect -1483 208567 -1173 208609
rect -1483 208449 -1467 208567
rect -1349 208449 -1307 208567
rect -1189 208449 -1173 208567
rect -1483 190727 -1173 208449
rect -1483 190609 -1467 190727
rect -1349 190609 -1307 190727
rect -1189 190609 -1173 190727
rect -1483 190567 -1173 190609
rect -1483 190449 -1467 190567
rect -1349 190449 -1307 190567
rect -1189 190449 -1173 190567
rect -1483 172727 -1173 190449
rect -1483 172609 -1467 172727
rect -1349 172609 -1307 172727
rect -1189 172609 -1173 172727
rect -1483 172567 -1173 172609
rect -1483 172449 -1467 172567
rect -1349 172449 -1307 172567
rect -1189 172449 -1173 172567
rect -1483 154727 -1173 172449
rect -1483 154609 -1467 154727
rect -1349 154609 -1307 154727
rect -1189 154609 -1173 154727
rect -1483 154567 -1173 154609
rect -1483 154449 -1467 154567
rect -1349 154449 -1307 154567
rect -1189 154449 -1173 154567
rect -1483 136727 -1173 154449
rect -1483 136609 -1467 136727
rect -1349 136609 -1307 136727
rect -1189 136609 -1173 136727
rect -1483 136567 -1173 136609
rect -1483 136449 -1467 136567
rect -1349 136449 -1307 136567
rect -1189 136449 -1173 136567
rect -1483 118727 -1173 136449
rect -1483 118609 -1467 118727
rect -1349 118609 -1307 118727
rect -1189 118609 -1173 118727
rect -1483 118567 -1173 118609
rect -1483 118449 -1467 118567
rect -1349 118449 -1307 118567
rect -1189 118449 -1173 118567
rect -1483 100727 -1173 118449
rect -1483 100609 -1467 100727
rect -1349 100609 -1307 100727
rect -1189 100609 -1173 100727
rect -1483 100567 -1173 100609
rect -1483 100449 -1467 100567
rect -1349 100449 -1307 100567
rect -1189 100449 -1173 100567
rect -1483 82727 -1173 100449
rect -1483 82609 -1467 82727
rect -1349 82609 -1307 82727
rect -1189 82609 -1173 82727
rect -1483 82567 -1173 82609
rect -1483 82449 -1467 82567
rect -1349 82449 -1307 82567
rect -1189 82449 -1173 82567
rect -1483 64727 -1173 82449
rect -1483 64609 -1467 64727
rect -1349 64609 -1307 64727
rect -1189 64609 -1173 64727
rect -1483 64567 -1173 64609
rect -1483 64449 -1467 64567
rect -1349 64449 -1307 64567
rect -1189 64449 -1173 64567
rect -1483 46727 -1173 64449
rect -1483 46609 -1467 46727
rect -1349 46609 -1307 46727
rect -1189 46609 -1173 46727
rect -1483 46567 -1173 46609
rect -1483 46449 -1467 46567
rect -1349 46449 -1307 46567
rect -1189 46449 -1173 46567
rect -1483 28727 -1173 46449
rect -1483 28609 -1467 28727
rect -1349 28609 -1307 28727
rect -1189 28609 -1173 28727
rect -1483 28567 -1173 28609
rect -1483 28449 -1467 28567
rect -1349 28449 -1307 28567
rect -1189 28449 -1173 28567
rect -1483 10727 -1173 28449
rect -1483 10609 -1467 10727
rect -1349 10609 -1307 10727
rect -1189 10609 -1173 10727
rect -1483 10567 -1173 10609
rect -1483 10449 -1467 10567
rect -1349 10449 -1307 10567
rect -1189 10449 -1173 10567
rect -1483 -653 -1173 10449
rect -1003 352419 -693 352435
rect -1003 352301 -987 352419
rect -869 352301 -827 352419
rect -709 352301 -693 352419
rect -1003 352259 -693 352301
rect -1003 352141 -987 352259
rect -869 352141 -827 352259
rect -709 352141 -693 352259
rect -1003 343727 -693 352141
rect -1003 343609 -987 343727
rect -869 343609 -827 343727
rect -709 343609 -693 343727
rect -1003 343567 -693 343609
rect -1003 343449 -987 343567
rect -869 343449 -827 343567
rect -709 343449 -693 343567
rect -1003 325727 -693 343449
rect -1003 325609 -987 325727
rect -869 325609 -827 325727
rect -709 325609 -693 325727
rect -1003 325567 -693 325609
rect -1003 325449 -987 325567
rect -869 325449 -827 325567
rect -709 325449 -693 325567
rect -1003 307727 -693 325449
rect -1003 307609 -987 307727
rect -869 307609 -827 307727
rect -709 307609 -693 307727
rect -1003 307567 -693 307609
rect -1003 307449 -987 307567
rect -869 307449 -827 307567
rect -709 307449 -693 307567
rect -1003 289727 -693 307449
rect -1003 289609 -987 289727
rect -869 289609 -827 289727
rect -709 289609 -693 289727
rect -1003 289567 -693 289609
rect -1003 289449 -987 289567
rect -869 289449 -827 289567
rect -709 289449 -693 289567
rect -1003 271727 -693 289449
rect -1003 271609 -987 271727
rect -869 271609 -827 271727
rect -709 271609 -693 271727
rect -1003 271567 -693 271609
rect -1003 271449 -987 271567
rect -869 271449 -827 271567
rect -709 271449 -693 271567
rect -1003 253727 -693 271449
rect -1003 253609 -987 253727
rect -869 253609 -827 253727
rect -709 253609 -693 253727
rect -1003 253567 -693 253609
rect -1003 253449 -987 253567
rect -869 253449 -827 253567
rect -709 253449 -693 253567
rect -1003 235727 -693 253449
rect -1003 235609 -987 235727
rect -869 235609 -827 235727
rect -709 235609 -693 235727
rect -1003 235567 -693 235609
rect -1003 235449 -987 235567
rect -869 235449 -827 235567
rect -709 235449 -693 235567
rect -1003 217727 -693 235449
rect -1003 217609 -987 217727
rect -869 217609 -827 217727
rect -709 217609 -693 217727
rect -1003 217567 -693 217609
rect -1003 217449 -987 217567
rect -869 217449 -827 217567
rect -709 217449 -693 217567
rect -1003 199727 -693 217449
rect -1003 199609 -987 199727
rect -869 199609 -827 199727
rect -709 199609 -693 199727
rect -1003 199567 -693 199609
rect -1003 199449 -987 199567
rect -869 199449 -827 199567
rect -709 199449 -693 199567
rect -1003 181727 -693 199449
rect -1003 181609 -987 181727
rect -869 181609 -827 181727
rect -709 181609 -693 181727
rect -1003 181567 -693 181609
rect -1003 181449 -987 181567
rect -869 181449 -827 181567
rect -709 181449 -693 181567
rect -1003 163727 -693 181449
rect -1003 163609 -987 163727
rect -869 163609 -827 163727
rect -709 163609 -693 163727
rect -1003 163567 -693 163609
rect -1003 163449 -987 163567
rect -869 163449 -827 163567
rect -709 163449 -693 163567
rect -1003 145727 -693 163449
rect -1003 145609 -987 145727
rect -869 145609 -827 145727
rect -709 145609 -693 145727
rect -1003 145567 -693 145609
rect -1003 145449 -987 145567
rect -869 145449 -827 145567
rect -709 145449 -693 145567
rect -1003 127727 -693 145449
rect -1003 127609 -987 127727
rect -869 127609 -827 127727
rect -709 127609 -693 127727
rect -1003 127567 -693 127609
rect -1003 127449 -987 127567
rect -869 127449 -827 127567
rect -709 127449 -693 127567
rect -1003 109727 -693 127449
rect -1003 109609 -987 109727
rect -869 109609 -827 109727
rect -709 109609 -693 109727
rect -1003 109567 -693 109609
rect -1003 109449 -987 109567
rect -869 109449 -827 109567
rect -709 109449 -693 109567
rect -1003 91727 -693 109449
rect -1003 91609 -987 91727
rect -869 91609 -827 91727
rect -709 91609 -693 91727
rect -1003 91567 -693 91609
rect -1003 91449 -987 91567
rect -869 91449 -827 91567
rect -709 91449 -693 91567
rect -1003 73727 -693 91449
rect -1003 73609 -987 73727
rect -869 73609 -827 73727
rect -709 73609 -693 73727
rect -1003 73567 -693 73609
rect -1003 73449 -987 73567
rect -869 73449 -827 73567
rect -709 73449 -693 73567
rect -1003 55727 -693 73449
rect -1003 55609 -987 55727
rect -869 55609 -827 55727
rect -709 55609 -693 55727
rect -1003 55567 -693 55609
rect -1003 55449 -987 55567
rect -869 55449 -827 55567
rect -709 55449 -693 55567
rect -1003 37727 -693 55449
rect -1003 37609 -987 37727
rect -869 37609 -827 37727
rect -709 37609 -693 37727
rect -1003 37567 -693 37609
rect -1003 37449 -987 37567
rect -869 37449 -827 37567
rect -709 37449 -693 37567
rect -1003 19727 -693 37449
rect -1003 19609 -987 19727
rect -869 19609 -827 19727
rect -709 19609 -693 19727
rect -1003 19567 -693 19609
rect -1003 19449 -987 19567
rect -869 19449 -827 19567
rect -709 19449 -693 19567
rect -1003 1727 -693 19449
rect -1003 1609 -987 1727
rect -869 1609 -827 1727
rect -709 1609 -693 1727
rect -1003 1567 -693 1609
rect -1003 1449 -987 1567
rect -869 1449 -827 1567
rect -709 1449 -693 1567
rect -1003 -173 -693 1449
rect -1003 -291 -987 -173
rect -869 -291 -827 -173
rect -709 -291 -693 -173
rect -1003 -333 -693 -291
rect -1003 -451 -987 -333
rect -869 -451 -827 -333
rect -709 -451 -693 -333
rect -1003 -467 -693 -451
rect 897 352419 1207 352915
rect 897 352301 913 352419
rect 1031 352301 1073 352419
rect 1191 352301 1207 352419
rect 897 352259 1207 352301
rect 897 352141 913 352259
rect 1031 352141 1073 352259
rect 1191 352141 1207 352259
rect 897 343727 1207 352141
rect 897 343609 913 343727
rect 1031 343609 1073 343727
rect 1191 343609 1207 343727
rect 897 343567 1207 343609
rect 897 343449 913 343567
rect 1031 343449 1073 343567
rect 1191 343449 1207 343567
rect 897 325727 1207 343449
rect 897 325609 913 325727
rect 1031 325609 1073 325727
rect 1191 325609 1207 325727
rect 897 325567 1207 325609
rect 897 325449 913 325567
rect 1031 325449 1073 325567
rect 1191 325449 1207 325567
rect 897 307727 1207 325449
rect 897 307609 913 307727
rect 1031 307609 1073 307727
rect 1191 307609 1207 307727
rect 897 307567 1207 307609
rect 897 307449 913 307567
rect 1031 307449 1073 307567
rect 1191 307449 1207 307567
rect 897 289727 1207 307449
rect 897 289609 913 289727
rect 1031 289609 1073 289727
rect 1191 289609 1207 289727
rect 897 289567 1207 289609
rect 897 289449 913 289567
rect 1031 289449 1073 289567
rect 1191 289449 1207 289567
rect 897 271727 1207 289449
rect 897 271609 913 271727
rect 1031 271609 1073 271727
rect 1191 271609 1207 271727
rect 897 271567 1207 271609
rect 897 271449 913 271567
rect 1031 271449 1073 271567
rect 1191 271449 1207 271567
rect 897 253727 1207 271449
rect 897 253609 913 253727
rect 1031 253609 1073 253727
rect 1191 253609 1207 253727
rect 897 253567 1207 253609
rect 897 253449 913 253567
rect 1031 253449 1073 253567
rect 1191 253449 1207 253567
rect 897 235727 1207 253449
rect 897 235609 913 235727
rect 1031 235609 1073 235727
rect 1191 235609 1207 235727
rect 897 235567 1207 235609
rect 897 235449 913 235567
rect 1031 235449 1073 235567
rect 1191 235449 1207 235567
rect 897 217727 1207 235449
rect 897 217609 913 217727
rect 1031 217609 1073 217727
rect 1191 217609 1207 217727
rect 897 217567 1207 217609
rect 897 217449 913 217567
rect 1031 217449 1073 217567
rect 1191 217449 1207 217567
rect 897 199727 1207 217449
rect 897 199609 913 199727
rect 1031 199609 1073 199727
rect 1191 199609 1207 199727
rect 897 199567 1207 199609
rect 897 199449 913 199567
rect 1031 199449 1073 199567
rect 1191 199449 1207 199567
rect 897 181727 1207 199449
rect 897 181609 913 181727
rect 1031 181609 1073 181727
rect 1191 181609 1207 181727
rect 897 181567 1207 181609
rect 897 181449 913 181567
rect 1031 181449 1073 181567
rect 1191 181449 1207 181567
rect 897 163727 1207 181449
rect 897 163609 913 163727
rect 1031 163609 1073 163727
rect 1191 163609 1207 163727
rect 897 163567 1207 163609
rect 897 163449 913 163567
rect 1031 163449 1073 163567
rect 1191 163449 1207 163567
rect 897 145727 1207 163449
rect 897 145609 913 145727
rect 1031 145609 1073 145727
rect 1191 145609 1207 145727
rect 897 145567 1207 145609
rect 897 145449 913 145567
rect 1031 145449 1073 145567
rect 1191 145449 1207 145567
rect 897 127727 1207 145449
rect 897 127609 913 127727
rect 1031 127609 1073 127727
rect 1191 127609 1207 127727
rect 897 127567 1207 127609
rect 897 127449 913 127567
rect 1031 127449 1073 127567
rect 1191 127449 1207 127567
rect 897 109727 1207 127449
rect 897 109609 913 109727
rect 1031 109609 1073 109727
rect 1191 109609 1207 109727
rect 897 109567 1207 109609
rect 897 109449 913 109567
rect 1031 109449 1073 109567
rect 1191 109449 1207 109567
rect 897 91727 1207 109449
rect 897 91609 913 91727
rect 1031 91609 1073 91727
rect 1191 91609 1207 91727
rect 897 91567 1207 91609
rect 897 91449 913 91567
rect 1031 91449 1073 91567
rect 1191 91449 1207 91567
rect 897 73727 1207 91449
rect 897 73609 913 73727
rect 1031 73609 1073 73727
rect 1191 73609 1207 73727
rect 897 73567 1207 73609
rect 897 73449 913 73567
rect 1031 73449 1073 73567
rect 1191 73449 1207 73567
rect 897 55727 1207 73449
rect 897 55609 913 55727
rect 1031 55609 1073 55727
rect 1191 55609 1207 55727
rect 897 55567 1207 55609
rect 897 55449 913 55567
rect 1031 55449 1073 55567
rect 1191 55449 1207 55567
rect 897 37727 1207 55449
rect 897 37609 913 37727
rect 1031 37609 1073 37727
rect 1191 37609 1207 37727
rect 897 37567 1207 37609
rect 897 37449 913 37567
rect 1031 37449 1073 37567
rect 1191 37449 1207 37567
rect 897 19727 1207 37449
rect 897 19609 913 19727
rect 1031 19609 1073 19727
rect 1191 19609 1207 19727
rect 897 19567 1207 19609
rect 897 19449 913 19567
rect 1031 19449 1073 19567
rect 1191 19449 1207 19567
rect 897 1727 1207 19449
rect 897 1609 913 1727
rect 1031 1609 1073 1727
rect 1191 1609 1207 1727
rect 897 1567 1207 1609
rect 897 1449 913 1567
rect 1031 1449 1073 1567
rect 1191 1449 1207 1567
rect 897 -173 1207 1449
rect 897 -291 913 -173
rect 1031 -291 1073 -173
rect 1191 -291 1207 -173
rect 897 -333 1207 -291
rect 897 -451 913 -333
rect 1031 -451 1073 -333
rect 1191 -451 1207 -333
rect -1483 -771 -1467 -653
rect -1349 -771 -1307 -653
rect -1189 -771 -1173 -653
rect -1483 -813 -1173 -771
rect -1483 -931 -1467 -813
rect -1349 -931 -1307 -813
rect -1189 -931 -1173 -813
rect -1483 -947 -1173 -931
rect 897 -947 1207 -451
rect 2757 345587 3067 353101
rect 2757 345469 2773 345587
rect 2891 345469 2933 345587
rect 3051 345469 3067 345587
rect 2757 345427 3067 345469
rect 2757 345309 2773 345427
rect 2891 345309 2933 345427
rect 3051 345309 3067 345427
rect 2757 327587 3067 345309
rect 2757 327469 2773 327587
rect 2891 327469 2933 327587
rect 3051 327469 3067 327587
rect 2757 327427 3067 327469
rect 2757 327309 2773 327427
rect 2891 327309 2933 327427
rect 3051 327309 3067 327427
rect 2757 309587 3067 327309
rect 2757 309469 2773 309587
rect 2891 309469 2933 309587
rect 3051 309469 3067 309587
rect 2757 309427 3067 309469
rect 2757 309309 2773 309427
rect 2891 309309 2933 309427
rect 3051 309309 3067 309427
rect 2757 291587 3067 309309
rect 2757 291469 2773 291587
rect 2891 291469 2933 291587
rect 3051 291469 3067 291587
rect 2757 291427 3067 291469
rect 2757 291309 2773 291427
rect 2891 291309 2933 291427
rect 3051 291309 3067 291427
rect 2757 273587 3067 291309
rect 2757 273469 2773 273587
rect 2891 273469 2933 273587
rect 3051 273469 3067 273587
rect 2757 273427 3067 273469
rect 2757 273309 2773 273427
rect 2891 273309 2933 273427
rect 3051 273309 3067 273427
rect 2757 255587 3067 273309
rect 2757 255469 2773 255587
rect 2891 255469 2933 255587
rect 3051 255469 3067 255587
rect 2757 255427 3067 255469
rect 2757 255309 2773 255427
rect 2891 255309 2933 255427
rect 3051 255309 3067 255427
rect 2757 237587 3067 255309
rect 2757 237469 2773 237587
rect 2891 237469 2933 237587
rect 3051 237469 3067 237587
rect 2757 237427 3067 237469
rect 2757 237309 2773 237427
rect 2891 237309 2933 237427
rect 3051 237309 3067 237427
rect 2757 219587 3067 237309
rect 2757 219469 2773 219587
rect 2891 219469 2933 219587
rect 3051 219469 3067 219587
rect 2757 219427 3067 219469
rect 2757 219309 2773 219427
rect 2891 219309 2933 219427
rect 3051 219309 3067 219427
rect 2757 201587 3067 219309
rect 2757 201469 2773 201587
rect 2891 201469 2933 201587
rect 3051 201469 3067 201587
rect 2757 201427 3067 201469
rect 2757 201309 2773 201427
rect 2891 201309 2933 201427
rect 3051 201309 3067 201427
rect 2757 183587 3067 201309
rect 2757 183469 2773 183587
rect 2891 183469 2933 183587
rect 3051 183469 3067 183587
rect 2757 183427 3067 183469
rect 2757 183309 2773 183427
rect 2891 183309 2933 183427
rect 3051 183309 3067 183427
rect 2757 165587 3067 183309
rect 2757 165469 2773 165587
rect 2891 165469 2933 165587
rect 3051 165469 3067 165587
rect 2757 165427 3067 165469
rect 2757 165309 2773 165427
rect 2891 165309 2933 165427
rect 3051 165309 3067 165427
rect 2757 147587 3067 165309
rect 2757 147469 2773 147587
rect 2891 147469 2933 147587
rect 3051 147469 3067 147587
rect 2757 147427 3067 147469
rect 2757 147309 2773 147427
rect 2891 147309 2933 147427
rect 3051 147309 3067 147427
rect 2757 129587 3067 147309
rect 2757 129469 2773 129587
rect 2891 129469 2933 129587
rect 3051 129469 3067 129587
rect 2757 129427 3067 129469
rect 2757 129309 2773 129427
rect 2891 129309 2933 129427
rect 3051 129309 3067 129427
rect 2757 111587 3067 129309
rect 2757 111469 2773 111587
rect 2891 111469 2933 111587
rect 3051 111469 3067 111587
rect 2757 111427 3067 111469
rect 2757 111309 2773 111427
rect 2891 111309 2933 111427
rect 3051 111309 3067 111427
rect 2757 93587 3067 111309
rect 2757 93469 2773 93587
rect 2891 93469 2933 93587
rect 3051 93469 3067 93587
rect 2757 93427 3067 93469
rect 2757 93309 2773 93427
rect 2891 93309 2933 93427
rect 3051 93309 3067 93427
rect 2757 75587 3067 93309
rect 2757 75469 2773 75587
rect 2891 75469 2933 75587
rect 3051 75469 3067 75587
rect 2757 75427 3067 75469
rect 2757 75309 2773 75427
rect 2891 75309 2933 75427
rect 3051 75309 3067 75427
rect 2757 57587 3067 75309
rect 2757 57469 2773 57587
rect 2891 57469 2933 57587
rect 3051 57469 3067 57587
rect 2757 57427 3067 57469
rect 2757 57309 2773 57427
rect 2891 57309 2933 57427
rect 3051 57309 3067 57427
rect 2757 39587 3067 57309
rect 2757 39469 2773 39587
rect 2891 39469 2933 39587
rect 3051 39469 3067 39587
rect 2757 39427 3067 39469
rect 2757 39309 2773 39427
rect 2891 39309 2933 39427
rect 3051 39309 3067 39427
rect 2757 21587 3067 39309
rect 2757 21469 2773 21587
rect 2891 21469 2933 21587
rect 3051 21469 3067 21587
rect 2757 21427 3067 21469
rect 2757 21309 2773 21427
rect 2891 21309 2933 21427
rect 3051 21309 3067 21427
rect 2757 3587 3067 21309
rect 2757 3469 2773 3587
rect 2891 3469 2933 3587
rect 3051 3469 3067 3587
rect 2757 3427 3067 3469
rect 2757 3309 2773 3427
rect 2891 3309 2933 3427
rect 3051 3309 3067 3427
rect -1963 -1251 -1947 -1133
rect -1829 -1251 -1787 -1133
rect -1669 -1251 -1653 -1133
rect -1963 -1293 -1653 -1251
rect -1963 -1411 -1947 -1293
rect -1829 -1411 -1787 -1293
rect -1669 -1411 -1653 -1293
rect -1963 -1427 -1653 -1411
rect 2757 -1133 3067 3309
rect 2757 -1251 2773 -1133
rect 2891 -1251 2933 -1133
rect 3051 -1251 3067 -1133
rect 2757 -1293 3067 -1251
rect 2757 -1411 2773 -1293
rect 2891 -1411 2933 -1293
rect 3051 -1411 3067 -1293
rect -2443 -1731 -2427 -1613
rect -2309 -1731 -2267 -1613
rect -2149 -1731 -2133 -1613
rect -2443 -1773 -2133 -1731
rect -2443 -1891 -2427 -1773
rect -2309 -1891 -2267 -1773
rect -2149 -1891 -2133 -1773
rect -2443 -1907 -2133 -1891
rect 2757 -1907 3067 -1411
rect 4617 347447 4927 354061
rect 4617 347329 4633 347447
rect 4751 347329 4793 347447
rect 4911 347329 4927 347447
rect 4617 347287 4927 347329
rect 4617 347169 4633 347287
rect 4751 347169 4793 347287
rect 4911 347169 4927 347287
rect 4617 329447 4927 347169
rect 4617 329329 4633 329447
rect 4751 329329 4793 329447
rect 4911 329329 4927 329447
rect 4617 329287 4927 329329
rect 4617 329169 4633 329287
rect 4751 329169 4793 329287
rect 4911 329169 4927 329287
rect 4617 311447 4927 329169
rect 4617 311329 4633 311447
rect 4751 311329 4793 311447
rect 4911 311329 4927 311447
rect 4617 311287 4927 311329
rect 4617 311169 4633 311287
rect 4751 311169 4793 311287
rect 4911 311169 4927 311287
rect 4617 293447 4927 311169
rect 4617 293329 4633 293447
rect 4751 293329 4793 293447
rect 4911 293329 4927 293447
rect 4617 293287 4927 293329
rect 4617 293169 4633 293287
rect 4751 293169 4793 293287
rect 4911 293169 4927 293287
rect 4617 275447 4927 293169
rect 4617 275329 4633 275447
rect 4751 275329 4793 275447
rect 4911 275329 4927 275447
rect 4617 275287 4927 275329
rect 4617 275169 4633 275287
rect 4751 275169 4793 275287
rect 4911 275169 4927 275287
rect 4617 257447 4927 275169
rect 4617 257329 4633 257447
rect 4751 257329 4793 257447
rect 4911 257329 4927 257447
rect 4617 257287 4927 257329
rect 4617 257169 4633 257287
rect 4751 257169 4793 257287
rect 4911 257169 4927 257287
rect 4617 239447 4927 257169
rect 4617 239329 4633 239447
rect 4751 239329 4793 239447
rect 4911 239329 4927 239447
rect 4617 239287 4927 239329
rect 4617 239169 4633 239287
rect 4751 239169 4793 239287
rect 4911 239169 4927 239287
rect 4617 221447 4927 239169
rect 4617 221329 4633 221447
rect 4751 221329 4793 221447
rect 4911 221329 4927 221447
rect 4617 221287 4927 221329
rect 4617 221169 4633 221287
rect 4751 221169 4793 221287
rect 4911 221169 4927 221287
rect 4617 203447 4927 221169
rect 4617 203329 4633 203447
rect 4751 203329 4793 203447
rect 4911 203329 4927 203447
rect 4617 203287 4927 203329
rect 4617 203169 4633 203287
rect 4751 203169 4793 203287
rect 4911 203169 4927 203287
rect 4617 185447 4927 203169
rect 4617 185329 4633 185447
rect 4751 185329 4793 185447
rect 4911 185329 4927 185447
rect 4617 185287 4927 185329
rect 4617 185169 4633 185287
rect 4751 185169 4793 185287
rect 4911 185169 4927 185287
rect 4617 167447 4927 185169
rect 4617 167329 4633 167447
rect 4751 167329 4793 167447
rect 4911 167329 4927 167447
rect 4617 167287 4927 167329
rect 4617 167169 4633 167287
rect 4751 167169 4793 167287
rect 4911 167169 4927 167287
rect 4617 149447 4927 167169
rect 4617 149329 4633 149447
rect 4751 149329 4793 149447
rect 4911 149329 4927 149447
rect 4617 149287 4927 149329
rect 4617 149169 4633 149287
rect 4751 149169 4793 149287
rect 4911 149169 4927 149287
rect 4617 131447 4927 149169
rect 4617 131329 4633 131447
rect 4751 131329 4793 131447
rect 4911 131329 4927 131447
rect 4617 131287 4927 131329
rect 4617 131169 4633 131287
rect 4751 131169 4793 131287
rect 4911 131169 4927 131287
rect 4617 113447 4927 131169
rect 4617 113329 4633 113447
rect 4751 113329 4793 113447
rect 4911 113329 4927 113447
rect 4617 113287 4927 113329
rect 4617 113169 4633 113287
rect 4751 113169 4793 113287
rect 4911 113169 4927 113287
rect 4617 95447 4927 113169
rect 4617 95329 4633 95447
rect 4751 95329 4793 95447
rect 4911 95329 4927 95447
rect 4617 95287 4927 95329
rect 4617 95169 4633 95287
rect 4751 95169 4793 95287
rect 4911 95169 4927 95287
rect 4617 77447 4927 95169
rect 4617 77329 4633 77447
rect 4751 77329 4793 77447
rect 4911 77329 4927 77447
rect 4617 77287 4927 77329
rect 4617 77169 4633 77287
rect 4751 77169 4793 77287
rect 4911 77169 4927 77287
rect 4617 59447 4927 77169
rect 4617 59329 4633 59447
rect 4751 59329 4793 59447
rect 4911 59329 4927 59447
rect 4617 59287 4927 59329
rect 4617 59169 4633 59287
rect 4751 59169 4793 59287
rect 4911 59169 4927 59287
rect 4617 41447 4927 59169
rect 4617 41329 4633 41447
rect 4751 41329 4793 41447
rect 4911 41329 4927 41447
rect 4617 41287 4927 41329
rect 4617 41169 4633 41287
rect 4751 41169 4793 41287
rect 4911 41169 4927 41287
rect 4617 23447 4927 41169
rect 4617 23329 4633 23447
rect 4751 23329 4793 23447
rect 4911 23329 4927 23447
rect 4617 23287 4927 23329
rect 4617 23169 4633 23287
rect 4751 23169 4793 23287
rect 4911 23169 4927 23287
rect 4617 5447 4927 23169
rect 4617 5329 4633 5447
rect 4751 5329 4793 5447
rect 4911 5329 4927 5447
rect 4617 5287 4927 5329
rect 4617 5169 4633 5287
rect 4751 5169 4793 5287
rect 4911 5169 4927 5287
rect -2923 -2211 -2907 -2093
rect -2789 -2211 -2747 -2093
rect -2629 -2211 -2613 -2093
rect -2923 -2253 -2613 -2211
rect -2923 -2371 -2907 -2253
rect -2789 -2371 -2747 -2253
rect -2629 -2371 -2613 -2253
rect -2923 -2387 -2613 -2371
rect 4617 -2093 4927 5169
rect 4617 -2211 4633 -2093
rect 4751 -2211 4793 -2093
rect 4911 -2211 4927 -2093
rect 4617 -2253 4927 -2211
rect 4617 -2371 4633 -2253
rect 4751 -2371 4793 -2253
rect 4911 -2371 4927 -2253
rect -3403 -2691 -3387 -2573
rect -3269 -2691 -3227 -2573
rect -3109 -2691 -3093 -2573
rect -3403 -2733 -3093 -2691
rect -3403 -2851 -3387 -2733
rect -3269 -2851 -3227 -2733
rect -3109 -2851 -3093 -2733
rect -3403 -2867 -3093 -2851
rect 4617 -2867 4927 -2371
rect 6477 349307 6787 355021
rect 15477 355779 15787 355795
rect 15477 355661 15493 355779
rect 15611 355661 15653 355779
rect 15771 355661 15787 355779
rect 15477 355619 15787 355661
rect 15477 355501 15493 355619
rect 15611 355501 15653 355619
rect 15771 355501 15787 355619
rect 13617 354819 13927 354835
rect 13617 354701 13633 354819
rect 13751 354701 13793 354819
rect 13911 354701 13927 354819
rect 13617 354659 13927 354701
rect 13617 354541 13633 354659
rect 13751 354541 13793 354659
rect 13911 354541 13927 354659
rect 11757 353859 12067 353875
rect 11757 353741 11773 353859
rect 11891 353741 11933 353859
rect 12051 353741 12067 353859
rect 11757 353699 12067 353741
rect 11757 353581 11773 353699
rect 11891 353581 11933 353699
rect 12051 353581 12067 353699
rect 6477 349189 6493 349307
rect 6611 349189 6653 349307
rect 6771 349189 6787 349307
rect 6477 349147 6787 349189
rect 6477 349029 6493 349147
rect 6611 349029 6653 349147
rect 6771 349029 6787 349147
rect 6477 331307 6787 349029
rect 6477 331189 6493 331307
rect 6611 331189 6653 331307
rect 6771 331189 6787 331307
rect 6477 331147 6787 331189
rect 6477 331029 6493 331147
rect 6611 331029 6653 331147
rect 6771 331029 6787 331147
rect 6477 313307 6787 331029
rect 6477 313189 6493 313307
rect 6611 313189 6653 313307
rect 6771 313189 6787 313307
rect 6477 313147 6787 313189
rect 6477 313029 6493 313147
rect 6611 313029 6653 313147
rect 6771 313029 6787 313147
rect 6477 295307 6787 313029
rect 6477 295189 6493 295307
rect 6611 295189 6653 295307
rect 6771 295189 6787 295307
rect 6477 295147 6787 295189
rect 6477 295029 6493 295147
rect 6611 295029 6653 295147
rect 6771 295029 6787 295147
rect 6477 277307 6787 295029
rect 6477 277189 6493 277307
rect 6611 277189 6653 277307
rect 6771 277189 6787 277307
rect 6477 277147 6787 277189
rect 6477 277029 6493 277147
rect 6611 277029 6653 277147
rect 6771 277029 6787 277147
rect 6477 259307 6787 277029
rect 6477 259189 6493 259307
rect 6611 259189 6653 259307
rect 6771 259189 6787 259307
rect 6477 259147 6787 259189
rect 6477 259029 6493 259147
rect 6611 259029 6653 259147
rect 6771 259029 6787 259147
rect 6477 241307 6787 259029
rect 6477 241189 6493 241307
rect 6611 241189 6653 241307
rect 6771 241189 6787 241307
rect 6477 241147 6787 241189
rect 6477 241029 6493 241147
rect 6611 241029 6653 241147
rect 6771 241029 6787 241147
rect 6477 223307 6787 241029
rect 6477 223189 6493 223307
rect 6611 223189 6653 223307
rect 6771 223189 6787 223307
rect 6477 223147 6787 223189
rect 6477 223029 6493 223147
rect 6611 223029 6653 223147
rect 6771 223029 6787 223147
rect 6477 205307 6787 223029
rect 6477 205189 6493 205307
rect 6611 205189 6653 205307
rect 6771 205189 6787 205307
rect 6477 205147 6787 205189
rect 6477 205029 6493 205147
rect 6611 205029 6653 205147
rect 6771 205029 6787 205147
rect 6477 187307 6787 205029
rect 6477 187189 6493 187307
rect 6611 187189 6653 187307
rect 6771 187189 6787 187307
rect 6477 187147 6787 187189
rect 6477 187029 6493 187147
rect 6611 187029 6653 187147
rect 6771 187029 6787 187147
rect 6477 169307 6787 187029
rect 6477 169189 6493 169307
rect 6611 169189 6653 169307
rect 6771 169189 6787 169307
rect 6477 169147 6787 169189
rect 6477 169029 6493 169147
rect 6611 169029 6653 169147
rect 6771 169029 6787 169147
rect 6477 151307 6787 169029
rect 6477 151189 6493 151307
rect 6611 151189 6653 151307
rect 6771 151189 6787 151307
rect 6477 151147 6787 151189
rect 6477 151029 6493 151147
rect 6611 151029 6653 151147
rect 6771 151029 6787 151147
rect 6477 133307 6787 151029
rect 6477 133189 6493 133307
rect 6611 133189 6653 133307
rect 6771 133189 6787 133307
rect 6477 133147 6787 133189
rect 6477 133029 6493 133147
rect 6611 133029 6653 133147
rect 6771 133029 6787 133147
rect 6477 115307 6787 133029
rect 6477 115189 6493 115307
rect 6611 115189 6653 115307
rect 6771 115189 6787 115307
rect 6477 115147 6787 115189
rect 6477 115029 6493 115147
rect 6611 115029 6653 115147
rect 6771 115029 6787 115147
rect 6477 97307 6787 115029
rect 6477 97189 6493 97307
rect 6611 97189 6653 97307
rect 6771 97189 6787 97307
rect 6477 97147 6787 97189
rect 6477 97029 6493 97147
rect 6611 97029 6653 97147
rect 6771 97029 6787 97147
rect 6477 79307 6787 97029
rect 6477 79189 6493 79307
rect 6611 79189 6653 79307
rect 6771 79189 6787 79307
rect 6477 79147 6787 79189
rect 6477 79029 6493 79147
rect 6611 79029 6653 79147
rect 6771 79029 6787 79147
rect 6477 61307 6787 79029
rect 6477 61189 6493 61307
rect 6611 61189 6653 61307
rect 6771 61189 6787 61307
rect 6477 61147 6787 61189
rect 6477 61029 6493 61147
rect 6611 61029 6653 61147
rect 6771 61029 6787 61147
rect 6477 43307 6787 61029
rect 6477 43189 6493 43307
rect 6611 43189 6653 43307
rect 6771 43189 6787 43307
rect 6477 43147 6787 43189
rect 6477 43029 6493 43147
rect 6611 43029 6653 43147
rect 6771 43029 6787 43147
rect 6477 25307 6787 43029
rect 6477 25189 6493 25307
rect 6611 25189 6653 25307
rect 6771 25189 6787 25307
rect 6477 25147 6787 25189
rect 6477 25029 6493 25147
rect 6611 25029 6653 25147
rect 6771 25029 6787 25147
rect 6477 7307 6787 25029
rect 6477 7189 6493 7307
rect 6611 7189 6653 7307
rect 6771 7189 6787 7307
rect 6477 7147 6787 7189
rect 6477 7029 6493 7147
rect 6611 7029 6653 7147
rect 6771 7029 6787 7147
rect -3883 -3171 -3867 -3053
rect -3749 -3171 -3707 -3053
rect -3589 -3171 -3573 -3053
rect -3883 -3213 -3573 -3171
rect -3883 -3331 -3867 -3213
rect -3749 -3331 -3707 -3213
rect -3589 -3331 -3573 -3213
rect -3883 -3347 -3573 -3331
rect 6477 -3053 6787 7029
rect 9897 352899 10207 352915
rect 9897 352781 9913 352899
rect 10031 352781 10073 352899
rect 10191 352781 10207 352899
rect 9897 352739 10207 352781
rect 9897 352621 9913 352739
rect 10031 352621 10073 352739
rect 10191 352621 10207 352739
rect 9897 334727 10207 352621
rect 9897 334609 9913 334727
rect 10031 334609 10073 334727
rect 10191 334609 10207 334727
rect 9897 334567 10207 334609
rect 9897 334449 9913 334567
rect 10031 334449 10073 334567
rect 10191 334449 10207 334567
rect 9897 316727 10207 334449
rect 9897 316609 9913 316727
rect 10031 316609 10073 316727
rect 10191 316609 10207 316727
rect 9897 316567 10207 316609
rect 9897 316449 9913 316567
rect 10031 316449 10073 316567
rect 10191 316449 10207 316567
rect 9897 298727 10207 316449
rect 9897 298609 9913 298727
rect 10031 298609 10073 298727
rect 10191 298609 10207 298727
rect 9897 298567 10207 298609
rect 9897 298449 9913 298567
rect 10031 298449 10073 298567
rect 10191 298449 10207 298567
rect 9897 280727 10207 298449
rect 9897 280609 9913 280727
rect 10031 280609 10073 280727
rect 10191 280609 10207 280727
rect 9897 280567 10207 280609
rect 9897 280449 9913 280567
rect 10031 280449 10073 280567
rect 10191 280449 10207 280567
rect 9897 262727 10207 280449
rect 9897 262609 9913 262727
rect 10031 262609 10073 262727
rect 10191 262609 10207 262727
rect 9897 262567 10207 262609
rect 9897 262449 9913 262567
rect 10031 262449 10073 262567
rect 10191 262449 10207 262567
rect 9897 244727 10207 262449
rect 9897 244609 9913 244727
rect 10031 244609 10073 244727
rect 10191 244609 10207 244727
rect 9897 244567 10207 244609
rect 9897 244449 9913 244567
rect 10031 244449 10073 244567
rect 10191 244449 10207 244567
rect 9897 226727 10207 244449
rect 9897 226609 9913 226727
rect 10031 226609 10073 226727
rect 10191 226609 10207 226727
rect 9897 226567 10207 226609
rect 9897 226449 9913 226567
rect 10031 226449 10073 226567
rect 10191 226449 10207 226567
rect 9897 208727 10207 226449
rect 9897 208609 9913 208727
rect 10031 208609 10073 208727
rect 10191 208609 10207 208727
rect 9897 208567 10207 208609
rect 9897 208449 9913 208567
rect 10031 208449 10073 208567
rect 10191 208449 10207 208567
rect 9897 190727 10207 208449
rect 9897 190609 9913 190727
rect 10031 190609 10073 190727
rect 10191 190609 10207 190727
rect 9897 190567 10207 190609
rect 9897 190449 9913 190567
rect 10031 190449 10073 190567
rect 10191 190449 10207 190567
rect 9897 172727 10207 190449
rect 9897 172609 9913 172727
rect 10031 172609 10073 172727
rect 10191 172609 10207 172727
rect 9897 172567 10207 172609
rect 9897 172449 9913 172567
rect 10031 172449 10073 172567
rect 10191 172449 10207 172567
rect 9897 154727 10207 172449
rect 9897 154609 9913 154727
rect 10031 154609 10073 154727
rect 10191 154609 10207 154727
rect 9897 154567 10207 154609
rect 9897 154449 9913 154567
rect 10031 154449 10073 154567
rect 10191 154449 10207 154567
rect 9897 136727 10207 154449
rect 9897 136609 9913 136727
rect 10031 136609 10073 136727
rect 10191 136609 10207 136727
rect 9897 136567 10207 136609
rect 9897 136449 9913 136567
rect 10031 136449 10073 136567
rect 10191 136449 10207 136567
rect 9897 118727 10207 136449
rect 9897 118609 9913 118727
rect 10031 118609 10073 118727
rect 10191 118609 10207 118727
rect 9897 118567 10207 118609
rect 9897 118449 9913 118567
rect 10031 118449 10073 118567
rect 10191 118449 10207 118567
rect 9897 100727 10207 118449
rect 9897 100609 9913 100727
rect 10031 100609 10073 100727
rect 10191 100609 10207 100727
rect 9897 100567 10207 100609
rect 9897 100449 9913 100567
rect 10031 100449 10073 100567
rect 10191 100449 10207 100567
rect 9897 82727 10207 100449
rect 9897 82609 9913 82727
rect 10031 82609 10073 82727
rect 10191 82609 10207 82727
rect 9897 82567 10207 82609
rect 9897 82449 9913 82567
rect 10031 82449 10073 82567
rect 10191 82449 10207 82567
rect 9897 64727 10207 82449
rect 9897 64609 9913 64727
rect 10031 64609 10073 64727
rect 10191 64609 10207 64727
rect 9897 64567 10207 64609
rect 9897 64449 9913 64567
rect 10031 64449 10073 64567
rect 10191 64449 10207 64567
rect 9897 46727 10207 64449
rect 9897 46609 9913 46727
rect 10031 46609 10073 46727
rect 10191 46609 10207 46727
rect 9897 46567 10207 46609
rect 9897 46449 9913 46567
rect 10031 46449 10073 46567
rect 10191 46449 10207 46567
rect 9897 28727 10207 46449
rect 9897 28609 9913 28727
rect 10031 28609 10073 28727
rect 10191 28609 10207 28727
rect 9897 28567 10207 28609
rect 9897 28449 9913 28567
rect 10031 28449 10073 28567
rect 10191 28449 10207 28567
rect 9897 10727 10207 28449
rect 9897 10609 9913 10727
rect 10031 10609 10073 10727
rect 10191 10609 10207 10727
rect 9897 10567 10207 10609
rect 9897 10449 9913 10567
rect 10031 10449 10073 10567
rect 10191 10449 10207 10567
rect 9897 -653 10207 10449
rect 9897 -771 9913 -653
rect 10031 -771 10073 -653
rect 10191 -771 10207 -653
rect 9897 -813 10207 -771
rect 9897 -931 9913 -813
rect 10031 -931 10073 -813
rect 10191 -931 10207 -813
rect 9897 -947 10207 -931
rect 11757 336587 12067 353581
rect 11757 336469 11773 336587
rect 11891 336469 11933 336587
rect 12051 336469 12067 336587
rect 11757 336427 12067 336469
rect 11757 336309 11773 336427
rect 11891 336309 11933 336427
rect 12051 336309 12067 336427
rect 11757 318587 12067 336309
rect 11757 318469 11773 318587
rect 11891 318469 11933 318587
rect 12051 318469 12067 318587
rect 11757 318427 12067 318469
rect 11757 318309 11773 318427
rect 11891 318309 11933 318427
rect 12051 318309 12067 318427
rect 11757 300587 12067 318309
rect 11757 300469 11773 300587
rect 11891 300469 11933 300587
rect 12051 300469 12067 300587
rect 11757 300427 12067 300469
rect 11757 300309 11773 300427
rect 11891 300309 11933 300427
rect 12051 300309 12067 300427
rect 11757 282587 12067 300309
rect 11757 282469 11773 282587
rect 11891 282469 11933 282587
rect 12051 282469 12067 282587
rect 11757 282427 12067 282469
rect 11757 282309 11773 282427
rect 11891 282309 11933 282427
rect 12051 282309 12067 282427
rect 11757 264587 12067 282309
rect 11757 264469 11773 264587
rect 11891 264469 11933 264587
rect 12051 264469 12067 264587
rect 11757 264427 12067 264469
rect 11757 264309 11773 264427
rect 11891 264309 11933 264427
rect 12051 264309 12067 264427
rect 11757 246587 12067 264309
rect 11757 246469 11773 246587
rect 11891 246469 11933 246587
rect 12051 246469 12067 246587
rect 11757 246427 12067 246469
rect 11757 246309 11773 246427
rect 11891 246309 11933 246427
rect 12051 246309 12067 246427
rect 11757 228587 12067 246309
rect 11757 228469 11773 228587
rect 11891 228469 11933 228587
rect 12051 228469 12067 228587
rect 11757 228427 12067 228469
rect 11757 228309 11773 228427
rect 11891 228309 11933 228427
rect 12051 228309 12067 228427
rect 11757 210587 12067 228309
rect 11757 210469 11773 210587
rect 11891 210469 11933 210587
rect 12051 210469 12067 210587
rect 11757 210427 12067 210469
rect 11757 210309 11773 210427
rect 11891 210309 11933 210427
rect 12051 210309 12067 210427
rect 11757 192587 12067 210309
rect 11757 192469 11773 192587
rect 11891 192469 11933 192587
rect 12051 192469 12067 192587
rect 11757 192427 12067 192469
rect 11757 192309 11773 192427
rect 11891 192309 11933 192427
rect 12051 192309 12067 192427
rect 11757 174587 12067 192309
rect 11757 174469 11773 174587
rect 11891 174469 11933 174587
rect 12051 174469 12067 174587
rect 11757 174427 12067 174469
rect 11757 174309 11773 174427
rect 11891 174309 11933 174427
rect 12051 174309 12067 174427
rect 11757 156587 12067 174309
rect 11757 156469 11773 156587
rect 11891 156469 11933 156587
rect 12051 156469 12067 156587
rect 11757 156427 12067 156469
rect 11757 156309 11773 156427
rect 11891 156309 11933 156427
rect 12051 156309 12067 156427
rect 11757 138587 12067 156309
rect 11757 138469 11773 138587
rect 11891 138469 11933 138587
rect 12051 138469 12067 138587
rect 11757 138427 12067 138469
rect 11757 138309 11773 138427
rect 11891 138309 11933 138427
rect 12051 138309 12067 138427
rect 11757 120587 12067 138309
rect 11757 120469 11773 120587
rect 11891 120469 11933 120587
rect 12051 120469 12067 120587
rect 11757 120427 12067 120469
rect 11757 120309 11773 120427
rect 11891 120309 11933 120427
rect 12051 120309 12067 120427
rect 11757 102587 12067 120309
rect 11757 102469 11773 102587
rect 11891 102469 11933 102587
rect 12051 102469 12067 102587
rect 11757 102427 12067 102469
rect 11757 102309 11773 102427
rect 11891 102309 11933 102427
rect 12051 102309 12067 102427
rect 11757 84587 12067 102309
rect 11757 84469 11773 84587
rect 11891 84469 11933 84587
rect 12051 84469 12067 84587
rect 11757 84427 12067 84469
rect 11757 84309 11773 84427
rect 11891 84309 11933 84427
rect 12051 84309 12067 84427
rect 11757 66587 12067 84309
rect 11757 66469 11773 66587
rect 11891 66469 11933 66587
rect 12051 66469 12067 66587
rect 11757 66427 12067 66469
rect 11757 66309 11773 66427
rect 11891 66309 11933 66427
rect 12051 66309 12067 66427
rect 11757 48587 12067 66309
rect 11757 48469 11773 48587
rect 11891 48469 11933 48587
rect 12051 48469 12067 48587
rect 11757 48427 12067 48469
rect 11757 48309 11773 48427
rect 11891 48309 11933 48427
rect 12051 48309 12067 48427
rect 11757 30587 12067 48309
rect 11757 30469 11773 30587
rect 11891 30469 11933 30587
rect 12051 30469 12067 30587
rect 11757 30427 12067 30469
rect 11757 30309 11773 30427
rect 11891 30309 11933 30427
rect 12051 30309 12067 30427
rect 11757 12587 12067 30309
rect 11757 12469 11773 12587
rect 11891 12469 11933 12587
rect 12051 12469 12067 12587
rect 11757 12427 12067 12469
rect 11757 12309 11773 12427
rect 11891 12309 11933 12427
rect 12051 12309 12067 12427
rect 11757 -1613 12067 12309
rect 11757 -1731 11773 -1613
rect 11891 -1731 11933 -1613
rect 12051 -1731 12067 -1613
rect 11757 -1773 12067 -1731
rect 11757 -1891 11773 -1773
rect 11891 -1891 11933 -1773
rect 12051 -1891 12067 -1773
rect 11757 -1907 12067 -1891
rect 13617 338447 13927 354541
rect 13617 338329 13633 338447
rect 13751 338329 13793 338447
rect 13911 338329 13927 338447
rect 13617 338287 13927 338329
rect 13617 338169 13633 338287
rect 13751 338169 13793 338287
rect 13911 338169 13927 338287
rect 13617 320447 13927 338169
rect 13617 320329 13633 320447
rect 13751 320329 13793 320447
rect 13911 320329 13927 320447
rect 13617 320287 13927 320329
rect 13617 320169 13633 320287
rect 13751 320169 13793 320287
rect 13911 320169 13927 320287
rect 13617 302447 13927 320169
rect 13617 302329 13633 302447
rect 13751 302329 13793 302447
rect 13911 302329 13927 302447
rect 13617 302287 13927 302329
rect 13617 302169 13633 302287
rect 13751 302169 13793 302287
rect 13911 302169 13927 302287
rect 13617 284447 13927 302169
rect 13617 284329 13633 284447
rect 13751 284329 13793 284447
rect 13911 284329 13927 284447
rect 13617 284287 13927 284329
rect 13617 284169 13633 284287
rect 13751 284169 13793 284287
rect 13911 284169 13927 284287
rect 13617 266447 13927 284169
rect 13617 266329 13633 266447
rect 13751 266329 13793 266447
rect 13911 266329 13927 266447
rect 13617 266287 13927 266329
rect 13617 266169 13633 266287
rect 13751 266169 13793 266287
rect 13911 266169 13927 266287
rect 13617 248447 13927 266169
rect 13617 248329 13633 248447
rect 13751 248329 13793 248447
rect 13911 248329 13927 248447
rect 13617 248287 13927 248329
rect 13617 248169 13633 248287
rect 13751 248169 13793 248287
rect 13911 248169 13927 248287
rect 13617 230447 13927 248169
rect 13617 230329 13633 230447
rect 13751 230329 13793 230447
rect 13911 230329 13927 230447
rect 13617 230287 13927 230329
rect 13617 230169 13633 230287
rect 13751 230169 13793 230287
rect 13911 230169 13927 230287
rect 13617 212447 13927 230169
rect 13617 212329 13633 212447
rect 13751 212329 13793 212447
rect 13911 212329 13927 212447
rect 13617 212287 13927 212329
rect 13617 212169 13633 212287
rect 13751 212169 13793 212287
rect 13911 212169 13927 212287
rect 13617 194447 13927 212169
rect 13617 194329 13633 194447
rect 13751 194329 13793 194447
rect 13911 194329 13927 194447
rect 13617 194287 13927 194329
rect 13617 194169 13633 194287
rect 13751 194169 13793 194287
rect 13911 194169 13927 194287
rect 13617 176447 13927 194169
rect 13617 176329 13633 176447
rect 13751 176329 13793 176447
rect 13911 176329 13927 176447
rect 13617 176287 13927 176329
rect 13617 176169 13633 176287
rect 13751 176169 13793 176287
rect 13911 176169 13927 176287
rect 13617 158447 13927 176169
rect 13617 158329 13633 158447
rect 13751 158329 13793 158447
rect 13911 158329 13927 158447
rect 13617 158287 13927 158329
rect 13617 158169 13633 158287
rect 13751 158169 13793 158287
rect 13911 158169 13927 158287
rect 13617 140447 13927 158169
rect 13617 140329 13633 140447
rect 13751 140329 13793 140447
rect 13911 140329 13927 140447
rect 13617 140287 13927 140329
rect 13617 140169 13633 140287
rect 13751 140169 13793 140287
rect 13911 140169 13927 140287
rect 13617 122447 13927 140169
rect 13617 122329 13633 122447
rect 13751 122329 13793 122447
rect 13911 122329 13927 122447
rect 13617 122287 13927 122329
rect 13617 122169 13633 122287
rect 13751 122169 13793 122287
rect 13911 122169 13927 122287
rect 13617 104447 13927 122169
rect 13617 104329 13633 104447
rect 13751 104329 13793 104447
rect 13911 104329 13927 104447
rect 13617 104287 13927 104329
rect 13617 104169 13633 104287
rect 13751 104169 13793 104287
rect 13911 104169 13927 104287
rect 13617 86447 13927 104169
rect 13617 86329 13633 86447
rect 13751 86329 13793 86447
rect 13911 86329 13927 86447
rect 13617 86287 13927 86329
rect 13617 86169 13633 86287
rect 13751 86169 13793 86287
rect 13911 86169 13927 86287
rect 13617 68447 13927 86169
rect 13617 68329 13633 68447
rect 13751 68329 13793 68447
rect 13911 68329 13927 68447
rect 13617 68287 13927 68329
rect 13617 68169 13633 68287
rect 13751 68169 13793 68287
rect 13911 68169 13927 68287
rect 13617 50447 13927 68169
rect 13617 50329 13633 50447
rect 13751 50329 13793 50447
rect 13911 50329 13927 50447
rect 13617 50287 13927 50329
rect 13617 50169 13633 50287
rect 13751 50169 13793 50287
rect 13911 50169 13927 50287
rect 13617 32447 13927 50169
rect 13617 32329 13633 32447
rect 13751 32329 13793 32447
rect 13911 32329 13927 32447
rect 13617 32287 13927 32329
rect 13617 32169 13633 32287
rect 13751 32169 13793 32287
rect 13911 32169 13927 32287
rect 13617 14447 13927 32169
rect 13617 14329 13633 14447
rect 13751 14329 13793 14447
rect 13911 14329 13927 14447
rect 13617 14287 13927 14329
rect 13617 14169 13633 14287
rect 13751 14169 13793 14287
rect 13911 14169 13927 14287
rect 13617 -2573 13927 14169
rect 13617 -2691 13633 -2573
rect 13751 -2691 13793 -2573
rect 13911 -2691 13927 -2573
rect 13617 -2733 13927 -2691
rect 13617 -2851 13633 -2733
rect 13751 -2851 13793 -2733
rect 13911 -2851 13927 -2733
rect 13617 -2867 13927 -2851
rect 15477 340307 15787 355501
rect 24477 355299 24787 355795
rect 24477 355181 24493 355299
rect 24611 355181 24653 355299
rect 24771 355181 24787 355299
rect 24477 355139 24787 355181
rect 24477 355021 24493 355139
rect 24611 355021 24653 355139
rect 24771 355021 24787 355139
rect 22617 354339 22927 354835
rect 22617 354221 22633 354339
rect 22751 354221 22793 354339
rect 22911 354221 22927 354339
rect 22617 354179 22927 354221
rect 22617 354061 22633 354179
rect 22751 354061 22793 354179
rect 22911 354061 22927 354179
rect 20757 353379 21067 353875
rect 20757 353261 20773 353379
rect 20891 353261 20933 353379
rect 21051 353261 21067 353379
rect 20757 353219 21067 353261
rect 20757 353101 20773 353219
rect 20891 353101 20933 353219
rect 21051 353101 21067 353219
rect 15477 340189 15493 340307
rect 15611 340189 15653 340307
rect 15771 340189 15787 340307
rect 15477 340147 15787 340189
rect 15477 340029 15493 340147
rect 15611 340029 15653 340147
rect 15771 340029 15787 340147
rect 15477 322307 15787 340029
rect 15477 322189 15493 322307
rect 15611 322189 15653 322307
rect 15771 322189 15787 322307
rect 15477 322147 15787 322189
rect 15477 322029 15493 322147
rect 15611 322029 15653 322147
rect 15771 322029 15787 322147
rect 15477 304307 15787 322029
rect 15477 304189 15493 304307
rect 15611 304189 15653 304307
rect 15771 304189 15787 304307
rect 15477 304147 15787 304189
rect 15477 304029 15493 304147
rect 15611 304029 15653 304147
rect 15771 304029 15787 304147
rect 15477 286307 15787 304029
rect 15477 286189 15493 286307
rect 15611 286189 15653 286307
rect 15771 286189 15787 286307
rect 15477 286147 15787 286189
rect 15477 286029 15493 286147
rect 15611 286029 15653 286147
rect 15771 286029 15787 286147
rect 15477 268307 15787 286029
rect 15477 268189 15493 268307
rect 15611 268189 15653 268307
rect 15771 268189 15787 268307
rect 15477 268147 15787 268189
rect 15477 268029 15493 268147
rect 15611 268029 15653 268147
rect 15771 268029 15787 268147
rect 15477 250307 15787 268029
rect 15477 250189 15493 250307
rect 15611 250189 15653 250307
rect 15771 250189 15787 250307
rect 15477 250147 15787 250189
rect 15477 250029 15493 250147
rect 15611 250029 15653 250147
rect 15771 250029 15787 250147
rect 15477 232307 15787 250029
rect 15477 232189 15493 232307
rect 15611 232189 15653 232307
rect 15771 232189 15787 232307
rect 15477 232147 15787 232189
rect 15477 232029 15493 232147
rect 15611 232029 15653 232147
rect 15771 232029 15787 232147
rect 15477 214307 15787 232029
rect 15477 214189 15493 214307
rect 15611 214189 15653 214307
rect 15771 214189 15787 214307
rect 15477 214147 15787 214189
rect 15477 214029 15493 214147
rect 15611 214029 15653 214147
rect 15771 214029 15787 214147
rect 15477 196307 15787 214029
rect 15477 196189 15493 196307
rect 15611 196189 15653 196307
rect 15771 196189 15787 196307
rect 15477 196147 15787 196189
rect 15477 196029 15493 196147
rect 15611 196029 15653 196147
rect 15771 196029 15787 196147
rect 15477 178307 15787 196029
rect 15477 178189 15493 178307
rect 15611 178189 15653 178307
rect 15771 178189 15787 178307
rect 15477 178147 15787 178189
rect 15477 178029 15493 178147
rect 15611 178029 15653 178147
rect 15771 178029 15787 178147
rect 15477 160307 15787 178029
rect 15477 160189 15493 160307
rect 15611 160189 15653 160307
rect 15771 160189 15787 160307
rect 15477 160147 15787 160189
rect 15477 160029 15493 160147
rect 15611 160029 15653 160147
rect 15771 160029 15787 160147
rect 15477 142307 15787 160029
rect 15477 142189 15493 142307
rect 15611 142189 15653 142307
rect 15771 142189 15787 142307
rect 15477 142147 15787 142189
rect 15477 142029 15493 142147
rect 15611 142029 15653 142147
rect 15771 142029 15787 142147
rect 15477 124307 15787 142029
rect 15477 124189 15493 124307
rect 15611 124189 15653 124307
rect 15771 124189 15787 124307
rect 15477 124147 15787 124189
rect 15477 124029 15493 124147
rect 15611 124029 15653 124147
rect 15771 124029 15787 124147
rect 15477 106307 15787 124029
rect 15477 106189 15493 106307
rect 15611 106189 15653 106307
rect 15771 106189 15787 106307
rect 15477 106147 15787 106189
rect 15477 106029 15493 106147
rect 15611 106029 15653 106147
rect 15771 106029 15787 106147
rect 15477 88307 15787 106029
rect 15477 88189 15493 88307
rect 15611 88189 15653 88307
rect 15771 88189 15787 88307
rect 15477 88147 15787 88189
rect 15477 88029 15493 88147
rect 15611 88029 15653 88147
rect 15771 88029 15787 88147
rect 15477 70307 15787 88029
rect 15477 70189 15493 70307
rect 15611 70189 15653 70307
rect 15771 70189 15787 70307
rect 15477 70147 15787 70189
rect 15477 70029 15493 70147
rect 15611 70029 15653 70147
rect 15771 70029 15787 70147
rect 15477 52307 15787 70029
rect 15477 52189 15493 52307
rect 15611 52189 15653 52307
rect 15771 52189 15787 52307
rect 15477 52147 15787 52189
rect 15477 52029 15493 52147
rect 15611 52029 15653 52147
rect 15771 52029 15787 52147
rect 15477 34307 15787 52029
rect 15477 34189 15493 34307
rect 15611 34189 15653 34307
rect 15771 34189 15787 34307
rect 15477 34147 15787 34189
rect 15477 34029 15493 34147
rect 15611 34029 15653 34147
rect 15771 34029 15787 34147
rect 15477 16307 15787 34029
rect 15477 16189 15493 16307
rect 15611 16189 15653 16307
rect 15771 16189 15787 16307
rect 15477 16147 15787 16189
rect 15477 16029 15493 16147
rect 15611 16029 15653 16147
rect 15771 16029 15787 16147
rect 6477 -3171 6493 -3053
rect 6611 -3171 6653 -3053
rect 6771 -3171 6787 -3053
rect 6477 -3213 6787 -3171
rect 6477 -3331 6493 -3213
rect 6611 -3331 6653 -3213
rect 6771 -3331 6787 -3213
rect -4363 -3651 -4347 -3533
rect -4229 -3651 -4187 -3533
rect -4069 -3651 -4053 -3533
rect -4363 -3693 -4053 -3651
rect -4363 -3811 -4347 -3693
rect -4229 -3811 -4187 -3693
rect -4069 -3811 -4053 -3693
rect -4363 -3827 -4053 -3811
rect 6477 -3827 6787 -3331
rect 15477 -3533 15787 16029
rect 18897 352419 19207 352915
rect 18897 352301 18913 352419
rect 19031 352301 19073 352419
rect 19191 352301 19207 352419
rect 18897 352259 19207 352301
rect 18897 352141 18913 352259
rect 19031 352141 19073 352259
rect 19191 352141 19207 352259
rect 18897 343727 19207 352141
rect 18897 343609 18913 343727
rect 19031 343609 19073 343727
rect 19191 343609 19207 343727
rect 18897 343567 19207 343609
rect 18897 343449 18913 343567
rect 19031 343449 19073 343567
rect 19191 343449 19207 343567
rect 18897 325727 19207 343449
rect 18897 325609 18913 325727
rect 19031 325609 19073 325727
rect 19191 325609 19207 325727
rect 18897 325567 19207 325609
rect 18897 325449 18913 325567
rect 19031 325449 19073 325567
rect 19191 325449 19207 325567
rect 18897 307727 19207 325449
rect 18897 307609 18913 307727
rect 19031 307609 19073 307727
rect 19191 307609 19207 307727
rect 18897 307567 19207 307609
rect 18897 307449 18913 307567
rect 19031 307449 19073 307567
rect 19191 307449 19207 307567
rect 18897 289727 19207 307449
rect 18897 289609 18913 289727
rect 19031 289609 19073 289727
rect 19191 289609 19207 289727
rect 18897 289567 19207 289609
rect 18897 289449 18913 289567
rect 19031 289449 19073 289567
rect 19191 289449 19207 289567
rect 18897 271727 19207 289449
rect 18897 271609 18913 271727
rect 19031 271609 19073 271727
rect 19191 271609 19207 271727
rect 18897 271567 19207 271609
rect 18897 271449 18913 271567
rect 19031 271449 19073 271567
rect 19191 271449 19207 271567
rect 18897 253727 19207 271449
rect 18897 253609 18913 253727
rect 19031 253609 19073 253727
rect 19191 253609 19207 253727
rect 18897 253567 19207 253609
rect 18897 253449 18913 253567
rect 19031 253449 19073 253567
rect 19191 253449 19207 253567
rect 18897 235727 19207 253449
rect 18897 235609 18913 235727
rect 19031 235609 19073 235727
rect 19191 235609 19207 235727
rect 18897 235567 19207 235609
rect 18897 235449 18913 235567
rect 19031 235449 19073 235567
rect 19191 235449 19207 235567
rect 18897 217727 19207 235449
rect 18897 217609 18913 217727
rect 19031 217609 19073 217727
rect 19191 217609 19207 217727
rect 18897 217567 19207 217609
rect 18897 217449 18913 217567
rect 19031 217449 19073 217567
rect 19191 217449 19207 217567
rect 18897 199727 19207 217449
rect 18897 199609 18913 199727
rect 19031 199609 19073 199727
rect 19191 199609 19207 199727
rect 18897 199567 19207 199609
rect 18897 199449 18913 199567
rect 19031 199449 19073 199567
rect 19191 199449 19207 199567
rect 18897 181727 19207 199449
rect 18897 181609 18913 181727
rect 19031 181609 19073 181727
rect 19191 181609 19207 181727
rect 18897 181567 19207 181609
rect 18897 181449 18913 181567
rect 19031 181449 19073 181567
rect 19191 181449 19207 181567
rect 18897 163727 19207 181449
rect 18897 163609 18913 163727
rect 19031 163609 19073 163727
rect 19191 163609 19207 163727
rect 18897 163567 19207 163609
rect 18897 163449 18913 163567
rect 19031 163449 19073 163567
rect 19191 163449 19207 163567
rect 18897 145727 19207 163449
rect 18897 145609 18913 145727
rect 19031 145609 19073 145727
rect 19191 145609 19207 145727
rect 18897 145567 19207 145609
rect 18897 145449 18913 145567
rect 19031 145449 19073 145567
rect 19191 145449 19207 145567
rect 18897 127727 19207 145449
rect 18897 127609 18913 127727
rect 19031 127609 19073 127727
rect 19191 127609 19207 127727
rect 18897 127567 19207 127609
rect 18897 127449 18913 127567
rect 19031 127449 19073 127567
rect 19191 127449 19207 127567
rect 18897 109727 19207 127449
rect 18897 109609 18913 109727
rect 19031 109609 19073 109727
rect 19191 109609 19207 109727
rect 18897 109567 19207 109609
rect 18897 109449 18913 109567
rect 19031 109449 19073 109567
rect 19191 109449 19207 109567
rect 18897 91727 19207 109449
rect 18897 91609 18913 91727
rect 19031 91609 19073 91727
rect 19191 91609 19207 91727
rect 18897 91567 19207 91609
rect 18897 91449 18913 91567
rect 19031 91449 19073 91567
rect 19191 91449 19207 91567
rect 18897 73727 19207 91449
rect 18897 73609 18913 73727
rect 19031 73609 19073 73727
rect 19191 73609 19207 73727
rect 18897 73567 19207 73609
rect 18897 73449 18913 73567
rect 19031 73449 19073 73567
rect 19191 73449 19207 73567
rect 18897 55727 19207 73449
rect 18897 55609 18913 55727
rect 19031 55609 19073 55727
rect 19191 55609 19207 55727
rect 18897 55567 19207 55609
rect 18897 55449 18913 55567
rect 19031 55449 19073 55567
rect 19191 55449 19207 55567
rect 18897 37727 19207 55449
rect 18897 37609 18913 37727
rect 19031 37609 19073 37727
rect 19191 37609 19207 37727
rect 18897 37567 19207 37609
rect 18897 37449 18913 37567
rect 19031 37449 19073 37567
rect 19191 37449 19207 37567
rect 18897 19727 19207 37449
rect 18897 19609 18913 19727
rect 19031 19609 19073 19727
rect 19191 19609 19207 19727
rect 18897 19567 19207 19609
rect 18897 19449 18913 19567
rect 19031 19449 19073 19567
rect 19191 19449 19207 19567
rect 18897 1727 19207 19449
rect 18897 1609 18913 1727
rect 19031 1609 19073 1727
rect 19191 1609 19207 1727
rect 18897 1567 19207 1609
rect 18897 1449 18913 1567
rect 19031 1449 19073 1567
rect 19191 1449 19207 1567
rect 18897 -173 19207 1449
rect 18897 -291 18913 -173
rect 19031 -291 19073 -173
rect 19191 -291 19207 -173
rect 18897 -333 19207 -291
rect 18897 -451 18913 -333
rect 19031 -451 19073 -333
rect 19191 -451 19207 -333
rect 18897 -947 19207 -451
rect 20757 345587 21067 353101
rect 20757 345469 20773 345587
rect 20891 345469 20933 345587
rect 21051 345469 21067 345587
rect 20757 345427 21067 345469
rect 20757 345309 20773 345427
rect 20891 345309 20933 345427
rect 21051 345309 21067 345427
rect 20757 327587 21067 345309
rect 20757 327469 20773 327587
rect 20891 327469 20933 327587
rect 21051 327469 21067 327587
rect 20757 327427 21067 327469
rect 20757 327309 20773 327427
rect 20891 327309 20933 327427
rect 21051 327309 21067 327427
rect 20757 309587 21067 327309
rect 20757 309469 20773 309587
rect 20891 309469 20933 309587
rect 21051 309469 21067 309587
rect 20757 309427 21067 309469
rect 20757 309309 20773 309427
rect 20891 309309 20933 309427
rect 21051 309309 21067 309427
rect 20757 291587 21067 309309
rect 20757 291469 20773 291587
rect 20891 291469 20933 291587
rect 21051 291469 21067 291587
rect 20757 291427 21067 291469
rect 20757 291309 20773 291427
rect 20891 291309 20933 291427
rect 21051 291309 21067 291427
rect 20757 273587 21067 291309
rect 20757 273469 20773 273587
rect 20891 273469 20933 273587
rect 21051 273469 21067 273587
rect 20757 273427 21067 273469
rect 20757 273309 20773 273427
rect 20891 273309 20933 273427
rect 21051 273309 21067 273427
rect 20757 255587 21067 273309
rect 20757 255469 20773 255587
rect 20891 255469 20933 255587
rect 21051 255469 21067 255587
rect 20757 255427 21067 255469
rect 20757 255309 20773 255427
rect 20891 255309 20933 255427
rect 21051 255309 21067 255427
rect 20757 237587 21067 255309
rect 20757 237469 20773 237587
rect 20891 237469 20933 237587
rect 21051 237469 21067 237587
rect 20757 237427 21067 237469
rect 20757 237309 20773 237427
rect 20891 237309 20933 237427
rect 21051 237309 21067 237427
rect 20757 219587 21067 237309
rect 20757 219469 20773 219587
rect 20891 219469 20933 219587
rect 21051 219469 21067 219587
rect 20757 219427 21067 219469
rect 20757 219309 20773 219427
rect 20891 219309 20933 219427
rect 21051 219309 21067 219427
rect 20757 201587 21067 219309
rect 20757 201469 20773 201587
rect 20891 201469 20933 201587
rect 21051 201469 21067 201587
rect 20757 201427 21067 201469
rect 20757 201309 20773 201427
rect 20891 201309 20933 201427
rect 21051 201309 21067 201427
rect 20757 183587 21067 201309
rect 20757 183469 20773 183587
rect 20891 183469 20933 183587
rect 21051 183469 21067 183587
rect 20757 183427 21067 183469
rect 20757 183309 20773 183427
rect 20891 183309 20933 183427
rect 21051 183309 21067 183427
rect 20757 165587 21067 183309
rect 20757 165469 20773 165587
rect 20891 165469 20933 165587
rect 21051 165469 21067 165587
rect 20757 165427 21067 165469
rect 20757 165309 20773 165427
rect 20891 165309 20933 165427
rect 21051 165309 21067 165427
rect 20757 147587 21067 165309
rect 20757 147469 20773 147587
rect 20891 147469 20933 147587
rect 21051 147469 21067 147587
rect 20757 147427 21067 147469
rect 20757 147309 20773 147427
rect 20891 147309 20933 147427
rect 21051 147309 21067 147427
rect 20757 129587 21067 147309
rect 20757 129469 20773 129587
rect 20891 129469 20933 129587
rect 21051 129469 21067 129587
rect 20757 129427 21067 129469
rect 20757 129309 20773 129427
rect 20891 129309 20933 129427
rect 21051 129309 21067 129427
rect 20757 111587 21067 129309
rect 20757 111469 20773 111587
rect 20891 111469 20933 111587
rect 21051 111469 21067 111587
rect 20757 111427 21067 111469
rect 20757 111309 20773 111427
rect 20891 111309 20933 111427
rect 21051 111309 21067 111427
rect 20757 93587 21067 111309
rect 20757 93469 20773 93587
rect 20891 93469 20933 93587
rect 21051 93469 21067 93587
rect 20757 93427 21067 93469
rect 20757 93309 20773 93427
rect 20891 93309 20933 93427
rect 21051 93309 21067 93427
rect 20757 75587 21067 93309
rect 20757 75469 20773 75587
rect 20891 75469 20933 75587
rect 21051 75469 21067 75587
rect 20757 75427 21067 75469
rect 20757 75309 20773 75427
rect 20891 75309 20933 75427
rect 21051 75309 21067 75427
rect 20757 57587 21067 75309
rect 20757 57469 20773 57587
rect 20891 57469 20933 57587
rect 21051 57469 21067 57587
rect 20757 57427 21067 57469
rect 20757 57309 20773 57427
rect 20891 57309 20933 57427
rect 21051 57309 21067 57427
rect 20757 39587 21067 57309
rect 20757 39469 20773 39587
rect 20891 39469 20933 39587
rect 21051 39469 21067 39587
rect 20757 39427 21067 39469
rect 20757 39309 20773 39427
rect 20891 39309 20933 39427
rect 21051 39309 21067 39427
rect 20757 21587 21067 39309
rect 20757 21469 20773 21587
rect 20891 21469 20933 21587
rect 21051 21469 21067 21587
rect 20757 21427 21067 21469
rect 20757 21309 20773 21427
rect 20891 21309 20933 21427
rect 21051 21309 21067 21427
rect 20757 3587 21067 21309
rect 20757 3469 20773 3587
rect 20891 3469 20933 3587
rect 21051 3469 21067 3587
rect 20757 3427 21067 3469
rect 20757 3309 20773 3427
rect 20891 3309 20933 3427
rect 21051 3309 21067 3427
rect 20757 -1133 21067 3309
rect 20757 -1251 20773 -1133
rect 20891 -1251 20933 -1133
rect 21051 -1251 21067 -1133
rect 20757 -1293 21067 -1251
rect 20757 -1411 20773 -1293
rect 20891 -1411 20933 -1293
rect 21051 -1411 21067 -1293
rect 20757 -1907 21067 -1411
rect 22617 347447 22927 354061
rect 22617 347329 22633 347447
rect 22751 347329 22793 347447
rect 22911 347329 22927 347447
rect 22617 347287 22927 347329
rect 22617 347169 22633 347287
rect 22751 347169 22793 347287
rect 22911 347169 22927 347287
rect 22617 329447 22927 347169
rect 22617 329329 22633 329447
rect 22751 329329 22793 329447
rect 22911 329329 22927 329447
rect 22617 329287 22927 329329
rect 22617 329169 22633 329287
rect 22751 329169 22793 329287
rect 22911 329169 22927 329287
rect 22617 311447 22927 329169
rect 22617 311329 22633 311447
rect 22751 311329 22793 311447
rect 22911 311329 22927 311447
rect 22617 311287 22927 311329
rect 22617 311169 22633 311287
rect 22751 311169 22793 311287
rect 22911 311169 22927 311287
rect 22617 293447 22927 311169
rect 22617 293329 22633 293447
rect 22751 293329 22793 293447
rect 22911 293329 22927 293447
rect 22617 293287 22927 293329
rect 22617 293169 22633 293287
rect 22751 293169 22793 293287
rect 22911 293169 22927 293287
rect 22617 275447 22927 293169
rect 22617 275329 22633 275447
rect 22751 275329 22793 275447
rect 22911 275329 22927 275447
rect 22617 275287 22927 275329
rect 22617 275169 22633 275287
rect 22751 275169 22793 275287
rect 22911 275169 22927 275287
rect 22617 257447 22927 275169
rect 22617 257329 22633 257447
rect 22751 257329 22793 257447
rect 22911 257329 22927 257447
rect 22617 257287 22927 257329
rect 22617 257169 22633 257287
rect 22751 257169 22793 257287
rect 22911 257169 22927 257287
rect 22617 239447 22927 257169
rect 22617 239329 22633 239447
rect 22751 239329 22793 239447
rect 22911 239329 22927 239447
rect 22617 239287 22927 239329
rect 22617 239169 22633 239287
rect 22751 239169 22793 239287
rect 22911 239169 22927 239287
rect 22617 221447 22927 239169
rect 22617 221329 22633 221447
rect 22751 221329 22793 221447
rect 22911 221329 22927 221447
rect 22617 221287 22927 221329
rect 22617 221169 22633 221287
rect 22751 221169 22793 221287
rect 22911 221169 22927 221287
rect 22617 203447 22927 221169
rect 22617 203329 22633 203447
rect 22751 203329 22793 203447
rect 22911 203329 22927 203447
rect 22617 203287 22927 203329
rect 22617 203169 22633 203287
rect 22751 203169 22793 203287
rect 22911 203169 22927 203287
rect 22617 185447 22927 203169
rect 22617 185329 22633 185447
rect 22751 185329 22793 185447
rect 22911 185329 22927 185447
rect 22617 185287 22927 185329
rect 22617 185169 22633 185287
rect 22751 185169 22793 185287
rect 22911 185169 22927 185287
rect 22617 167447 22927 185169
rect 22617 167329 22633 167447
rect 22751 167329 22793 167447
rect 22911 167329 22927 167447
rect 22617 167287 22927 167329
rect 22617 167169 22633 167287
rect 22751 167169 22793 167287
rect 22911 167169 22927 167287
rect 22617 149447 22927 167169
rect 22617 149329 22633 149447
rect 22751 149329 22793 149447
rect 22911 149329 22927 149447
rect 22617 149287 22927 149329
rect 22617 149169 22633 149287
rect 22751 149169 22793 149287
rect 22911 149169 22927 149287
rect 22617 131447 22927 149169
rect 22617 131329 22633 131447
rect 22751 131329 22793 131447
rect 22911 131329 22927 131447
rect 22617 131287 22927 131329
rect 22617 131169 22633 131287
rect 22751 131169 22793 131287
rect 22911 131169 22927 131287
rect 22617 113447 22927 131169
rect 22617 113329 22633 113447
rect 22751 113329 22793 113447
rect 22911 113329 22927 113447
rect 22617 113287 22927 113329
rect 22617 113169 22633 113287
rect 22751 113169 22793 113287
rect 22911 113169 22927 113287
rect 22617 95447 22927 113169
rect 22617 95329 22633 95447
rect 22751 95329 22793 95447
rect 22911 95329 22927 95447
rect 22617 95287 22927 95329
rect 22617 95169 22633 95287
rect 22751 95169 22793 95287
rect 22911 95169 22927 95287
rect 22617 77447 22927 95169
rect 22617 77329 22633 77447
rect 22751 77329 22793 77447
rect 22911 77329 22927 77447
rect 22617 77287 22927 77329
rect 22617 77169 22633 77287
rect 22751 77169 22793 77287
rect 22911 77169 22927 77287
rect 22617 59447 22927 77169
rect 22617 59329 22633 59447
rect 22751 59329 22793 59447
rect 22911 59329 22927 59447
rect 22617 59287 22927 59329
rect 22617 59169 22633 59287
rect 22751 59169 22793 59287
rect 22911 59169 22927 59287
rect 22617 41447 22927 59169
rect 22617 41329 22633 41447
rect 22751 41329 22793 41447
rect 22911 41329 22927 41447
rect 22617 41287 22927 41329
rect 22617 41169 22633 41287
rect 22751 41169 22793 41287
rect 22911 41169 22927 41287
rect 22617 23447 22927 41169
rect 22617 23329 22633 23447
rect 22751 23329 22793 23447
rect 22911 23329 22927 23447
rect 22617 23287 22927 23329
rect 22617 23169 22633 23287
rect 22751 23169 22793 23287
rect 22911 23169 22927 23287
rect 22617 5447 22927 23169
rect 22617 5329 22633 5447
rect 22751 5329 22793 5447
rect 22911 5329 22927 5447
rect 22617 5287 22927 5329
rect 22617 5169 22633 5287
rect 22751 5169 22793 5287
rect 22911 5169 22927 5287
rect 22617 -2093 22927 5169
rect 22617 -2211 22633 -2093
rect 22751 -2211 22793 -2093
rect 22911 -2211 22927 -2093
rect 22617 -2253 22927 -2211
rect 22617 -2371 22633 -2253
rect 22751 -2371 22793 -2253
rect 22911 -2371 22927 -2253
rect 22617 -2867 22927 -2371
rect 24477 349307 24787 355021
rect 33477 355779 33787 355795
rect 33477 355661 33493 355779
rect 33611 355661 33653 355779
rect 33771 355661 33787 355779
rect 33477 355619 33787 355661
rect 33477 355501 33493 355619
rect 33611 355501 33653 355619
rect 33771 355501 33787 355619
rect 31617 354819 31927 354835
rect 31617 354701 31633 354819
rect 31751 354701 31793 354819
rect 31911 354701 31927 354819
rect 31617 354659 31927 354701
rect 31617 354541 31633 354659
rect 31751 354541 31793 354659
rect 31911 354541 31927 354659
rect 29757 353859 30067 353875
rect 29757 353741 29773 353859
rect 29891 353741 29933 353859
rect 30051 353741 30067 353859
rect 29757 353699 30067 353741
rect 29757 353581 29773 353699
rect 29891 353581 29933 353699
rect 30051 353581 30067 353699
rect 24477 349189 24493 349307
rect 24611 349189 24653 349307
rect 24771 349189 24787 349307
rect 24477 349147 24787 349189
rect 24477 349029 24493 349147
rect 24611 349029 24653 349147
rect 24771 349029 24787 349147
rect 24477 331307 24787 349029
rect 24477 331189 24493 331307
rect 24611 331189 24653 331307
rect 24771 331189 24787 331307
rect 24477 331147 24787 331189
rect 24477 331029 24493 331147
rect 24611 331029 24653 331147
rect 24771 331029 24787 331147
rect 24477 313307 24787 331029
rect 24477 313189 24493 313307
rect 24611 313189 24653 313307
rect 24771 313189 24787 313307
rect 24477 313147 24787 313189
rect 24477 313029 24493 313147
rect 24611 313029 24653 313147
rect 24771 313029 24787 313147
rect 24477 295307 24787 313029
rect 24477 295189 24493 295307
rect 24611 295189 24653 295307
rect 24771 295189 24787 295307
rect 24477 295147 24787 295189
rect 24477 295029 24493 295147
rect 24611 295029 24653 295147
rect 24771 295029 24787 295147
rect 24477 277307 24787 295029
rect 24477 277189 24493 277307
rect 24611 277189 24653 277307
rect 24771 277189 24787 277307
rect 24477 277147 24787 277189
rect 24477 277029 24493 277147
rect 24611 277029 24653 277147
rect 24771 277029 24787 277147
rect 24477 259307 24787 277029
rect 24477 259189 24493 259307
rect 24611 259189 24653 259307
rect 24771 259189 24787 259307
rect 24477 259147 24787 259189
rect 24477 259029 24493 259147
rect 24611 259029 24653 259147
rect 24771 259029 24787 259147
rect 24477 241307 24787 259029
rect 24477 241189 24493 241307
rect 24611 241189 24653 241307
rect 24771 241189 24787 241307
rect 24477 241147 24787 241189
rect 24477 241029 24493 241147
rect 24611 241029 24653 241147
rect 24771 241029 24787 241147
rect 24477 223307 24787 241029
rect 24477 223189 24493 223307
rect 24611 223189 24653 223307
rect 24771 223189 24787 223307
rect 24477 223147 24787 223189
rect 24477 223029 24493 223147
rect 24611 223029 24653 223147
rect 24771 223029 24787 223147
rect 24477 205307 24787 223029
rect 24477 205189 24493 205307
rect 24611 205189 24653 205307
rect 24771 205189 24787 205307
rect 24477 205147 24787 205189
rect 24477 205029 24493 205147
rect 24611 205029 24653 205147
rect 24771 205029 24787 205147
rect 24477 187307 24787 205029
rect 24477 187189 24493 187307
rect 24611 187189 24653 187307
rect 24771 187189 24787 187307
rect 24477 187147 24787 187189
rect 24477 187029 24493 187147
rect 24611 187029 24653 187147
rect 24771 187029 24787 187147
rect 24477 169307 24787 187029
rect 24477 169189 24493 169307
rect 24611 169189 24653 169307
rect 24771 169189 24787 169307
rect 24477 169147 24787 169189
rect 24477 169029 24493 169147
rect 24611 169029 24653 169147
rect 24771 169029 24787 169147
rect 24477 151307 24787 169029
rect 24477 151189 24493 151307
rect 24611 151189 24653 151307
rect 24771 151189 24787 151307
rect 24477 151147 24787 151189
rect 24477 151029 24493 151147
rect 24611 151029 24653 151147
rect 24771 151029 24787 151147
rect 24477 133307 24787 151029
rect 24477 133189 24493 133307
rect 24611 133189 24653 133307
rect 24771 133189 24787 133307
rect 24477 133147 24787 133189
rect 24477 133029 24493 133147
rect 24611 133029 24653 133147
rect 24771 133029 24787 133147
rect 24477 115307 24787 133029
rect 24477 115189 24493 115307
rect 24611 115189 24653 115307
rect 24771 115189 24787 115307
rect 24477 115147 24787 115189
rect 24477 115029 24493 115147
rect 24611 115029 24653 115147
rect 24771 115029 24787 115147
rect 24477 97307 24787 115029
rect 24477 97189 24493 97307
rect 24611 97189 24653 97307
rect 24771 97189 24787 97307
rect 24477 97147 24787 97189
rect 24477 97029 24493 97147
rect 24611 97029 24653 97147
rect 24771 97029 24787 97147
rect 24477 79307 24787 97029
rect 24477 79189 24493 79307
rect 24611 79189 24653 79307
rect 24771 79189 24787 79307
rect 24477 79147 24787 79189
rect 24477 79029 24493 79147
rect 24611 79029 24653 79147
rect 24771 79029 24787 79147
rect 24477 61307 24787 79029
rect 24477 61189 24493 61307
rect 24611 61189 24653 61307
rect 24771 61189 24787 61307
rect 24477 61147 24787 61189
rect 24477 61029 24493 61147
rect 24611 61029 24653 61147
rect 24771 61029 24787 61147
rect 24477 43307 24787 61029
rect 24477 43189 24493 43307
rect 24611 43189 24653 43307
rect 24771 43189 24787 43307
rect 24477 43147 24787 43189
rect 24477 43029 24493 43147
rect 24611 43029 24653 43147
rect 24771 43029 24787 43147
rect 24477 25307 24787 43029
rect 24477 25189 24493 25307
rect 24611 25189 24653 25307
rect 24771 25189 24787 25307
rect 24477 25147 24787 25189
rect 24477 25029 24493 25147
rect 24611 25029 24653 25147
rect 24771 25029 24787 25147
rect 24477 7307 24787 25029
rect 24477 7189 24493 7307
rect 24611 7189 24653 7307
rect 24771 7189 24787 7307
rect 24477 7147 24787 7189
rect 24477 7029 24493 7147
rect 24611 7029 24653 7147
rect 24771 7029 24787 7147
rect 15477 -3651 15493 -3533
rect 15611 -3651 15653 -3533
rect 15771 -3651 15787 -3533
rect 15477 -3693 15787 -3651
rect 15477 -3811 15493 -3693
rect 15611 -3811 15653 -3693
rect 15771 -3811 15787 -3693
rect 15477 -3827 15787 -3811
rect 24477 -3053 24787 7029
rect 27897 352899 28207 352915
rect 27897 352781 27913 352899
rect 28031 352781 28073 352899
rect 28191 352781 28207 352899
rect 27897 352739 28207 352781
rect 27897 352621 27913 352739
rect 28031 352621 28073 352739
rect 28191 352621 28207 352739
rect 27897 334727 28207 352621
rect 27897 334609 27913 334727
rect 28031 334609 28073 334727
rect 28191 334609 28207 334727
rect 27897 334567 28207 334609
rect 27897 334449 27913 334567
rect 28031 334449 28073 334567
rect 28191 334449 28207 334567
rect 27897 316727 28207 334449
rect 27897 316609 27913 316727
rect 28031 316609 28073 316727
rect 28191 316609 28207 316727
rect 27897 316567 28207 316609
rect 27897 316449 27913 316567
rect 28031 316449 28073 316567
rect 28191 316449 28207 316567
rect 27897 298727 28207 316449
rect 27897 298609 27913 298727
rect 28031 298609 28073 298727
rect 28191 298609 28207 298727
rect 27897 298567 28207 298609
rect 27897 298449 27913 298567
rect 28031 298449 28073 298567
rect 28191 298449 28207 298567
rect 27897 280727 28207 298449
rect 27897 280609 27913 280727
rect 28031 280609 28073 280727
rect 28191 280609 28207 280727
rect 27897 280567 28207 280609
rect 27897 280449 27913 280567
rect 28031 280449 28073 280567
rect 28191 280449 28207 280567
rect 27897 262727 28207 280449
rect 27897 262609 27913 262727
rect 28031 262609 28073 262727
rect 28191 262609 28207 262727
rect 27897 262567 28207 262609
rect 27897 262449 27913 262567
rect 28031 262449 28073 262567
rect 28191 262449 28207 262567
rect 27897 244727 28207 262449
rect 27897 244609 27913 244727
rect 28031 244609 28073 244727
rect 28191 244609 28207 244727
rect 27897 244567 28207 244609
rect 27897 244449 27913 244567
rect 28031 244449 28073 244567
rect 28191 244449 28207 244567
rect 27897 226727 28207 244449
rect 27897 226609 27913 226727
rect 28031 226609 28073 226727
rect 28191 226609 28207 226727
rect 27897 226567 28207 226609
rect 27897 226449 27913 226567
rect 28031 226449 28073 226567
rect 28191 226449 28207 226567
rect 27897 208727 28207 226449
rect 27897 208609 27913 208727
rect 28031 208609 28073 208727
rect 28191 208609 28207 208727
rect 27897 208567 28207 208609
rect 27897 208449 27913 208567
rect 28031 208449 28073 208567
rect 28191 208449 28207 208567
rect 27897 190727 28207 208449
rect 27897 190609 27913 190727
rect 28031 190609 28073 190727
rect 28191 190609 28207 190727
rect 27897 190567 28207 190609
rect 27897 190449 27913 190567
rect 28031 190449 28073 190567
rect 28191 190449 28207 190567
rect 27897 172727 28207 190449
rect 27897 172609 27913 172727
rect 28031 172609 28073 172727
rect 28191 172609 28207 172727
rect 27897 172567 28207 172609
rect 27897 172449 27913 172567
rect 28031 172449 28073 172567
rect 28191 172449 28207 172567
rect 27897 154727 28207 172449
rect 27897 154609 27913 154727
rect 28031 154609 28073 154727
rect 28191 154609 28207 154727
rect 27897 154567 28207 154609
rect 27897 154449 27913 154567
rect 28031 154449 28073 154567
rect 28191 154449 28207 154567
rect 27897 136727 28207 154449
rect 27897 136609 27913 136727
rect 28031 136609 28073 136727
rect 28191 136609 28207 136727
rect 27897 136567 28207 136609
rect 27897 136449 27913 136567
rect 28031 136449 28073 136567
rect 28191 136449 28207 136567
rect 27897 118727 28207 136449
rect 27897 118609 27913 118727
rect 28031 118609 28073 118727
rect 28191 118609 28207 118727
rect 27897 118567 28207 118609
rect 27897 118449 27913 118567
rect 28031 118449 28073 118567
rect 28191 118449 28207 118567
rect 27897 100727 28207 118449
rect 27897 100609 27913 100727
rect 28031 100609 28073 100727
rect 28191 100609 28207 100727
rect 27897 100567 28207 100609
rect 27897 100449 27913 100567
rect 28031 100449 28073 100567
rect 28191 100449 28207 100567
rect 27897 82727 28207 100449
rect 27897 82609 27913 82727
rect 28031 82609 28073 82727
rect 28191 82609 28207 82727
rect 27897 82567 28207 82609
rect 27897 82449 27913 82567
rect 28031 82449 28073 82567
rect 28191 82449 28207 82567
rect 27897 64727 28207 82449
rect 27897 64609 27913 64727
rect 28031 64609 28073 64727
rect 28191 64609 28207 64727
rect 27897 64567 28207 64609
rect 27897 64449 27913 64567
rect 28031 64449 28073 64567
rect 28191 64449 28207 64567
rect 27897 46727 28207 64449
rect 27897 46609 27913 46727
rect 28031 46609 28073 46727
rect 28191 46609 28207 46727
rect 27897 46567 28207 46609
rect 27897 46449 27913 46567
rect 28031 46449 28073 46567
rect 28191 46449 28207 46567
rect 27897 28727 28207 46449
rect 27897 28609 27913 28727
rect 28031 28609 28073 28727
rect 28191 28609 28207 28727
rect 27897 28567 28207 28609
rect 27897 28449 27913 28567
rect 28031 28449 28073 28567
rect 28191 28449 28207 28567
rect 27897 10727 28207 28449
rect 27897 10609 27913 10727
rect 28031 10609 28073 10727
rect 28191 10609 28207 10727
rect 27897 10567 28207 10609
rect 27897 10449 27913 10567
rect 28031 10449 28073 10567
rect 28191 10449 28207 10567
rect 27897 -653 28207 10449
rect 27897 -771 27913 -653
rect 28031 -771 28073 -653
rect 28191 -771 28207 -653
rect 27897 -813 28207 -771
rect 27897 -931 27913 -813
rect 28031 -931 28073 -813
rect 28191 -931 28207 -813
rect 27897 -947 28207 -931
rect 29757 336587 30067 353581
rect 29757 336469 29773 336587
rect 29891 336469 29933 336587
rect 30051 336469 30067 336587
rect 29757 336427 30067 336469
rect 29757 336309 29773 336427
rect 29891 336309 29933 336427
rect 30051 336309 30067 336427
rect 29757 318587 30067 336309
rect 29757 318469 29773 318587
rect 29891 318469 29933 318587
rect 30051 318469 30067 318587
rect 29757 318427 30067 318469
rect 29757 318309 29773 318427
rect 29891 318309 29933 318427
rect 30051 318309 30067 318427
rect 29757 300587 30067 318309
rect 29757 300469 29773 300587
rect 29891 300469 29933 300587
rect 30051 300469 30067 300587
rect 29757 300427 30067 300469
rect 29757 300309 29773 300427
rect 29891 300309 29933 300427
rect 30051 300309 30067 300427
rect 29757 282587 30067 300309
rect 29757 282469 29773 282587
rect 29891 282469 29933 282587
rect 30051 282469 30067 282587
rect 29757 282427 30067 282469
rect 29757 282309 29773 282427
rect 29891 282309 29933 282427
rect 30051 282309 30067 282427
rect 29757 264587 30067 282309
rect 29757 264469 29773 264587
rect 29891 264469 29933 264587
rect 30051 264469 30067 264587
rect 29757 264427 30067 264469
rect 29757 264309 29773 264427
rect 29891 264309 29933 264427
rect 30051 264309 30067 264427
rect 29757 246587 30067 264309
rect 29757 246469 29773 246587
rect 29891 246469 29933 246587
rect 30051 246469 30067 246587
rect 29757 246427 30067 246469
rect 29757 246309 29773 246427
rect 29891 246309 29933 246427
rect 30051 246309 30067 246427
rect 29757 228587 30067 246309
rect 29757 228469 29773 228587
rect 29891 228469 29933 228587
rect 30051 228469 30067 228587
rect 29757 228427 30067 228469
rect 29757 228309 29773 228427
rect 29891 228309 29933 228427
rect 30051 228309 30067 228427
rect 29757 210587 30067 228309
rect 29757 210469 29773 210587
rect 29891 210469 29933 210587
rect 30051 210469 30067 210587
rect 29757 210427 30067 210469
rect 29757 210309 29773 210427
rect 29891 210309 29933 210427
rect 30051 210309 30067 210427
rect 29757 192587 30067 210309
rect 29757 192469 29773 192587
rect 29891 192469 29933 192587
rect 30051 192469 30067 192587
rect 29757 192427 30067 192469
rect 29757 192309 29773 192427
rect 29891 192309 29933 192427
rect 30051 192309 30067 192427
rect 29757 174587 30067 192309
rect 29757 174469 29773 174587
rect 29891 174469 29933 174587
rect 30051 174469 30067 174587
rect 29757 174427 30067 174469
rect 29757 174309 29773 174427
rect 29891 174309 29933 174427
rect 30051 174309 30067 174427
rect 29757 156587 30067 174309
rect 29757 156469 29773 156587
rect 29891 156469 29933 156587
rect 30051 156469 30067 156587
rect 29757 156427 30067 156469
rect 29757 156309 29773 156427
rect 29891 156309 29933 156427
rect 30051 156309 30067 156427
rect 29757 138587 30067 156309
rect 29757 138469 29773 138587
rect 29891 138469 29933 138587
rect 30051 138469 30067 138587
rect 29757 138427 30067 138469
rect 29757 138309 29773 138427
rect 29891 138309 29933 138427
rect 30051 138309 30067 138427
rect 29757 120587 30067 138309
rect 29757 120469 29773 120587
rect 29891 120469 29933 120587
rect 30051 120469 30067 120587
rect 29757 120427 30067 120469
rect 29757 120309 29773 120427
rect 29891 120309 29933 120427
rect 30051 120309 30067 120427
rect 29757 102587 30067 120309
rect 29757 102469 29773 102587
rect 29891 102469 29933 102587
rect 30051 102469 30067 102587
rect 29757 102427 30067 102469
rect 29757 102309 29773 102427
rect 29891 102309 29933 102427
rect 30051 102309 30067 102427
rect 29757 84587 30067 102309
rect 29757 84469 29773 84587
rect 29891 84469 29933 84587
rect 30051 84469 30067 84587
rect 29757 84427 30067 84469
rect 29757 84309 29773 84427
rect 29891 84309 29933 84427
rect 30051 84309 30067 84427
rect 29757 66587 30067 84309
rect 29757 66469 29773 66587
rect 29891 66469 29933 66587
rect 30051 66469 30067 66587
rect 29757 66427 30067 66469
rect 29757 66309 29773 66427
rect 29891 66309 29933 66427
rect 30051 66309 30067 66427
rect 29757 48587 30067 66309
rect 29757 48469 29773 48587
rect 29891 48469 29933 48587
rect 30051 48469 30067 48587
rect 29757 48427 30067 48469
rect 29757 48309 29773 48427
rect 29891 48309 29933 48427
rect 30051 48309 30067 48427
rect 29757 30587 30067 48309
rect 29757 30469 29773 30587
rect 29891 30469 29933 30587
rect 30051 30469 30067 30587
rect 29757 30427 30067 30469
rect 29757 30309 29773 30427
rect 29891 30309 29933 30427
rect 30051 30309 30067 30427
rect 29757 12587 30067 30309
rect 29757 12469 29773 12587
rect 29891 12469 29933 12587
rect 30051 12469 30067 12587
rect 29757 12427 30067 12469
rect 29757 12309 29773 12427
rect 29891 12309 29933 12427
rect 30051 12309 30067 12427
rect 29757 -1613 30067 12309
rect 29757 -1731 29773 -1613
rect 29891 -1731 29933 -1613
rect 30051 -1731 30067 -1613
rect 29757 -1773 30067 -1731
rect 29757 -1891 29773 -1773
rect 29891 -1891 29933 -1773
rect 30051 -1891 30067 -1773
rect 29757 -1907 30067 -1891
rect 31617 338447 31927 354541
rect 31617 338329 31633 338447
rect 31751 338329 31793 338447
rect 31911 338329 31927 338447
rect 31617 338287 31927 338329
rect 31617 338169 31633 338287
rect 31751 338169 31793 338287
rect 31911 338169 31927 338287
rect 31617 320447 31927 338169
rect 31617 320329 31633 320447
rect 31751 320329 31793 320447
rect 31911 320329 31927 320447
rect 31617 320287 31927 320329
rect 31617 320169 31633 320287
rect 31751 320169 31793 320287
rect 31911 320169 31927 320287
rect 31617 302447 31927 320169
rect 31617 302329 31633 302447
rect 31751 302329 31793 302447
rect 31911 302329 31927 302447
rect 31617 302287 31927 302329
rect 31617 302169 31633 302287
rect 31751 302169 31793 302287
rect 31911 302169 31927 302287
rect 31617 284447 31927 302169
rect 31617 284329 31633 284447
rect 31751 284329 31793 284447
rect 31911 284329 31927 284447
rect 31617 284287 31927 284329
rect 31617 284169 31633 284287
rect 31751 284169 31793 284287
rect 31911 284169 31927 284287
rect 31617 266447 31927 284169
rect 31617 266329 31633 266447
rect 31751 266329 31793 266447
rect 31911 266329 31927 266447
rect 31617 266287 31927 266329
rect 31617 266169 31633 266287
rect 31751 266169 31793 266287
rect 31911 266169 31927 266287
rect 31617 248447 31927 266169
rect 31617 248329 31633 248447
rect 31751 248329 31793 248447
rect 31911 248329 31927 248447
rect 31617 248287 31927 248329
rect 31617 248169 31633 248287
rect 31751 248169 31793 248287
rect 31911 248169 31927 248287
rect 31617 230447 31927 248169
rect 31617 230329 31633 230447
rect 31751 230329 31793 230447
rect 31911 230329 31927 230447
rect 31617 230287 31927 230329
rect 31617 230169 31633 230287
rect 31751 230169 31793 230287
rect 31911 230169 31927 230287
rect 31617 212447 31927 230169
rect 31617 212329 31633 212447
rect 31751 212329 31793 212447
rect 31911 212329 31927 212447
rect 31617 212287 31927 212329
rect 31617 212169 31633 212287
rect 31751 212169 31793 212287
rect 31911 212169 31927 212287
rect 31617 194447 31927 212169
rect 31617 194329 31633 194447
rect 31751 194329 31793 194447
rect 31911 194329 31927 194447
rect 31617 194287 31927 194329
rect 31617 194169 31633 194287
rect 31751 194169 31793 194287
rect 31911 194169 31927 194287
rect 31617 176447 31927 194169
rect 31617 176329 31633 176447
rect 31751 176329 31793 176447
rect 31911 176329 31927 176447
rect 31617 176287 31927 176329
rect 31617 176169 31633 176287
rect 31751 176169 31793 176287
rect 31911 176169 31927 176287
rect 31617 158447 31927 176169
rect 31617 158329 31633 158447
rect 31751 158329 31793 158447
rect 31911 158329 31927 158447
rect 31617 158287 31927 158329
rect 31617 158169 31633 158287
rect 31751 158169 31793 158287
rect 31911 158169 31927 158287
rect 31617 140447 31927 158169
rect 31617 140329 31633 140447
rect 31751 140329 31793 140447
rect 31911 140329 31927 140447
rect 31617 140287 31927 140329
rect 31617 140169 31633 140287
rect 31751 140169 31793 140287
rect 31911 140169 31927 140287
rect 31617 122447 31927 140169
rect 31617 122329 31633 122447
rect 31751 122329 31793 122447
rect 31911 122329 31927 122447
rect 31617 122287 31927 122329
rect 31617 122169 31633 122287
rect 31751 122169 31793 122287
rect 31911 122169 31927 122287
rect 31617 104447 31927 122169
rect 31617 104329 31633 104447
rect 31751 104329 31793 104447
rect 31911 104329 31927 104447
rect 31617 104287 31927 104329
rect 31617 104169 31633 104287
rect 31751 104169 31793 104287
rect 31911 104169 31927 104287
rect 31617 86447 31927 104169
rect 31617 86329 31633 86447
rect 31751 86329 31793 86447
rect 31911 86329 31927 86447
rect 31617 86287 31927 86329
rect 31617 86169 31633 86287
rect 31751 86169 31793 86287
rect 31911 86169 31927 86287
rect 31617 68447 31927 86169
rect 31617 68329 31633 68447
rect 31751 68329 31793 68447
rect 31911 68329 31927 68447
rect 31617 68287 31927 68329
rect 31617 68169 31633 68287
rect 31751 68169 31793 68287
rect 31911 68169 31927 68287
rect 31617 50447 31927 68169
rect 31617 50329 31633 50447
rect 31751 50329 31793 50447
rect 31911 50329 31927 50447
rect 31617 50287 31927 50329
rect 31617 50169 31633 50287
rect 31751 50169 31793 50287
rect 31911 50169 31927 50287
rect 31617 32447 31927 50169
rect 31617 32329 31633 32447
rect 31751 32329 31793 32447
rect 31911 32329 31927 32447
rect 31617 32287 31927 32329
rect 31617 32169 31633 32287
rect 31751 32169 31793 32287
rect 31911 32169 31927 32287
rect 31617 14447 31927 32169
rect 31617 14329 31633 14447
rect 31751 14329 31793 14447
rect 31911 14329 31927 14447
rect 31617 14287 31927 14329
rect 31617 14169 31633 14287
rect 31751 14169 31793 14287
rect 31911 14169 31927 14287
rect 31617 -2573 31927 14169
rect 31617 -2691 31633 -2573
rect 31751 -2691 31793 -2573
rect 31911 -2691 31927 -2573
rect 31617 -2733 31927 -2691
rect 31617 -2851 31633 -2733
rect 31751 -2851 31793 -2733
rect 31911 -2851 31927 -2733
rect 31617 -2867 31927 -2851
rect 33477 340307 33787 355501
rect 42477 355299 42787 355795
rect 42477 355181 42493 355299
rect 42611 355181 42653 355299
rect 42771 355181 42787 355299
rect 42477 355139 42787 355181
rect 42477 355021 42493 355139
rect 42611 355021 42653 355139
rect 42771 355021 42787 355139
rect 40617 354339 40927 354835
rect 40617 354221 40633 354339
rect 40751 354221 40793 354339
rect 40911 354221 40927 354339
rect 40617 354179 40927 354221
rect 40617 354061 40633 354179
rect 40751 354061 40793 354179
rect 40911 354061 40927 354179
rect 38757 353379 39067 353875
rect 38757 353261 38773 353379
rect 38891 353261 38933 353379
rect 39051 353261 39067 353379
rect 38757 353219 39067 353261
rect 38757 353101 38773 353219
rect 38891 353101 38933 353219
rect 39051 353101 39067 353219
rect 33477 340189 33493 340307
rect 33611 340189 33653 340307
rect 33771 340189 33787 340307
rect 33477 340147 33787 340189
rect 33477 340029 33493 340147
rect 33611 340029 33653 340147
rect 33771 340029 33787 340147
rect 33477 322307 33787 340029
rect 33477 322189 33493 322307
rect 33611 322189 33653 322307
rect 33771 322189 33787 322307
rect 33477 322147 33787 322189
rect 33477 322029 33493 322147
rect 33611 322029 33653 322147
rect 33771 322029 33787 322147
rect 33477 304307 33787 322029
rect 33477 304189 33493 304307
rect 33611 304189 33653 304307
rect 33771 304189 33787 304307
rect 33477 304147 33787 304189
rect 33477 304029 33493 304147
rect 33611 304029 33653 304147
rect 33771 304029 33787 304147
rect 33477 286307 33787 304029
rect 33477 286189 33493 286307
rect 33611 286189 33653 286307
rect 33771 286189 33787 286307
rect 33477 286147 33787 286189
rect 33477 286029 33493 286147
rect 33611 286029 33653 286147
rect 33771 286029 33787 286147
rect 33477 268307 33787 286029
rect 33477 268189 33493 268307
rect 33611 268189 33653 268307
rect 33771 268189 33787 268307
rect 33477 268147 33787 268189
rect 33477 268029 33493 268147
rect 33611 268029 33653 268147
rect 33771 268029 33787 268147
rect 33477 250307 33787 268029
rect 33477 250189 33493 250307
rect 33611 250189 33653 250307
rect 33771 250189 33787 250307
rect 33477 250147 33787 250189
rect 33477 250029 33493 250147
rect 33611 250029 33653 250147
rect 33771 250029 33787 250147
rect 33477 232307 33787 250029
rect 33477 232189 33493 232307
rect 33611 232189 33653 232307
rect 33771 232189 33787 232307
rect 33477 232147 33787 232189
rect 33477 232029 33493 232147
rect 33611 232029 33653 232147
rect 33771 232029 33787 232147
rect 33477 214307 33787 232029
rect 33477 214189 33493 214307
rect 33611 214189 33653 214307
rect 33771 214189 33787 214307
rect 33477 214147 33787 214189
rect 33477 214029 33493 214147
rect 33611 214029 33653 214147
rect 33771 214029 33787 214147
rect 33477 196307 33787 214029
rect 33477 196189 33493 196307
rect 33611 196189 33653 196307
rect 33771 196189 33787 196307
rect 33477 196147 33787 196189
rect 33477 196029 33493 196147
rect 33611 196029 33653 196147
rect 33771 196029 33787 196147
rect 33477 178307 33787 196029
rect 33477 178189 33493 178307
rect 33611 178189 33653 178307
rect 33771 178189 33787 178307
rect 33477 178147 33787 178189
rect 33477 178029 33493 178147
rect 33611 178029 33653 178147
rect 33771 178029 33787 178147
rect 33477 160307 33787 178029
rect 33477 160189 33493 160307
rect 33611 160189 33653 160307
rect 33771 160189 33787 160307
rect 33477 160147 33787 160189
rect 33477 160029 33493 160147
rect 33611 160029 33653 160147
rect 33771 160029 33787 160147
rect 33477 142307 33787 160029
rect 33477 142189 33493 142307
rect 33611 142189 33653 142307
rect 33771 142189 33787 142307
rect 33477 142147 33787 142189
rect 33477 142029 33493 142147
rect 33611 142029 33653 142147
rect 33771 142029 33787 142147
rect 33477 124307 33787 142029
rect 33477 124189 33493 124307
rect 33611 124189 33653 124307
rect 33771 124189 33787 124307
rect 33477 124147 33787 124189
rect 33477 124029 33493 124147
rect 33611 124029 33653 124147
rect 33771 124029 33787 124147
rect 33477 106307 33787 124029
rect 33477 106189 33493 106307
rect 33611 106189 33653 106307
rect 33771 106189 33787 106307
rect 33477 106147 33787 106189
rect 33477 106029 33493 106147
rect 33611 106029 33653 106147
rect 33771 106029 33787 106147
rect 33477 88307 33787 106029
rect 33477 88189 33493 88307
rect 33611 88189 33653 88307
rect 33771 88189 33787 88307
rect 33477 88147 33787 88189
rect 33477 88029 33493 88147
rect 33611 88029 33653 88147
rect 33771 88029 33787 88147
rect 33477 70307 33787 88029
rect 33477 70189 33493 70307
rect 33611 70189 33653 70307
rect 33771 70189 33787 70307
rect 33477 70147 33787 70189
rect 33477 70029 33493 70147
rect 33611 70029 33653 70147
rect 33771 70029 33787 70147
rect 33477 52307 33787 70029
rect 33477 52189 33493 52307
rect 33611 52189 33653 52307
rect 33771 52189 33787 52307
rect 33477 52147 33787 52189
rect 33477 52029 33493 52147
rect 33611 52029 33653 52147
rect 33771 52029 33787 52147
rect 33477 34307 33787 52029
rect 33477 34189 33493 34307
rect 33611 34189 33653 34307
rect 33771 34189 33787 34307
rect 33477 34147 33787 34189
rect 33477 34029 33493 34147
rect 33611 34029 33653 34147
rect 33771 34029 33787 34147
rect 33477 16307 33787 34029
rect 33477 16189 33493 16307
rect 33611 16189 33653 16307
rect 33771 16189 33787 16307
rect 33477 16147 33787 16189
rect 33477 16029 33493 16147
rect 33611 16029 33653 16147
rect 33771 16029 33787 16147
rect 24477 -3171 24493 -3053
rect 24611 -3171 24653 -3053
rect 24771 -3171 24787 -3053
rect 24477 -3213 24787 -3171
rect 24477 -3331 24493 -3213
rect 24611 -3331 24653 -3213
rect 24771 -3331 24787 -3213
rect 24477 -3827 24787 -3331
rect 33477 -3533 33787 16029
rect 36897 352419 37207 352915
rect 36897 352301 36913 352419
rect 37031 352301 37073 352419
rect 37191 352301 37207 352419
rect 36897 352259 37207 352301
rect 36897 352141 36913 352259
rect 37031 352141 37073 352259
rect 37191 352141 37207 352259
rect 36897 343727 37207 352141
rect 36897 343609 36913 343727
rect 37031 343609 37073 343727
rect 37191 343609 37207 343727
rect 36897 343567 37207 343609
rect 36897 343449 36913 343567
rect 37031 343449 37073 343567
rect 37191 343449 37207 343567
rect 36897 325727 37207 343449
rect 36897 325609 36913 325727
rect 37031 325609 37073 325727
rect 37191 325609 37207 325727
rect 36897 325567 37207 325609
rect 36897 325449 36913 325567
rect 37031 325449 37073 325567
rect 37191 325449 37207 325567
rect 36897 307727 37207 325449
rect 36897 307609 36913 307727
rect 37031 307609 37073 307727
rect 37191 307609 37207 307727
rect 36897 307567 37207 307609
rect 36897 307449 36913 307567
rect 37031 307449 37073 307567
rect 37191 307449 37207 307567
rect 36897 289727 37207 307449
rect 36897 289609 36913 289727
rect 37031 289609 37073 289727
rect 37191 289609 37207 289727
rect 36897 289567 37207 289609
rect 36897 289449 36913 289567
rect 37031 289449 37073 289567
rect 37191 289449 37207 289567
rect 36897 271727 37207 289449
rect 36897 271609 36913 271727
rect 37031 271609 37073 271727
rect 37191 271609 37207 271727
rect 36897 271567 37207 271609
rect 36897 271449 36913 271567
rect 37031 271449 37073 271567
rect 37191 271449 37207 271567
rect 36897 253727 37207 271449
rect 36897 253609 36913 253727
rect 37031 253609 37073 253727
rect 37191 253609 37207 253727
rect 36897 253567 37207 253609
rect 36897 253449 36913 253567
rect 37031 253449 37073 253567
rect 37191 253449 37207 253567
rect 36897 235727 37207 253449
rect 36897 235609 36913 235727
rect 37031 235609 37073 235727
rect 37191 235609 37207 235727
rect 36897 235567 37207 235609
rect 36897 235449 36913 235567
rect 37031 235449 37073 235567
rect 37191 235449 37207 235567
rect 36897 217727 37207 235449
rect 36897 217609 36913 217727
rect 37031 217609 37073 217727
rect 37191 217609 37207 217727
rect 36897 217567 37207 217609
rect 36897 217449 36913 217567
rect 37031 217449 37073 217567
rect 37191 217449 37207 217567
rect 36897 199727 37207 217449
rect 36897 199609 36913 199727
rect 37031 199609 37073 199727
rect 37191 199609 37207 199727
rect 36897 199567 37207 199609
rect 36897 199449 36913 199567
rect 37031 199449 37073 199567
rect 37191 199449 37207 199567
rect 36897 181727 37207 199449
rect 36897 181609 36913 181727
rect 37031 181609 37073 181727
rect 37191 181609 37207 181727
rect 36897 181567 37207 181609
rect 36897 181449 36913 181567
rect 37031 181449 37073 181567
rect 37191 181449 37207 181567
rect 36897 163727 37207 181449
rect 36897 163609 36913 163727
rect 37031 163609 37073 163727
rect 37191 163609 37207 163727
rect 36897 163567 37207 163609
rect 36897 163449 36913 163567
rect 37031 163449 37073 163567
rect 37191 163449 37207 163567
rect 36897 145727 37207 163449
rect 36897 145609 36913 145727
rect 37031 145609 37073 145727
rect 37191 145609 37207 145727
rect 36897 145567 37207 145609
rect 36897 145449 36913 145567
rect 37031 145449 37073 145567
rect 37191 145449 37207 145567
rect 36897 127727 37207 145449
rect 36897 127609 36913 127727
rect 37031 127609 37073 127727
rect 37191 127609 37207 127727
rect 36897 127567 37207 127609
rect 36897 127449 36913 127567
rect 37031 127449 37073 127567
rect 37191 127449 37207 127567
rect 36897 109727 37207 127449
rect 36897 109609 36913 109727
rect 37031 109609 37073 109727
rect 37191 109609 37207 109727
rect 36897 109567 37207 109609
rect 36897 109449 36913 109567
rect 37031 109449 37073 109567
rect 37191 109449 37207 109567
rect 36897 91727 37207 109449
rect 36897 91609 36913 91727
rect 37031 91609 37073 91727
rect 37191 91609 37207 91727
rect 36897 91567 37207 91609
rect 36897 91449 36913 91567
rect 37031 91449 37073 91567
rect 37191 91449 37207 91567
rect 36897 73727 37207 91449
rect 36897 73609 36913 73727
rect 37031 73609 37073 73727
rect 37191 73609 37207 73727
rect 36897 73567 37207 73609
rect 36897 73449 36913 73567
rect 37031 73449 37073 73567
rect 37191 73449 37207 73567
rect 36897 55727 37207 73449
rect 36897 55609 36913 55727
rect 37031 55609 37073 55727
rect 37191 55609 37207 55727
rect 36897 55567 37207 55609
rect 36897 55449 36913 55567
rect 37031 55449 37073 55567
rect 37191 55449 37207 55567
rect 36897 37727 37207 55449
rect 36897 37609 36913 37727
rect 37031 37609 37073 37727
rect 37191 37609 37207 37727
rect 36897 37567 37207 37609
rect 36897 37449 36913 37567
rect 37031 37449 37073 37567
rect 37191 37449 37207 37567
rect 36897 19727 37207 37449
rect 36897 19609 36913 19727
rect 37031 19609 37073 19727
rect 37191 19609 37207 19727
rect 36897 19567 37207 19609
rect 36897 19449 36913 19567
rect 37031 19449 37073 19567
rect 37191 19449 37207 19567
rect 36897 1727 37207 19449
rect 36897 1609 36913 1727
rect 37031 1609 37073 1727
rect 37191 1609 37207 1727
rect 36897 1567 37207 1609
rect 36897 1449 36913 1567
rect 37031 1449 37073 1567
rect 37191 1449 37207 1567
rect 36897 -173 37207 1449
rect 36897 -291 36913 -173
rect 37031 -291 37073 -173
rect 37191 -291 37207 -173
rect 36897 -333 37207 -291
rect 36897 -451 36913 -333
rect 37031 -451 37073 -333
rect 37191 -451 37207 -333
rect 36897 -947 37207 -451
rect 38757 345587 39067 353101
rect 38757 345469 38773 345587
rect 38891 345469 38933 345587
rect 39051 345469 39067 345587
rect 38757 345427 39067 345469
rect 38757 345309 38773 345427
rect 38891 345309 38933 345427
rect 39051 345309 39067 345427
rect 38757 327587 39067 345309
rect 38757 327469 38773 327587
rect 38891 327469 38933 327587
rect 39051 327469 39067 327587
rect 38757 327427 39067 327469
rect 38757 327309 38773 327427
rect 38891 327309 38933 327427
rect 39051 327309 39067 327427
rect 38757 309587 39067 327309
rect 38757 309469 38773 309587
rect 38891 309469 38933 309587
rect 39051 309469 39067 309587
rect 38757 309427 39067 309469
rect 38757 309309 38773 309427
rect 38891 309309 38933 309427
rect 39051 309309 39067 309427
rect 38757 291587 39067 309309
rect 38757 291469 38773 291587
rect 38891 291469 38933 291587
rect 39051 291469 39067 291587
rect 38757 291427 39067 291469
rect 38757 291309 38773 291427
rect 38891 291309 38933 291427
rect 39051 291309 39067 291427
rect 38757 273587 39067 291309
rect 38757 273469 38773 273587
rect 38891 273469 38933 273587
rect 39051 273469 39067 273587
rect 38757 273427 39067 273469
rect 38757 273309 38773 273427
rect 38891 273309 38933 273427
rect 39051 273309 39067 273427
rect 38757 255587 39067 273309
rect 38757 255469 38773 255587
rect 38891 255469 38933 255587
rect 39051 255469 39067 255587
rect 38757 255427 39067 255469
rect 38757 255309 38773 255427
rect 38891 255309 38933 255427
rect 39051 255309 39067 255427
rect 38757 237587 39067 255309
rect 38757 237469 38773 237587
rect 38891 237469 38933 237587
rect 39051 237469 39067 237587
rect 38757 237427 39067 237469
rect 38757 237309 38773 237427
rect 38891 237309 38933 237427
rect 39051 237309 39067 237427
rect 38757 219587 39067 237309
rect 38757 219469 38773 219587
rect 38891 219469 38933 219587
rect 39051 219469 39067 219587
rect 38757 219427 39067 219469
rect 38757 219309 38773 219427
rect 38891 219309 38933 219427
rect 39051 219309 39067 219427
rect 38757 201587 39067 219309
rect 38757 201469 38773 201587
rect 38891 201469 38933 201587
rect 39051 201469 39067 201587
rect 38757 201427 39067 201469
rect 38757 201309 38773 201427
rect 38891 201309 38933 201427
rect 39051 201309 39067 201427
rect 38757 183587 39067 201309
rect 38757 183469 38773 183587
rect 38891 183469 38933 183587
rect 39051 183469 39067 183587
rect 38757 183427 39067 183469
rect 38757 183309 38773 183427
rect 38891 183309 38933 183427
rect 39051 183309 39067 183427
rect 38757 165587 39067 183309
rect 38757 165469 38773 165587
rect 38891 165469 38933 165587
rect 39051 165469 39067 165587
rect 38757 165427 39067 165469
rect 38757 165309 38773 165427
rect 38891 165309 38933 165427
rect 39051 165309 39067 165427
rect 38757 147587 39067 165309
rect 38757 147469 38773 147587
rect 38891 147469 38933 147587
rect 39051 147469 39067 147587
rect 38757 147427 39067 147469
rect 38757 147309 38773 147427
rect 38891 147309 38933 147427
rect 39051 147309 39067 147427
rect 38757 129587 39067 147309
rect 38757 129469 38773 129587
rect 38891 129469 38933 129587
rect 39051 129469 39067 129587
rect 38757 129427 39067 129469
rect 38757 129309 38773 129427
rect 38891 129309 38933 129427
rect 39051 129309 39067 129427
rect 38757 111587 39067 129309
rect 38757 111469 38773 111587
rect 38891 111469 38933 111587
rect 39051 111469 39067 111587
rect 38757 111427 39067 111469
rect 38757 111309 38773 111427
rect 38891 111309 38933 111427
rect 39051 111309 39067 111427
rect 38757 93587 39067 111309
rect 38757 93469 38773 93587
rect 38891 93469 38933 93587
rect 39051 93469 39067 93587
rect 38757 93427 39067 93469
rect 38757 93309 38773 93427
rect 38891 93309 38933 93427
rect 39051 93309 39067 93427
rect 38757 75587 39067 93309
rect 38757 75469 38773 75587
rect 38891 75469 38933 75587
rect 39051 75469 39067 75587
rect 38757 75427 39067 75469
rect 38757 75309 38773 75427
rect 38891 75309 38933 75427
rect 39051 75309 39067 75427
rect 38757 57587 39067 75309
rect 38757 57469 38773 57587
rect 38891 57469 38933 57587
rect 39051 57469 39067 57587
rect 38757 57427 39067 57469
rect 38757 57309 38773 57427
rect 38891 57309 38933 57427
rect 39051 57309 39067 57427
rect 38757 39587 39067 57309
rect 38757 39469 38773 39587
rect 38891 39469 38933 39587
rect 39051 39469 39067 39587
rect 38757 39427 39067 39469
rect 38757 39309 38773 39427
rect 38891 39309 38933 39427
rect 39051 39309 39067 39427
rect 38757 21587 39067 39309
rect 38757 21469 38773 21587
rect 38891 21469 38933 21587
rect 39051 21469 39067 21587
rect 38757 21427 39067 21469
rect 38757 21309 38773 21427
rect 38891 21309 38933 21427
rect 39051 21309 39067 21427
rect 38757 3587 39067 21309
rect 38757 3469 38773 3587
rect 38891 3469 38933 3587
rect 39051 3469 39067 3587
rect 38757 3427 39067 3469
rect 38757 3309 38773 3427
rect 38891 3309 38933 3427
rect 39051 3309 39067 3427
rect 38757 -1133 39067 3309
rect 38757 -1251 38773 -1133
rect 38891 -1251 38933 -1133
rect 39051 -1251 39067 -1133
rect 38757 -1293 39067 -1251
rect 38757 -1411 38773 -1293
rect 38891 -1411 38933 -1293
rect 39051 -1411 39067 -1293
rect 38757 -1907 39067 -1411
rect 40617 347447 40927 354061
rect 40617 347329 40633 347447
rect 40751 347329 40793 347447
rect 40911 347329 40927 347447
rect 40617 347287 40927 347329
rect 40617 347169 40633 347287
rect 40751 347169 40793 347287
rect 40911 347169 40927 347287
rect 40617 329447 40927 347169
rect 40617 329329 40633 329447
rect 40751 329329 40793 329447
rect 40911 329329 40927 329447
rect 40617 329287 40927 329329
rect 40617 329169 40633 329287
rect 40751 329169 40793 329287
rect 40911 329169 40927 329287
rect 40617 311447 40927 329169
rect 40617 311329 40633 311447
rect 40751 311329 40793 311447
rect 40911 311329 40927 311447
rect 40617 311287 40927 311329
rect 40617 311169 40633 311287
rect 40751 311169 40793 311287
rect 40911 311169 40927 311287
rect 40617 293447 40927 311169
rect 40617 293329 40633 293447
rect 40751 293329 40793 293447
rect 40911 293329 40927 293447
rect 40617 293287 40927 293329
rect 40617 293169 40633 293287
rect 40751 293169 40793 293287
rect 40911 293169 40927 293287
rect 40617 275447 40927 293169
rect 40617 275329 40633 275447
rect 40751 275329 40793 275447
rect 40911 275329 40927 275447
rect 40617 275287 40927 275329
rect 40617 275169 40633 275287
rect 40751 275169 40793 275287
rect 40911 275169 40927 275287
rect 40617 257447 40927 275169
rect 40617 257329 40633 257447
rect 40751 257329 40793 257447
rect 40911 257329 40927 257447
rect 40617 257287 40927 257329
rect 40617 257169 40633 257287
rect 40751 257169 40793 257287
rect 40911 257169 40927 257287
rect 40617 239447 40927 257169
rect 40617 239329 40633 239447
rect 40751 239329 40793 239447
rect 40911 239329 40927 239447
rect 40617 239287 40927 239329
rect 40617 239169 40633 239287
rect 40751 239169 40793 239287
rect 40911 239169 40927 239287
rect 40617 221447 40927 239169
rect 40617 221329 40633 221447
rect 40751 221329 40793 221447
rect 40911 221329 40927 221447
rect 40617 221287 40927 221329
rect 40617 221169 40633 221287
rect 40751 221169 40793 221287
rect 40911 221169 40927 221287
rect 40617 203447 40927 221169
rect 40617 203329 40633 203447
rect 40751 203329 40793 203447
rect 40911 203329 40927 203447
rect 40617 203287 40927 203329
rect 40617 203169 40633 203287
rect 40751 203169 40793 203287
rect 40911 203169 40927 203287
rect 40617 185447 40927 203169
rect 40617 185329 40633 185447
rect 40751 185329 40793 185447
rect 40911 185329 40927 185447
rect 40617 185287 40927 185329
rect 40617 185169 40633 185287
rect 40751 185169 40793 185287
rect 40911 185169 40927 185287
rect 40617 167447 40927 185169
rect 40617 167329 40633 167447
rect 40751 167329 40793 167447
rect 40911 167329 40927 167447
rect 40617 167287 40927 167329
rect 40617 167169 40633 167287
rect 40751 167169 40793 167287
rect 40911 167169 40927 167287
rect 40617 149447 40927 167169
rect 40617 149329 40633 149447
rect 40751 149329 40793 149447
rect 40911 149329 40927 149447
rect 40617 149287 40927 149329
rect 40617 149169 40633 149287
rect 40751 149169 40793 149287
rect 40911 149169 40927 149287
rect 40617 131447 40927 149169
rect 40617 131329 40633 131447
rect 40751 131329 40793 131447
rect 40911 131329 40927 131447
rect 40617 131287 40927 131329
rect 40617 131169 40633 131287
rect 40751 131169 40793 131287
rect 40911 131169 40927 131287
rect 40617 113447 40927 131169
rect 40617 113329 40633 113447
rect 40751 113329 40793 113447
rect 40911 113329 40927 113447
rect 40617 113287 40927 113329
rect 40617 113169 40633 113287
rect 40751 113169 40793 113287
rect 40911 113169 40927 113287
rect 40617 95447 40927 113169
rect 40617 95329 40633 95447
rect 40751 95329 40793 95447
rect 40911 95329 40927 95447
rect 40617 95287 40927 95329
rect 40617 95169 40633 95287
rect 40751 95169 40793 95287
rect 40911 95169 40927 95287
rect 40617 77447 40927 95169
rect 40617 77329 40633 77447
rect 40751 77329 40793 77447
rect 40911 77329 40927 77447
rect 40617 77287 40927 77329
rect 40617 77169 40633 77287
rect 40751 77169 40793 77287
rect 40911 77169 40927 77287
rect 40617 59447 40927 77169
rect 40617 59329 40633 59447
rect 40751 59329 40793 59447
rect 40911 59329 40927 59447
rect 40617 59287 40927 59329
rect 40617 59169 40633 59287
rect 40751 59169 40793 59287
rect 40911 59169 40927 59287
rect 40617 41447 40927 59169
rect 40617 41329 40633 41447
rect 40751 41329 40793 41447
rect 40911 41329 40927 41447
rect 40617 41287 40927 41329
rect 40617 41169 40633 41287
rect 40751 41169 40793 41287
rect 40911 41169 40927 41287
rect 40617 23447 40927 41169
rect 40617 23329 40633 23447
rect 40751 23329 40793 23447
rect 40911 23329 40927 23447
rect 40617 23287 40927 23329
rect 40617 23169 40633 23287
rect 40751 23169 40793 23287
rect 40911 23169 40927 23287
rect 40617 5447 40927 23169
rect 40617 5329 40633 5447
rect 40751 5329 40793 5447
rect 40911 5329 40927 5447
rect 40617 5287 40927 5329
rect 40617 5169 40633 5287
rect 40751 5169 40793 5287
rect 40911 5169 40927 5287
rect 40617 -2093 40927 5169
rect 40617 -2211 40633 -2093
rect 40751 -2211 40793 -2093
rect 40911 -2211 40927 -2093
rect 40617 -2253 40927 -2211
rect 40617 -2371 40633 -2253
rect 40751 -2371 40793 -2253
rect 40911 -2371 40927 -2253
rect 40617 -2867 40927 -2371
rect 42477 349307 42787 355021
rect 51477 355779 51787 355795
rect 51477 355661 51493 355779
rect 51611 355661 51653 355779
rect 51771 355661 51787 355779
rect 51477 355619 51787 355661
rect 51477 355501 51493 355619
rect 51611 355501 51653 355619
rect 51771 355501 51787 355619
rect 49617 354819 49927 354835
rect 49617 354701 49633 354819
rect 49751 354701 49793 354819
rect 49911 354701 49927 354819
rect 49617 354659 49927 354701
rect 49617 354541 49633 354659
rect 49751 354541 49793 354659
rect 49911 354541 49927 354659
rect 47757 353859 48067 353875
rect 47757 353741 47773 353859
rect 47891 353741 47933 353859
rect 48051 353741 48067 353859
rect 47757 353699 48067 353741
rect 47757 353581 47773 353699
rect 47891 353581 47933 353699
rect 48051 353581 48067 353699
rect 42477 349189 42493 349307
rect 42611 349189 42653 349307
rect 42771 349189 42787 349307
rect 42477 349147 42787 349189
rect 42477 349029 42493 349147
rect 42611 349029 42653 349147
rect 42771 349029 42787 349147
rect 42477 331307 42787 349029
rect 42477 331189 42493 331307
rect 42611 331189 42653 331307
rect 42771 331189 42787 331307
rect 42477 331147 42787 331189
rect 42477 331029 42493 331147
rect 42611 331029 42653 331147
rect 42771 331029 42787 331147
rect 42477 313307 42787 331029
rect 42477 313189 42493 313307
rect 42611 313189 42653 313307
rect 42771 313189 42787 313307
rect 42477 313147 42787 313189
rect 42477 313029 42493 313147
rect 42611 313029 42653 313147
rect 42771 313029 42787 313147
rect 42477 295307 42787 313029
rect 42477 295189 42493 295307
rect 42611 295189 42653 295307
rect 42771 295189 42787 295307
rect 42477 295147 42787 295189
rect 42477 295029 42493 295147
rect 42611 295029 42653 295147
rect 42771 295029 42787 295147
rect 42477 277307 42787 295029
rect 42477 277189 42493 277307
rect 42611 277189 42653 277307
rect 42771 277189 42787 277307
rect 42477 277147 42787 277189
rect 42477 277029 42493 277147
rect 42611 277029 42653 277147
rect 42771 277029 42787 277147
rect 42477 259307 42787 277029
rect 42477 259189 42493 259307
rect 42611 259189 42653 259307
rect 42771 259189 42787 259307
rect 42477 259147 42787 259189
rect 42477 259029 42493 259147
rect 42611 259029 42653 259147
rect 42771 259029 42787 259147
rect 42477 241307 42787 259029
rect 42477 241189 42493 241307
rect 42611 241189 42653 241307
rect 42771 241189 42787 241307
rect 42477 241147 42787 241189
rect 42477 241029 42493 241147
rect 42611 241029 42653 241147
rect 42771 241029 42787 241147
rect 42477 223307 42787 241029
rect 42477 223189 42493 223307
rect 42611 223189 42653 223307
rect 42771 223189 42787 223307
rect 42477 223147 42787 223189
rect 42477 223029 42493 223147
rect 42611 223029 42653 223147
rect 42771 223029 42787 223147
rect 42477 205307 42787 223029
rect 42477 205189 42493 205307
rect 42611 205189 42653 205307
rect 42771 205189 42787 205307
rect 42477 205147 42787 205189
rect 42477 205029 42493 205147
rect 42611 205029 42653 205147
rect 42771 205029 42787 205147
rect 42477 187307 42787 205029
rect 42477 187189 42493 187307
rect 42611 187189 42653 187307
rect 42771 187189 42787 187307
rect 42477 187147 42787 187189
rect 42477 187029 42493 187147
rect 42611 187029 42653 187147
rect 42771 187029 42787 187147
rect 42477 169307 42787 187029
rect 42477 169189 42493 169307
rect 42611 169189 42653 169307
rect 42771 169189 42787 169307
rect 42477 169147 42787 169189
rect 42477 169029 42493 169147
rect 42611 169029 42653 169147
rect 42771 169029 42787 169147
rect 42477 151307 42787 169029
rect 42477 151189 42493 151307
rect 42611 151189 42653 151307
rect 42771 151189 42787 151307
rect 42477 151147 42787 151189
rect 42477 151029 42493 151147
rect 42611 151029 42653 151147
rect 42771 151029 42787 151147
rect 42477 133307 42787 151029
rect 42477 133189 42493 133307
rect 42611 133189 42653 133307
rect 42771 133189 42787 133307
rect 42477 133147 42787 133189
rect 42477 133029 42493 133147
rect 42611 133029 42653 133147
rect 42771 133029 42787 133147
rect 42477 115307 42787 133029
rect 42477 115189 42493 115307
rect 42611 115189 42653 115307
rect 42771 115189 42787 115307
rect 42477 115147 42787 115189
rect 42477 115029 42493 115147
rect 42611 115029 42653 115147
rect 42771 115029 42787 115147
rect 42477 97307 42787 115029
rect 42477 97189 42493 97307
rect 42611 97189 42653 97307
rect 42771 97189 42787 97307
rect 42477 97147 42787 97189
rect 42477 97029 42493 97147
rect 42611 97029 42653 97147
rect 42771 97029 42787 97147
rect 42477 79307 42787 97029
rect 42477 79189 42493 79307
rect 42611 79189 42653 79307
rect 42771 79189 42787 79307
rect 42477 79147 42787 79189
rect 42477 79029 42493 79147
rect 42611 79029 42653 79147
rect 42771 79029 42787 79147
rect 42477 61307 42787 79029
rect 42477 61189 42493 61307
rect 42611 61189 42653 61307
rect 42771 61189 42787 61307
rect 42477 61147 42787 61189
rect 42477 61029 42493 61147
rect 42611 61029 42653 61147
rect 42771 61029 42787 61147
rect 42477 43307 42787 61029
rect 42477 43189 42493 43307
rect 42611 43189 42653 43307
rect 42771 43189 42787 43307
rect 42477 43147 42787 43189
rect 42477 43029 42493 43147
rect 42611 43029 42653 43147
rect 42771 43029 42787 43147
rect 42477 25307 42787 43029
rect 42477 25189 42493 25307
rect 42611 25189 42653 25307
rect 42771 25189 42787 25307
rect 42477 25147 42787 25189
rect 42477 25029 42493 25147
rect 42611 25029 42653 25147
rect 42771 25029 42787 25147
rect 42477 7307 42787 25029
rect 42477 7189 42493 7307
rect 42611 7189 42653 7307
rect 42771 7189 42787 7307
rect 42477 7147 42787 7189
rect 42477 7029 42493 7147
rect 42611 7029 42653 7147
rect 42771 7029 42787 7147
rect 33477 -3651 33493 -3533
rect 33611 -3651 33653 -3533
rect 33771 -3651 33787 -3533
rect 33477 -3693 33787 -3651
rect 33477 -3811 33493 -3693
rect 33611 -3811 33653 -3693
rect 33771 -3811 33787 -3693
rect 33477 -3827 33787 -3811
rect 42477 -3053 42787 7029
rect 45897 352899 46207 352915
rect 45897 352781 45913 352899
rect 46031 352781 46073 352899
rect 46191 352781 46207 352899
rect 45897 352739 46207 352781
rect 45897 352621 45913 352739
rect 46031 352621 46073 352739
rect 46191 352621 46207 352739
rect 45897 334727 46207 352621
rect 45897 334609 45913 334727
rect 46031 334609 46073 334727
rect 46191 334609 46207 334727
rect 45897 334567 46207 334609
rect 45897 334449 45913 334567
rect 46031 334449 46073 334567
rect 46191 334449 46207 334567
rect 45897 316727 46207 334449
rect 45897 316609 45913 316727
rect 46031 316609 46073 316727
rect 46191 316609 46207 316727
rect 45897 316567 46207 316609
rect 45897 316449 45913 316567
rect 46031 316449 46073 316567
rect 46191 316449 46207 316567
rect 45897 298727 46207 316449
rect 45897 298609 45913 298727
rect 46031 298609 46073 298727
rect 46191 298609 46207 298727
rect 45897 298567 46207 298609
rect 45897 298449 45913 298567
rect 46031 298449 46073 298567
rect 46191 298449 46207 298567
rect 45897 280727 46207 298449
rect 45897 280609 45913 280727
rect 46031 280609 46073 280727
rect 46191 280609 46207 280727
rect 45897 280567 46207 280609
rect 45897 280449 45913 280567
rect 46031 280449 46073 280567
rect 46191 280449 46207 280567
rect 45897 262727 46207 280449
rect 45897 262609 45913 262727
rect 46031 262609 46073 262727
rect 46191 262609 46207 262727
rect 45897 262567 46207 262609
rect 45897 262449 45913 262567
rect 46031 262449 46073 262567
rect 46191 262449 46207 262567
rect 45897 244727 46207 262449
rect 45897 244609 45913 244727
rect 46031 244609 46073 244727
rect 46191 244609 46207 244727
rect 45897 244567 46207 244609
rect 45897 244449 45913 244567
rect 46031 244449 46073 244567
rect 46191 244449 46207 244567
rect 45897 226727 46207 244449
rect 45897 226609 45913 226727
rect 46031 226609 46073 226727
rect 46191 226609 46207 226727
rect 45897 226567 46207 226609
rect 45897 226449 45913 226567
rect 46031 226449 46073 226567
rect 46191 226449 46207 226567
rect 45897 208727 46207 226449
rect 45897 208609 45913 208727
rect 46031 208609 46073 208727
rect 46191 208609 46207 208727
rect 45897 208567 46207 208609
rect 45897 208449 45913 208567
rect 46031 208449 46073 208567
rect 46191 208449 46207 208567
rect 45897 190727 46207 208449
rect 45897 190609 45913 190727
rect 46031 190609 46073 190727
rect 46191 190609 46207 190727
rect 45897 190567 46207 190609
rect 45897 190449 45913 190567
rect 46031 190449 46073 190567
rect 46191 190449 46207 190567
rect 45897 172727 46207 190449
rect 45897 172609 45913 172727
rect 46031 172609 46073 172727
rect 46191 172609 46207 172727
rect 45897 172567 46207 172609
rect 45897 172449 45913 172567
rect 46031 172449 46073 172567
rect 46191 172449 46207 172567
rect 45897 154727 46207 172449
rect 45897 154609 45913 154727
rect 46031 154609 46073 154727
rect 46191 154609 46207 154727
rect 45897 154567 46207 154609
rect 45897 154449 45913 154567
rect 46031 154449 46073 154567
rect 46191 154449 46207 154567
rect 45897 136727 46207 154449
rect 45897 136609 45913 136727
rect 46031 136609 46073 136727
rect 46191 136609 46207 136727
rect 45897 136567 46207 136609
rect 45897 136449 45913 136567
rect 46031 136449 46073 136567
rect 46191 136449 46207 136567
rect 45897 118727 46207 136449
rect 45897 118609 45913 118727
rect 46031 118609 46073 118727
rect 46191 118609 46207 118727
rect 45897 118567 46207 118609
rect 45897 118449 45913 118567
rect 46031 118449 46073 118567
rect 46191 118449 46207 118567
rect 45897 100727 46207 118449
rect 45897 100609 45913 100727
rect 46031 100609 46073 100727
rect 46191 100609 46207 100727
rect 45897 100567 46207 100609
rect 45897 100449 45913 100567
rect 46031 100449 46073 100567
rect 46191 100449 46207 100567
rect 45897 82727 46207 100449
rect 45897 82609 45913 82727
rect 46031 82609 46073 82727
rect 46191 82609 46207 82727
rect 45897 82567 46207 82609
rect 45897 82449 45913 82567
rect 46031 82449 46073 82567
rect 46191 82449 46207 82567
rect 45897 64727 46207 82449
rect 45897 64609 45913 64727
rect 46031 64609 46073 64727
rect 46191 64609 46207 64727
rect 45897 64567 46207 64609
rect 45897 64449 45913 64567
rect 46031 64449 46073 64567
rect 46191 64449 46207 64567
rect 45897 46727 46207 64449
rect 45897 46609 45913 46727
rect 46031 46609 46073 46727
rect 46191 46609 46207 46727
rect 45897 46567 46207 46609
rect 45897 46449 45913 46567
rect 46031 46449 46073 46567
rect 46191 46449 46207 46567
rect 45897 28727 46207 46449
rect 45897 28609 45913 28727
rect 46031 28609 46073 28727
rect 46191 28609 46207 28727
rect 45897 28567 46207 28609
rect 45897 28449 45913 28567
rect 46031 28449 46073 28567
rect 46191 28449 46207 28567
rect 45897 10727 46207 28449
rect 45897 10609 45913 10727
rect 46031 10609 46073 10727
rect 46191 10609 46207 10727
rect 45897 10567 46207 10609
rect 45897 10449 45913 10567
rect 46031 10449 46073 10567
rect 46191 10449 46207 10567
rect 45897 -653 46207 10449
rect 45897 -771 45913 -653
rect 46031 -771 46073 -653
rect 46191 -771 46207 -653
rect 45897 -813 46207 -771
rect 45897 -931 45913 -813
rect 46031 -931 46073 -813
rect 46191 -931 46207 -813
rect 45897 -947 46207 -931
rect 47757 336587 48067 353581
rect 47757 336469 47773 336587
rect 47891 336469 47933 336587
rect 48051 336469 48067 336587
rect 47757 336427 48067 336469
rect 47757 336309 47773 336427
rect 47891 336309 47933 336427
rect 48051 336309 48067 336427
rect 47757 318587 48067 336309
rect 47757 318469 47773 318587
rect 47891 318469 47933 318587
rect 48051 318469 48067 318587
rect 47757 318427 48067 318469
rect 47757 318309 47773 318427
rect 47891 318309 47933 318427
rect 48051 318309 48067 318427
rect 47757 300587 48067 318309
rect 47757 300469 47773 300587
rect 47891 300469 47933 300587
rect 48051 300469 48067 300587
rect 47757 300427 48067 300469
rect 47757 300309 47773 300427
rect 47891 300309 47933 300427
rect 48051 300309 48067 300427
rect 47757 282587 48067 300309
rect 47757 282469 47773 282587
rect 47891 282469 47933 282587
rect 48051 282469 48067 282587
rect 47757 282427 48067 282469
rect 47757 282309 47773 282427
rect 47891 282309 47933 282427
rect 48051 282309 48067 282427
rect 47757 264587 48067 282309
rect 47757 264469 47773 264587
rect 47891 264469 47933 264587
rect 48051 264469 48067 264587
rect 47757 264427 48067 264469
rect 47757 264309 47773 264427
rect 47891 264309 47933 264427
rect 48051 264309 48067 264427
rect 47757 246587 48067 264309
rect 47757 246469 47773 246587
rect 47891 246469 47933 246587
rect 48051 246469 48067 246587
rect 47757 246427 48067 246469
rect 47757 246309 47773 246427
rect 47891 246309 47933 246427
rect 48051 246309 48067 246427
rect 47757 228587 48067 246309
rect 47757 228469 47773 228587
rect 47891 228469 47933 228587
rect 48051 228469 48067 228587
rect 47757 228427 48067 228469
rect 47757 228309 47773 228427
rect 47891 228309 47933 228427
rect 48051 228309 48067 228427
rect 47757 210587 48067 228309
rect 47757 210469 47773 210587
rect 47891 210469 47933 210587
rect 48051 210469 48067 210587
rect 47757 210427 48067 210469
rect 47757 210309 47773 210427
rect 47891 210309 47933 210427
rect 48051 210309 48067 210427
rect 47757 192587 48067 210309
rect 47757 192469 47773 192587
rect 47891 192469 47933 192587
rect 48051 192469 48067 192587
rect 47757 192427 48067 192469
rect 47757 192309 47773 192427
rect 47891 192309 47933 192427
rect 48051 192309 48067 192427
rect 47757 174587 48067 192309
rect 47757 174469 47773 174587
rect 47891 174469 47933 174587
rect 48051 174469 48067 174587
rect 47757 174427 48067 174469
rect 47757 174309 47773 174427
rect 47891 174309 47933 174427
rect 48051 174309 48067 174427
rect 47757 156587 48067 174309
rect 47757 156469 47773 156587
rect 47891 156469 47933 156587
rect 48051 156469 48067 156587
rect 47757 156427 48067 156469
rect 47757 156309 47773 156427
rect 47891 156309 47933 156427
rect 48051 156309 48067 156427
rect 47757 138587 48067 156309
rect 47757 138469 47773 138587
rect 47891 138469 47933 138587
rect 48051 138469 48067 138587
rect 47757 138427 48067 138469
rect 47757 138309 47773 138427
rect 47891 138309 47933 138427
rect 48051 138309 48067 138427
rect 47757 120587 48067 138309
rect 47757 120469 47773 120587
rect 47891 120469 47933 120587
rect 48051 120469 48067 120587
rect 47757 120427 48067 120469
rect 47757 120309 47773 120427
rect 47891 120309 47933 120427
rect 48051 120309 48067 120427
rect 47757 102587 48067 120309
rect 47757 102469 47773 102587
rect 47891 102469 47933 102587
rect 48051 102469 48067 102587
rect 47757 102427 48067 102469
rect 47757 102309 47773 102427
rect 47891 102309 47933 102427
rect 48051 102309 48067 102427
rect 47757 84587 48067 102309
rect 47757 84469 47773 84587
rect 47891 84469 47933 84587
rect 48051 84469 48067 84587
rect 47757 84427 48067 84469
rect 47757 84309 47773 84427
rect 47891 84309 47933 84427
rect 48051 84309 48067 84427
rect 47757 66587 48067 84309
rect 47757 66469 47773 66587
rect 47891 66469 47933 66587
rect 48051 66469 48067 66587
rect 47757 66427 48067 66469
rect 47757 66309 47773 66427
rect 47891 66309 47933 66427
rect 48051 66309 48067 66427
rect 47757 48587 48067 66309
rect 47757 48469 47773 48587
rect 47891 48469 47933 48587
rect 48051 48469 48067 48587
rect 47757 48427 48067 48469
rect 47757 48309 47773 48427
rect 47891 48309 47933 48427
rect 48051 48309 48067 48427
rect 47757 30587 48067 48309
rect 47757 30469 47773 30587
rect 47891 30469 47933 30587
rect 48051 30469 48067 30587
rect 47757 30427 48067 30469
rect 47757 30309 47773 30427
rect 47891 30309 47933 30427
rect 48051 30309 48067 30427
rect 47757 12587 48067 30309
rect 47757 12469 47773 12587
rect 47891 12469 47933 12587
rect 48051 12469 48067 12587
rect 47757 12427 48067 12469
rect 47757 12309 47773 12427
rect 47891 12309 47933 12427
rect 48051 12309 48067 12427
rect 47757 -1613 48067 12309
rect 47757 -1731 47773 -1613
rect 47891 -1731 47933 -1613
rect 48051 -1731 48067 -1613
rect 47757 -1773 48067 -1731
rect 47757 -1891 47773 -1773
rect 47891 -1891 47933 -1773
rect 48051 -1891 48067 -1773
rect 47757 -1907 48067 -1891
rect 49617 338447 49927 354541
rect 49617 338329 49633 338447
rect 49751 338329 49793 338447
rect 49911 338329 49927 338447
rect 49617 338287 49927 338329
rect 49617 338169 49633 338287
rect 49751 338169 49793 338287
rect 49911 338169 49927 338287
rect 49617 320447 49927 338169
rect 49617 320329 49633 320447
rect 49751 320329 49793 320447
rect 49911 320329 49927 320447
rect 49617 320287 49927 320329
rect 49617 320169 49633 320287
rect 49751 320169 49793 320287
rect 49911 320169 49927 320287
rect 49617 302447 49927 320169
rect 49617 302329 49633 302447
rect 49751 302329 49793 302447
rect 49911 302329 49927 302447
rect 49617 302287 49927 302329
rect 49617 302169 49633 302287
rect 49751 302169 49793 302287
rect 49911 302169 49927 302287
rect 49617 284447 49927 302169
rect 49617 284329 49633 284447
rect 49751 284329 49793 284447
rect 49911 284329 49927 284447
rect 49617 284287 49927 284329
rect 49617 284169 49633 284287
rect 49751 284169 49793 284287
rect 49911 284169 49927 284287
rect 49617 266447 49927 284169
rect 49617 266329 49633 266447
rect 49751 266329 49793 266447
rect 49911 266329 49927 266447
rect 49617 266287 49927 266329
rect 49617 266169 49633 266287
rect 49751 266169 49793 266287
rect 49911 266169 49927 266287
rect 49617 248447 49927 266169
rect 49617 248329 49633 248447
rect 49751 248329 49793 248447
rect 49911 248329 49927 248447
rect 49617 248287 49927 248329
rect 49617 248169 49633 248287
rect 49751 248169 49793 248287
rect 49911 248169 49927 248287
rect 49617 230447 49927 248169
rect 49617 230329 49633 230447
rect 49751 230329 49793 230447
rect 49911 230329 49927 230447
rect 49617 230287 49927 230329
rect 49617 230169 49633 230287
rect 49751 230169 49793 230287
rect 49911 230169 49927 230287
rect 49617 212447 49927 230169
rect 49617 212329 49633 212447
rect 49751 212329 49793 212447
rect 49911 212329 49927 212447
rect 49617 212287 49927 212329
rect 49617 212169 49633 212287
rect 49751 212169 49793 212287
rect 49911 212169 49927 212287
rect 49617 194447 49927 212169
rect 49617 194329 49633 194447
rect 49751 194329 49793 194447
rect 49911 194329 49927 194447
rect 49617 194287 49927 194329
rect 49617 194169 49633 194287
rect 49751 194169 49793 194287
rect 49911 194169 49927 194287
rect 49617 176447 49927 194169
rect 49617 176329 49633 176447
rect 49751 176329 49793 176447
rect 49911 176329 49927 176447
rect 49617 176287 49927 176329
rect 49617 176169 49633 176287
rect 49751 176169 49793 176287
rect 49911 176169 49927 176287
rect 49617 158447 49927 176169
rect 49617 158329 49633 158447
rect 49751 158329 49793 158447
rect 49911 158329 49927 158447
rect 49617 158287 49927 158329
rect 49617 158169 49633 158287
rect 49751 158169 49793 158287
rect 49911 158169 49927 158287
rect 49617 140447 49927 158169
rect 49617 140329 49633 140447
rect 49751 140329 49793 140447
rect 49911 140329 49927 140447
rect 49617 140287 49927 140329
rect 49617 140169 49633 140287
rect 49751 140169 49793 140287
rect 49911 140169 49927 140287
rect 49617 122447 49927 140169
rect 49617 122329 49633 122447
rect 49751 122329 49793 122447
rect 49911 122329 49927 122447
rect 49617 122287 49927 122329
rect 49617 122169 49633 122287
rect 49751 122169 49793 122287
rect 49911 122169 49927 122287
rect 49617 104447 49927 122169
rect 49617 104329 49633 104447
rect 49751 104329 49793 104447
rect 49911 104329 49927 104447
rect 49617 104287 49927 104329
rect 49617 104169 49633 104287
rect 49751 104169 49793 104287
rect 49911 104169 49927 104287
rect 49617 86447 49927 104169
rect 49617 86329 49633 86447
rect 49751 86329 49793 86447
rect 49911 86329 49927 86447
rect 49617 86287 49927 86329
rect 49617 86169 49633 86287
rect 49751 86169 49793 86287
rect 49911 86169 49927 86287
rect 49617 68447 49927 86169
rect 49617 68329 49633 68447
rect 49751 68329 49793 68447
rect 49911 68329 49927 68447
rect 49617 68287 49927 68329
rect 49617 68169 49633 68287
rect 49751 68169 49793 68287
rect 49911 68169 49927 68287
rect 49617 50447 49927 68169
rect 49617 50329 49633 50447
rect 49751 50329 49793 50447
rect 49911 50329 49927 50447
rect 49617 50287 49927 50329
rect 49617 50169 49633 50287
rect 49751 50169 49793 50287
rect 49911 50169 49927 50287
rect 49617 32447 49927 50169
rect 49617 32329 49633 32447
rect 49751 32329 49793 32447
rect 49911 32329 49927 32447
rect 49617 32287 49927 32329
rect 49617 32169 49633 32287
rect 49751 32169 49793 32287
rect 49911 32169 49927 32287
rect 49617 14447 49927 32169
rect 49617 14329 49633 14447
rect 49751 14329 49793 14447
rect 49911 14329 49927 14447
rect 49617 14287 49927 14329
rect 49617 14169 49633 14287
rect 49751 14169 49793 14287
rect 49911 14169 49927 14287
rect 49617 -2573 49927 14169
rect 49617 -2691 49633 -2573
rect 49751 -2691 49793 -2573
rect 49911 -2691 49927 -2573
rect 49617 -2733 49927 -2691
rect 49617 -2851 49633 -2733
rect 49751 -2851 49793 -2733
rect 49911 -2851 49927 -2733
rect 49617 -2867 49927 -2851
rect 51477 340307 51787 355501
rect 60477 355299 60787 355795
rect 60477 355181 60493 355299
rect 60611 355181 60653 355299
rect 60771 355181 60787 355299
rect 60477 355139 60787 355181
rect 60477 355021 60493 355139
rect 60611 355021 60653 355139
rect 60771 355021 60787 355139
rect 58617 354339 58927 354835
rect 58617 354221 58633 354339
rect 58751 354221 58793 354339
rect 58911 354221 58927 354339
rect 58617 354179 58927 354221
rect 58617 354061 58633 354179
rect 58751 354061 58793 354179
rect 58911 354061 58927 354179
rect 56757 353379 57067 353875
rect 56757 353261 56773 353379
rect 56891 353261 56933 353379
rect 57051 353261 57067 353379
rect 56757 353219 57067 353261
rect 56757 353101 56773 353219
rect 56891 353101 56933 353219
rect 57051 353101 57067 353219
rect 51477 340189 51493 340307
rect 51611 340189 51653 340307
rect 51771 340189 51787 340307
rect 51477 340147 51787 340189
rect 51477 340029 51493 340147
rect 51611 340029 51653 340147
rect 51771 340029 51787 340147
rect 51477 322307 51787 340029
rect 51477 322189 51493 322307
rect 51611 322189 51653 322307
rect 51771 322189 51787 322307
rect 51477 322147 51787 322189
rect 51477 322029 51493 322147
rect 51611 322029 51653 322147
rect 51771 322029 51787 322147
rect 51477 304307 51787 322029
rect 51477 304189 51493 304307
rect 51611 304189 51653 304307
rect 51771 304189 51787 304307
rect 51477 304147 51787 304189
rect 51477 304029 51493 304147
rect 51611 304029 51653 304147
rect 51771 304029 51787 304147
rect 51477 286307 51787 304029
rect 51477 286189 51493 286307
rect 51611 286189 51653 286307
rect 51771 286189 51787 286307
rect 51477 286147 51787 286189
rect 51477 286029 51493 286147
rect 51611 286029 51653 286147
rect 51771 286029 51787 286147
rect 51477 268307 51787 286029
rect 51477 268189 51493 268307
rect 51611 268189 51653 268307
rect 51771 268189 51787 268307
rect 51477 268147 51787 268189
rect 51477 268029 51493 268147
rect 51611 268029 51653 268147
rect 51771 268029 51787 268147
rect 51477 250307 51787 268029
rect 51477 250189 51493 250307
rect 51611 250189 51653 250307
rect 51771 250189 51787 250307
rect 51477 250147 51787 250189
rect 51477 250029 51493 250147
rect 51611 250029 51653 250147
rect 51771 250029 51787 250147
rect 51477 232307 51787 250029
rect 51477 232189 51493 232307
rect 51611 232189 51653 232307
rect 51771 232189 51787 232307
rect 51477 232147 51787 232189
rect 51477 232029 51493 232147
rect 51611 232029 51653 232147
rect 51771 232029 51787 232147
rect 51477 214307 51787 232029
rect 51477 214189 51493 214307
rect 51611 214189 51653 214307
rect 51771 214189 51787 214307
rect 51477 214147 51787 214189
rect 51477 214029 51493 214147
rect 51611 214029 51653 214147
rect 51771 214029 51787 214147
rect 51477 196307 51787 214029
rect 51477 196189 51493 196307
rect 51611 196189 51653 196307
rect 51771 196189 51787 196307
rect 51477 196147 51787 196189
rect 51477 196029 51493 196147
rect 51611 196029 51653 196147
rect 51771 196029 51787 196147
rect 51477 178307 51787 196029
rect 51477 178189 51493 178307
rect 51611 178189 51653 178307
rect 51771 178189 51787 178307
rect 51477 178147 51787 178189
rect 51477 178029 51493 178147
rect 51611 178029 51653 178147
rect 51771 178029 51787 178147
rect 51477 160307 51787 178029
rect 51477 160189 51493 160307
rect 51611 160189 51653 160307
rect 51771 160189 51787 160307
rect 51477 160147 51787 160189
rect 51477 160029 51493 160147
rect 51611 160029 51653 160147
rect 51771 160029 51787 160147
rect 51477 142307 51787 160029
rect 51477 142189 51493 142307
rect 51611 142189 51653 142307
rect 51771 142189 51787 142307
rect 51477 142147 51787 142189
rect 51477 142029 51493 142147
rect 51611 142029 51653 142147
rect 51771 142029 51787 142147
rect 51477 124307 51787 142029
rect 51477 124189 51493 124307
rect 51611 124189 51653 124307
rect 51771 124189 51787 124307
rect 51477 124147 51787 124189
rect 51477 124029 51493 124147
rect 51611 124029 51653 124147
rect 51771 124029 51787 124147
rect 51477 106307 51787 124029
rect 51477 106189 51493 106307
rect 51611 106189 51653 106307
rect 51771 106189 51787 106307
rect 51477 106147 51787 106189
rect 51477 106029 51493 106147
rect 51611 106029 51653 106147
rect 51771 106029 51787 106147
rect 51477 88307 51787 106029
rect 51477 88189 51493 88307
rect 51611 88189 51653 88307
rect 51771 88189 51787 88307
rect 51477 88147 51787 88189
rect 51477 88029 51493 88147
rect 51611 88029 51653 88147
rect 51771 88029 51787 88147
rect 51477 70307 51787 88029
rect 51477 70189 51493 70307
rect 51611 70189 51653 70307
rect 51771 70189 51787 70307
rect 51477 70147 51787 70189
rect 51477 70029 51493 70147
rect 51611 70029 51653 70147
rect 51771 70029 51787 70147
rect 51477 52307 51787 70029
rect 51477 52189 51493 52307
rect 51611 52189 51653 52307
rect 51771 52189 51787 52307
rect 51477 52147 51787 52189
rect 51477 52029 51493 52147
rect 51611 52029 51653 52147
rect 51771 52029 51787 52147
rect 51477 34307 51787 52029
rect 51477 34189 51493 34307
rect 51611 34189 51653 34307
rect 51771 34189 51787 34307
rect 51477 34147 51787 34189
rect 51477 34029 51493 34147
rect 51611 34029 51653 34147
rect 51771 34029 51787 34147
rect 51477 16307 51787 34029
rect 51477 16189 51493 16307
rect 51611 16189 51653 16307
rect 51771 16189 51787 16307
rect 51477 16147 51787 16189
rect 51477 16029 51493 16147
rect 51611 16029 51653 16147
rect 51771 16029 51787 16147
rect 42477 -3171 42493 -3053
rect 42611 -3171 42653 -3053
rect 42771 -3171 42787 -3053
rect 42477 -3213 42787 -3171
rect 42477 -3331 42493 -3213
rect 42611 -3331 42653 -3213
rect 42771 -3331 42787 -3213
rect 42477 -3827 42787 -3331
rect 51477 -3533 51787 16029
rect 54897 352419 55207 352915
rect 54897 352301 54913 352419
rect 55031 352301 55073 352419
rect 55191 352301 55207 352419
rect 54897 352259 55207 352301
rect 54897 352141 54913 352259
rect 55031 352141 55073 352259
rect 55191 352141 55207 352259
rect 54897 343727 55207 352141
rect 54897 343609 54913 343727
rect 55031 343609 55073 343727
rect 55191 343609 55207 343727
rect 54897 343567 55207 343609
rect 54897 343449 54913 343567
rect 55031 343449 55073 343567
rect 55191 343449 55207 343567
rect 54897 325727 55207 343449
rect 54897 325609 54913 325727
rect 55031 325609 55073 325727
rect 55191 325609 55207 325727
rect 54897 325567 55207 325609
rect 54897 325449 54913 325567
rect 55031 325449 55073 325567
rect 55191 325449 55207 325567
rect 54897 307727 55207 325449
rect 54897 307609 54913 307727
rect 55031 307609 55073 307727
rect 55191 307609 55207 307727
rect 54897 307567 55207 307609
rect 54897 307449 54913 307567
rect 55031 307449 55073 307567
rect 55191 307449 55207 307567
rect 54897 289727 55207 307449
rect 54897 289609 54913 289727
rect 55031 289609 55073 289727
rect 55191 289609 55207 289727
rect 54897 289567 55207 289609
rect 54897 289449 54913 289567
rect 55031 289449 55073 289567
rect 55191 289449 55207 289567
rect 54897 271727 55207 289449
rect 54897 271609 54913 271727
rect 55031 271609 55073 271727
rect 55191 271609 55207 271727
rect 54897 271567 55207 271609
rect 54897 271449 54913 271567
rect 55031 271449 55073 271567
rect 55191 271449 55207 271567
rect 54897 253727 55207 271449
rect 54897 253609 54913 253727
rect 55031 253609 55073 253727
rect 55191 253609 55207 253727
rect 54897 253567 55207 253609
rect 54897 253449 54913 253567
rect 55031 253449 55073 253567
rect 55191 253449 55207 253567
rect 54897 235727 55207 253449
rect 54897 235609 54913 235727
rect 55031 235609 55073 235727
rect 55191 235609 55207 235727
rect 54897 235567 55207 235609
rect 54897 235449 54913 235567
rect 55031 235449 55073 235567
rect 55191 235449 55207 235567
rect 54897 217727 55207 235449
rect 54897 217609 54913 217727
rect 55031 217609 55073 217727
rect 55191 217609 55207 217727
rect 54897 217567 55207 217609
rect 54897 217449 54913 217567
rect 55031 217449 55073 217567
rect 55191 217449 55207 217567
rect 54897 199727 55207 217449
rect 54897 199609 54913 199727
rect 55031 199609 55073 199727
rect 55191 199609 55207 199727
rect 54897 199567 55207 199609
rect 54897 199449 54913 199567
rect 55031 199449 55073 199567
rect 55191 199449 55207 199567
rect 54897 181727 55207 199449
rect 54897 181609 54913 181727
rect 55031 181609 55073 181727
rect 55191 181609 55207 181727
rect 54897 181567 55207 181609
rect 54897 181449 54913 181567
rect 55031 181449 55073 181567
rect 55191 181449 55207 181567
rect 54897 163727 55207 181449
rect 54897 163609 54913 163727
rect 55031 163609 55073 163727
rect 55191 163609 55207 163727
rect 54897 163567 55207 163609
rect 54897 163449 54913 163567
rect 55031 163449 55073 163567
rect 55191 163449 55207 163567
rect 54897 145727 55207 163449
rect 54897 145609 54913 145727
rect 55031 145609 55073 145727
rect 55191 145609 55207 145727
rect 54897 145567 55207 145609
rect 54897 145449 54913 145567
rect 55031 145449 55073 145567
rect 55191 145449 55207 145567
rect 54897 127727 55207 145449
rect 54897 127609 54913 127727
rect 55031 127609 55073 127727
rect 55191 127609 55207 127727
rect 54897 127567 55207 127609
rect 54897 127449 54913 127567
rect 55031 127449 55073 127567
rect 55191 127449 55207 127567
rect 54897 109727 55207 127449
rect 54897 109609 54913 109727
rect 55031 109609 55073 109727
rect 55191 109609 55207 109727
rect 54897 109567 55207 109609
rect 54897 109449 54913 109567
rect 55031 109449 55073 109567
rect 55191 109449 55207 109567
rect 54897 91727 55207 109449
rect 54897 91609 54913 91727
rect 55031 91609 55073 91727
rect 55191 91609 55207 91727
rect 54897 91567 55207 91609
rect 54897 91449 54913 91567
rect 55031 91449 55073 91567
rect 55191 91449 55207 91567
rect 54897 73727 55207 91449
rect 54897 73609 54913 73727
rect 55031 73609 55073 73727
rect 55191 73609 55207 73727
rect 54897 73567 55207 73609
rect 54897 73449 54913 73567
rect 55031 73449 55073 73567
rect 55191 73449 55207 73567
rect 54897 55727 55207 73449
rect 54897 55609 54913 55727
rect 55031 55609 55073 55727
rect 55191 55609 55207 55727
rect 54897 55567 55207 55609
rect 54897 55449 54913 55567
rect 55031 55449 55073 55567
rect 55191 55449 55207 55567
rect 54897 37727 55207 55449
rect 54897 37609 54913 37727
rect 55031 37609 55073 37727
rect 55191 37609 55207 37727
rect 54897 37567 55207 37609
rect 54897 37449 54913 37567
rect 55031 37449 55073 37567
rect 55191 37449 55207 37567
rect 54897 19727 55207 37449
rect 54897 19609 54913 19727
rect 55031 19609 55073 19727
rect 55191 19609 55207 19727
rect 54897 19567 55207 19609
rect 54897 19449 54913 19567
rect 55031 19449 55073 19567
rect 55191 19449 55207 19567
rect 54897 1727 55207 19449
rect 54897 1609 54913 1727
rect 55031 1609 55073 1727
rect 55191 1609 55207 1727
rect 54897 1567 55207 1609
rect 54897 1449 54913 1567
rect 55031 1449 55073 1567
rect 55191 1449 55207 1567
rect 54897 -173 55207 1449
rect 54897 -291 54913 -173
rect 55031 -291 55073 -173
rect 55191 -291 55207 -173
rect 54897 -333 55207 -291
rect 54897 -451 54913 -333
rect 55031 -451 55073 -333
rect 55191 -451 55207 -333
rect 54897 -947 55207 -451
rect 56757 345587 57067 353101
rect 56757 345469 56773 345587
rect 56891 345469 56933 345587
rect 57051 345469 57067 345587
rect 56757 345427 57067 345469
rect 56757 345309 56773 345427
rect 56891 345309 56933 345427
rect 57051 345309 57067 345427
rect 56757 327587 57067 345309
rect 56757 327469 56773 327587
rect 56891 327469 56933 327587
rect 57051 327469 57067 327587
rect 56757 327427 57067 327469
rect 56757 327309 56773 327427
rect 56891 327309 56933 327427
rect 57051 327309 57067 327427
rect 56757 309587 57067 327309
rect 56757 309469 56773 309587
rect 56891 309469 56933 309587
rect 57051 309469 57067 309587
rect 56757 309427 57067 309469
rect 56757 309309 56773 309427
rect 56891 309309 56933 309427
rect 57051 309309 57067 309427
rect 56757 291587 57067 309309
rect 56757 291469 56773 291587
rect 56891 291469 56933 291587
rect 57051 291469 57067 291587
rect 56757 291427 57067 291469
rect 56757 291309 56773 291427
rect 56891 291309 56933 291427
rect 57051 291309 57067 291427
rect 56757 273587 57067 291309
rect 56757 273469 56773 273587
rect 56891 273469 56933 273587
rect 57051 273469 57067 273587
rect 56757 273427 57067 273469
rect 56757 273309 56773 273427
rect 56891 273309 56933 273427
rect 57051 273309 57067 273427
rect 56757 255587 57067 273309
rect 56757 255469 56773 255587
rect 56891 255469 56933 255587
rect 57051 255469 57067 255587
rect 56757 255427 57067 255469
rect 56757 255309 56773 255427
rect 56891 255309 56933 255427
rect 57051 255309 57067 255427
rect 56757 237587 57067 255309
rect 56757 237469 56773 237587
rect 56891 237469 56933 237587
rect 57051 237469 57067 237587
rect 56757 237427 57067 237469
rect 56757 237309 56773 237427
rect 56891 237309 56933 237427
rect 57051 237309 57067 237427
rect 56757 219587 57067 237309
rect 56757 219469 56773 219587
rect 56891 219469 56933 219587
rect 57051 219469 57067 219587
rect 56757 219427 57067 219469
rect 56757 219309 56773 219427
rect 56891 219309 56933 219427
rect 57051 219309 57067 219427
rect 56757 201587 57067 219309
rect 56757 201469 56773 201587
rect 56891 201469 56933 201587
rect 57051 201469 57067 201587
rect 56757 201427 57067 201469
rect 56757 201309 56773 201427
rect 56891 201309 56933 201427
rect 57051 201309 57067 201427
rect 56757 183587 57067 201309
rect 56757 183469 56773 183587
rect 56891 183469 56933 183587
rect 57051 183469 57067 183587
rect 56757 183427 57067 183469
rect 56757 183309 56773 183427
rect 56891 183309 56933 183427
rect 57051 183309 57067 183427
rect 56757 165587 57067 183309
rect 56757 165469 56773 165587
rect 56891 165469 56933 165587
rect 57051 165469 57067 165587
rect 56757 165427 57067 165469
rect 56757 165309 56773 165427
rect 56891 165309 56933 165427
rect 57051 165309 57067 165427
rect 56757 147587 57067 165309
rect 56757 147469 56773 147587
rect 56891 147469 56933 147587
rect 57051 147469 57067 147587
rect 56757 147427 57067 147469
rect 56757 147309 56773 147427
rect 56891 147309 56933 147427
rect 57051 147309 57067 147427
rect 56757 129587 57067 147309
rect 56757 129469 56773 129587
rect 56891 129469 56933 129587
rect 57051 129469 57067 129587
rect 56757 129427 57067 129469
rect 56757 129309 56773 129427
rect 56891 129309 56933 129427
rect 57051 129309 57067 129427
rect 56757 111587 57067 129309
rect 56757 111469 56773 111587
rect 56891 111469 56933 111587
rect 57051 111469 57067 111587
rect 56757 111427 57067 111469
rect 56757 111309 56773 111427
rect 56891 111309 56933 111427
rect 57051 111309 57067 111427
rect 56757 93587 57067 111309
rect 56757 93469 56773 93587
rect 56891 93469 56933 93587
rect 57051 93469 57067 93587
rect 56757 93427 57067 93469
rect 56757 93309 56773 93427
rect 56891 93309 56933 93427
rect 57051 93309 57067 93427
rect 56757 75587 57067 93309
rect 56757 75469 56773 75587
rect 56891 75469 56933 75587
rect 57051 75469 57067 75587
rect 56757 75427 57067 75469
rect 56757 75309 56773 75427
rect 56891 75309 56933 75427
rect 57051 75309 57067 75427
rect 56757 57587 57067 75309
rect 56757 57469 56773 57587
rect 56891 57469 56933 57587
rect 57051 57469 57067 57587
rect 56757 57427 57067 57469
rect 56757 57309 56773 57427
rect 56891 57309 56933 57427
rect 57051 57309 57067 57427
rect 56757 39587 57067 57309
rect 56757 39469 56773 39587
rect 56891 39469 56933 39587
rect 57051 39469 57067 39587
rect 56757 39427 57067 39469
rect 56757 39309 56773 39427
rect 56891 39309 56933 39427
rect 57051 39309 57067 39427
rect 56757 21587 57067 39309
rect 56757 21469 56773 21587
rect 56891 21469 56933 21587
rect 57051 21469 57067 21587
rect 56757 21427 57067 21469
rect 56757 21309 56773 21427
rect 56891 21309 56933 21427
rect 57051 21309 57067 21427
rect 56757 3587 57067 21309
rect 56757 3469 56773 3587
rect 56891 3469 56933 3587
rect 57051 3469 57067 3587
rect 56757 3427 57067 3469
rect 56757 3309 56773 3427
rect 56891 3309 56933 3427
rect 57051 3309 57067 3427
rect 56757 -1133 57067 3309
rect 56757 -1251 56773 -1133
rect 56891 -1251 56933 -1133
rect 57051 -1251 57067 -1133
rect 56757 -1293 57067 -1251
rect 56757 -1411 56773 -1293
rect 56891 -1411 56933 -1293
rect 57051 -1411 57067 -1293
rect 56757 -1907 57067 -1411
rect 58617 347447 58927 354061
rect 58617 347329 58633 347447
rect 58751 347329 58793 347447
rect 58911 347329 58927 347447
rect 58617 347287 58927 347329
rect 58617 347169 58633 347287
rect 58751 347169 58793 347287
rect 58911 347169 58927 347287
rect 58617 329447 58927 347169
rect 58617 329329 58633 329447
rect 58751 329329 58793 329447
rect 58911 329329 58927 329447
rect 58617 329287 58927 329329
rect 58617 329169 58633 329287
rect 58751 329169 58793 329287
rect 58911 329169 58927 329287
rect 58617 311447 58927 329169
rect 58617 311329 58633 311447
rect 58751 311329 58793 311447
rect 58911 311329 58927 311447
rect 58617 311287 58927 311329
rect 58617 311169 58633 311287
rect 58751 311169 58793 311287
rect 58911 311169 58927 311287
rect 58617 293447 58927 311169
rect 58617 293329 58633 293447
rect 58751 293329 58793 293447
rect 58911 293329 58927 293447
rect 58617 293287 58927 293329
rect 58617 293169 58633 293287
rect 58751 293169 58793 293287
rect 58911 293169 58927 293287
rect 58617 275447 58927 293169
rect 58617 275329 58633 275447
rect 58751 275329 58793 275447
rect 58911 275329 58927 275447
rect 58617 275287 58927 275329
rect 58617 275169 58633 275287
rect 58751 275169 58793 275287
rect 58911 275169 58927 275287
rect 58617 257447 58927 275169
rect 58617 257329 58633 257447
rect 58751 257329 58793 257447
rect 58911 257329 58927 257447
rect 58617 257287 58927 257329
rect 58617 257169 58633 257287
rect 58751 257169 58793 257287
rect 58911 257169 58927 257287
rect 58617 239447 58927 257169
rect 58617 239329 58633 239447
rect 58751 239329 58793 239447
rect 58911 239329 58927 239447
rect 58617 239287 58927 239329
rect 58617 239169 58633 239287
rect 58751 239169 58793 239287
rect 58911 239169 58927 239287
rect 58617 221447 58927 239169
rect 58617 221329 58633 221447
rect 58751 221329 58793 221447
rect 58911 221329 58927 221447
rect 58617 221287 58927 221329
rect 58617 221169 58633 221287
rect 58751 221169 58793 221287
rect 58911 221169 58927 221287
rect 58617 203447 58927 221169
rect 58617 203329 58633 203447
rect 58751 203329 58793 203447
rect 58911 203329 58927 203447
rect 58617 203287 58927 203329
rect 58617 203169 58633 203287
rect 58751 203169 58793 203287
rect 58911 203169 58927 203287
rect 58617 185447 58927 203169
rect 58617 185329 58633 185447
rect 58751 185329 58793 185447
rect 58911 185329 58927 185447
rect 58617 185287 58927 185329
rect 58617 185169 58633 185287
rect 58751 185169 58793 185287
rect 58911 185169 58927 185287
rect 58617 167447 58927 185169
rect 58617 167329 58633 167447
rect 58751 167329 58793 167447
rect 58911 167329 58927 167447
rect 58617 167287 58927 167329
rect 58617 167169 58633 167287
rect 58751 167169 58793 167287
rect 58911 167169 58927 167287
rect 58617 149447 58927 167169
rect 58617 149329 58633 149447
rect 58751 149329 58793 149447
rect 58911 149329 58927 149447
rect 58617 149287 58927 149329
rect 58617 149169 58633 149287
rect 58751 149169 58793 149287
rect 58911 149169 58927 149287
rect 58617 131447 58927 149169
rect 58617 131329 58633 131447
rect 58751 131329 58793 131447
rect 58911 131329 58927 131447
rect 58617 131287 58927 131329
rect 58617 131169 58633 131287
rect 58751 131169 58793 131287
rect 58911 131169 58927 131287
rect 58617 113447 58927 131169
rect 58617 113329 58633 113447
rect 58751 113329 58793 113447
rect 58911 113329 58927 113447
rect 58617 113287 58927 113329
rect 58617 113169 58633 113287
rect 58751 113169 58793 113287
rect 58911 113169 58927 113287
rect 58617 95447 58927 113169
rect 58617 95329 58633 95447
rect 58751 95329 58793 95447
rect 58911 95329 58927 95447
rect 58617 95287 58927 95329
rect 58617 95169 58633 95287
rect 58751 95169 58793 95287
rect 58911 95169 58927 95287
rect 58617 77447 58927 95169
rect 58617 77329 58633 77447
rect 58751 77329 58793 77447
rect 58911 77329 58927 77447
rect 58617 77287 58927 77329
rect 58617 77169 58633 77287
rect 58751 77169 58793 77287
rect 58911 77169 58927 77287
rect 58617 59447 58927 77169
rect 58617 59329 58633 59447
rect 58751 59329 58793 59447
rect 58911 59329 58927 59447
rect 58617 59287 58927 59329
rect 58617 59169 58633 59287
rect 58751 59169 58793 59287
rect 58911 59169 58927 59287
rect 58617 41447 58927 59169
rect 58617 41329 58633 41447
rect 58751 41329 58793 41447
rect 58911 41329 58927 41447
rect 58617 41287 58927 41329
rect 58617 41169 58633 41287
rect 58751 41169 58793 41287
rect 58911 41169 58927 41287
rect 58617 23447 58927 41169
rect 58617 23329 58633 23447
rect 58751 23329 58793 23447
rect 58911 23329 58927 23447
rect 58617 23287 58927 23329
rect 58617 23169 58633 23287
rect 58751 23169 58793 23287
rect 58911 23169 58927 23287
rect 58617 5447 58927 23169
rect 58617 5329 58633 5447
rect 58751 5329 58793 5447
rect 58911 5329 58927 5447
rect 58617 5287 58927 5329
rect 58617 5169 58633 5287
rect 58751 5169 58793 5287
rect 58911 5169 58927 5287
rect 58617 -2093 58927 5169
rect 58617 -2211 58633 -2093
rect 58751 -2211 58793 -2093
rect 58911 -2211 58927 -2093
rect 58617 -2253 58927 -2211
rect 58617 -2371 58633 -2253
rect 58751 -2371 58793 -2253
rect 58911 -2371 58927 -2253
rect 58617 -2867 58927 -2371
rect 60477 349307 60787 355021
rect 69477 355779 69787 355795
rect 69477 355661 69493 355779
rect 69611 355661 69653 355779
rect 69771 355661 69787 355779
rect 69477 355619 69787 355661
rect 69477 355501 69493 355619
rect 69611 355501 69653 355619
rect 69771 355501 69787 355619
rect 67617 354819 67927 354835
rect 67617 354701 67633 354819
rect 67751 354701 67793 354819
rect 67911 354701 67927 354819
rect 67617 354659 67927 354701
rect 67617 354541 67633 354659
rect 67751 354541 67793 354659
rect 67911 354541 67927 354659
rect 65757 353859 66067 353875
rect 65757 353741 65773 353859
rect 65891 353741 65933 353859
rect 66051 353741 66067 353859
rect 65757 353699 66067 353741
rect 65757 353581 65773 353699
rect 65891 353581 65933 353699
rect 66051 353581 66067 353699
rect 60477 349189 60493 349307
rect 60611 349189 60653 349307
rect 60771 349189 60787 349307
rect 60477 349147 60787 349189
rect 60477 349029 60493 349147
rect 60611 349029 60653 349147
rect 60771 349029 60787 349147
rect 60477 331307 60787 349029
rect 60477 331189 60493 331307
rect 60611 331189 60653 331307
rect 60771 331189 60787 331307
rect 60477 331147 60787 331189
rect 60477 331029 60493 331147
rect 60611 331029 60653 331147
rect 60771 331029 60787 331147
rect 60477 313307 60787 331029
rect 60477 313189 60493 313307
rect 60611 313189 60653 313307
rect 60771 313189 60787 313307
rect 60477 313147 60787 313189
rect 60477 313029 60493 313147
rect 60611 313029 60653 313147
rect 60771 313029 60787 313147
rect 60477 295307 60787 313029
rect 60477 295189 60493 295307
rect 60611 295189 60653 295307
rect 60771 295189 60787 295307
rect 60477 295147 60787 295189
rect 60477 295029 60493 295147
rect 60611 295029 60653 295147
rect 60771 295029 60787 295147
rect 60477 277307 60787 295029
rect 60477 277189 60493 277307
rect 60611 277189 60653 277307
rect 60771 277189 60787 277307
rect 60477 277147 60787 277189
rect 60477 277029 60493 277147
rect 60611 277029 60653 277147
rect 60771 277029 60787 277147
rect 60477 259307 60787 277029
rect 60477 259189 60493 259307
rect 60611 259189 60653 259307
rect 60771 259189 60787 259307
rect 60477 259147 60787 259189
rect 60477 259029 60493 259147
rect 60611 259029 60653 259147
rect 60771 259029 60787 259147
rect 60477 241307 60787 259029
rect 60477 241189 60493 241307
rect 60611 241189 60653 241307
rect 60771 241189 60787 241307
rect 60477 241147 60787 241189
rect 60477 241029 60493 241147
rect 60611 241029 60653 241147
rect 60771 241029 60787 241147
rect 60477 223307 60787 241029
rect 60477 223189 60493 223307
rect 60611 223189 60653 223307
rect 60771 223189 60787 223307
rect 60477 223147 60787 223189
rect 60477 223029 60493 223147
rect 60611 223029 60653 223147
rect 60771 223029 60787 223147
rect 60477 205307 60787 223029
rect 60477 205189 60493 205307
rect 60611 205189 60653 205307
rect 60771 205189 60787 205307
rect 60477 205147 60787 205189
rect 60477 205029 60493 205147
rect 60611 205029 60653 205147
rect 60771 205029 60787 205147
rect 60477 187307 60787 205029
rect 60477 187189 60493 187307
rect 60611 187189 60653 187307
rect 60771 187189 60787 187307
rect 60477 187147 60787 187189
rect 60477 187029 60493 187147
rect 60611 187029 60653 187147
rect 60771 187029 60787 187147
rect 60477 169307 60787 187029
rect 60477 169189 60493 169307
rect 60611 169189 60653 169307
rect 60771 169189 60787 169307
rect 60477 169147 60787 169189
rect 60477 169029 60493 169147
rect 60611 169029 60653 169147
rect 60771 169029 60787 169147
rect 60477 151307 60787 169029
rect 60477 151189 60493 151307
rect 60611 151189 60653 151307
rect 60771 151189 60787 151307
rect 60477 151147 60787 151189
rect 60477 151029 60493 151147
rect 60611 151029 60653 151147
rect 60771 151029 60787 151147
rect 60477 133307 60787 151029
rect 60477 133189 60493 133307
rect 60611 133189 60653 133307
rect 60771 133189 60787 133307
rect 60477 133147 60787 133189
rect 60477 133029 60493 133147
rect 60611 133029 60653 133147
rect 60771 133029 60787 133147
rect 60477 115307 60787 133029
rect 60477 115189 60493 115307
rect 60611 115189 60653 115307
rect 60771 115189 60787 115307
rect 60477 115147 60787 115189
rect 60477 115029 60493 115147
rect 60611 115029 60653 115147
rect 60771 115029 60787 115147
rect 60477 97307 60787 115029
rect 60477 97189 60493 97307
rect 60611 97189 60653 97307
rect 60771 97189 60787 97307
rect 60477 97147 60787 97189
rect 60477 97029 60493 97147
rect 60611 97029 60653 97147
rect 60771 97029 60787 97147
rect 60477 79307 60787 97029
rect 60477 79189 60493 79307
rect 60611 79189 60653 79307
rect 60771 79189 60787 79307
rect 60477 79147 60787 79189
rect 60477 79029 60493 79147
rect 60611 79029 60653 79147
rect 60771 79029 60787 79147
rect 60477 61307 60787 79029
rect 60477 61189 60493 61307
rect 60611 61189 60653 61307
rect 60771 61189 60787 61307
rect 60477 61147 60787 61189
rect 60477 61029 60493 61147
rect 60611 61029 60653 61147
rect 60771 61029 60787 61147
rect 60477 43307 60787 61029
rect 60477 43189 60493 43307
rect 60611 43189 60653 43307
rect 60771 43189 60787 43307
rect 60477 43147 60787 43189
rect 60477 43029 60493 43147
rect 60611 43029 60653 43147
rect 60771 43029 60787 43147
rect 60477 25307 60787 43029
rect 60477 25189 60493 25307
rect 60611 25189 60653 25307
rect 60771 25189 60787 25307
rect 60477 25147 60787 25189
rect 60477 25029 60493 25147
rect 60611 25029 60653 25147
rect 60771 25029 60787 25147
rect 60477 7307 60787 25029
rect 60477 7189 60493 7307
rect 60611 7189 60653 7307
rect 60771 7189 60787 7307
rect 60477 7147 60787 7189
rect 60477 7029 60493 7147
rect 60611 7029 60653 7147
rect 60771 7029 60787 7147
rect 51477 -3651 51493 -3533
rect 51611 -3651 51653 -3533
rect 51771 -3651 51787 -3533
rect 51477 -3693 51787 -3651
rect 51477 -3811 51493 -3693
rect 51611 -3811 51653 -3693
rect 51771 -3811 51787 -3693
rect 51477 -3827 51787 -3811
rect 60477 -3053 60787 7029
rect 63897 352899 64207 352915
rect 63897 352781 63913 352899
rect 64031 352781 64073 352899
rect 64191 352781 64207 352899
rect 63897 352739 64207 352781
rect 63897 352621 63913 352739
rect 64031 352621 64073 352739
rect 64191 352621 64207 352739
rect 63897 334727 64207 352621
rect 63897 334609 63913 334727
rect 64031 334609 64073 334727
rect 64191 334609 64207 334727
rect 63897 334567 64207 334609
rect 63897 334449 63913 334567
rect 64031 334449 64073 334567
rect 64191 334449 64207 334567
rect 63897 316727 64207 334449
rect 63897 316609 63913 316727
rect 64031 316609 64073 316727
rect 64191 316609 64207 316727
rect 63897 316567 64207 316609
rect 63897 316449 63913 316567
rect 64031 316449 64073 316567
rect 64191 316449 64207 316567
rect 63897 298727 64207 316449
rect 63897 298609 63913 298727
rect 64031 298609 64073 298727
rect 64191 298609 64207 298727
rect 63897 298567 64207 298609
rect 63897 298449 63913 298567
rect 64031 298449 64073 298567
rect 64191 298449 64207 298567
rect 63897 280727 64207 298449
rect 63897 280609 63913 280727
rect 64031 280609 64073 280727
rect 64191 280609 64207 280727
rect 63897 280567 64207 280609
rect 63897 280449 63913 280567
rect 64031 280449 64073 280567
rect 64191 280449 64207 280567
rect 63897 262727 64207 280449
rect 63897 262609 63913 262727
rect 64031 262609 64073 262727
rect 64191 262609 64207 262727
rect 63897 262567 64207 262609
rect 63897 262449 63913 262567
rect 64031 262449 64073 262567
rect 64191 262449 64207 262567
rect 63897 244727 64207 262449
rect 63897 244609 63913 244727
rect 64031 244609 64073 244727
rect 64191 244609 64207 244727
rect 63897 244567 64207 244609
rect 63897 244449 63913 244567
rect 64031 244449 64073 244567
rect 64191 244449 64207 244567
rect 63897 226727 64207 244449
rect 63897 226609 63913 226727
rect 64031 226609 64073 226727
rect 64191 226609 64207 226727
rect 63897 226567 64207 226609
rect 63897 226449 63913 226567
rect 64031 226449 64073 226567
rect 64191 226449 64207 226567
rect 63897 208727 64207 226449
rect 63897 208609 63913 208727
rect 64031 208609 64073 208727
rect 64191 208609 64207 208727
rect 63897 208567 64207 208609
rect 63897 208449 63913 208567
rect 64031 208449 64073 208567
rect 64191 208449 64207 208567
rect 63897 190727 64207 208449
rect 63897 190609 63913 190727
rect 64031 190609 64073 190727
rect 64191 190609 64207 190727
rect 63897 190567 64207 190609
rect 63897 190449 63913 190567
rect 64031 190449 64073 190567
rect 64191 190449 64207 190567
rect 63897 172727 64207 190449
rect 63897 172609 63913 172727
rect 64031 172609 64073 172727
rect 64191 172609 64207 172727
rect 63897 172567 64207 172609
rect 63897 172449 63913 172567
rect 64031 172449 64073 172567
rect 64191 172449 64207 172567
rect 63897 154727 64207 172449
rect 63897 154609 63913 154727
rect 64031 154609 64073 154727
rect 64191 154609 64207 154727
rect 63897 154567 64207 154609
rect 63897 154449 63913 154567
rect 64031 154449 64073 154567
rect 64191 154449 64207 154567
rect 63897 136727 64207 154449
rect 63897 136609 63913 136727
rect 64031 136609 64073 136727
rect 64191 136609 64207 136727
rect 63897 136567 64207 136609
rect 63897 136449 63913 136567
rect 64031 136449 64073 136567
rect 64191 136449 64207 136567
rect 63897 118727 64207 136449
rect 63897 118609 63913 118727
rect 64031 118609 64073 118727
rect 64191 118609 64207 118727
rect 63897 118567 64207 118609
rect 63897 118449 63913 118567
rect 64031 118449 64073 118567
rect 64191 118449 64207 118567
rect 63897 100727 64207 118449
rect 63897 100609 63913 100727
rect 64031 100609 64073 100727
rect 64191 100609 64207 100727
rect 63897 100567 64207 100609
rect 63897 100449 63913 100567
rect 64031 100449 64073 100567
rect 64191 100449 64207 100567
rect 63897 82727 64207 100449
rect 63897 82609 63913 82727
rect 64031 82609 64073 82727
rect 64191 82609 64207 82727
rect 63897 82567 64207 82609
rect 63897 82449 63913 82567
rect 64031 82449 64073 82567
rect 64191 82449 64207 82567
rect 63897 64727 64207 82449
rect 63897 64609 63913 64727
rect 64031 64609 64073 64727
rect 64191 64609 64207 64727
rect 63897 64567 64207 64609
rect 63897 64449 63913 64567
rect 64031 64449 64073 64567
rect 64191 64449 64207 64567
rect 63897 46727 64207 64449
rect 63897 46609 63913 46727
rect 64031 46609 64073 46727
rect 64191 46609 64207 46727
rect 63897 46567 64207 46609
rect 63897 46449 63913 46567
rect 64031 46449 64073 46567
rect 64191 46449 64207 46567
rect 63897 28727 64207 46449
rect 63897 28609 63913 28727
rect 64031 28609 64073 28727
rect 64191 28609 64207 28727
rect 63897 28567 64207 28609
rect 63897 28449 63913 28567
rect 64031 28449 64073 28567
rect 64191 28449 64207 28567
rect 63897 10727 64207 28449
rect 63897 10609 63913 10727
rect 64031 10609 64073 10727
rect 64191 10609 64207 10727
rect 63897 10567 64207 10609
rect 63897 10449 63913 10567
rect 64031 10449 64073 10567
rect 64191 10449 64207 10567
rect 63897 -653 64207 10449
rect 63897 -771 63913 -653
rect 64031 -771 64073 -653
rect 64191 -771 64207 -653
rect 63897 -813 64207 -771
rect 63897 -931 63913 -813
rect 64031 -931 64073 -813
rect 64191 -931 64207 -813
rect 63897 -947 64207 -931
rect 65757 336587 66067 353581
rect 65757 336469 65773 336587
rect 65891 336469 65933 336587
rect 66051 336469 66067 336587
rect 65757 336427 66067 336469
rect 65757 336309 65773 336427
rect 65891 336309 65933 336427
rect 66051 336309 66067 336427
rect 65757 318587 66067 336309
rect 65757 318469 65773 318587
rect 65891 318469 65933 318587
rect 66051 318469 66067 318587
rect 65757 318427 66067 318469
rect 65757 318309 65773 318427
rect 65891 318309 65933 318427
rect 66051 318309 66067 318427
rect 65757 300587 66067 318309
rect 65757 300469 65773 300587
rect 65891 300469 65933 300587
rect 66051 300469 66067 300587
rect 65757 300427 66067 300469
rect 65757 300309 65773 300427
rect 65891 300309 65933 300427
rect 66051 300309 66067 300427
rect 65757 282587 66067 300309
rect 65757 282469 65773 282587
rect 65891 282469 65933 282587
rect 66051 282469 66067 282587
rect 65757 282427 66067 282469
rect 65757 282309 65773 282427
rect 65891 282309 65933 282427
rect 66051 282309 66067 282427
rect 65757 264587 66067 282309
rect 65757 264469 65773 264587
rect 65891 264469 65933 264587
rect 66051 264469 66067 264587
rect 65757 264427 66067 264469
rect 65757 264309 65773 264427
rect 65891 264309 65933 264427
rect 66051 264309 66067 264427
rect 65757 246587 66067 264309
rect 65757 246469 65773 246587
rect 65891 246469 65933 246587
rect 66051 246469 66067 246587
rect 65757 246427 66067 246469
rect 65757 246309 65773 246427
rect 65891 246309 65933 246427
rect 66051 246309 66067 246427
rect 65757 228587 66067 246309
rect 65757 228469 65773 228587
rect 65891 228469 65933 228587
rect 66051 228469 66067 228587
rect 65757 228427 66067 228469
rect 65757 228309 65773 228427
rect 65891 228309 65933 228427
rect 66051 228309 66067 228427
rect 65757 210587 66067 228309
rect 65757 210469 65773 210587
rect 65891 210469 65933 210587
rect 66051 210469 66067 210587
rect 65757 210427 66067 210469
rect 65757 210309 65773 210427
rect 65891 210309 65933 210427
rect 66051 210309 66067 210427
rect 65757 192587 66067 210309
rect 65757 192469 65773 192587
rect 65891 192469 65933 192587
rect 66051 192469 66067 192587
rect 65757 192427 66067 192469
rect 65757 192309 65773 192427
rect 65891 192309 65933 192427
rect 66051 192309 66067 192427
rect 65757 174587 66067 192309
rect 65757 174469 65773 174587
rect 65891 174469 65933 174587
rect 66051 174469 66067 174587
rect 65757 174427 66067 174469
rect 65757 174309 65773 174427
rect 65891 174309 65933 174427
rect 66051 174309 66067 174427
rect 65757 156587 66067 174309
rect 65757 156469 65773 156587
rect 65891 156469 65933 156587
rect 66051 156469 66067 156587
rect 65757 156427 66067 156469
rect 65757 156309 65773 156427
rect 65891 156309 65933 156427
rect 66051 156309 66067 156427
rect 65757 138587 66067 156309
rect 65757 138469 65773 138587
rect 65891 138469 65933 138587
rect 66051 138469 66067 138587
rect 65757 138427 66067 138469
rect 65757 138309 65773 138427
rect 65891 138309 65933 138427
rect 66051 138309 66067 138427
rect 65757 120587 66067 138309
rect 65757 120469 65773 120587
rect 65891 120469 65933 120587
rect 66051 120469 66067 120587
rect 65757 120427 66067 120469
rect 65757 120309 65773 120427
rect 65891 120309 65933 120427
rect 66051 120309 66067 120427
rect 65757 102587 66067 120309
rect 65757 102469 65773 102587
rect 65891 102469 65933 102587
rect 66051 102469 66067 102587
rect 65757 102427 66067 102469
rect 65757 102309 65773 102427
rect 65891 102309 65933 102427
rect 66051 102309 66067 102427
rect 65757 84587 66067 102309
rect 65757 84469 65773 84587
rect 65891 84469 65933 84587
rect 66051 84469 66067 84587
rect 65757 84427 66067 84469
rect 65757 84309 65773 84427
rect 65891 84309 65933 84427
rect 66051 84309 66067 84427
rect 65757 66587 66067 84309
rect 65757 66469 65773 66587
rect 65891 66469 65933 66587
rect 66051 66469 66067 66587
rect 65757 66427 66067 66469
rect 65757 66309 65773 66427
rect 65891 66309 65933 66427
rect 66051 66309 66067 66427
rect 65757 48587 66067 66309
rect 65757 48469 65773 48587
rect 65891 48469 65933 48587
rect 66051 48469 66067 48587
rect 65757 48427 66067 48469
rect 65757 48309 65773 48427
rect 65891 48309 65933 48427
rect 66051 48309 66067 48427
rect 65757 30587 66067 48309
rect 65757 30469 65773 30587
rect 65891 30469 65933 30587
rect 66051 30469 66067 30587
rect 65757 30427 66067 30469
rect 65757 30309 65773 30427
rect 65891 30309 65933 30427
rect 66051 30309 66067 30427
rect 65757 12587 66067 30309
rect 65757 12469 65773 12587
rect 65891 12469 65933 12587
rect 66051 12469 66067 12587
rect 65757 12427 66067 12469
rect 65757 12309 65773 12427
rect 65891 12309 65933 12427
rect 66051 12309 66067 12427
rect 65757 -1613 66067 12309
rect 65757 -1731 65773 -1613
rect 65891 -1731 65933 -1613
rect 66051 -1731 66067 -1613
rect 65757 -1773 66067 -1731
rect 65757 -1891 65773 -1773
rect 65891 -1891 65933 -1773
rect 66051 -1891 66067 -1773
rect 65757 -1907 66067 -1891
rect 67617 338447 67927 354541
rect 67617 338329 67633 338447
rect 67751 338329 67793 338447
rect 67911 338329 67927 338447
rect 67617 338287 67927 338329
rect 67617 338169 67633 338287
rect 67751 338169 67793 338287
rect 67911 338169 67927 338287
rect 67617 320447 67927 338169
rect 67617 320329 67633 320447
rect 67751 320329 67793 320447
rect 67911 320329 67927 320447
rect 67617 320287 67927 320329
rect 67617 320169 67633 320287
rect 67751 320169 67793 320287
rect 67911 320169 67927 320287
rect 67617 302447 67927 320169
rect 67617 302329 67633 302447
rect 67751 302329 67793 302447
rect 67911 302329 67927 302447
rect 67617 302287 67927 302329
rect 67617 302169 67633 302287
rect 67751 302169 67793 302287
rect 67911 302169 67927 302287
rect 67617 284447 67927 302169
rect 67617 284329 67633 284447
rect 67751 284329 67793 284447
rect 67911 284329 67927 284447
rect 67617 284287 67927 284329
rect 67617 284169 67633 284287
rect 67751 284169 67793 284287
rect 67911 284169 67927 284287
rect 67617 266447 67927 284169
rect 67617 266329 67633 266447
rect 67751 266329 67793 266447
rect 67911 266329 67927 266447
rect 67617 266287 67927 266329
rect 67617 266169 67633 266287
rect 67751 266169 67793 266287
rect 67911 266169 67927 266287
rect 67617 248447 67927 266169
rect 67617 248329 67633 248447
rect 67751 248329 67793 248447
rect 67911 248329 67927 248447
rect 67617 248287 67927 248329
rect 67617 248169 67633 248287
rect 67751 248169 67793 248287
rect 67911 248169 67927 248287
rect 67617 230447 67927 248169
rect 67617 230329 67633 230447
rect 67751 230329 67793 230447
rect 67911 230329 67927 230447
rect 67617 230287 67927 230329
rect 67617 230169 67633 230287
rect 67751 230169 67793 230287
rect 67911 230169 67927 230287
rect 67617 212447 67927 230169
rect 67617 212329 67633 212447
rect 67751 212329 67793 212447
rect 67911 212329 67927 212447
rect 67617 212287 67927 212329
rect 67617 212169 67633 212287
rect 67751 212169 67793 212287
rect 67911 212169 67927 212287
rect 67617 194447 67927 212169
rect 67617 194329 67633 194447
rect 67751 194329 67793 194447
rect 67911 194329 67927 194447
rect 67617 194287 67927 194329
rect 67617 194169 67633 194287
rect 67751 194169 67793 194287
rect 67911 194169 67927 194287
rect 67617 176447 67927 194169
rect 67617 176329 67633 176447
rect 67751 176329 67793 176447
rect 67911 176329 67927 176447
rect 67617 176287 67927 176329
rect 67617 176169 67633 176287
rect 67751 176169 67793 176287
rect 67911 176169 67927 176287
rect 67617 158447 67927 176169
rect 67617 158329 67633 158447
rect 67751 158329 67793 158447
rect 67911 158329 67927 158447
rect 67617 158287 67927 158329
rect 67617 158169 67633 158287
rect 67751 158169 67793 158287
rect 67911 158169 67927 158287
rect 67617 140447 67927 158169
rect 67617 140329 67633 140447
rect 67751 140329 67793 140447
rect 67911 140329 67927 140447
rect 67617 140287 67927 140329
rect 67617 140169 67633 140287
rect 67751 140169 67793 140287
rect 67911 140169 67927 140287
rect 67617 122447 67927 140169
rect 67617 122329 67633 122447
rect 67751 122329 67793 122447
rect 67911 122329 67927 122447
rect 67617 122287 67927 122329
rect 67617 122169 67633 122287
rect 67751 122169 67793 122287
rect 67911 122169 67927 122287
rect 67617 104447 67927 122169
rect 67617 104329 67633 104447
rect 67751 104329 67793 104447
rect 67911 104329 67927 104447
rect 67617 104287 67927 104329
rect 67617 104169 67633 104287
rect 67751 104169 67793 104287
rect 67911 104169 67927 104287
rect 67617 86447 67927 104169
rect 67617 86329 67633 86447
rect 67751 86329 67793 86447
rect 67911 86329 67927 86447
rect 67617 86287 67927 86329
rect 67617 86169 67633 86287
rect 67751 86169 67793 86287
rect 67911 86169 67927 86287
rect 67617 68447 67927 86169
rect 67617 68329 67633 68447
rect 67751 68329 67793 68447
rect 67911 68329 67927 68447
rect 67617 68287 67927 68329
rect 67617 68169 67633 68287
rect 67751 68169 67793 68287
rect 67911 68169 67927 68287
rect 67617 50447 67927 68169
rect 67617 50329 67633 50447
rect 67751 50329 67793 50447
rect 67911 50329 67927 50447
rect 67617 50287 67927 50329
rect 67617 50169 67633 50287
rect 67751 50169 67793 50287
rect 67911 50169 67927 50287
rect 67617 32447 67927 50169
rect 67617 32329 67633 32447
rect 67751 32329 67793 32447
rect 67911 32329 67927 32447
rect 67617 32287 67927 32329
rect 67617 32169 67633 32287
rect 67751 32169 67793 32287
rect 67911 32169 67927 32287
rect 67617 14447 67927 32169
rect 67617 14329 67633 14447
rect 67751 14329 67793 14447
rect 67911 14329 67927 14447
rect 67617 14287 67927 14329
rect 67617 14169 67633 14287
rect 67751 14169 67793 14287
rect 67911 14169 67927 14287
rect 67617 -2573 67927 14169
rect 67617 -2691 67633 -2573
rect 67751 -2691 67793 -2573
rect 67911 -2691 67927 -2573
rect 67617 -2733 67927 -2691
rect 67617 -2851 67633 -2733
rect 67751 -2851 67793 -2733
rect 67911 -2851 67927 -2733
rect 67617 -2867 67927 -2851
rect 69477 340307 69787 355501
rect 78477 355299 78787 355795
rect 78477 355181 78493 355299
rect 78611 355181 78653 355299
rect 78771 355181 78787 355299
rect 78477 355139 78787 355181
rect 78477 355021 78493 355139
rect 78611 355021 78653 355139
rect 78771 355021 78787 355139
rect 76617 354339 76927 354835
rect 76617 354221 76633 354339
rect 76751 354221 76793 354339
rect 76911 354221 76927 354339
rect 76617 354179 76927 354221
rect 76617 354061 76633 354179
rect 76751 354061 76793 354179
rect 76911 354061 76927 354179
rect 74757 353379 75067 353875
rect 74757 353261 74773 353379
rect 74891 353261 74933 353379
rect 75051 353261 75067 353379
rect 74757 353219 75067 353261
rect 74757 353101 74773 353219
rect 74891 353101 74933 353219
rect 75051 353101 75067 353219
rect 69477 340189 69493 340307
rect 69611 340189 69653 340307
rect 69771 340189 69787 340307
rect 69477 340147 69787 340189
rect 69477 340029 69493 340147
rect 69611 340029 69653 340147
rect 69771 340029 69787 340147
rect 69477 322307 69787 340029
rect 69477 322189 69493 322307
rect 69611 322189 69653 322307
rect 69771 322189 69787 322307
rect 69477 322147 69787 322189
rect 69477 322029 69493 322147
rect 69611 322029 69653 322147
rect 69771 322029 69787 322147
rect 69477 304307 69787 322029
rect 69477 304189 69493 304307
rect 69611 304189 69653 304307
rect 69771 304189 69787 304307
rect 69477 304147 69787 304189
rect 69477 304029 69493 304147
rect 69611 304029 69653 304147
rect 69771 304029 69787 304147
rect 69477 286307 69787 304029
rect 69477 286189 69493 286307
rect 69611 286189 69653 286307
rect 69771 286189 69787 286307
rect 69477 286147 69787 286189
rect 69477 286029 69493 286147
rect 69611 286029 69653 286147
rect 69771 286029 69787 286147
rect 69477 268307 69787 286029
rect 69477 268189 69493 268307
rect 69611 268189 69653 268307
rect 69771 268189 69787 268307
rect 69477 268147 69787 268189
rect 69477 268029 69493 268147
rect 69611 268029 69653 268147
rect 69771 268029 69787 268147
rect 69477 250307 69787 268029
rect 69477 250189 69493 250307
rect 69611 250189 69653 250307
rect 69771 250189 69787 250307
rect 69477 250147 69787 250189
rect 69477 250029 69493 250147
rect 69611 250029 69653 250147
rect 69771 250029 69787 250147
rect 69477 232307 69787 250029
rect 69477 232189 69493 232307
rect 69611 232189 69653 232307
rect 69771 232189 69787 232307
rect 69477 232147 69787 232189
rect 69477 232029 69493 232147
rect 69611 232029 69653 232147
rect 69771 232029 69787 232147
rect 69477 214307 69787 232029
rect 69477 214189 69493 214307
rect 69611 214189 69653 214307
rect 69771 214189 69787 214307
rect 69477 214147 69787 214189
rect 69477 214029 69493 214147
rect 69611 214029 69653 214147
rect 69771 214029 69787 214147
rect 69477 196307 69787 214029
rect 69477 196189 69493 196307
rect 69611 196189 69653 196307
rect 69771 196189 69787 196307
rect 69477 196147 69787 196189
rect 69477 196029 69493 196147
rect 69611 196029 69653 196147
rect 69771 196029 69787 196147
rect 69477 178307 69787 196029
rect 69477 178189 69493 178307
rect 69611 178189 69653 178307
rect 69771 178189 69787 178307
rect 69477 178147 69787 178189
rect 69477 178029 69493 178147
rect 69611 178029 69653 178147
rect 69771 178029 69787 178147
rect 69477 160307 69787 178029
rect 69477 160189 69493 160307
rect 69611 160189 69653 160307
rect 69771 160189 69787 160307
rect 69477 160147 69787 160189
rect 69477 160029 69493 160147
rect 69611 160029 69653 160147
rect 69771 160029 69787 160147
rect 69477 142307 69787 160029
rect 69477 142189 69493 142307
rect 69611 142189 69653 142307
rect 69771 142189 69787 142307
rect 69477 142147 69787 142189
rect 69477 142029 69493 142147
rect 69611 142029 69653 142147
rect 69771 142029 69787 142147
rect 69477 124307 69787 142029
rect 69477 124189 69493 124307
rect 69611 124189 69653 124307
rect 69771 124189 69787 124307
rect 69477 124147 69787 124189
rect 69477 124029 69493 124147
rect 69611 124029 69653 124147
rect 69771 124029 69787 124147
rect 69477 106307 69787 124029
rect 69477 106189 69493 106307
rect 69611 106189 69653 106307
rect 69771 106189 69787 106307
rect 69477 106147 69787 106189
rect 69477 106029 69493 106147
rect 69611 106029 69653 106147
rect 69771 106029 69787 106147
rect 69477 88307 69787 106029
rect 69477 88189 69493 88307
rect 69611 88189 69653 88307
rect 69771 88189 69787 88307
rect 69477 88147 69787 88189
rect 69477 88029 69493 88147
rect 69611 88029 69653 88147
rect 69771 88029 69787 88147
rect 69477 70307 69787 88029
rect 69477 70189 69493 70307
rect 69611 70189 69653 70307
rect 69771 70189 69787 70307
rect 69477 70147 69787 70189
rect 69477 70029 69493 70147
rect 69611 70029 69653 70147
rect 69771 70029 69787 70147
rect 69477 52307 69787 70029
rect 69477 52189 69493 52307
rect 69611 52189 69653 52307
rect 69771 52189 69787 52307
rect 69477 52147 69787 52189
rect 69477 52029 69493 52147
rect 69611 52029 69653 52147
rect 69771 52029 69787 52147
rect 69477 34307 69787 52029
rect 69477 34189 69493 34307
rect 69611 34189 69653 34307
rect 69771 34189 69787 34307
rect 69477 34147 69787 34189
rect 69477 34029 69493 34147
rect 69611 34029 69653 34147
rect 69771 34029 69787 34147
rect 69477 16307 69787 34029
rect 69477 16189 69493 16307
rect 69611 16189 69653 16307
rect 69771 16189 69787 16307
rect 69477 16147 69787 16189
rect 69477 16029 69493 16147
rect 69611 16029 69653 16147
rect 69771 16029 69787 16147
rect 60477 -3171 60493 -3053
rect 60611 -3171 60653 -3053
rect 60771 -3171 60787 -3053
rect 60477 -3213 60787 -3171
rect 60477 -3331 60493 -3213
rect 60611 -3331 60653 -3213
rect 60771 -3331 60787 -3213
rect 60477 -3827 60787 -3331
rect 69477 -3533 69787 16029
rect 72897 352419 73207 352915
rect 72897 352301 72913 352419
rect 73031 352301 73073 352419
rect 73191 352301 73207 352419
rect 72897 352259 73207 352301
rect 72897 352141 72913 352259
rect 73031 352141 73073 352259
rect 73191 352141 73207 352259
rect 72897 343727 73207 352141
rect 72897 343609 72913 343727
rect 73031 343609 73073 343727
rect 73191 343609 73207 343727
rect 72897 343567 73207 343609
rect 72897 343449 72913 343567
rect 73031 343449 73073 343567
rect 73191 343449 73207 343567
rect 72897 325727 73207 343449
rect 72897 325609 72913 325727
rect 73031 325609 73073 325727
rect 73191 325609 73207 325727
rect 72897 325567 73207 325609
rect 72897 325449 72913 325567
rect 73031 325449 73073 325567
rect 73191 325449 73207 325567
rect 72897 307727 73207 325449
rect 72897 307609 72913 307727
rect 73031 307609 73073 307727
rect 73191 307609 73207 307727
rect 72897 307567 73207 307609
rect 72897 307449 72913 307567
rect 73031 307449 73073 307567
rect 73191 307449 73207 307567
rect 72897 289727 73207 307449
rect 72897 289609 72913 289727
rect 73031 289609 73073 289727
rect 73191 289609 73207 289727
rect 72897 289567 73207 289609
rect 72897 289449 72913 289567
rect 73031 289449 73073 289567
rect 73191 289449 73207 289567
rect 72897 271727 73207 289449
rect 72897 271609 72913 271727
rect 73031 271609 73073 271727
rect 73191 271609 73207 271727
rect 72897 271567 73207 271609
rect 72897 271449 72913 271567
rect 73031 271449 73073 271567
rect 73191 271449 73207 271567
rect 72897 253727 73207 271449
rect 72897 253609 72913 253727
rect 73031 253609 73073 253727
rect 73191 253609 73207 253727
rect 72897 253567 73207 253609
rect 72897 253449 72913 253567
rect 73031 253449 73073 253567
rect 73191 253449 73207 253567
rect 72897 235727 73207 253449
rect 72897 235609 72913 235727
rect 73031 235609 73073 235727
rect 73191 235609 73207 235727
rect 72897 235567 73207 235609
rect 72897 235449 72913 235567
rect 73031 235449 73073 235567
rect 73191 235449 73207 235567
rect 72897 217727 73207 235449
rect 72897 217609 72913 217727
rect 73031 217609 73073 217727
rect 73191 217609 73207 217727
rect 72897 217567 73207 217609
rect 72897 217449 72913 217567
rect 73031 217449 73073 217567
rect 73191 217449 73207 217567
rect 72897 199727 73207 217449
rect 72897 199609 72913 199727
rect 73031 199609 73073 199727
rect 73191 199609 73207 199727
rect 72897 199567 73207 199609
rect 72897 199449 72913 199567
rect 73031 199449 73073 199567
rect 73191 199449 73207 199567
rect 72897 181727 73207 199449
rect 72897 181609 72913 181727
rect 73031 181609 73073 181727
rect 73191 181609 73207 181727
rect 72897 181567 73207 181609
rect 72897 181449 72913 181567
rect 73031 181449 73073 181567
rect 73191 181449 73207 181567
rect 72897 163727 73207 181449
rect 72897 163609 72913 163727
rect 73031 163609 73073 163727
rect 73191 163609 73207 163727
rect 72897 163567 73207 163609
rect 72897 163449 72913 163567
rect 73031 163449 73073 163567
rect 73191 163449 73207 163567
rect 72897 145727 73207 163449
rect 72897 145609 72913 145727
rect 73031 145609 73073 145727
rect 73191 145609 73207 145727
rect 72897 145567 73207 145609
rect 72897 145449 72913 145567
rect 73031 145449 73073 145567
rect 73191 145449 73207 145567
rect 72897 127727 73207 145449
rect 72897 127609 72913 127727
rect 73031 127609 73073 127727
rect 73191 127609 73207 127727
rect 72897 127567 73207 127609
rect 72897 127449 72913 127567
rect 73031 127449 73073 127567
rect 73191 127449 73207 127567
rect 72897 109727 73207 127449
rect 72897 109609 72913 109727
rect 73031 109609 73073 109727
rect 73191 109609 73207 109727
rect 72897 109567 73207 109609
rect 72897 109449 72913 109567
rect 73031 109449 73073 109567
rect 73191 109449 73207 109567
rect 72897 91727 73207 109449
rect 72897 91609 72913 91727
rect 73031 91609 73073 91727
rect 73191 91609 73207 91727
rect 72897 91567 73207 91609
rect 72897 91449 72913 91567
rect 73031 91449 73073 91567
rect 73191 91449 73207 91567
rect 72897 73727 73207 91449
rect 72897 73609 72913 73727
rect 73031 73609 73073 73727
rect 73191 73609 73207 73727
rect 72897 73567 73207 73609
rect 72897 73449 72913 73567
rect 73031 73449 73073 73567
rect 73191 73449 73207 73567
rect 72897 55727 73207 73449
rect 72897 55609 72913 55727
rect 73031 55609 73073 55727
rect 73191 55609 73207 55727
rect 72897 55567 73207 55609
rect 72897 55449 72913 55567
rect 73031 55449 73073 55567
rect 73191 55449 73207 55567
rect 72897 37727 73207 55449
rect 72897 37609 72913 37727
rect 73031 37609 73073 37727
rect 73191 37609 73207 37727
rect 72897 37567 73207 37609
rect 72897 37449 72913 37567
rect 73031 37449 73073 37567
rect 73191 37449 73207 37567
rect 72897 19727 73207 37449
rect 72897 19609 72913 19727
rect 73031 19609 73073 19727
rect 73191 19609 73207 19727
rect 72897 19567 73207 19609
rect 72897 19449 72913 19567
rect 73031 19449 73073 19567
rect 73191 19449 73207 19567
rect 72897 1727 73207 19449
rect 72897 1609 72913 1727
rect 73031 1609 73073 1727
rect 73191 1609 73207 1727
rect 72897 1567 73207 1609
rect 72897 1449 72913 1567
rect 73031 1449 73073 1567
rect 73191 1449 73207 1567
rect 72897 -173 73207 1449
rect 72897 -291 72913 -173
rect 73031 -291 73073 -173
rect 73191 -291 73207 -173
rect 72897 -333 73207 -291
rect 72897 -451 72913 -333
rect 73031 -451 73073 -333
rect 73191 -451 73207 -333
rect 72897 -947 73207 -451
rect 74757 345587 75067 353101
rect 74757 345469 74773 345587
rect 74891 345469 74933 345587
rect 75051 345469 75067 345587
rect 74757 345427 75067 345469
rect 74757 345309 74773 345427
rect 74891 345309 74933 345427
rect 75051 345309 75067 345427
rect 74757 327587 75067 345309
rect 74757 327469 74773 327587
rect 74891 327469 74933 327587
rect 75051 327469 75067 327587
rect 74757 327427 75067 327469
rect 74757 327309 74773 327427
rect 74891 327309 74933 327427
rect 75051 327309 75067 327427
rect 74757 309587 75067 327309
rect 74757 309469 74773 309587
rect 74891 309469 74933 309587
rect 75051 309469 75067 309587
rect 74757 309427 75067 309469
rect 74757 309309 74773 309427
rect 74891 309309 74933 309427
rect 75051 309309 75067 309427
rect 74757 291587 75067 309309
rect 74757 291469 74773 291587
rect 74891 291469 74933 291587
rect 75051 291469 75067 291587
rect 74757 291427 75067 291469
rect 74757 291309 74773 291427
rect 74891 291309 74933 291427
rect 75051 291309 75067 291427
rect 74757 273587 75067 291309
rect 74757 273469 74773 273587
rect 74891 273469 74933 273587
rect 75051 273469 75067 273587
rect 74757 273427 75067 273469
rect 74757 273309 74773 273427
rect 74891 273309 74933 273427
rect 75051 273309 75067 273427
rect 74757 255587 75067 273309
rect 74757 255469 74773 255587
rect 74891 255469 74933 255587
rect 75051 255469 75067 255587
rect 74757 255427 75067 255469
rect 74757 255309 74773 255427
rect 74891 255309 74933 255427
rect 75051 255309 75067 255427
rect 74757 237587 75067 255309
rect 74757 237469 74773 237587
rect 74891 237469 74933 237587
rect 75051 237469 75067 237587
rect 74757 237427 75067 237469
rect 74757 237309 74773 237427
rect 74891 237309 74933 237427
rect 75051 237309 75067 237427
rect 74757 219587 75067 237309
rect 74757 219469 74773 219587
rect 74891 219469 74933 219587
rect 75051 219469 75067 219587
rect 74757 219427 75067 219469
rect 74757 219309 74773 219427
rect 74891 219309 74933 219427
rect 75051 219309 75067 219427
rect 74757 201587 75067 219309
rect 74757 201469 74773 201587
rect 74891 201469 74933 201587
rect 75051 201469 75067 201587
rect 74757 201427 75067 201469
rect 74757 201309 74773 201427
rect 74891 201309 74933 201427
rect 75051 201309 75067 201427
rect 74757 183587 75067 201309
rect 74757 183469 74773 183587
rect 74891 183469 74933 183587
rect 75051 183469 75067 183587
rect 74757 183427 75067 183469
rect 74757 183309 74773 183427
rect 74891 183309 74933 183427
rect 75051 183309 75067 183427
rect 74757 165587 75067 183309
rect 74757 165469 74773 165587
rect 74891 165469 74933 165587
rect 75051 165469 75067 165587
rect 74757 165427 75067 165469
rect 74757 165309 74773 165427
rect 74891 165309 74933 165427
rect 75051 165309 75067 165427
rect 74757 147587 75067 165309
rect 74757 147469 74773 147587
rect 74891 147469 74933 147587
rect 75051 147469 75067 147587
rect 74757 147427 75067 147469
rect 74757 147309 74773 147427
rect 74891 147309 74933 147427
rect 75051 147309 75067 147427
rect 74757 129587 75067 147309
rect 74757 129469 74773 129587
rect 74891 129469 74933 129587
rect 75051 129469 75067 129587
rect 74757 129427 75067 129469
rect 74757 129309 74773 129427
rect 74891 129309 74933 129427
rect 75051 129309 75067 129427
rect 74757 111587 75067 129309
rect 74757 111469 74773 111587
rect 74891 111469 74933 111587
rect 75051 111469 75067 111587
rect 74757 111427 75067 111469
rect 74757 111309 74773 111427
rect 74891 111309 74933 111427
rect 75051 111309 75067 111427
rect 74757 93587 75067 111309
rect 74757 93469 74773 93587
rect 74891 93469 74933 93587
rect 75051 93469 75067 93587
rect 74757 93427 75067 93469
rect 74757 93309 74773 93427
rect 74891 93309 74933 93427
rect 75051 93309 75067 93427
rect 74757 75587 75067 93309
rect 74757 75469 74773 75587
rect 74891 75469 74933 75587
rect 75051 75469 75067 75587
rect 74757 75427 75067 75469
rect 74757 75309 74773 75427
rect 74891 75309 74933 75427
rect 75051 75309 75067 75427
rect 74757 57587 75067 75309
rect 74757 57469 74773 57587
rect 74891 57469 74933 57587
rect 75051 57469 75067 57587
rect 74757 57427 75067 57469
rect 74757 57309 74773 57427
rect 74891 57309 74933 57427
rect 75051 57309 75067 57427
rect 74757 39587 75067 57309
rect 74757 39469 74773 39587
rect 74891 39469 74933 39587
rect 75051 39469 75067 39587
rect 74757 39427 75067 39469
rect 74757 39309 74773 39427
rect 74891 39309 74933 39427
rect 75051 39309 75067 39427
rect 74757 21587 75067 39309
rect 74757 21469 74773 21587
rect 74891 21469 74933 21587
rect 75051 21469 75067 21587
rect 74757 21427 75067 21469
rect 74757 21309 74773 21427
rect 74891 21309 74933 21427
rect 75051 21309 75067 21427
rect 74757 3587 75067 21309
rect 74757 3469 74773 3587
rect 74891 3469 74933 3587
rect 75051 3469 75067 3587
rect 74757 3427 75067 3469
rect 74757 3309 74773 3427
rect 74891 3309 74933 3427
rect 75051 3309 75067 3427
rect 74757 -1133 75067 3309
rect 74757 -1251 74773 -1133
rect 74891 -1251 74933 -1133
rect 75051 -1251 75067 -1133
rect 74757 -1293 75067 -1251
rect 74757 -1411 74773 -1293
rect 74891 -1411 74933 -1293
rect 75051 -1411 75067 -1293
rect 74757 -1907 75067 -1411
rect 76617 347447 76927 354061
rect 76617 347329 76633 347447
rect 76751 347329 76793 347447
rect 76911 347329 76927 347447
rect 76617 347287 76927 347329
rect 76617 347169 76633 347287
rect 76751 347169 76793 347287
rect 76911 347169 76927 347287
rect 76617 329447 76927 347169
rect 76617 329329 76633 329447
rect 76751 329329 76793 329447
rect 76911 329329 76927 329447
rect 76617 329287 76927 329329
rect 76617 329169 76633 329287
rect 76751 329169 76793 329287
rect 76911 329169 76927 329287
rect 76617 311447 76927 329169
rect 76617 311329 76633 311447
rect 76751 311329 76793 311447
rect 76911 311329 76927 311447
rect 76617 311287 76927 311329
rect 76617 311169 76633 311287
rect 76751 311169 76793 311287
rect 76911 311169 76927 311287
rect 76617 293447 76927 311169
rect 76617 293329 76633 293447
rect 76751 293329 76793 293447
rect 76911 293329 76927 293447
rect 76617 293287 76927 293329
rect 76617 293169 76633 293287
rect 76751 293169 76793 293287
rect 76911 293169 76927 293287
rect 76617 275447 76927 293169
rect 76617 275329 76633 275447
rect 76751 275329 76793 275447
rect 76911 275329 76927 275447
rect 76617 275287 76927 275329
rect 76617 275169 76633 275287
rect 76751 275169 76793 275287
rect 76911 275169 76927 275287
rect 76617 257447 76927 275169
rect 76617 257329 76633 257447
rect 76751 257329 76793 257447
rect 76911 257329 76927 257447
rect 76617 257287 76927 257329
rect 76617 257169 76633 257287
rect 76751 257169 76793 257287
rect 76911 257169 76927 257287
rect 76617 239447 76927 257169
rect 76617 239329 76633 239447
rect 76751 239329 76793 239447
rect 76911 239329 76927 239447
rect 76617 239287 76927 239329
rect 76617 239169 76633 239287
rect 76751 239169 76793 239287
rect 76911 239169 76927 239287
rect 76617 221447 76927 239169
rect 76617 221329 76633 221447
rect 76751 221329 76793 221447
rect 76911 221329 76927 221447
rect 76617 221287 76927 221329
rect 76617 221169 76633 221287
rect 76751 221169 76793 221287
rect 76911 221169 76927 221287
rect 76617 203447 76927 221169
rect 76617 203329 76633 203447
rect 76751 203329 76793 203447
rect 76911 203329 76927 203447
rect 76617 203287 76927 203329
rect 76617 203169 76633 203287
rect 76751 203169 76793 203287
rect 76911 203169 76927 203287
rect 76617 185447 76927 203169
rect 76617 185329 76633 185447
rect 76751 185329 76793 185447
rect 76911 185329 76927 185447
rect 76617 185287 76927 185329
rect 76617 185169 76633 185287
rect 76751 185169 76793 185287
rect 76911 185169 76927 185287
rect 76617 167447 76927 185169
rect 76617 167329 76633 167447
rect 76751 167329 76793 167447
rect 76911 167329 76927 167447
rect 76617 167287 76927 167329
rect 76617 167169 76633 167287
rect 76751 167169 76793 167287
rect 76911 167169 76927 167287
rect 76617 149447 76927 167169
rect 76617 149329 76633 149447
rect 76751 149329 76793 149447
rect 76911 149329 76927 149447
rect 76617 149287 76927 149329
rect 76617 149169 76633 149287
rect 76751 149169 76793 149287
rect 76911 149169 76927 149287
rect 76617 131447 76927 149169
rect 76617 131329 76633 131447
rect 76751 131329 76793 131447
rect 76911 131329 76927 131447
rect 76617 131287 76927 131329
rect 76617 131169 76633 131287
rect 76751 131169 76793 131287
rect 76911 131169 76927 131287
rect 76617 113447 76927 131169
rect 76617 113329 76633 113447
rect 76751 113329 76793 113447
rect 76911 113329 76927 113447
rect 76617 113287 76927 113329
rect 76617 113169 76633 113287
rect 76751 113169 76793 113287
rect 76911 113169 76927 113287
rect 76617 95447 76927 113169
rect 76617 95329 76633 95447
rect 76751 95329 76793 95447
rect 76911 95329 76927 95447
rect 76617 95287 76927 95329
rect 76617 95169 76633 95287
rect 76751 95169 76793 95287
rect 76911 95169 76927 95287
rect 76617 77447 76927 95169
rect 76617 77329 76633 77447
rect 76751 77329 76793 77447
rect 76911 77329 76927 77447
rect 76617 77287 76927 77329
rect 76617 77169 76633 77287
rect 76751 77169 76793 77287
rect 76911 77169 76927 77287
rect 76617 59447 76927 77169
rect 76617 59329 76633 59447
rect 76751 59329 76793 59447
rect 76911 59329 76927 59447
rect 76617 59287 76927 59329
rect 76617 59169 76633 59287
rect 76751 59169 76793 59287
rect 76911 59169 76927 59287
rect 76617 41447 76927 59169
rect 76617 41329 76633 41447
rect 76751 41329 76793 41447
rect 76911 41329 76927 41447
rect 76617 41287 76927 41329
rect 76617 41169 76633 41287
rect 76751 41169 76793 41287
rect 76911 41169 76927 41287
rect 76617 23447 76927 41169
rect 76617 23329 76633 23447
rect 76751 23329 76793 23447
rect 76911 23329 76927 23447
rect 76617 23287 76927 23329
rect 76617 23169 76633 23287
rect 76751 23169 76793 23287
rect 76911 23169 76927 23287
rect 76617 5447 76927 23169
rect 76617 5329 76633 5447
rect 76751 5329 76793 5447
rect 76911 5329 76927 5447
rect 76617 5287 76927 5329
rect 76617 5169 76633 5287
rect 76751 5169 76793 5287
rect 76911 5169 76927 5287
rect 76617 -2093 76927 5169
rect 76617 -2211 76633 -2093
rect 76751 -2211 76793 -2093
rect 76911 -2211 76927 -2093
rect 76617 -2253 76927 -2211
rect 76617 -2371 76633 -2253
rect 76751 -2371 76793 -2253
rect 76911 -2371 76927 -2253
rect 76617 -2867 76927 -2371
rect 78477 349307 78787 355021
rect 87477 355779 87787 355795
rect 87477 355661 87493 355779
rect 87611 355661 87653 355779
rect 87771 355661 87787 355779
rect 87477 355619 87787 355661
rect 87477 355501 87493 355619
rect 87611 355501 87653 355619
rect 87771 355501 87787 355619
rect 85617 354819 85927 354835
rect 85617 354701 85633 354819
rect 85751 354701 85793 354819
rect 85911 354701 85927 354819
rect 85617 354659 85927 354701
rect 85617 354541 85633 354659
rect 85751 354541 85793 354659
rect 85911 354541 85927 354659
rect 83757 353859 84067 353875
rect 83757 353741 83773 353859
rect 83891 353741 83933 353859
rect 84051 353741 84067 353859
rect 83757 353699 84067 353741
rect 83757 353581 83773 353699
rect 83891 353581 83933 353699
rect 84051 353581 84067 353699
rect 78477 349189 78493 349307
rect 78611 349189 78653 349307
rect 78771 349189 78787 349307
rect 78477 349147 78787 349189
rect 78477 349029 78493 349147
rect 78611 349029 78653 349147
rect 78771 349029 78787 349147
rect 78477 331307 78787 349029
rect 78477 331189 78493 331307
rect 78611 331189 78653 331307
rect 78771 331189 78787 331307
rect 78477 331147 78787 331189
rect 78477 331029 78493 331147
rect 78611 331029 78653 331147
rect 78771 331029 78787 331147
rect 78477 313307 78787 331029
rect 78477 313189 78493 313307
rect 78611 313189 78653 313307
rect 78771 313189 78787 313307
rect 78477 313147 78787 313189
rect 78477 313029 78493 313147
rect 78611 313029 78653 313147
rect 78771 313029 78787 313147
rect 78477 295307 78787 313029
rect 78477 295189 78493 295307
rect 78611 295189 78653 295307
rect 78771 295189 78787 295307
rect 78477 295147 78787 295189
rect 78477 295029 78493 295147
rect 78611 295029 78653 295147
rect 78771 295029 78787 295147
rect 78477 277307 78787 295029
rect 78477 277189 78493 277307
rect 78611 277189 78653 277307
rect 78771 277189 78787 277307
rect 78477 277147 78787 277189
rect 78477 277029 78493 277147
rect 78611 277029 78653 277147
rect 78771 277029 78787 277147
rect 78477 259307 78787 277029
rect 78477 259189 78493 259307
rect 78611 259189 78653 259307
rect 78771 259189 78787 259307
rect 78477 259147 78787 259189
rect 78477 259029 78493 259147
rect 78611 259029 78653 259147
rect 78771 259029 78787 259147
rect 78477 241307 78787 259029
rect 78477 241189 78493 241307
rect 78611 241189 78653 241307
rect 78771 241189 78787 241307
rect 78477 241147 78787 241189
rect 78477 241029 78493 241147
rect 78611 241029 78653 241147
rect 78771 241029 78787 241147
rect 78477 223307 78787 241029
rect 78477 223189 78493 223307
rect 78611 223189 78653 223307
rect 78771 223189 78787 223307
rect 78477 223147 78787 223189
rect 78477 223029 78493 223147
rect 78611 223029 78653 223147
rect 78771 223029 78787 223147
rect 78477 205307 78787 223029
rect 78477 205189 78493 205307
rect 78611 205189 78653 205307
rect 78771 205189 78787 205307
rect 78477 205147 78787 205189
rect 78477 205029 78493 205147
rect 78611 205029 78653 205147
rect 78771 205029 78787 205147
rect 78477 187307 78787 205029
rect 78477 187189 78493 187307
rect 78611 187189 78653 187307
rect 78771 187189 78787 187307
rect 78477 187147 78787 187189
rect 78477 187029 78493 187147
rect 78611 187029 78653 187147
rect 78771 187029 78787 187147
rect 78477 169307 78787 187029
rect 78477 169189 78493 169307
rect 78611 169189 78653 169307
rect 78771 169189 78787 169307
rect 78477 169147 78787 169189
rect 78477 169029 78493 169147
rect 78611 169029 78653 169147
rect 78771 169029 78787 169147
rect 78477 151307 78787 169029
rect 78477 151189 78493 151307
rect 78611 151189 78653 151307
rect 78771 151189 78787 151307
rect 78477 151147 78787 151189
rect 78477 151029 78493 151147
rect 78611 151029 78653 151147
rect 78771 151029 78787 151147
rect 78477 133307 78787 151029
rect 78477 133189 78493 133307
rect 78611 133189 78653 133307
rect 78771 133189 78787 133307
rect 78477 133147 78787 133189
rect 78477 133029 78493 133147
rect 78611 133029 78653 133147
rect 78771 133029 78787 133147
rect 78477 115307 78787 133029
rect 78477 115189 78493 115307
rect 78611 115189 78653 115307
rect 78771 115189 78787 115307
rect 78477 115147 78787 115189
rect 78477 115029 78493 115147
rect 78611 115029 78653 115147
rect 78771 115029 78787 115147
rect 78477 97307 78787 115029
rect 78477 97189 78493 97307
rect 78611 97189 78653 97307
rect 78771 97189 78787 97307
rect 78477 97147 78787 97189
rect 78477 97029 78493 97147
rect 78611 97029 78653 97147
rect 78771 97029 78787 97147
rect 78477 79307 78787 97029
rect 78477 79189 78493 79307
rect 78611 79189 78653 79307
rect 78771 79189 78787 79307
rect 78477 79147 78787 79189
rect 78477 79029 78493 79147
rect 78611 79029 78653 79147
rect 78771 79029 78787 79147
rect 78477 61307 78787 79029
rect 78477 61189 78493 61307
rect 78611 61189 78653 61307
rect 78771 61189 78787 61307
rect 78477 61147 78787 61189
rect 78477 61029 78493 61147
rect 78611 61029 78653 61147
rect 78771 61029 78787 61147
rect 78477 43307 78787 61029
rect 78477 43189 78493 43307
rect 78611 43189 78653 43307
rect 78771 43189 78787 43307
rect 78477 43147 78787 43189
rect 78477 43029 78493 43147
rect 78611 43029 78653 43147
rect 78771 43029 78787 43147
rect 78477 25307 78787 43029
rect 78477 25189 78493 25307
rect 78611 25189 78653 25307
rect 78771 25189 78787 25307
rect 78477 25147 78787 25189
rect 78477 25029 78493 25147
rect 78611 25029 78653 25147
rect 78771 25029 78787 25147
rect 78477 7307 78787 25029
rect 78477 7189 78493 7307
rect 78611 7189 78653 7307
rect 78771 7189 78787 7307
rect 78477 7147 78787 7189
rect 78477 7029 78493 7147
rect 78611 7029 78653 7147
rect 78771 7029 78787 7147
rect 69477 -3651 69493 -3533
rect 69611 -3651 69653 -3533
rect 69771 -3651 69787 -3533
rect 69477 -3693 69787 -3651
rect 69477 -3811 69493 -3693
rect 69611 -3811 69653 -3693
rect 69771 -3811 69787 -3693
rect 69477 -3827 69787 -3811
rect 78477 -3053 78787 7029
rect 81897 352899 82207 352915
rect 81897 352781 81913 352899
rect 82031 352781 82073 352899
rect 82191 352781 82207 352899
rect 81897 352739 82207 352781
rect 81897 352621 81913 352739
rect 82031 352621 82073 352739
rect 82191 352621 82207 352739
rect 81897 334727 82207 352621
rect 81897 334609 81913 334727
rect 82031 334609 82073 334727
rect 82191 334609 82207 334727
rect 81897 334567 82207 334609
rect 81897 334449 81913 334567
rect 82031 334449 82073 334567
rect 82191 334449 82207 334567
rect 81897 316727 82207 334449
rect 81897 316609 81913 316727
rect 82031 316609 82073 316727
rect 82191 316609 82207 316727
rect 81897 316567 82207 316609
rect 81897 316449 81913 316567
rect 82031 316449 82073 316567
rect 82191 316449 82207 316567
rect 81897 298727 82207 316449
rect 81897 298609 81913 298727
rect 82031 298609 82073 298727
rect 82191 298609 82207 298727
rect 81897 298567 82207 298609
rect 81897 298449 81913 298567
rect 82031 298449 82073 298567
rect 82191 298449 82207 298567
rect 81897 280727 82207 298449
rect 81897 280609 81913 280727
rect 82031 280609 82073 280727
rect 82191 280609 82207 280727
rect 81897 280567 82207 280609
rect 81897 280449 81913 280567
rect 82031 280449 82073 280567
rect 82191 280449 82207 280567
rect 81897 262727 82207 280449
rect 81897 262609 81913 262727
rect 82031 262609 82073 262727
rect 82191 262609 82207 262727
rect 81897 262567 82207 262609
rect 81897 262449 81913 262567
rect 82031 262449 82073 262567
rect 82191 262449 82207 262567
rect 81897 244727 82207 262449
rect 81897 244609 81913 244727
rect 82031 244609 82073 244727
rect 82191 244609 82207 244727
rect 81897 244567 82207 244609
rect 81897 244449 81913 244567
rect 82031 244449 82073 244567
rect 82191 244449 82207 244567
rect 81897 226727 82207 244449
rect 81897 226609 81913 226727
rect 82031 226609 82073 226727
rect 82191 226609 82207 226727
rect 81897 226567 82207 226609
rect 81897 226449 81913 226567
rect 82031 226449 82073 226567
rect 82191 226449 82207 226567
rect 81897 208727 82207 226449
rect 81897 208609 81913 208727
rect 82031 208609 82073 208727
rect 82191 208609 82207 208727
rect 81897 208567 82207 208609
rect 81897 208449 81913 208567
rect 82031 208449 82073 208567
rect 82191 208449 82207 208567
rect 81897 190727 82207 208449
rect 81897 190609 81913 190727
rect 82031 190609 82073 190727
rect 82191 190609 82207 190727
rect 81897 190567 82207 190609
rect 81897 190449 81913 190567
rect 82031 190449 82073 190567
rect 82191 190449 82207 190567
rect 81897 172727 82207 190449
rect 81897 172609 81913 172727
rect 82031 172609 82073 172727
rect 82191 172609 82207 172727
rect 81897 172567 82207 172609
rect 81897 172449 81913 172567
rect 82031 172449 82073 172567
rect 82191 172449 82207 172567
rect 81897 154727 82207 172449
rect 81897 154609 81913 154727
rect 82031 154609 82073 154727
rect 82191 154609 82207 154727
rect 81897 154567 82207 154609
rect 81897 154449 81913 154567
rect 82031 154449 82073 154567
rect 82191 154449 82207 154567
rect 81897 136727 82207 154449
rect 81897 136609 81913 136727
rect 82031 136609 82073 136727
rect 82191 136609 82207 136727
rect 81897 136567 82207 136609
rect 81897 136449 81913 136567
rect 82031 136449 82073 136567
rect 82191 136449 82207 136567
rect 81897 118727 82207 136449
rect 81897 118609 81913 118727
rect 82031 118609 82073 118727
rect 82191 118609 82207 118727
rect 81897 118567 82207 118609
rect 81897 118449 81913 118567
rect 82031 118449 82073 118567
rect 82191 118449 82207 118567
rect 81897 100727 82207 118449
rect 81897 100609 81913 100727
rect 82031 100609 82073 100727
rect 82191 100609 82207 100727
rect 81897 100567 82207 100609
rect 81897 100449 81913 100567
rect 82031 100449 82073 100567
rect 82191 100449 82207 100567
rect 81897 82727 82207 100449
rect 81897 82609 81913 82727
rect 82031 82609 82073 82727
rect 82191 82609 82207 82727
rect 81897 82567 82207 82609
rect 81897 82449 81913 82567
rect 82031 82449 82073 82567
rect 82191 82449 82207 82567
rect 81897 64727 82207 82449
rect 81897 64609 81913 64727
rect 82031 64609 82073 64727
rect 82191 64609 82207 64727
rect 81897 64567 82207 64609
rect 81897 64449 81913 64567
rect 82031 64449 82073 64567
rect 82191 64449 82207 64567
rect 81897 46727 82207 64449
rect 81897 46609 81913 46727
rect 82031 46609 82073 46727
rect 82191 46609 82207 46727
rect 81897 46567 82207 46609
rect 81897 46449 81913 46567
rect 82031 46449 82073 46567
rect 82191 46449 82207 46567
rect 81897 28727 82207 46449
rect 81897 28609 81913 28727
rect 82031 28609 82073 28727
rect 82191 28609 82207 28727
rect 81897 28567 82207 28609
rect 81897 28449 81913 28567
rect 82031 28449 82073 28567
rect 82191 28449 82207 28567
rect 81897 10727 82207 28449
rect 81897 10609 81913 10727
rect 82031 10609 82073 10727
rect 82191 10609 82207 10727
rect 81897 10567 82207 10609
rect 81897 10449 81913 10567
rect 82031 10449 82073 10567
rect 82191 10449 82207 10567
rect 81897 -653 82207 10449
rect 81897 -771 81913 -653
rect 82031 -771 82073 -653
rect 82191 -771 82207 -653
rect 81897 -813 82207 -771
rect 81897 -931 81913 -813
rect 82031 -931 82073 -813
rect 82191 -931 82207 -813
rect 81897 -947 82207 -931
rect 83757 336587 84067 353581
rect 83757 336469 83773 336587
rect 83891 336469 83933 336587
rect 84051 336469 84067 336587
rect 83757 336427 84067 336469
rect 83757 336309 83773 336427
rect 83891 336309 83933 336427
rect 84051 336309 84067 336427
rect 83757 318587 84067 336309
rect 83757 318469 83773 318587
rect 83891 318469 83933 318587
rect 84051 318469 84067 318587
rect 83757 318427 84067 318469
rect 83757 318309 83773 318427
rect 83891 318309 83933 318427
rect 84051 318309 84067 318427
rect 83757 300587 84067 318309
rect 83757 300469 83773 300587
rect 83891 300469 83933 300587
rect 84051 300469 84067 300587
rect 83757 300427 84067 300469
rect 83757 300309 83773 300427
rect 83891 300309 83933 300427
rect 84051 300309 84067 300427
rect 83757 282587 84067 300309
rect 83757 282469 83773 282587
rect 83891 282469 83933 282587
rect 84051 282469 84067 282587
rect 83757 282427 84067 282469
rect 83757 282309 83773 282427
rect 83891 282309 83933 282427
rect 84051 282309 84067 282427
rect 83757 264587 84067 282309
rect 83757 264469 83773 264587
rect 83891 264469 83933 264587
rect 84051 264469 84067 264587
rect 83757 264427 84067 264469
rect 83757 264309 83773 264427
rect 83891 264309 83933 264427
rect 84051 264309 84067 264427
rect 83757 246587 84067 264309
rect 83757 246469 83773 246587
rect 83891 246469 83933 246587
rect 84051 246469 84067 246587
rect 83757 246427 84067 246469
rect 83757 246309 83773 246427
rect 83891 246309 83933 246427
rect 84051 246309 84067 246427
rect 83757 228587 84067 246309
rect 83757 228469 83773 228587
rect 83891 228469 83933 228587
rect 84051 228469 84067 228587
rect 83757 228427 84067 228469
rect 83757 228309 83773 228427
rect 83891 228309 83933 228427
rect 84051 228309 84067 228427
rect 83757 210587 84067 228309
rect 83757 210469 83773 210587
rect 83891 210469 83933 210587
rect 84051 210469 84067 210587
rect 83757 210427 84067 210469
rect 83757 210309 83773 210427
rect 83891 210309 83933 210427
rect 84051 210309 84067 210427
rect 83757 192587 84067 210309
rect 83757 192469 83773 192587
rect 83891 192469 83933 192587
rect 84051 192469 84067 192587
rect 83757 192427 84067 192469
rect 83757 192309 83773 192427
rect 83891 192309 83933 192427
rect 84051 192309 84067 192427
rect 83757 174587 84067 192309
rect 83757 174469 83773 174587
rect 83891 174469 83933 174587
rect 84051 174469 84067 174587
rect 83757 174427 84067 174469
rect 83757 174309 83773 174427
rect 83891 174309 83933 174427
rect 84051 174309 84067 174427
rect 83757 156587 84067 174309
rect 83757 156469 83773 156587
rect 83891 156469 83933 156587
rect 84051 156469 84067 156587
rect 83757 156427 84067 156469
rect 83757 156309 83773 156427
rect 83891 156309 83933 156427
rect 84051 156309 84067 156427
rect 83757 138587 84067 156309
rect 83757 138469 83773 138587
rect 83891 138469 83933 138587
rect 84051 138469 84067 138587
rect 83757 138427 84067 138469
rect 83757 138309 83773 138427
rect 83891 138309 83933 138427
rect 84051 138309 84067 138427
rect 83757 120587 84067 138309
rect 83757 120469 83773 120587
rect 83891 120469 83933 120587
rect 84051 120469 84067 120587
rect 83757 120427 84067 120469
rect 83757 120309 83773 120427
rect 83891 120309 83933 120427
rect 84051 120309 84067 120427
rect 83757 102587 84067 120309
rect 83757 102469 83773 102587
rect 83891 102469 83933 102587
rect 84051 102469 84067 102587
rect 83757 102427 84067 102469
rect 83757 102309 83773 102427
rect 83891 102309 83933 102427
rect 84051 102309 84067 102427
rect 83757 84587 84067 102309
rect 83757 84469 83773 84587
rect 83891 84469 83933 84587
rect 84051 84469 84067 84587
rect 83757 84427 84067 84469
rect 83757 84309 83773 84427
rect 83891 84309 83933 84427
rect 84051 84309 84067 84427
rect 83757 66587 84067 84309
rect 83757 66469 83773 66587
rect 83891 66469 83933 66587
rect 84051 66469 84067 66587
rect 83757 66427 84067 66469
rect 83757 66309 83773 66427
rect 83891 66309 83933 66427
rect 84051 66309 84067 66427
rect 83757 48587 84067 66309
rect 83757 48469 83773 48587
rect 83891 48469 83933 48587
rect 84051 48469 84067 48587
rect 83757 48427 84067 48469
rect 83757 48309 83773 48427
rect 83891 48309 83933 48427
rect 84051 48309 84067 48427
rect 83757 30587 84067 48309
rect 83757 30469 83773 30587
rect 83891 30469 83933 30587
rect 84051 30469 84067 30587
rect 83757 30427 84067 30469
rect 83757 30309 83773 30427
rect 83891 30309 83933 30427
rect 84051 30309 84067 30427
rect 83757 12587 84067 30309
rect 83757 12469 83773 12587
rect 83891 12469 83933 12587
rect 84051 12469 84067 12587
rect 83757 12427 84067 12469
rect 83757 12309 83773 12427
rect 83891 12309 83933 12427
rect 84051 12309 84067 12427
rect 83757 -1613 84067 12309
rect 83757 -1731 83773 -1613
rect 83891 -1731 83933 -1613
rect 84051 -1731 84067 -1613
rect 83757 -1773 84067 -1731
rect 83757 -1891 83773 -1773
rect 83891 -1891 83933 -1773
rect 84051 -1891 84067 -1773
rect 83757 -1907 84067 -1891
rect 85617 338447 85927 354541
rect 85617 338329 85633 338447
rect 85751 338329 85793 338447
rect 85911 338329 85927 338447
rect 85617 338287 85927 338329
rect 85617 338169 85633 338287
rect 85751 338169 85793 338287
rect 85911 338169 85927 338287
rect 85617 320447 85927 338169
rect 85617 320329 85633 320447
rect 85751 320329 85793 320447
rect 85911 320329 85927 320447
rect 85617 320287 85927 320329
rect 85617 320169 85633 320287
rect 85751 320169 85793 320287
rect 85911 320169 85927 320287
rect 85617 302447 85927 320169
rect 85617 302329 85633 302447
rect 85751 302329 85793 302447
rect 85911 302329 85927 302447
rect 85617 302287 85927 302329
rect 85617 302169 85633 302287
rect 85751 302169 85793 302287
rect 85911 302169 85927 302287
rect 85617 284447 85927 302169
rect 85617 284329 85633 284447
rect 85751 284329 85793 284447
rect 85911 284329 85927 284447
rect 85617 284287 85927 284329
rect 85617 284169 85633 284287
rect 85751 284169 85793 284287
rect 85911 284169 85927 284287
rect 85617 266447 85927 284169
rect 85617 266329 85633 266447
rect 85751 266329 85793 266447
rect 85911 266329 85927 266447
rect 85617 266287 85927 266329
rect 85617 266169 85633 266287
rect 85751 266169 85793 266287
rect 85911 266169 85927 266287
rect 85617 248447 85927 266169
rect 85617 248329 85633 248447
rect 85751 248329 85793 248447
rect 85911 248329 85927 248447
rect 85617 248287 85927 248329
rect 85617 248169 85633 248287
rect 85751 248169 85793 248287
rect 85911 248169 85927 248287
rect 85617 230447 85927 248169
rect 85617 230329 85633 230447
rect 85751 230329 85793 230447
rect 85911 230329 85927 230447
rect 85617 230287 85927 230329
rect 85617 230169 85633 230287
rect 85751 230169 85793 230287
rect 85911 230169 85927 230287
rect 85617 212447 85927 230169
rect 85617 212329 85633 212447
rect 85751 212329 85793 212447
rect 85911 212329 85927 212447
rect 85617 212287 85927 212329
rect 85617 212169 85633 212287
rect 85751 212169 85793 212287
rect 85911 212169 85927 212287
rect 85617 194447 85927 212169
rect 85617 194329 85633 194447
rect 85751 194329 85793 194447
rect 85911 194329 85927 194447
rect 85617 194287 85927 194329
rect 85617 194169 85633 194287
rect 85751 194169 85793 194287
rect 85911 194169 85927 194287
rect 85617 176447 85927 194169
rect 85617 176329 85633 176447
rect 85751 176329 85793 176447
rect 85911 176329 85927 176447
rect 85617 176287 85927 176329
rect 85617 176169 85633 176287
rect 85751 176169 85793 176287
rect 85911 176169 85927 176287
rect 85617 158447 85927 176169
rect 85617 158329 85633 158447
rect 85751 158329 85793 158447
rect 85911 158329 85927 158447
rect 85617 158287 85927 158329
rect 85617 158169 85633 158287
rect 85751 158169 85793 158287
rect 85911 158169 85927 158287
rect 85617 140447 85927 158169
rect 85617 140329 85633 140447
rect 85751 140329 85793 140447
rect 85911 140329 85927 140447
rect 85617 140287 85927 140329
rect 85617 140169 85633 140287
rect 85751 140169 85793 140287
rect 85911 140169 85927 140287
rect 85617 122447 85927 140169
rect 85617 122329 85633 122447
rect 85751 122329 85793 122447
rect 85911 122329 85927 122447
rect 85617 122287 85927 122329
rect 85617 122169 85633 122287
rect 85751 122169 85793 122287
rect 85911 122169 85927 122287
rect 85617 104447 85927 122169
rect 85617 104329 85633 104447
rect 85751 104329 85793 104447
rect 85911 104329 85927 104447
rect 85617 104287 85927 104329
rect 85617 104169 85633 104287
rect 85751 104169 85793 104287
rect 85911 104169 85927 104287
rect 85617 86447 85927 104169
rect 85617 86329 85633 86447
rect 85751 86329 85793 86447
rect 85911 86329 85927 86447
rect 85617 86287 85927 86329
rect 85617 86169 85633 86287
rect 85751 86169 85793 86287
rect 85911 86169 85927 86287
rect 85617 68447 85927 86169
rect 85617 68329 85633 68447
rect 85751 68329 85793 68447
rect 85911 68329 85927 68447
rect 85617 68287 85927 68329
rect 85617 68169 85633 68287
rect 85751 68169 85793 68287
rect 85911 68169 85927 68287
rect 85617 50447 85927 68169
rect 85617 50329 85633 50447
rect 85751 50329 85793 50447
rect 85911 50329 85927 50447
rect 85617 50287 85927 50329
rect 85617 50169 85633 50287
rect 85751 50169 85793 50287
rect 85911 50169 85927 50287
rect 85617 32447 85927 50169
rect 85617 32329 85633 32447
rect 85751 32329 85793 32447
rect 85911 32329 85927 32447
rect 85617 32287 85927 32329
rect 85617 32169 85633 32287
rect 85751 32169 85793 32287
rect 85911 32169 85927 32287
rect 85617 14447 85927 32169
rect 85617 14329 85633 14447
rect 85751 14329 85793 14447
rect 85911 14329 85927 14447
rect 85617 14287 85927 14329
rect 85617 14169 85633 14287
rect 85751 14169 85793 14287
rect 85911 14169 85927 14287
rect 85617 -2573 85927 14169
rect 85617 -2691 85633 -2573
rect 85751 -2691 85793 -2573
rect 85911 -2691 85927 -2573
rect 85617 -2733 85927 -2691
rect 85617 -2851 85633 -2733
rect 85751 -2851 85793 -2733
rect 85911 -2851 85927 -2733
rect 85617 -2867 85927 -2851
rect 87477 340307 87787 355501
rect 96477 355299 96787 355795
rect 96477 355181 96493 355299
rect 96611 355181 96653 355299
rect 96771 355181 96787 355299
rect 96477 355139 96787 355181
rect 96477 355021 96493 355139
rect 96611 355021 96653 355139
rect 96771 355021 96787 355139
rect 94617 354339 94927 354835
rect 94617 354221 94633 354339
rect 94751 354221 94793 354339
rect 94911 354221 94927 354339
rect 94617 354179 94927 354221
rect 94617 354061 94633 354179
rect 94751 354061 94793 354179
rect 94911 354061 94927 354179
rect 92757 353379 93067 353875
rect 92757 353261 92773 353379
rect 92891 353261 92933 353379
rect 93051 353261 93067 353379
rect 92757 353219 93067 353261
rect 92757 353101 92773 353219
rect 92891 353101 92933 353219
rect 93051 353101 93067 353219
rect 87477 340189 87493 340307
rect 87611 340189 87653 340307
rect 87771 340189 87787 340307
rect 87477 340147 87787 340189
rect 87477 340029 87493 340147
rect 87611 340029 87653 340147
rect 87771 340029 87787 340147
rect 87477 322307 87787 340029
rect 87477 322189 87493 322307
rect 87611 322189 87653 322307
rect 87771 322189 87787 322307
rect 87477 322147 87787 322189
rect 87477 322029 87493 322147
rect 87611 322029 87653 322147
rect 87771 322029 87787 322147
rect 87477 304307 87787 322029
rect 87477 304189 87493 304307
rect 87611 304189 87653 304307
rect 87771 304189 87787 304307
rect 87477 304147 87787 304189
rect 87477 304029 87493 304147
rect 87611 304029 87653 304147
rect 87771 304029 87787 304147
rect 87477 286307 87787 304029
rect 87477 286189 87493 286307
rect 87611 286189 87653 286307
rect 87771 286189 87787 286307
rect 87477 286147 87787 286189
rect 87477 286029 87493 286147
rect 87611 286029 87653 286147
rect 87771 286029 87787 286147
rect 87477 268307 87787 286029
rect 87477 268189 87493 268307
rect 87611 268189 87653 268307
rect 87771 268189 87787 268307
rect 87477 268147 87787 268189
rect 87477 268029 87493 268147
rect 87611 268029 87653 268147
rect 87771 268029 87787 268147
rect 87477 250307 87787 268029
rect 87477 250189 87493 250307
rect 87611 250189 87653 250307
rect 87771 250189 87787 250307
rect 87477 250147 87787 250189
rect 87477 250029 87493 250147
rect 87611 250029 87653 250147
rect 87771 250029 87787 250147
rect 87477 232307 87787 250029
rect 87477 232189 87493 232307
rect 87611 232189 87653 232307
rect 87771 232189 87787 232307
rect 87477 232147 87787 232189
rect 87477 232029 87493 232147
rect 87611 232029 87653 232147
rect 87771 232029 87787 232147
rect 87477 214307 87787 232029
rect 87477 214189 87493 214307
rect 87611 214189 87653 214307
rect 87771 214189 87787 214307
rect 87477 214147 87787 214189
rect 87477 214029 87493 214147
rect 87611 214029 87653 214147
rect 87771 214029 87787 214147
rect 87477 196307 87787 214029
rect 87477 196189 87493 196307
rect 87611 196189 87653 196307
rect 87771 196189 87787 196307
rect 87477 196147 87787 196189
rect 87477 196029 87493 196147
rect 87611 196029 87653 196147
rect 87771 196029 87787 196147
rect 87477 178307 87787 196029
rect 87477 178189 87493 178307
rect 87611 178189 87653 178307
rect 87771 178189 87787 178307
rect 87477 178147 87787 178189
rect 87477 178029 87493 178147
rect 87611 178029 87653 178147
rect 87771 178029 87787 178147
rect 87477 160307 87787 178029
rect 87477 160189 87493 160307
rect 87611 160189 87653 160307
rect 87771 160189 87787 160307
rect 87477 160147 87787 160189
rect 87477 160029 87493 160147
rect 87611 160029 87653 160147
rect 87771 160029 87787 160147
rect 87477 142307 87787 160029
rect 87477 142189 87493 142307
rect 87611 142189 87653 142307
rect 87771 142189 87787 142307
rect 87477 142147 87787 142189
rect 87477 142029 87493 142147
rect 87611 142029 87653 142147
rect 87771 142029 87787 142147
rect 87477 124307 87787 142029
rect 87477 124189 87493 124307
rect 87611 124189 87653 124307
rect 87771 124189 87787 124307
rect 87477 124147 87787 124189
rect 87477 124029 87493 124147
rect 87611 124029 87653 124147
rect 87771 124029 87787 124147
rect 87477 106307 87787 124029
rect 87477 106189 87493 106307
rect 87611 106189 87653 106307
rect 87771 106189 87787 106307
rect 87477 106147 87787 106189
rect 87477 106029 87493 106147
rect 87611 106029 87653 106147
rect 87771 106029 87787 106147
rect 87477 88307 87787 106029
rect 87477 88189 87493 88307
rect 87611 88189 87653 88307
rect 87771 88189 87787 88307
rect 87477 88147 87787 88189
rect 87477 88029 87493 88147
rect 87611 88029 87653 88147
rect 87771 88029 87787 88147
rect 87477 70307 87787 88029
rect 87477 70189 87493 70307
rect 87611 70189 87653 70307
rect 87771 70189 87787 70307
rect 87477 70147 87787 70189
rect 87477 70029 87493 70147
rect 87611 70029 87653 70147
rect 87771 70029 87787 70147
rect 87477 52307 87787 70029
rect 87477 52189 87493 52307
rect 87611 52189 87653 52307
rect 87771 52189 87787 52307
rect 87477 52147 87787 52189
rect 87477 52029 87493 52147
rect 87611 52029 87653 52147
rect 87771 52029 87787 52147
rect 87477 34307 87787 52029
rect 87477 34189 87493 34307
rect 87611 34189 87653 34307
rect 87771 34189 87787 34307
rect 87477 34147 87787 34189
rect 87477 34029 87493 34147
rect 87611 34029 87653 34147
rect 87771 34029 87787 34147
rect 87477 16307 87787 34029
rect 87477 16189 87493 16307
rect 87611 16189 87653 16307
rect 87771 16189 87787 16307
rect 87477 16147 87787 16189
rect 87477 16029 87493 16147
rect 87611 16029 87653 16147
rect 87771 16029 87787 16147
rect 78477 -3171 78493 -3053
rect 78611 -3171 78653 -3053
rect 78771 -3171 78787 -3053
rect 78477 -3213 78787 -3171
rect 78477 -3331 78493 -3213
rect 78611 -3331 78653 -3213
rect 78771 -3331 78787 -3213
rect 78477 -3827 78787 -3331
rect 87477 -3533 87787 16029
rect 90897 352419 91207 352915
rect 90897 352301 90913 352419
rect 91031 352301 91073 352419
rect 91191 352301 91207 352419
rect 90897 352259 91207 352301
rect 90897 352141 90913 352259
rect 91031 352141 91073 352259
rect 91191 352141 91207 352259
rect 90897 343727 91207 352141
rect 90897 343609 90913 343727
rect 91031 343609 91073 343727
rect 91191 343609 91207 343727
rect 90897 343567 91207 343609
rect 90897 343449 90913 343567
rect 91031 343449 91073 343567
rect 91191 343449 91207 343567
rect 90897 325727 91207 343449
rect 90897 325609 90913 325727
rect 91031 325609 91073 325727
rect 91191 325609 91207 325727
rect 90897 325567 91207 325609
rect 90897 325449 90913 325567
rect 91031 325449 91073 325567
rect 91191 325449 91207 325567
rect 90897 307727 91207 325449
rect 90897 307609 90913 307727
rect 91031 307609 91073 307727
rect 91191 307609 91207 307727
rect 90897 307567 91207 307609
rect 90897 307449 90913 307567
rect 91031 307449 91073 307567
rect 91191 307449 91207 307567
rect 90897 289727 91207 307449
rect 90897 289609 90913 289727
rect 91031 289609 91073 289727
rect 91191 289609 91207 289727
rect 90897 289567 91207 289609
rect 90897 289449 90913 289567
rect 91031 289449 91073 289567
rect 91191 289449 91207 289567
rect 90897 271727 91207 289449
rect 90897 271609 90913 271727
rect 91031 271609 91073 271727
rect 91191 271609 91207 271727
rect 90897 271567 91207 271609
rect 90897 271449 90913 271567
rect 91031 271449 91073 271567
rect 91191 271449 91207 271567
rect 90897 253727 91207 271449
rect 90897 253609 90913 253727
rect 91031 253609 91073 253727
rect 91191 253609 91207 253727
rect 90897 253567 91207 253609
rect 90897 253449 90913 253567
rect 91031 253449 91073 253567
rect 91191 253449 91207 253567
rect 90897 235727 91207 253449
rect 90897 235609 90913 235727
rect 91031 235609 91073 235727
rect 91191 235609 91207 235727
rect 90897 235567 91207 235609
rect 90897 235449 90913 235567
rect 91031 235449 91073 235567
rect 91191 235449 91207 235567
rect 90897 217727 91207 235449
rect 90897 217609 90913 217727
rect 91031 217609 91073 217727
rect 91191 217609 91207 217727
rect 90897 217567 91207 217609
rect 90897 217449 90913 217567
rect 91031 217449 91073 217567
rect 91191 217449 91207 217567
rect 90897 199727 91207 217449
rect 90897 199609 90913 199727
rect 91031 199609 91073 199727
rect 91191 199609 91207 199727
rect 90897 199567 91207 199609
rect 90897 199449 90913 199567
rect 91031 199449 91073 199567
rect 91191 199449 91207 199567
rect 90897 181727 91207 199449
rect 90897 181609 90913 181727
rect 91031 181609 91073 181727
rect 91191 181609 91207 181727
rect 90897 181567 91207 181609
rect 90897 181449 90913 181567
rect 91031 181449 91073 181567
rect 91191 181449 91207 181567
rect 90897 163727 91207 181449
rect 90897 163609 90913 163727
rect 91031 163609 91073 163727
rect 91191 163609 91207 163727
rect 90897 163567 91207 163609
rect 90897 163449 90913 163567
rect 91031 163449 91073 163567
rect 91191 163449 91207 163567
rect 90897 145727 91207 163449
rect 90897 145609 90913 145727
rect 91031 145609 91073 145727
rect 91191 145609 91207 145727
rect 90897 145567 91207 145609
rect 90897 145449 90913 145567
rect 91031 145449 91073 145567
rect 91191 145449 91207 145567
rect 90897 127727 91207 145449
rect 90897 127609 90913 127727
rect 91031 127609 91073 127727
rect 91191 127609 91207 127727
rect 90897 127567 91207 127609
rect 90897 127449 90913 127567
rect 91031 127449 91073 127567
rect 91191 127449 91207 127567
rect 90897 109727 91207 127449
rect 90897 109609 90913 109727
rect 91031 109609 91073 109727
rect 91191 109609 91207 109727
rect 90897 109567 91207 109609
rect 90897 109449 90913 109567
rect 91031 109449 91073 109567
rect 91191 109449 91207 109567
rect 90897 91727 91207 109449
rect 90897 91609 90913 91727
rect 91031 91609 91073 91727
rect 91191 91609 91207 91727
rect 90897 91567 91207 91609
rect 90897 91449 90913 91567
rect 91031 91449 91073 91567
rect 91191 91449 91207 91567
rect 90897 73727 91207 91449
rect 90897 73609 90913 73727
rect 91031 73609 91073 73727
rect 91191 73609 91207 73727
rect 90897 73567 91207 73609
rect 90897 73449 90913 73567
rect 91031 73449 91073 73567
rect 91191 73449 91207 73567
rect 90897 55727 91207 73449
rect 90897 55609 90913 55727
rect 91031 55609 91073 55727
rect 91191 55609 91207 55727
rect 90897 55567 91207 55609
rect 90897 55449 90913 55567
rect 91031 55449 91073 55567
rect 91191 55449 91207 55567
rect 90897 37727 91207 55449
rect 90897 37609 90913 37727
rect 91031 37609 91073 37727
rect 91191 37609 91207 37727
rect 90897 37567 91207 37609
rect 90897 37449 90913 37567
rect 91031 37449 91073 37567
rect 91191 37449 91207 37567
rect 90897 19727 91207 37449
rect 90897 19609 90913 19727
rect 91031 19609 91073 19727
rect 91191 19609 91207 19727
rect 90897 19567 91207 19609
rect 90897 19449 90913 19567
rect 91031 19449 91073 19567
rect 91191 19449 91207 19567
rect 90897 1727 91207 19449
rect 90897 1609 90913 1727
rect 91031 1609 91073 1727
rect 91191 1609 91207 1727
rect 90897 1567 91207 1609
rect 90897 1449 90913 1567
rect 91031 1449 91073 1567
rect 91191 1449 91207 1567
rect 90897 -173 91207 1449
rect 90897 -291 90913 -173
rect 91031 -291 91073 -173
rect 91191 -291 91207 -173
rect 90897 -333 91207 -291
rect 90897 -451 90913 -333
rect 91031 -451 91073 -333
rect 91191 -451 91207 -333
rect 90897 -947 91207 -451
rect 92757 345587 93067 353101
rect 92757 345469 92773 345587
rect 92891 345469 92933 345587
rect 93051 345469 93067 345587
rect 92757 345427 93067 345469
rect 92757 345309 92773 345427
rect 92891 345309 92933 345427
rect 93051 345309 93067 345427
rect 92757 327587 93067 345309
rect 92757 327469 92773 327587
rect 92891 327469 92933 327587
rect 93051 327469 93067 327587
rect 92757 327427 93067 327469
rect 92757 327309 92773 327427
rect 92891 327309 92933 327427
rect 93051 327309 93067 327427
rect 92757 309587 93067 327309
rect 92757 309469 92773 309587
rect 92891 309469 92933 309587
rect 93051 309469 93067 309587
rect 92757 309427 93067 309469
rect 92757 309309 92773 309427
rect 92891 309309 92933 309427
rect 93051 309309 93067 309427
rect 92757 291587 93067 309309
rect 92757 291469 92773 291587
rect 92891 291469 92933 291587
rect 93051 291469 93067 291587
rect 92757 291427 93067 291469
rect 92757 291309 92773 291427
rect 92891 291309 92933 291427
rect 93051 291309 93067 291427
rect 92757 273587 93067 291309
rect 92757 273469 92773 273587
rect 92891 273469 92933 273587
rect 93051 273469 93067 273587
rect 92757 273427 93067 273469
rect 92757 273309 92773 273427
rect 92891 273309 92933 273427
rect 93051 273309 93067 273427
rect 92757 255587 93067 273309
rect 92757 255469 92773 255587
rect 92891 255469 92933 255587
rect 93051 255469 93067 255587
rect 92757 255427 93067 255469
rect 92757 255309 92773 255427
rect 92891 255309 92933 255427
rect 93051 255309 93067 255427
rect 92757 237587 93067 255309
rect 92757 237469 92773 237587
rect 92891 237469 92933 237587
rect 93051 237469 93067 237587
rect 92757 237427 93067 237469
rect 92757 237309 92773 237427
rect 92891 237309 92933 237427
rect 93051 237309 93067 237427
rect 92757 219587 93067 237309
rect 92757 219469 92773 219587
rect 92891 219469 92933 219587
rect 93051 219469 93067 219587
rect 92757 219427 93067 219469
rect 92757 219309 92773 219427
rect 92891 219309 92933 219427
rect 93051 219309 93067 219427
rect 92757 201587 93067 219309
rect 92757 201469 92773 201587
rect 92891 201469 92933 201587
rect 93051 201469 93067 201587
rect 92757 201427 93067 201469
rect 92757 201309 92773 201427
rect 92891 201309 92933 201427
rect 93051 201309 93067 201427
rect 92757 183587 93067 201309
rect 92757 183469 92773 183587
rect 92891 183469 92933 183587
rect 93051 183469 93067 183587
rect 92757 183427 93067 183469
rect 92757 183309 92773 183427
rect 92891 183309 92933 183427
rect 93051 183309 93067 183427
rect 92757 165587 93067 183309
rect 92757 165469 92773 165587
rect 92891 165469 92933 165587
rect 93051 165469 93067 165587
rect 92757 165427 93067 165469
rect 92757 165309 92773 165427
rect 92891 165309 92933 165427
rect 93051 165309 93067 165427
rect 92757 147587 93067 165309
rect 92757 147469 92773 147587
rect 92891 147469 92933 147587
rect 93051 147469 93067 147587
rect 92757 147427 93067 147469
rect 92757 147309 92773 147427
rect 92891 147309 92933 147427
rect 93051 147309 93067 147427
rect 92757 129587 93067 147309
rect 92757 129469 92773 129587
rect 92891 129469 92933 129587
rect 93051 129469 93067 129587
rect 92757 129427 93067 129469
rect 92757 129309 92773 129427
rect 92891 129309 92933 129427
rect 93051 129309 93067 129427
rect 92757 111587 93067 129309
rect 92757 111469 92773 111587
rect 92891 111469 92933 111587
rect 93051 111469 93067 111587
rect 92757 111427 93067 111469
rect 92757 111309 92773 111427
rect 92891 111309 92933 111427
rect 93051 111309 93067 111427
rect 92757 93587 93067 111309
rect 92757 93469 92773 93587
rect 92891 93469 92933 93587
rect 93051 93469 93067 93587
rect 92757 93427 93067 93469
rect 92757 93309 92773 93427
rect 92891 93309 92933 93427
rect 93051 93309 93067 93427
rect 92757 75587 93067 93309
rect 92757 75469 92773 75587
rect 92891 75469 92933 75587
rect 93051 75469 93067 75587
rect 92757 75427 93067 75469
rect 92757 75309 92773 75427
rect 92891 75309 92933 75427
rect 93051 75309 93067 75427
rect 92757 57587 93067 75309
rect 92757 57469 92773 57587
rect 92891 57469 92933 57587
rect 93051 57469 93067 57587
rect 92757 57427 93067 57469
rect 92757 57309 92773 57427
rect 92891 57309 92933 57427
rect 93051 57309 93067 57427
rect 92757 39587 93067 57309
rect 92757 39469 92773 39587
rect 92891 39469 92933 39587
rect 93051 39469 93067 39587
rect 92757 39427 93067 39469
rect 92757 39309 92773 39427
rect 92891 39309 92933 39427
rect 93051 39309 93067 39427
rect 92757 21587 93067 39309
rect 92757 21469 92773 21587
rect 92891 21469 92933 21587
rect 93051 21469 93067 21587
rect 92757 21427 93067 21469
rect 92757 21309 92773 21427
rect 92891 21309 92933 21427
rect 93051 21309 93067 21427
rect 92757 3587 93067 21309
rect 92757 3469 92773 3587
rect 92891 3469 92933 3587
rect 93051 3469 93067 3587
rect 92757 3427 93067 3469
rect 92757 3309 92773 3427
rect 92891 3309 92933 3427
rect 93051 3309 93067 3427
rect 92757 -1133 93067 3309
rect 92757 -1251 92773 -1133
rect 92891 -1251 92933 -1133
rect 93051 -1251 93067 -1133
rect 92757 -1293 93067 -1251
rect 92757 -1411 92773 -1293
rect 92891 -1411 92933 -1293
rect 93051 -1411 93067 -1293
rect 92757 -1907 93067 -1411
rect 94617 347447 94927 354061
rect 94617 347329 94633 347447
rect 94751 347329 94793 347447
rect 94911 347329 94927 347447
rect 94617 347287 94927 347329
rect 94617 347169 94633 347287
rect 94751 347169 94793 347287
rect 94911 347169 94927 347287
rect 94617 329447 94927 347169
rect 94617 329329 94633 329447
rect 94751 329329 94793 329447
rect 94911 329329 94927 329447
rect 94617 329287 94927 329329
rect 94617 329169 94633 329287
rect 94751 329169 94793 329287
rect 94911 329169 94927 329287
rect 94617 311447 94927 329169
rect 94617 311329 94633 311447
rect 94751 311329 94793 311447
rect 94911 311329 94927 311447
rect 94617 311287 94927 311329
rect 94617 311169 94633 311287
rect 94751 311169 94793 311287
rect 94911 311169 94927 311287
rect 94617 293447 94927 311169
rect 94617 293329 94633 293447
rect 94751 293329 94793 293447
rect 94911 293329 94927 293447
rect 94617 293287 94927 293329
rect 94617 293169 94633 293287
rect 94751 293169 94793 293287
rect 94911 293169 94927 293287
rect 94617 275447 94927 293169
rect 94617 275329 94633 275447
rect 94751 275329 94793 275447
rect 94911 275329 94927 275447
rect 94617 275287 94927 275329
rect 94617 275169 94633 275287
rect 94751 275169 94793 275287
rect 94911 275169 94927 275287
rect 94617 257447 94927 275169
rect 94617 257329 94633 257447
rect 94751 257329 94793 257447
rect 94911 257329 94927 257447
rect 94617 257287 94927 257329
rect 94617 257169 94633 257287
rect 94751 257169 94793 257287
rect 94911 257169 94927 257287
rect 94617 239447 94927 257169
rect 94617 239329 94633 239447
rect 94751 239329 94793 239447
rect 94911 239329 94927 239447
rect 94617 239287 94927 239329
rect 94617 239169 94633 239287
rect 94751 239169 94793 239287
rect 94911 239169 94927 239287
rect 94617 221447 94927 239169
rect 94617 221329 94633 221447
rect 94751 221329 94793 221447
rect 94911 221329 94927 221447
rect 94617 221287 94927 221329
rect 94617 221169 94633 221287
rect 94751 221169 94793 221287
rect 94911 221169 94927 221287
rect 94617 203447 94927 221169
rect 94617 203329 94633 203447
rect 94751 203329 94793 203447
rect 94911 203329 94927 203447
rect 94617 203287 94927 203329
rect 94617 203169 94633 203287
rect 94751 203169 94793 203287
rect 94911 203169 94927 203287
rect 94617 185447 94927 203169
rect 94617 185329 94633 185447
rect 94751 185329 94793 185447
rect 94911 185329 94927 185447
rect 94617 185287 94927 185329
rect 94617 185169 94633 185287
rect 94751 185169 94793 185287
rect 94911 185169 94927 185287
rect 94617 167447 94927 185169
rect 94617 167329 94633 167447
rect 94751 167329 94793 167447
rect 94911 167329 94927 167447
rect 94617 167287 94927 167329
rect 94617 167169 94633 167287
rect 94751 167169 94793 167287
rect 94911 167169 94927 167287
rect 94617 149447 94927 167169
rect 94617 149329 94633 149447
rect 94751 149329 94793 149447
rect 94911 149329 94927 149447
rect 94617 149287 94927 149329
rect 94617 149169 94633 149287
rect 94751 149169 94793 149287
rect 94911 149169 94927 149287
rect 94617 131447 94927 149169
rect 94617 131329 94633 131447
rect 94751 131329 94793 131447
rect 94911 131329 94927 131447
rect 94617 131287 94927 131329
rect 94617 131169 94633 131287
rect 94751 131169 94793 131287
rect 94911 131169 94927 131287
rect 94617 113447 94927 131169
rect 94617 113329 94633 113447
rect 94751 113329 94793 113447
rect 94911 113329 94927 113447
rect 94617 113287 94927 113329
rect 94617 113169 94633 113287
rect 94751 113169 94793 113287
rect 94911 113169 94927 113287
rect 94617 95447 94927 113169
rect 94617 95329 94633 95447
rect 94751 95329 94793 95447
rect 94911 95329 94927 95447
rect 94617 95287 94927 95329
rect 94617 95169 94633 95287
rect 94751 95169 94793 95287
rect 94911 95169 94927 95287
rect 94617 77447 94927 95169
rect 94617 77329 94633 77447
rect 94751 77329 94793 77447
rect 94911 77329 94927 77447
rect 94617 77287 94927 77329
rect 94617 77169 94633 77287
rect 94751 77169 94793 77287
rect 94911 77169 94927 77287
rect 94617 59447 94927 77169
rect 94617 59329 94633 59447
rect 94751 59329 94793 59447
rect 94911 59329 94927 59447
rect 94617 59287 94927 59329
rect 94617 59169 94633 59287
rect 94751 59169 94793 59287
rect 94911 59169 94927 59287
rect 94617 41447 94927 59169
rect 94617 41329 94633 41447
rect 94751 41329 94793 41447
rect 94911 41329 94927 41447
rect 94617 41287 94927 41329
rect 94617 41169 94633 41287
rect 94751 41169 94793 41287
rect 94911 41169 94927 41287
rect 94617 23447 94927 41169
rect 94617 23329 94633 23447
rect 94751 23329 94793 23447
rect 94911 23329 94927 23447
rect 94617 23287 94927 23329
rect 94617 23169 94633 23287
rect 94751 23169 94793 23287
rect 94911 23169 94927 23287
rect 94617 5447 94927 23169
rect 94617 5329 94633 5447
rect 94751 5329 94793 5447
rect 94911 5329 94927 5447
rect 94617 5287 94927 5329
rect 94617 5169 94633 5287
rect 94751 5169 94793 5287
rect 94911 5169 94927 5287
rect 94617 -2093 94927 5169
rect 94617 -2211 94633 -2093
rect 94751 -2211 94793 -2093
rect 94911 -2211 94927 -2093
rect 94617 -2253 94927 -2211
rect 94617 -2371 94633 -2253
rect 94751 -2371 94793 -2253
rect 94911 -2371 94927 -2253
rect 94617 -2867 94927 -2371
rect 96477 349307 96787 355021
rect 105477 355779 105787 355795
rect 105477 355661 105493 355779
rect 105611 355661 105653 355779
rect 105771 355661 105787 355779
rect 105477 355619 105787 355661
rect 105477 355501 105493 355619
rect 105611 355501 105653 355619
rect 105771 355501 105787 355619
rect 103617 354819 103927 354835
rect 103617 354701 103633 354819
rect 103751 354701 103793 354819
rect 103911 354701 103927 354819
rect 103617 354659 103927 354701
rect 103617 354541 103633 354659
rect 103751 354541 103793 354659
rect 103911 354541 103927 354659
rect 101757 353859 102067 353875
rect 101757 353741 101773 353859
rect 101891 353741 101933 353859
rect 102051 353741 102067 353859
rect 101757 353699 102067 353741
rect 101757 353581 101773 353699
rect 101891 353581 101933 353699
rect 102051 353581 102067 353699
rect 96477 349189 96493 349307
rect 96611 349189 96653 349307
rect 96771 349189 96787 349307
rect 96477 349147 96787 349189
rect 96477 349029 96493 349147
rect 96611 349029 96653 349147
rect 96771 349029 96787 349147
rect 96477 331307 96787 349029
rect 96477 331189 96493 331307
rect 96611 331189 96653 331307
rect 96771 331189 96787 331307
rect 96477 331147 96787 331189
rect 96477 331029 96493 331147
rect 96611 331029 96653 331147
rect 96771 331029 96787 331147
rect 96477 313307 96787 331029
rect 96477 313189 96493 313307
rect 96611 313189 96653 313307
rect 96771 313189 96787 313307
rect 96477 313147 96787 313189
rect 96477 313029 96493 313147
rect 96611 313029 96653 313147
rect 96771 313029 96787 313147
rect 96477 295307 96787 313029
rect 96477 295189 96493 295307
rect 96611 295189 96653 295307
rect 96771 295189 96787 295307
rect 96477 295147 96787 295189
rect 96477 295029 96493 295147
rect 96611 295029 96653 295147
rect 96771 295029 96787 295147
rect 96477 277307 96787 295029
rect 96477 277189 96493 277307
rect 96611 277189 96653 277307
rect 96771 277189 96787 277307
rect 96477 277147 96787 277189
rect 96477 277029 96493 277147
rect 96611 277029 96653 277147
rect 96771 277029 96787 277147
rect 96477 259307 96787 277029
rect 96477 259189 96493 259307
rect 96611 259189 96653 259307
rect 96771 259189 96787 259307
rect 96477 259147 96787 259189
rect 96477 259029 96493 259147
rect 96611 259029 96653 259147
rect 96771 259029 96787 259147
rect 96477 241307 96787 259029
rect 96477 241189 96493 241307
rect 96611 241189 96653 241307
rect 96771 241189 96787 241307
rect 96477 241147 96787 241189
rect 96477 241029 96493 241147
rect 96611 241029 96653 241147
rect 96771 241029 96787 241147
rect 96477 223307 96787 241029
rect 96477 223189 96493 223307
rect 96611 223189 96653 223307
rect 96771 223189 96787 223307
rect 96477 223147 96787 223189
rect 96477 223029 96493 223147
rect 96611 223029 96653 223147
rect 96771 223029 96787 223147
rect 96477 205307 96787 223029
rect 96477 205189 96493 205307
rect 96611 205189 96653 205307
rect 96771 205189 96787 205307
rect 96477 205147 96787 205189
rect 96477 205029 96493 205147
rect 96611 205029 96653 205147
rect 96771 205029 96787 205147
rect 96477 187307 96787 205029
rect 96477 187189 96493 187307
rect 96611 187189 96653 187307
rect 96771 187189 96787 187307
rect 96477 187147 96787 187189
rect 96477 187029 96493 187147
rect 96611 187029 96653 187147
rect 96771 187029 96787 187147
rect 96477 169307 96787 187029
rect 96477 169189 96493 169307
rect 96611 169189 96653 169307
rect 96771 169189 96787 169307
rect 96477 169147 96787 169189
rect 96477 169029 96493 169147
rect 96611 169029 96653 169147
rect 96771 169029 96787 169147
rect 96477 151307 96787 169029
rect 96477 151189 96493 151307
rect 96611 151189 96653 151307
rect 96771 151189 96787 151307
rect 96477 151147 96787 151189
rect 96477 151029 96493 151147
rect 96611 151029 96653 151147
rect 96771 151029 96787 151147
rect 96477 133307 96787 151029
rect 96477 133189 96493 133307
rect 96611 133189 96653 133307
rect 96771 133189 96787 133307
rect 96477 133147 96787 133189
rect 96477 133029 96493 133147
rect 96611 133029 96653 133147
rect 96771 133029 96787 133147
rect 96477 115307 96787 133029
rect 96477 115189 96493 115307
rect 96611 115189 96653 115307
rect 96771 115189 96787 115307
rect 96477 115147 96787 115189
rect 96477 115029 96493 115147
rect 96611 115029 96653 115147
rect 96771 115029 96787 115147
rect 96477 97307 96787 115029
rect 96477 97189 96493 97307
rect 96611 97189 96653 97307
rect 96771 97189 96787 97307
rect 96477 97147 96787 97189
rect 96477 97029 96493 97147
rect 96611 97029 96653 97147
rect 96771 97029 96787 97147
rect 96477 79307 96787 97029
rect 96477 79189 96493 79307
rect 96611 79189 96653 79307
rect 96771 79189 96787 79307
rect 96477 79147 96787 79189
rect 96477 79029 96493 79147
rect 96611 79029 96653 79147
rect 96771 79029 96787 79147
rect 96477 61307 96787 79029
rect 96477 61189 96493 61307
rect 96611 61189 96653 61307
rect 96771 61189 96787 61307
rect 96477 61147 96787 61189
rect 96477 61029 96493 61147
rect 96611 61029 96653 61147
rect 96771 61029 96787 61147
rect 96477 43307 96787 61029
rect 96477 43189 96493 43307
rect 96611 43189 96653 43307
rect 96771 43189 96787 43307
rect 96477 43147 96787 43189
rect 96477 43029 96493 43147
rect 96611 43029 96653 43147
rect 96771 43029 96787 43147
rect 96477 25307 96787 43029
rect 96477 25189 96493 25307
rect 96611 25189 96653 25307
rect 96771 25189 96787 25307
rect 96477 25147 96787 25189
rect 96477 25029 96493 25147
rect 96611 25029 96653 25147
rect 96771 25029 96787 25147
rect 96477 7307 96787 25029
rect 96477 7189 96493 7307
rect 96611 7189 96653 7307
rect 96771 7189 96787 7307
rect 96477 7147 96787 7189
rect 96477 7029 96493 7147
rect 96611 7029 96653 7147
rect 96771 7029 96787 7147
rect 87477 -3651 87493 -3533
rect 87611 -3651 87653 -3533
rect 87771 -3651 87787 -3533
rect 87477 -3693 87787 -3651
rect 87477 -3811 87493 -3693
rect 87611 -3811 87653 -3693
rect 87771 -3811 87787 -3693
rect 87477 -3827 87787 -3811
rect 96477 -3053 96787 7029
rect 99897 352899 100207 352915
rect 99897 352781 99913 352899
rect 100031 352781 100073 352899
rect 100191 352781 100207 352899
rect 99897 352739 100207 352781
rect 99897 352621 99913 352739
rect 100031 352621 100073 352739
rect 100191 352621 100207 352739
rect 99897 334727 100207 352621
rect 99897 334609 99913 334727
rect 100031 334609 100073 334727
rect 100191 334609 100207 334727
rect 99897 334567 100207 334609
rect 99897 334449 99913 334567
rect 100031 334449 100073 334567
rect 100191 334449 100207 334567
rect 99897 316727 100207 334449
rect 99897 316609 99913 316727
rect 100031 316609 100073 316727
rect 100191 316609 100207 316727
rect 99897 316567 100207 316609
rect 99897 316449 99913 316567
rect 100031 316449 100073 316567
rect 100191 316449 100207 316567
rect 99897 298727 100207 316449
rect 99897 298609 99913 298727
rect 100031 298609 100073 298727
rect 100191 298609 100207 298727
rect 99897 298567 100207 298609
rect 99897 298449 99913 298567
rect 100031 298449 100073 298567
rect 100191 298449 100207 298567
rect 99897 280727 100207 298449
rect 99897 280609 99913 280727
rect 100031 280609 100073 280727
rect 100191 280609 100207 280727
rect 99897 280567 100207 280609
rect 99897 280449 99913 280567
rect 100031 280449 100073 280567
rect 100191 280449 100207 280567
rect 99897 262727 100207 280449
rect 99897 262609 99913 262727
rect 100031 262609 100073 262727
rect 100191 262609 100207 262727
rect 99897 262567 100207 262609
rect 99897 262449 99913 262567
rect 100031 262449 100073 262567
rect 100191 262449 100207 262567
rect 99897 244727 100207 262449
rect 99897 244609 99913 244727
rect 100031 244609 100073 244727
rect 100191 244609 100207 244727
rect 99897 244567 100207 244609
rect 99897 244449 99913 244567
rect 100031 244449 100073 244567
rect 100191 244449 100207 244567
rect 99897 226727 100207 244449
rect 99897 226609 99913 226727
rect 100031 226609 100073 226727
rect 100191 226609 100207 226727
rect 99897 226567 100207 226609
rect 99897 226449 99913 226567
rect 100031 226449 100073 226567
rect 100191 226449 100207 226567
rect 99897 208727 100207 226449
rect 99897 208609 99913 208727
rect 100031 208609 100073 208727
rect 100191 208609 100207 208727
rect 99897 208567 100207 208609
rect 99897 208449 99913 208567
rect 100031 208449 100073 208567
rect 100191 208449 100207 208567
rect 99897 190727 100207 208449
rect 99897 190609 99913 190727
rect 100031 190609 100073 190727
rect 100191 190609 100207 190727
rect 99897 190567 100207 190609
rect 99897 190449 99913 190567
rect 100031 190449 100073 190567
rect 100191 190449 100207 190567
rect 99897 172727 100207 190449
rect 99897 172609 99913 172727
rect 100031 172609 100073 172727
rect 100191 172609 100207 172727
rect 99897 172567 100207 172609
rect 99897 172449 99913 172567
rect 100031 172449 100073 172567
rect 100191 172449 100207 172567
rect 99897 154727 100207 172449
rect 99897 154609 99913 154727
rect 100031 154609 100073 154727
rect 100191 154609 100207 154727
rect 99897 154567 100207 154609
rect 99897 154449 99913 154567
rect 100031 154449 100073 154567
rect 100191 154449 100207 154567
rect 99897 136727 100207 154449
rect 99897 136609 99913 136727
rect 100031 136609 100073 136727
rect 100191 136609 100207 136727
rect 99897 136567 100207 136609
rect 99897 136449 99913 136567
rect 100031 136449 100073 136567
rect 100191 136449 100207 136567
rect 99897 118727 100207 136449
rect 99897 118609 99913 118727
rect 100031 118609 100073 118727
rect 100191 118609 100207 118727
rect 99897 118567 100207 118609
rect 99897 118449 99913 118567
rect 100031 118449 100073 118567
rect 100191 118449 100207 118567
rect 99897 100727 100207 118449
rect 99897 100609 99913 100727
rect 100031 100609 100073 100727
rect 100191 100609 100207 100727
rect 99897 100567 100207 100609
rect 99897 100449 99913 100567
rect 100031 100449 100073 100567
rect 100191 100449 100207 100567
rect 99897 82727 100207 100449
rect 99897 82609 99913 82727
rect 100031 82609 100073 82727
rect 100191 82609 100207 82727
rect 99897 82567 100207 82609
rect 99897 82449 99913 82567
rect 100031 82449 100073 82567
rect 100191 82449 100207 82567
rect 99897 64727 100207 82449
rect 99897 64609 99913 64727
rect 100031 64609 100073 64727
rect 100191 64609 100207 64727
rect 99897 64567 100207 64609
rect 99897 64449 99913 64567
rect 100031 64449 100073 64567
rect 100191 64449 100207 64567
rect 99897 46727 100207 64449
rect 99897 46609 99913 46727
rect 100031 46609 100073 46727
rect 100191 46609 100207 46727
rect 99897 46567 100207 46609
rect 99897 46449 99913 46567
rect 100031 46449 100073 46567
rect 100191 46449 100207 46567
rect 99897 28727 100207 46449
rect 99897 28609 99913 28727
rect 100031 28609 100073 28727
rect 100191 28609 100207 28727
rect 99897 28567 100207 28609
rect 99897 28449 99913 28567
rect 100031 28449 100073 28567
rect 100191 28449 100207 28567
rect 99897 10727 100207 28449
rect 99897 10609 99913 10727
rect 100031 10609 100073 10727
rect 100191 10609 100207 10727
rect 99897 10567 100207 10609
rect 99897 10449 99913 10567
rect 100031 10449 100073 10567
rect 100191 10449 100207 10567
rect 99897 -653 100207 10449
rect 99897 -771 99913 -653
rect 100031 -771 100073 -653
rect 100191 -771 100207 -653
rect 99897 -813 100207 -771
rect 99897 -931 99913 -813
rect 100031 -931 100073 -813
rect 100191 -931 100207 -813
rect 99897 -947 100207 -931
rect 101757 336587 102067 353581
rect 101757 336469 101773 336587
rect 101891 336469 101933 336587
rect 102051 336469 102067 336587
rect 101757 336427 102067 336469
rect 101757 336309 101773 336427
rect 101891 336309 101933 336427
rect 102051 336309 102067 336427
rect 101757 318587 102067 336309
rect 101757 318469 101773 318587
rect 101891 318469 101933 318587
rect 102051 318469 102067 318587
rect 101757 318427 102067 318469
rect 101757 318309 101773 318427
rect 101891 318309 101933 318427
rect 102051 318309 102067 318427
rect 101757 300587 102067 318309
rect 101757 300469 101773 300587
rect 101891 300469 101933 300587
rect 102051 300469 102067 300587
rect 101757 300427 102067 300469
rect 101757 300309 101773 300427
rect 101891 300309 101933 300427
rect 102051 300309 102067 300427
rect 101757 282587 102067 300309
rect 101757 282469 101773 282587
rect 101891 282469 101933 282587
rect 102051 282469 102067 282587
rect 101757 282427 102067 282469
rect 101757 282309 101773 282427
rect 101891 282309 101933 282427
rect 102051 282309 102067 282427
rect 101757 264587 102067 282309
rect 101757 264469 101773 264587
rect 101891 264469 101933 264587
rect 102051 264469 102067 264587
rect 101757 264427 102067 264469
rect 101757 264309 101773 264427
rect 101891 264309 101933 264427
rect 102051 264309 102067 264427
rect 101757 246587 102067 264309
rect 101757 246469 101773 246587
rect 101891 246469 101933 246587
rect 102051 246469 102067 246587
rect 101757 246427 102067 246469
rect 101757 246309 101773 246427
rect 101891 246309 101933 246427
rect 102051 246309 102067 246427
rect 101757 228587 102067 246309
rect 101757 228469 101773 228587
rect 101891 228469 101933 228587
rect 102051 228469 102067 228587
rect 101757 228427 102067 228469
rect 101757 228309 101773 228427
rect 101891 228309 101933 228427
rect 102051 228309 102067 228427
rect 101757 210587 102067 228309
rect 101757 210469 101773 210587
rect 101891 210469 101933 210587
rect 102051 210469 102067 210587
rect 101757 210427 102067 210469
rect 101757 210309 101773 210427
rect 101891 210309 101933 210427
rect 102051 210309 102067 210427
rect 101757 192587 102067 210309
rect 101757 192469 101773 192587
rect 101891 192469 101933 192587
rect 102051 192469 102067 192587
rect 101757 192427 102067 192469
rect 101757 192309 101773 192427
rect 101891 192309 101933 192427
rect 102051 192309 102067 192427
rect 101757 174587 102067 192309
rect 101757 174469 101773 174587
rect 101891 174469 101933 174587
rect 102051 174469 102067 174587
rect 101757 174427 102067 174469
rect 101757 174309 101773 174427
rect 101891 174309 101933 174427
rect 102051 174309 102067 174427
rect 101757 156587 102067 174309
rect 101757 156469 101773 156587
rect 101891 156469 101933 156587
rect 102051 156469 102067 156587
rect 101757 156427 102067 156469
rect 101757 156309 101773 156427
rect 101891 156309 101933 156427
rect 102051 156309 102067 156427
rect 101757 138587 102067 156309
rect 101757 138469 101773 138587
rect 101891 138469 101933 138587
rect 102051 138469 102067 138587
rect 101757 138427 102067 138469
rect 101757 138309 101773 138427
rect 101891 138309 101933 138427
rect 102051 138309 102067 138427
rect 101757 120587 102067 138309
rect 101757 120469 101773 120587
rect 101891 120469 101933 120587
rect 102051 120469 102067 120587
rect 101757 120427 102067 120469
rect 101757 120309 101773 120427
rect 101891 120309 101933 120427
rect 102051 120309 102067 120427
rect 101757 102587 102067 120309
rect 101757 102469 101773 102587
rect 101891 102469 101933 102587
rect 102051 102469 102067 102587
rect 101757 102427 102067 102469
rect 101757 102309 101773 102427
rect 101891 102309 101933 102427
rect 102051 102309 102067 102427
rect 101757 84587 102067 102309
rect 101757 84469 101773 84587
rect 101891 84469 101933 84587
rect 102051 84469 102067 84587
rect 101757 84427 102067 84469
rect 101757 84309 101773 84427
rect 101891 84309 101933 84427
rect 102051 84309 102067 84427
rect 101757 66587 102067 84309
rect 101757 66469 101773 66587
rect 101891 66469 101933 66587
rect 102051 66469 102067 66587
rect 101757 66427 102067 66469
rect 101757 66309 101773 66427
rect 101891 66309 101933 66427
rect 102051 66309 102067 66427
rect 101757 48587 102067 66309
rect 101757 48469 101773 48587
rect 101891 48469 101933 48587
rect 102051 48469 102067 48587
rect 101757 48427 102067 48469
rect 101757 48309 101773 48427
rect 101891 48309 101933 48427
rect 102051 48309 102067 48427
rect 101757 30587 102067 48309
rect 101757 30469 101773 30587
rect 101891 30469 101933 30587
rect 102051 30469 102067 30587
rect 101757 30427 102067 30469
rect 101757 30309 101773 30427
rect 101891 30309 101933 30427
rect 102051 30309 102067 30427
rect 101757 12587 102067 30309
rect 101757 12469 101773 12587
rect 101891 12469 101933 12587
rect 102051 12469 102067 12587
rect 101757 12427 102067 12469
rect 101757 12309 101773 12427
rect 101891 12309 101933 12427
rect 102051 12309 102067 12427
rect 101757 -1613 102067 12309
rect 101757 -1731 101773 -1613
rect 101891 -1731 101933 -1613
rect 102051 -1731 102067 -1613
rect 101757 -1773 102067 -1731
rect 101757 -1891 101773 -1773
rect 101891 -1891 101933 -1773
rect 102051 -1891 102067 -1773
rect 101757 -1907 102067 -1891
rect 103617 338447 103927 354541
rect 103617 338329 103633 338447
rect 103751 338329 103793 338447
rect 103911 338329 103927 338447
rect 103617 338287 103927 338329
rect 103617 338169 103633 338287
rect 103751 338169 103793 338287
rect 103911 338169 103927 338287
rect 103617 320447 103927 338169
rect 103617 320329 103633 320447
rect 103751 320329 103793 320447
rect 103911 320329 103927 320447
rect 103617 320287 103927 320329
rect 103617 320169 103633 320287
rect 103751 320169 103793 320287
rect 103911 320169 103927 320287
rect 103617 302447 103927 320169
rect 103617 302329 103633 302447
rect 103751 302329 103793 302447
rect 103911 302329 103927 302447
rect 103617 302287 103927 302329
rect 103617 302169 103633 302287
rect 103751 302169 103793 302287
rect 103911 302169 103927 302287
rect 103617 284447 103927 302169
rect 103617 284329 103633 284447
rect 103751 284329 103793 284447
rect 103911 284329 103927 284447
rect 103617 284287 103927 284329
rect 103617 284169 103633 284287
rect 103751 284169 103793 284287
rect 103911 284169 103927 284287
rect 103617 266447 103927 284169
rect 103617 266329 103633 266447
rect 103751 266329 103793 266447
rect 103911 266329 103927 266447
rect 103617 266287 103927 266329
rect 103617 266169 103633 266287
rect 103751 266169 103793 266287
rect 103911 266169 103927 266287
rect 103617 248447 103927 266169
rect 103617 248329 103633 248447
rect 103751 248329 103793 248447
rect 103911 248329 103927 248447
rect 103617 248287 103927 248329
rect 103617 248169 103633 248287
rect 103751 248169 103793 248287
rect 103911 248169 103927 248287
rect 103617 230447 103927 248169
rect 103617 230329 103633 230447
rect 103751 230329 103793 230447
rect 103911 230329 103927 230447
rect 103617 230287 103927 230329
rect 103617 230169 103633 230287
rect 103751 230169 103793 230287
rect 103911 230169 103927 230287
rect 103617 212447 103927 230169
rect 103617 212329 103633 212447
rect 103751 212329 103793 212447
rect 103911 212329 103927 212447
rect 103617 212287 103927 212329
rect 103617 212169 103633 212287
rect 103751 212169 103793 212287
rect 103911 212169 103927 212287
rect 103617 194447 103927 212169
rect 103617 194329 103633 194447
rect 103751 194329 103793 194447
rect 103911 194329 103927 194447
rect 103617 194287 103927 194329
rect 103617 194169 103633 194287
rect 103751 194169 103793 194287
rect 103911 194169 103927 194287
rect 103617 176447 103927 194169
rect 103617 176329 103633 176447
rect 103751 176329 103793 176447
rect 103911 176329 103927 176447
rect 103617 176287 103927 176329
rect 103617 176169 103633 176287
rect 103751 176169 103793 176287
rect 103911 176169 103927 176287
rect 103617 158447 103927 176169
rect 103617 158329 103633 158447
rect 103751 158329 103793 158447
rect 103911 158329 103927 158447
rect 103617 158287 103927 158329
rect 103617 158169 103633 158287
rect 103751 158169 103793 158287
rect 103911 158169 103927 158287
rect 103617 140447 103927 158169
rect 103617 140329 103633 140447
rect 103751 140329 103793 140447
rect 103911 140329 103927 140447
rect 103617 140287 103927 140329
rect 103617 140169 103633 140287
rect 103751 140169 103793 140287
rect 103911 140169 103927 140287
rect 103617 122447 103927 140169
rect 103617 122329 103633 122447
rect 103751 122329 103793 122447
rect 103911 122329 103927 122447
rect 103617 122287 103927 122329
rect 103617 122169 103633 122287
rect 103751 122169 103793 122287
rect 103911 122169 103927 122287
rect 103617 104447 103927 122169
rect 103617 104329 103633 104447
rect 103751 104329 103793 104447
rect 103911 104329 103927 104447
rect 103617 104287 103927 104329
rect 103617 104169 103633 104287
rect 103751 104169 103793 104287
rect 103911 104169 103927 104287
rect 103617 86447 103927 104169
rect 103617 86329 103633 86447
rect 103751 86329 103793 86447
rect 103911 86329 103927 86447
rect 103617 86287 103927 86329
rect 103617 86169 103633 86287
rect 103751 86169 103793 86287
rect 103911 86169 103927 86287
rect 103617 68447 103927 86169
rect 103617 68329 103633 68447
rect 103751 68329 103793 68447
rect 103911 68329 103927 68447
rect 103617 68287 103927 68329
rect 103617 68169 103633 68287
rect 103751 68169 103793 68287
rect 103911 68169 103927 68287
rect 103617 50447 103927 68169
rect 103617 50329 103633 50447
rect 103751 50329 103793 50447
rect 103911 50329 103927 50447
rect 103617 50287 103927 50329
rect 103617 50169 103633 50287
rect 103751 50169 103793 50287
rect 103911 50169 103927 50287
rect 103617 32447 103927 50169
rect 103617 32329 103633 32447
rect 103751 32329 103793 32447
rect 103911 32329 103927 32447
rect 103617 32287 103927 32329
rect 103617 32169 103633 32287
rect 103751 32169 103793 32287
rect 103911 32169 103927 32287
rect 103617 14447 103927 32169
rect 103617 14329 103633 14447
rect 103751 14329 103793 14447
rect 103911 14329 103927 14447
rect 103617 14287 103927 14329
rect 103617 14169 103633 14287
rect 103751 14169 103793 14287
rect 103911 14169 103927 14287
rect 103617 -2573 103927 14169
rect 103617 -2691 103633 -2573
rect 103751 -2691 103793 -2573
rect 103911 -2691 103927 -2573
rect 103617 -2733 103927 -2691
rect 103617 -2851 103633 -2733
rect 103751 -2851 103793 -2733
rect 103911 -2851 103927 -2733
rect 103617 -2867 103927 -2851
rect 105477 340307 105787 355501
rect 114477 355299 114787 355795
rect 114477 355181 114493 355299
rect 114611 355181 114653 355299
rect 114771 355181 114787 355299
rect 114477 355139 114787 355181
rect 114477 355021 114493 355139
rect 114611 355021 114653 355139
rect 114771 355021 114787 355139
rect 112617 354339 112927 354835
rect 112617 354221 112633 354339
rect 112751 354221 112793 354339
rect 112911 354221 112927 354339
rect 112617 354179 112927 354221
rect 112617 354061 112633 354179
rect 112751 354061 112793 354179
rect 112911 354061 112927 354179
rect 110757 353379 111067 353875
rect 110757 353261 110773 353379
rect 110891 353261 110933 353379
rect 111051 353261 111067 353379
rect 110757 353219 111067 353261
rect 110757 353101 110773 353219
rect 110891 353101 110933 353219
rect 111051 353101 111067 353219
rect 105477 340189 105493 340307
rect 105611 340189 105653 340307
rect 105771 340189 105787 340307
rect 105477 340147 105787 340189
rect 105477 340029 105493 340147
rect 105611 340029 105653 340147
rect 105771 340029 105787 340147
rect 105477 322307 105787 340029
rect 105477 322189 105493 322307
rect 105611 322189 105653 322307
rect 105771 322189 105787 322307
rect 105477 322147 105787 322189
rect 105477 322029 105493 322147
rect 105611 322029 105653 322147
rect 105771 322029 105787 322147
rect 105477 304307 105787 322029
rect 105477 304189 105493 304307
rect 105611 304189 105653 304307
rect 105771 304189 105787 304307
rect 105477 304147 105787 304189
rect 105477 304029 105493 304147
rect 105611 304029 105653 304147
rect 105771 304029 105787 304147
rect 105477 286307 105787 304029
rect 105477 286189 105493 286307
rect 105611 286189 105653 286307
rect 105771 286189 105787 286307
rect 105477 286147 105787 286189
rect 105477 286029 105493 286147
rect 105611 286029 105653 286147
rect 105771 286029 105787 286147
rect 105477 268307 105787 286029
rect 105477 268189 105493 268307
rect 105611 268189 105653 268307
rect 105771 268189 105787 268307
rect 105477 268147 105787 268189
rect 105477 268029 105493 268147
rect 105611 268029 105653 268147
rect 105771 268029 105787 268147
rect 105477 250307 105787 268029
rect 105477 250189 105493 250307
rect 105611 250189 105653 250307
rect 105771 250189 105787 250307
rect 105477 250147 105787 250189
rect 105477 250029 105493 250147
rect 105611 250029 105653 250147
rect 105771 250029 105787 250147
rect 105477 232307 105787 250029
rect 105477 232189 105493 232307
rect 105611 232189 105653 232307
rect 105771 232189 105787 232307
rect 105477 232147 105787 232189
rect 105477 232029 105493 232147
rect 105611 232029 105653 232147
rect 105771 232029 105787 232147
rect 105477 214307 105787 232029
rect 105477 214189 105493 214307
rect 105611 214189 105653 214307
rect 105771 214189 105787 214307
rect 105477 214147 105787 214189
rect 105477 214029 105493 214147
rect 105611 214029 105653 214147
rect 105771 214029 105787 214147
rect 105477 196307 105787 214029
rect 105477 196189 105493 196307
rect 105611 196189 105653 196307
rect 105771 196189 105787 196307
rect 105477 196147 105787 196189
rect 105477 196029 105493 196147
rect 105611 196029 105653 196147
rect 105771 196029 105787 196147
rect 105477 178307 105787 196029
rect 105477 178189 105493 178307
rect 105611 178189 105653 178307
rect 105771 178189 105787 178307
rect 105477 178147 105787 178189
rect 105477 178029 105493 178147
rect 105611 178029 105653 178147
rect 105771 178029 105787 178147
rect 105477 160307 105787 178029
rect 105477 160189 105493 160307
rect 105611 160189 105653 160307
rect 105771 160189 105787 160307
rect 105477 160147 105787 160189
rect 105477 160029 105493 160147
rect 105611 160029 105653 160147
rect 105771 160029 105787 160147
rect 105477 142307 105787 160029
rect 105477 142189 105493 142307
rect 105611 142189 105653 142307
rect 105771 142189 105787 142307
rect 105477 142147 105787 142189
rect 105477 142029 105493 142147
rect 105611 142029 105653 142147
rect 105771 142029 105787 142147
rect 105477 124307 105787 142029
rect 105477 124189 105493 124307
rect 105611 124189 105653 124307
rect 105771 124189 105787 124307
rect 105477 124147 105787 124189
rect 105477 124029 105493 124147
rect 105611 124029 105653 124147
rect 105771 124029 105787 124147
rect 105477 106307 105787 124029
rect 105477 106189 105493 106307
rect 105611 106189 105653 106307
rect 105771 106189 105787 106307
rect 105477 106147 105787 106189
rect 105477 106029 105493 106147
rect 105611 106029 105653 106147
rect 105771 106029 105787 106147
rect 105477 88307 105787 106029
rect 105477 88189 105493 88307
rect 105611 88189 105653 88307
rect 105771 88189 105787 88307
rect 105477 88147 105787 88189
rect 105477 88029 105493 88147
rect 105611 88029 105653 88147
rect 105771 88029 105787 88147
rect 105477 70307 105787 88029
rect 105477 70189 105493 70307
rect 105611 70189 105653 70307
rect 105771 70189 105787 70307
rect 105477 70147 105787 70189
rect 105477 70029 105493 70147
rect 105611 70029 105653 70147
rect 105771 70029 105787 70147
rect 105477 52307 105787 70029
rect 105477 52189 105493 52307
rect 105611 52189 105653 52307
rect 105771 52189 105787 52307
rect 105477 52147 105787 52189
rect 105477 52029 105493 52147
rect 105611 52029 105653 52147
rect 105771 52029 105787 52147
rect 105477 34307 105787 52029
rect 105477 34189 105493 34307
rect 105611 34189 105653 34307
rect 105771 34189 105787 34307
rect 105477 34147 105787 34189
rect 105477 34029 105493 34147
rect 105611 34029 105653 34147
rect 105771 34029 105787 34147
rect 105477 16307 105787 34029
rect 105477 16189 105493 16307
rect 105611 16189 105653 16307
rect 105771 16189 105787 16307
rect 105477 16147 105787 16189
rect 105477 16029 105493 16147
rect 105611 16029 105653 16147
rect 105771 16029 105787 16147
rect 96477 -3171 96493 -3053
rect 96611 -3171 96653 -3053
rect 96771 -3171 96787 -3053
rect 96477 -3213 96787 -3171
rect 96477 -3331 96493 -3213
rect 96611 -3331 96653 -3213
rect 96771 -3331 96787 -3213
rect 96477 -3827 96787 -3331
rect 105477 -3533 105787 16029
rect 108897 352419 109207 352915
rect 108897 352301 108913 352419
rect 109031 352301 109073 352419
rect 109191 352301 109207 352419
rect 108897 352259 109207 352301
rect 108897 352141 108913 352259
rect 109031 352141 109073 352259
rect 109191 352141 109207 352259
rect 108897 343727 109207 352141
rect 108897 343609 108913 343727
rect 109031 343609 109073 343727
rect 109191 343609 109207 343727
rect 108897 343567 109207 343609
rect 108897 343449 108913 343567
rect 109031 343449 109073 343567
rect 109191 343449 109207 343567
rect 108897 325727 109207 343449
rect 108897 325609 108913 325727
rect 109031 325609 109073 325727
rect 109191 325609 109207 325727
rect 108897 325567 109207 325609
rect 108897 325449 108913 325567
rect 109031 325449 109073 325567
rect 109191 325449 109207 325567
rect 108897 307727 109207 325449
rect 108897 307609 108913 307727
rect 109031 307609 109073 307727
rect 109191 307609 109207 307727
rect 108897 307567 109207 307609
rect 108897 307449 108913 307567
rect 109031 307449 109073 307567
rect 109191 307449 109207 307567
rect 108897 289727 109207 307449
rect 108897 289609 108913 289727
rect 109031 289609 109073 289727
rect 109191 289609 109207 289727
rect 108897 289567 109207 289609
rect 108897 289449 108913 289567
rect 109031 289449 109073 289567
rect 109191 289449 109207 289567
rect 108897 271727 109207 289449
rect 108897 271609 108913 271727
rect 109031 271609 109073 271727
rect 109191 271609 109207 271727
rect 108897 271567 109207 271609
rect 108897 271449 108913 271567
rect 109031 271449 109073 271567
rect 109191 271449 109207 271567
rect 108897 253727 109207 271449
rect 108897 253609 108913 253727
rect 109031 253609 109073 253727
rect 109191 253609 109207 253727
rect 108897 253567 109207 253609
rect 108897 253449 108913 253567
rect 109031 253449 109073 253567
rect 109191 253449 109207 253567
rect 108897 235727 109207 253449
rect 108897 235609 108913 235727
rect 109031 235609 109073 235727
rect 109191 235609 109207 235727
rect 108897 235567 109207 235609
rect 108897 235449 108913 235567
rect 109031 235449 109073 235567
rect 109191 235449 109207 235567
rect 108897 217727 109207 235449
rect 108897 217609 108913 217727
rect 109031 217609 109073 217727
rect 109191 217609 109207 217727
rect 108897 217567 109207 217609
rect 108897 217449 108913 217567
rect 109031 217449 109073 217567
rect 109191 217449 109207 217567
rect 108897 199727 109207 217449
rect 108897 199609 108913 199727
rect 109031 199609 109073 199727
rect 109191 199609 109207 199727
rect 108897 199567 109207 199609
rect 108897 199449 108913 199567
rect 109031 199449 109073 199567
rect 109191 199449 109207 199567
rect 108897 181727 109207 199449
rect 108897 181609 108913 181727
rect 109031 181609 109073 181727
rect 109191 181609 109207 181727
rect 108897 181567 109207 181609
rect 108897 181449 108913 181567
rect 109031 181449 109073 181567
rect 109191 181449 109207 181567
rect 108897 163727 109207 181449
rect 108897 163609 108913 163727
rect 109031 163609 109073 163727
rect 109191 163609 109207 163727
rect 108897 163567 109207 163609
rect 108897 163449 108913 163567
rect 109031 163449 109073 163567
rect 109191 163449 109207 163567
rect 108897 145727 109207 163449
rect 108897 145609 108913 145727
rect 109031 145609 109073 145727
rect 109191 145609 109207 145727
rect 108897 145567 109207 145609
rect 108897 145449 108913 145567
rect 109031 145449 109073 145567
rect 109191 145449 109207 145567
rect 108897 127727 109207 145449
rect 108897 127609 108913 127727
rect 109031 127609 109073 127727
rect 109191 127609 109207 127727
rect 108897 127567 109207 127609
rect 108897 127449 108913 127567
rect 109031 127449 109073 127567
rect 109191 127449 109207 127567
rect 108897 109727 109207 127449
rect 108897 109609 108913 109727
rect 109031 109609 109073 109727
rect 109191 109609 109207 109727
rect 108897 109567 109207 109609
rect 108897 109449 108913 109567
rect 109031 109449 109073 109567
rect 109191 109449 109207 109567
rect 108897 91727 109207 109449
rect 108897 91609 108913 91727
rect 109031 91609 109073 91727
rect 109191 91609 109207 91727
rect 108897 91567 109207 91609
rect 108897 91449 108913 91567
rect 109031 91449 109073 91567
rect 109191 91449 109207 91567
rect 108897 73727 109207 91449
rect 108897 73609 108913 73727
rect 109031 73609 109073 73727
rect 109191 73609 109207 73727
rect 108897 73567 109207 73609
rect 108897 73449 108913 73567
rect 109031 73449 109073 73567
rect 109191 73449 109207 73567
rect 108897 55727 109207 73449
rect 108897 55609 108913 55727
rect 109031 55609 109073 55727
rect 109191 55609 109207 55727
rect 108897 55567 109207 55609
rect 108897 55449 108913 55567
rect 109031 55449 109073 55567
rect 109191 55449 109207 55567
rect 108897 37727 109207 55449
rect 108897 37609 108913 37727
rect 109031 37609 109073 37727
rect 109191 37609 109207 37727
rect 108897 37567 109207 37609
rect 108897 37449 108913 37567
rect 109031 37449 109073 37567
rect 109191 37449 109207 37567
rect 108897 19727 109207 37449
rect 108897 19609 108913 19727
rect 109031 19609 109073 19727
rect 109191 19609 109207 19727
rect 108897 19567 109207 19609
rect 108897 19449 108913 19567
rect 109031 19449 109073 19567
rect 109191 19449 109207 19567
rect 108897 1727 109207 19449
rect 108897 1609 108913 1727
rect 109031 1609 109073 1727
rect 109191 1609 109207 1727
rect 108897 1567 109207 1609
rect 108897 1449 108913 1567
rect 109031 1449 109073 1567
rect 109191 1449 109207 1567
rect 108897 -173 109207 1449
rect 108897 -291 108913 -173
rect 109031 -291 109073 -173
rect 109191 -291 109207 -173
rect 108897 -333 109207 -291
rect 108897 -451 108913 -333
rect 109031 -451 109073 -333
rect 109191 -451 109207 -333
rect 108897 -947 109207 -451
rect 110757 345587 111067 353101
rect 110757 345469 110773 345587
rect 110891 345469 110933 345587
rect 111051 345469 111067 345587
rect 110757 345427 111067 345469
rect 110757 345309 110773 345427
rect 110891 345309 110933 345427
rect 111051 345309 111067 345427
rect 110757 327587 111067 345309
rect 110757 327469 110773 327587
rect 110891 327469 110933 327587
rect 111051 327469 111067 327587
rect 110757 327427 111067 327469
rect 110757 327309 110773 327427
rect 110891 327309 110933 327427
rect 111051 327309 111067 327427
rect 110757 309587 111067 327309
rect 110757 309469 110773 309587
rect 110891 309469 110933 309587
rect 111051 309469 111067 309587
rect 110757 309427 111067 309469
rect 110757 309309 110773 309427
rect 110891 309309 110933 309427
rect 111051 309309 111067 309427
rect 110757 291587 111067 309309
rect 110757 291469 110773 291587
rect 110891 291469 110933 291587
rect 111051 291469 111067 291587
rect 110757 291427 111067 291469
rect 110757 291309 110773 291427
rect 110891 291309 110933 291427
rect 111051 291309 111067 291427
rect 110757 273587 111067 291309
rect 110757 273469 110773 273587
rect 110891 273469 110933 273587
rect 111051 273469 111067 273587
rect 110757 273427 111067 273469
rect 110757 273309 110773 273427
rect 110891 273309 110933 273427
rect 111051 273309 111067 273427
rect 110757 255587 111067 273309
rect 110757 255469 110773 255587
rect 110891 255469 110933 255587
rect 111051 255469 111067 255587
rect 110757 255427 111067 255469
rect 110757 255309 110773 255427
rect 110891 255309 110933 255427
rect 111051 255309 111067 255427
rect 110757 237587 111067 255309
rect 110757 237469 110773 237587
rect 110891 237469 110933 237587
rect 111051 237469 111067 237587
rect 110757 237427 111067 237469
rect 110757 237309 110773 237427
rect 110891 237309 110933 237427
rect 111051 237309 111067 237427
rect 110757 219587 111067 237309
rect 110757 219469 110773 219587
rect 110891 219469 110933 219587
rect 111051 219469 111067 219587
rect 110757 219427 111067 219469
rect 110757 219309 110773 219427
rect 110891 219309 110933 219427
rect 111051 219309 111067 219427
rect 110757 201587 111067 219309
rect 110757 201469 110773 201587
rect 110891 201469 110933 201587
rect 111051 201469 111067 201587
rect 110757 201427 111067 201469
rect 110757 201309 110773 201427
rect 110891 201309 110933 201427
rect 111051 201309 111067 201427
rect 110757 183587 111067 201309
rect 110757 183469 110773 183587
rect 110891 183469 110933 183587
rect 111051 183469 111067 183587
rect 110757 183427 111067 183469
rect 110757 183309 110773 183427
rect 110891 183309 110933 183427
rect 111051 183309 111067 183427
rect 110757 165587 111067 183309
rect 110757 165469 110773 165587
rect 110891 165469 110933 165587
rect 111051 165469 111067 165587
rect 110757 165427 111067 165469
rect 110757 165309 110773 165427
rect 110891 165309 110933 165427
rect 111051 165309 111067 165427
rect 110757 147587 111067 165309
rect 110757 147469 110773 147587
rect 110891 147469 110933 147587
rect 111051 147469 111067 147587
rect 110757 147427 111067 147469
rect 110757 147309 110773 147427
rect 110891 147309 110933 147427
rect 111051 147309 111067 147427
rect 110757 129587 111067 147309
rect 110757 129469 110773 129587
rect 110891 129469 110933 129587
rect 111051 129469 111067 129587
rect 110757 129427 111067 129469
rect 110757 129309 110773 129427
rect 110891 129309 110933 129427
rect 111051 129309 111067 129427
rect 110757 111587 111067 129309
rect 110757 111469 110773 111587
rect 110891 111469 110933 111587
rect 111051 111469 111067 111587
rect 110757 111427 111067 111469
rect 110757 111309 110773 111427
rect 110891 111309 110933 111427
rect 111051 111309 111067 111427
rect 110757 93587 111067 111309
rect 110757 93469 110773 93587
rect 110891 93469 110933 93587
rect 111051 93469 111067 93587
rect 110757 93427 111067 93469
rect 110757 93309 110773 93427
rect 110891 93309 110933 93427
rect 111051 93309 111067 93427
rect 110757 75587 111067 93309
rect 110757 75469 110773 75587
rect 110891 75469 110933 75587
rect 111051 75469 111067 75587
rect 110757 75427 111067 75469
rect 110757 75309 110773 75427
rect 110891 75309 110933 75427
rect 111051 75309 111067 75427
rect 110757 57587 111067 75309
rect 110757 57469 110773 57587
rect 110891 57469 110933 57587
rect 111051 57469 111067 57587
rect 110757 57427 111067 57469
rect 110757 57309 110773 57427
rect 110891 57309 110933 57427
rect 111051 57309 111067 57427
rect 110757 39587 111067 57309
rect 110757 39469 110773 39587
rect 110891 39469 110933 39587
rect 111051 39469 111067 39587
rect 110757 39427 111067 39469
rect 110757 39309 110773 39427
rect 110891 39309 110933 39427
rect 111051 39309 111067 39427
rect 110757 21587 111067 39309
rect 110757 21469 110773 21587
rect 110891 21469 110933 21587
rect 111051 21469 111067 21587
rect 110757 21427 111067 21469
rect 110757 21309 110773 21427
rect 110891 21309 110933 21427
rect 111051 21309 111067 21427
rect 110757 3587 111067 21309
rect 110757 3469 110773 3587
rect 110891 3469 110933 3587
rect 111051 3469 111067 3587
rect 110757 3427 111067 3469
rect 110757 3309 110773 3427
rect 110891 3309 110933 3427
rect 111051 3309 111067 3427
rect 110757 -1133 111067 3309
rect 110757 -1251 110773 -1133
rect 110891 -1251 110933 -1133
rect 111051 -1251 111067 -1133
rect 110757 -1293 111067 -1251
rect 110757 -1411 110773 -1293
rect 110891 -1411 110933 -1293
rect 111051 -1411 111067 -1293
rect 110757 -1907 111067 -1411
rect 112617 347447 112927 354061
rect 112617 347329 112633 347447
rect 112751 347329 112793 347447
rect 112911 347329 112927 347447
rect 112617 347287 112927 347329
rect 112617 347169 112633 347287
rect 112751 347169 112793 347287
rect 112911 347169 112927 347287
rect 112617 329447 112927 347169
rect 112617 329329 112633 329447
rect 112751 329329 112793 329447
rect 112911 329329 112927 329447
rect 112617 329287 112927 329329
rect 112617 329169 112633 329287
rect 112751 329169 112793 329287
rect 112911 329169 112927 329287
rect 112617 311447 112927 329169
rect 112617 311329 112633 311447
rect 112751 311329 112793 311447
rect 112911 311329 112927 311447
rect 112617 311287 112927 311329
rect 112617 311169 112633 311287
rect 112751 311169 112793 311287
rect 112911 311169 112927 311287
rect 112617 293447 112927 311169
rect 112617 293329 112633 293447
rect 112751 293329 112793 293447
rect 112911 293329 112927 293447
rect 112617 293287 112927 293329
rect 112617 293169 112633 293287
rect 112751 293169 112793 293287
rect 112911 293169 112927 293287
rect 112617 275447 112927 293169
rect 112617 275329 112633 275447
rect 112751 275329 112793 275447
rect 112911 275329 112927 275447
rect 112617 275287 112927 275329
rect 112617 275169 112633 275287
rect 112751 275169 112793 275287
rect 112911 275169 112927 275287
rect 112617 257447 112927 275169
rect 112617 257329 112633 257447
rect 112751 257329 112793 257447
rect 112911 257329 112927 257447
rect 112617 257287 112927 257329
rect 112617 257169 112633 257287
rect 112751 257169 112793 257287
rect 112911 257169 112927 257287
rect 112617 239447 112927 257169
rect 112617 239329 112633 239447
rect 112751 239329 112793 239447
rect 112911 239329 112927 239447
rect 112617 239287 112927 239329
rect 112617 239169 112633 239287
rect 112751 239169 112793 239287
rect 112911 239169 112927 239287
rect 112617 221447 112927 239169
rect 112617 221329 112633 221447
rect 112751 221329 112793 221447
rect 112911 221329 112927 221447
rect 112617 221287 112927 221329
rect 112617 221169 112633 221287
rect 112751 221169 112793 221287
rect 112911 221169 112927 221287
rect 112617 203447 112927 221169
rect 112617 203329 112633 203447
rect 112751 203329 112793 203447
rect 112911 203329 112927 203447
rect 112617 203287 112927 203329
rect 112617 203169 112633 203287
rect 112751 203169 112793 203287
rect 112911 203169 112927 203287
rect 112617 185447 112927 203169
rect 112617 185329 112633 185447
rect 112751 185329 112793 185447
rect 112911 185329 112927 185447
rect 112617 185287 112927 185329
rect 112617 185169 112633 185287
rect 112751 185169 112793 185287
rect 112911 185169 112927 185287
rect 112617 167447 112927 185169
rect 112617 167329 112633 167447
rect 112751 167329 112793 167447
rect 112911 167329 112927 167447
rect 112617 167287 112927 167329
rect 112617 167169 112633 167287
rect 112751 167169 112793 167287
rect 112911 167169 112927 167287
rect 112617 149447 112927 167169
rect 112617 149329 112633 149447
rect 112751 149329 112793 149447
rect 112911 149329 112927 149447
rect 112617 149287 112927 149329
rect 112617 149169 112633 149287
rect 112751 149169 112793 149287
rect 112911 149169 112927 149287
rect 112617 131447 112927 149169
rect 112617 131329 112633 131447
rect 112751 131329 112793 131447
rect 112911 131329 112927 131447
rect 112617 131287 112927 131329
rect 112617 131169 112633 131287
rect 112751 131169 112793 131287
rect 112911 131169 112927 131287
rect 112617 113447 112927 131169
rect 112617 113329 112633 113447
rect 112751 113329 112793 113447
rect 112911 113329 112927 113447
rect 112617 113287 112927 113329
rect 112617 113169 112633 113287
rect 112751 113169 112793 113287
rect 112911 113169 112927 113287
rect 112617 95447 112927 113169
rect 112617 95329 112633 95447
rect 112751 95329 112793 95447
rect 112911 95329 112927 95447
rect 112617 95287 112927 95329
rect 112617 95169 112633 95287
rect 112751 95169 112793 95287
rect 112911 95169 112927 95287
rect 112617 77447 112927 95169
rect 112617 77329 112633 77447
rect 112751 77329 112793 77447
rect 112911 77329 112927 77447
rect 112617 77287 112927 77329
rect 112617 77169 112633 77287
rect 112751 77169 112793 77287
rect 112911 77169 112927 77287
rect 112617 59447 112927 77169
rect 112617 59329 112633 59447
rect 112751 59329 112793 59447
rect 112911 59329 112927 59447
rect 112617 59287 112927 59329
rect 112617 59169 112633 59287
rect 112751 59169 112793 59287
rect 112911 59169 112927 59287
rect 112617 41447 112927 59169
rect 112617 41329 112633 41447
rect 112751 41329 112793 41447
rect 112911 41329 112927 41447
rect 112617 41287 112927 41329
rect 112617 41169 112633 41287
rect 112751 41169 112793 41287
rect 112911 41169 112927 41287
rect 112617 23447 112927 41169
rect 112617 23329 112633 23447
rect 112751 23329 112793 23447
rect 112911 23329 112927 23447
rect 112617 23287 112927 23329
rect 112617 23169 112633 23287
rect 112751 23169 112793 23287
rect 112911 23169 112927 23287
rect 112617 5447 112927 23169
rect 112617 5329 112633 5447
rect 112751 5329 112793 5447
rect 112911 5329 112927 5447
rect 112617 5287 112927 5329
rect 112617 5169 112633 5287
rect 112751 5169 112793 5287
rect 112911 5169 112927 5287
rect 112617 -2093 112927 5169
rect 112617 -2211 112633 -2093
rect 112751 -2211 112793 -2093
rect 112911 -2211 112927 -2093
rect 112617 -2253 112927 -2211
rect 112617 -2371 112633 -2253
rect 112751 -2371 112793 -2253
rect 112911 -2371 112927 -2253
rect 112617 -2867 112927 -2371
rect 114477 349307 114787 355021
rect 123477 355779 123787 355795
rect 123477 355661 123493 355779
rect 123611 355661 123653 355779
rect 123771 355661 123787 355779
rect 123477 355619 123787 355661
rect 123477 355501 123493 355619
rect 123611 355501 123653 355619
rect 123771 355501 123787 355619
rect 121617 354819 121927 354835
rect 121617 354701 121633 354819
rect 121751 354701 121793 354819
rect 121911 354701 121927 354819
rect 121617 354659 121927 354701
rect 121617 354541 121633 354659
rect 121751 354541 121793 354659
rect 121911 354541 121927 354659
rect 119757 353859 120067 353875
rect 119757 353741 119773 353859
rect 119891 353741 119933 353859
rect 120051 353741 120067 353859
rect 119757 353699 120067 353741
rect 119757 353581 119773 353699
rect 119891 353581 119933 353699
rect 120051 353581 120067 353699
rect 114477 349189 114493 349307
rect 114611 349189 114653 349307
rect 114771 349189 114787 349307
rect 114477 349147 114787 349189
rect 114477 349029 114493 349147
rect 114611 349029 114653 349147
rect 114771 349029 114787 349147
rect 114477 331307 114787 349029
rect 114477 331189 114493 331307
rect 114611 331189 114653 331307
rect 114771 331189 114787 331307
rect 114477 331147 114787 331189
rect 114477 331029 114493 331147
rect 114611 331029 114653 331147
rect 114771 331029 114787 331147
rect 114477 313307 114787 331029
rect 114477 313189 114493 313307
rect 114611 313189 114653 313307
rect 114771 313189 114787 313307
rect 114477 313147 114787 313189
rect 114477 313029 114493 313147
rect 114611 313029 114653 313147
rect 114771 313029 114787 313147
rect 114477 295307 114787 313029
rect 114477 295189 114493 295307
rect 114611 295189 114653 295307
rect 114771 295189 114787 295307
rect 114477 295147 114787 295189
rect 114477 295029 114493 295147
rect 114611 295029 114653 295147
rect 114771 295029 114787 295147
rect 114477 277307 114787 295029
rect 114477 277189 114493 277307
rect 114611 277189 114653 277307
rect 114771 277189 114787 277307
rect 114477 277147 114787 277189
rect 114477 277029 114493 277147
rect 114611 277029 114653 277147
rect 114771 277029 114787 277147
rect 114477 259307 114787 277029
rect 114477 259189 114493 259307
rect 114611 259189 114653 259307
rect 114771 259189 114787 259307
rect 114477 259147 114787 259189
rect 114477 259029 114493 259147
rect 114611 259029 114653 259147
rect 114771 259029 114787 259147
rect 114477 241307 114787 259029
rect 114477 241189 114493 241307
rect 114611 241189 114653 241307
rect 114771 241189 114787 241307
rect 114477 241147 114787 241189
rect 114477 241029 114493 241147
rect 114611 241029 114653 241147
rect 114771 241029 114787 241147
rect 114477 223307 114787 241029
rect 114477 223189 114493 223307
rect 114611 223189 114653 223307
rect 114771 223189 114787 223307
rect 114477 223147 114787 223189
rect 114477 223029 114493 223147
rect 114611 223029 114653 223147
rect 114771 223029 114787 223147
rect 114477 205307 114787 223029
rect 114477 205189 114493 205307
rect 114611 205189 114653 205307
rect 114771 205189 114787 205307
rect 114477 205147 114787 205189
rect 114477 205029 114493 205147
rect 114611 205029 114653 205147
rect 114771 205029 114787 205147
rect 114477 187307 114787 205029
rect 114477 187189 114493 187307
rect 114611 187189 114653 187307
rect 114771 187189 114787 187307
rect 114477 187147 114787 187189
rect 114477 187029 114493 187147
rect 114611 187029 114653 187147
rect 114771 187029 114787 187147
rect 114477 169307 114787 187029
rect 114477 169189 114493 169307
rect 114611 169189 114653 169307
rect 114771 169189 114787 169307
rect 114477 169147 114787 169189
rect 114477 169029 114493 169147
rect 114611 169029 114653 169147
rect 114771 169029 114787 169147
rect 114477 151307 114787 169029
rect 114477 151189 114493 151307
rect 114611 151189 114653 151307
rect 114771 151189 114787 151307
rect 114477 151147 114787 151189
rect 114477 151029 114493 151147
rect 114611 151029 114653 151147
rect 114771 151029 114787 151147
rect 114477 133307 114787 151029
rect 114477 133189 114493 133307
rect 114611 133189 114653 133307
rect 114771 133189 114787 133307
rect 114477 133147 114787 133189
rect 114477 133029 114493 133147
rect 114611 133029 114653 133147
rect 114771 133029 114787 133147
rect 114477 115307 114787 133029
rect 114477 115189 114493 115307
rect 114611 115189 114653 115307
rect 114771 115189 114787 115307
rect 114477 115147 114787 115189
rect 114477 115029 114493 115147
rect 114611 115029 114653 115147
rect 114771 115029 114787 115147
rect 114477 97307 114787 115029
rect 114477 97189 114493 97307
rect 114611 97189 114653 97307
rect 114771 97189 114787 97307
rect 114477 97147 114787 97189
rect 114477 97029 114493 97147
rect 114611 97029 114653 97147
rect 114771 97029 114787 97147
rect 114477 79307 114787 97029
rect 114477 79189 114493 79307
rect 114611 79189 114653 79307
rect 114771 79189 114787 79307
rect 114477 79147 114787 79189
rect 114477 79029 114493 79147
rect 114611 79029 114653 79147
rect 114771 79029 114787 79147
rect 114477 61307 114787 79029
rect 114477 61189 114493 61307
rect 114611 61189 114653 61307
rect 114771 61189 114787 61307
rect 114477 61147 114787 61189
rect 114477 61029 114493 61147
rect 114611 61029 114653 61147
rect 114771 61029 114787 61147
rect 114477 43307 114787 61029
rect 114477 43189 114493 43307
rect 114611 43189 114653 43307
rect 114771 43189 114787 43307
rect 114477 43147 114787 43189
rect 114477 43029 114493 43147
rect 114611 43029 114653 43147
rect 114771 43029 114787 43147
rect 114477 25307 114787 43029
rect 114477 25189 114493 25307
rect 114611 25189 114653 25307
rect 114771 25189 114787 25307
rect 114477 25147 114787 25189
rect 114477 25029 114493 25147
rect 114611 25029 114653 25147
rect 114771 25029 114787 25147
rect 114477 7307 114787 25029
rect 114477 7189 114493 7307
rect 114611 7189 114653 7307
rect 114771 7189 114787 7307
rect 114477 7147 114787 7189
rect 114477 7029 114493 7147
rect 114611 7029 114653 7147
rect 114771 7029 114787 7147
rect 105477 -3651 105493 -3533
rect 105611 -3651 105653 -3533
rect 105771 -3651 105787 -3533
rect 105477 -3693 105787 -3651
rect 105477 -3811 105493 -3693
rect 105611 -3811 105653 -3693
rect 105771 -3811 105787 -3693
rect 105477 -3827 105787 -3811
rect 114477 -3053 114787 7029
rect 117897 352899 118207 352915
rect 117897 352781 117913 352899
rect 118031 352781 118073 352899
rect 118191 352781 118207 352899
rect 117897 352739 118207 352781
rect 117897 352621 117913 352739
rect 118031 352621 118073 352739
rect 118191 352621 118207 352739
rect 117897 334727 118207 352621
rect 117897 334609 117913 334727
rect 118031 334609 118073 334727
rect 118191 334609 118207 334727
rect 117897 334567 118207 334609
rect 117897 334449 117913 334567
rect 118031 334449 118073 334567
rect 118191 334449 118207 334567
rect 117897 316727 118207 334449
rect 117897 316609 117913 316727
rect 118031 316609 118073 316727
rect 118191 316609 118207 316727
rect 117897 316567 118207 316609
rect 117897 316449 117913 316567
rect 118031 316449 118073 316567
rect 118191 316449 118207 316567
rect 117897 298727 118207 316449
rect 117897 298609 117913 298727
rect 118031 298609 118073 298727
rect 118191 298609 118207 298727
rect 117897 298567 118207 298609
rect 117897 298449 117913 298567
rect 118031 298449 118073 298567
rect 118191 298449 118207 298567
rect 117897 280727 118207 298449
rect 117897 280609 117913 280727
rect 118031 280609 118073 280727
rect 118191 280609 118207 280727
rect 117897 280567 118207 280609
rect 117897 280449 117913 280567
rect 118031 280449 118073 280567
rect 118191 280449 118207 280567
rect 117897 262727 118207 280449
rect 117897 262609 117913 262727
rect 118031 262609 118073 262727
rect 118191 262609 118207 262727
rect 117897 262567 118207 262609
rect 117897 262449 117913 262567
rect 118031 262449 118073 262567
rect 118191 262449 118207 262567
rect 117897 244727 118207 262449
rect 117897 244609 117913 244727
rect 118031 244609 118073 244727
rect 118191 244609 118207 244727
rect 117897 244567 118207 244609
rect 117897 244449 117913 244567
rect 118031 244449 118073 244567
rect 118191 244449 118207 244567
rect 117897 226727 118207 244449
rect 117897 226609 117913 226727
rect 118031 226609 118073 226727
rect 118191 226609 118207 226727
rect 117897 226567 118207 226609
rect 117897 226449 117913 226567
rect 118031 226449 118073 226567
rect 118191 226449 118207 226567
rect 117897 208727 118207 226449
rect 117897 208609 117913 208727
rect 118031 208609 118073 208727
rect 118191 208609 118207 208727
rect 117897 208567 118207 208609
rect 117897 208449 117913 208567
rect 118031 208449 118073 208567
rect 118191 208449 118207 208567
rect 117897 190727 118207 208449
rect 117897 190609 117913 190727
rect 118031 190609 118073 190727
rect 118191 190609 118207 190727
rect 117897 190567 118207 190609
rect 117897 190449 117913 190567
rect 118031 190449 118073 190567
rect 118191 190449 118207 190567
rect 117897 172727 118207 190449
rect 117897 172609 117913 172727
rect 118031 172609 118073 172727
rect 118191 172609 118207 172727
rect 117897 172567 118207 172609
rect 117897 172449 117913 172567
rect 118031 172449 118073 172567
rect 118191 172449 118207 172567
rect 117897 154727 118207 172449
rect 117897 154609 117913 154727
rect 118031 154609 118073 154727
rect 118191 154609 118207 154727
rect 117897 154567 118207 154609
rect 117897 154449 117913 154567
rect 118031 154449 118073 154567
rect 118191 154449 118207 154567
rect 117897 136727 118207 154449
rect 117897 136609 117913 136727
rect 118031 136609 118073 136727
rect 118191 136609 118207 136727
rect 117897 136567 118207 136609
rect 117897 136449 117913 136567
rect 118031 136449 118073 136567
rect 118191 136449 118207 136567
rect 117897 118727 118207 136449
rect 117897 118609 117913 118727
rect 118031 118609 118073 118727
rect 118191 118609 118207 118727
rect 117897 118567 118207 118609
rect 117897 118449 117913 118567
rect 118031 118449 118073 118567
rect 118191 118449 118207 118567
rect 117897 100727 118207 118449
rect 117897 100609 117913 100727
rect 118031 100609 118073 100727
rect 118191 100609 118207 100727
rect 117897 100567 118207 100609
rect 117897 100449 117913 100567
rect 118031 100449 118073 100567
rect 118191 100449 118207 100567
rect 117897 82727 118207 100449
rect 117897 82609 117913 82727
rect 118031 82609 118073 82727
rect 118191 82609 118207 82727
rect 117897 82567 118207 82609
rect 117897 82449 117913 82567
rect 118031 82449 118073 82567
rect 118191 82449 118207 82567
rect 117897 64727 118207 82449
rect 117897 64609 117913 64727
rect 118031 64609 118073 64727
rect 118191 64609 118207 64727
rect 117897 64567 118207 64609
rect 117897 64449 117913 64567
rect 118031 64449 118073 64567
rect 118191 64449 118207 64567
rect 117897 46727 118207 64449
rect 117897 46609 117913 46727
rect 118031 46609 118073 46727
rect 118191 46609 118207 46727
rect 117897 46567 118207 46609
rect 117897 46449 117913 46567
rect 118031 46449 118073 46567
rect 118191 46449 118207 46567
rect 117897 28727 118207 46449
rect 117897 28609 117913 28727
rect 118031 28609 118073 28727
rect 118191 28609 118207 28727
rect 117897 28567 118207 28609
rect 117897 28449 117913 28567
rect 118031 28449 118073 28567
rect 118191 28449 118207 28567
rect 117897 10727 118207 28449
rect 117897 10609 117913 10727
rect 118031 10609 118073 10727
rect 118191 10609 118207 10727
rect 117897 10567 118207 10609
rect 117897 10449 117913 10567
rect 118031 10449 118073 10567
rect 118191 10449 118207 10567
rect 117897 -653 118207 10449
rect 117897 -771 117913 -653
rect 118031 -771 118073 -653
rect 118191 -771 118207 -653
rect 117897 -813 118207 -771
rect 117897 -931 117913 -813
rect 118031 -931 118073 -813
rect 118191 -931 118207 -813
rect 117897 -947 118207 -931
rect 119757 336587 120067 353581
rect 119757 336469 119773 336587
rect 119891 336469 119933 336587
rect 120051 336469 120067 336587
rect 119757 336427 120067 336469
rect 119757 336309 119773 336427
rect 119891 336309 119933 336427
rect 120051 336309 120067 336427
rect 119757 318587 120067 336309
rect 119757 318469 119773 318587
rect 119891 318469 119933 318587
rect 120051 318469 120067 318587
rect 119757 318427 120067 318469
rect 119757 318309 119773 318427
rect 119891 318309 119933 318427
rect 120051 318309 120067 318427
rect 119757 300587 120067 318309
rect 119757 300469 119773 300587
rect 119891 300469 119933 300587
rect 120051 300469 120067 300587
rect 119757 300427 120067 300469
rect 119757 300309 119773 300427
rect 119891 300309 119933 300427
rect 120051 300309 120067 300427
rect 119757 282587 120067 300309
rect 119757 282469 119773 282587
rect 119891 282469 119933 282587
rect 120051 282469 120067 282587
rect 119757 282427 120067 282469
rect 119757 282309 119773 282427
rect 119891 282309 119933 282427
rect 120051 282309 120067 282427
rect 119757 264587 120067 282309
rect 119757 264469 119773 264587
rect 119891 264469 119933 264587
rect 120051 264469 120067 264587
rect 119757 264427 120067 264469
rect 119757 264309 119773 264427
rect 119891 264309 119933 264427
rect 120051 264309 120067 264427
rect 119757 246587 120067 264309
rect 119757 246469 119773 246587
rect 119891 246469 119933 246587
rect 120051 246469 120067 246587
rect 119757 246427 120067 246469
rect 119757 246309 119773 246427
rect 119891 246309 119933 246427
rect 120051 246309 120067 246427
rect 119757 228587 120067 246309
rect 119757 228469 119773 228587
rect 119891 228469 119933 228587
rect 120051 228469 120067 228587
rect 119757 228427 120067 228469
rect 119757 228309 119773 228427
rect 119891 228309 119933 228427
rect 120051 228309 120067 228427
rect 119757 210587 120067 228309
rect 119757 210469 119773 210587
rect 119891 210469 119933 210587
rect 120051 210469 120067 210587
rect 119757 210427 120067 210469
rect 119757 210309 119773 210427
rect 119891 210309 119933 210427
rect 120051 210309 120067 210427
rect 119757 192587 120067 210309
rect 119757 192469 119773 192587
rect 119891 192469 119933 192587
rect 120051 192469 120067 192587
rect 119757 192427 120067 192469
rect 119757 192309 119773 192427
rect 119891 192309 119933 192427
rect 120051 192309 120067 192427
rect 119757 174587 120067 192309
rect 119757 174469 119773 174587
rect 119891 174469 119933 174587
rect 120051 174469 120067 174587
rect 119757 174427 120067 174469
rect 119757 174309 119773 174427
rect 119891 174309 119933 174427
rect 120051 174309 120067 174427
rect 119757 156587 120067 174309
rect 119757 156469 119773 156587
rect 119891 156469 119933 156587
rect 120051 156469 120067 156587
rect 119757 156427 120067 156469
rect 119757 156309 119773 156427
rect 119891 156309 119933 156427
rect 120051 156309 120067 156427
rect 119757 138587 120067 156309
rect 119757 138469 119773 138587
rect 119891 138469 119933 138587
rect 120051 138469 120067 138587
rect 119757 138427 120067 138469
rect 119757 138309 119773 138427
rect 119891 138309 119933 138427
rect 120051 138309 120067 138427
rect 119757 120587 120067 138309
rect 119757 120469 119773 120587
rect 119891 120469 119933 120587
rect 120051 120469 120067 120587
rect 119757 120427 120067 120469
rect 119757 120309 119773 120427
rect 119891 120309 119933 120427
rect 120051 120309 120067 120427
rect 119757 102587 120067 120309
rect 119757 102469 119773 102587
rect 119891 102469 119933 102587
rect 120051 102469 120067 102587
rect 119757 102427 120067 102469
rect 119757 102309 119773 102427
rect 119891 102309 119933 102427
rect 120051 102309 120067 102427
rect 119757 84587 120067 102309
rect 119757 84469 119773 84587
rect 119891 84469 119933 84587
rect 120051 84469 120067 84587
rect 119757 84427 120067 84469
rect 119757 84309 119773 84427
rect 119891 84309 119933 84427
rect 120051 84309 120067 84427
rect 119757 66587 120067 84309
rect 119757 66469 119773 66587
rect 119891 66469 119933 66587
rect 120051 66469 120067 66587
rect 119757 66427 120067 66469
rect 119757 66309 119773 66427
rect 119891 66309 119933 66427
rect 120051 66309 120067 66427
rect 119757 48587 120067 66309
rect 119757 48469 119773 48587
rect 119891 48469 119933 48587
rect 120051 48469 120067 48587
rect 119757 48427 120067 48469
rect 119757 48309 119773 48427
rect 119891 48309 119933 48427
rect 120051 48309 120067 48427
rect 119757 30587 120067 48309
rect 119757 30469 119773 30587
rect 119891 30469 119933 30587
rect 120051 30469 120067 30587
rect 119757 30427 120067 30469
rect 119757 30309 119773 30427
rect 119891 30309 119933 30427
rect 120051 30309 120067 30427
rect 119757 12587 120067 30309
rect 119757 12469 119773 12587
rect 119891 12469 119933 12587
rect 120051 12469 120067 12587
rect 119757 12427 120067 12469
rect 119757 12309 119773 12427
rect 119891 12309 119933 12427
rect 120051 12309 120067 12427
rect 119757 -1613 120067 12309
rect 119757 -1731 119773 -1613
rect 119891 -1731 119933 -1613
rect 120051 -1731 120067 -1613
rect 119757 -1773 120067 -1731
rect 119757 -1891 119773 -1773
rect 119891 -1891 119933 -1773
rect 120051 -1891 120067 -1773
rect 119757 -1907 120067 -1891
rect 121617 338447 121927 354541
rect 121617 338329 121633 338447
rect 121751 338329 121793 338447
rect 121911 338329 121927 338447
rect 121617 338287 121927 338329
rect 121617 338169 121633 338287
rect 121751 338169 121793 338287
rect 121911 338169 121927 338287
rect 121617 320447 121927 338169
rect 121617 320329 121633 320447
rect 121751 320329 121793 320447
rect 121911 320329 121927 320447
rect 121617 320287 121927 320329
rect 121617 320169 121633 320287
rect 121751 320169 121793 320287
rect 121911 320169 121927 320287
rect 121617 302447 121927 320169
rect 121617 302329 121633 302447
rect 121751 302329 121793 302447
rect 121911 302329 121927 302447
rect 121617 302287 121927 302329
rect 121617 302169 121633 302287
rect 121751 302169 121793 302287
rect 121911 302169 121927 302287
rect 121617 284447 121927 302169
rect 121617 284329 121633 284447
rect 121751 284329 121793 284447
rect 121911 284329 121927 284447
rect 121617 284287 121927 284329
rect 121617 284169 121633 284287
rect 121751 284169 121793 284287
rect 121911 284169 121927 284287
rect 121617 266447 121927 284169
rect 121617 266329 121633 266447
rect 121751 266329 121793 266447
rect 121911 266329 121927 266447
rect 121617 266287 121927 266329
rect 121617 266169 121633 266287
rect 121751 266169 121793 266287
rect 121911 266169 121927 266287
rect 121617 248447 121927 266169
rect 121617 248329 121633 248447
rect 121751 248329 121793 248447
rect 121911 248329 121927 248447
rect 121617 248287 121927 248329
rect 121617 248169 121633 248287
rect 121751 248169 121793 248287
rect 121911 248169 121927 248287
rect 121617 230447 121927 248169
rect 121617 230329 121633 230447
rect 121751 230329 121793 230447
rect 121911 230329 121927 230447
rect 121617 230287 121927 230329
rect 121617 230169 121633 230287
rect 121751 230169 121793 230287
rect 121911 230169 121927 230287
rect 121617 212447 121927 230169
rect 121617 212329 121633 212447
rect 121751 212329 121793 212447
rect 121911 212329 121927 212447
rect 121617 212287 121927 212329
rect 121617 212169 121633 212287
rect 121751 212169 121793 212287
rect 121911 212169 121927 212287
rect 121617 194447 121927 212169
rect 121617 194329 121633 194447
rect 121751 194329 121793 194447
rect 121911 194329 121927 194447
rect 121617 194287 121927 194329
rect 121617 194169 121633 194287
rect 121751 194169 121793 194287
rect 121911 194169 121927 194287
rect 121617 176447 121927 194169
rect 121617 176329 121633 176447
rect 121751 176329 121793 176447
rect 121911 176329 121927 176447
rect 121617 176287 121927 176329
rect 121617 176169 121633 176287
rect 121751 176169 121793 176287
rect 121911 176169 121927 176287
rect 121617 158447 121927 176169
rect 121617 158329 121633 158447
rect 121751 158329 121793 158447
rect 121911 158329 121927 158447
rect 121617 158287 121927 158329
rect 121617 158169 121633 158287
rect 121751 158169 121793 158287
rect 121911 158169 121927 158287
rect 121617 140447 121927 158169
rect 121617 140329 121633 140447
rect 121751 140329 121793 140447
rect 121911 140329 121927 140447
rect 121617 140287 121927 140329
rect 121617 140169 121633 140287
rect 121751 140169 121793 140287
rect 121911 140169 121927 140287
rect 121617 122447 121927 140169
rect 121617 122329 121633 122447
rect 121751 122329 121793 122447
rect 121911 122329 121927 122447
rect 121617 122287 121927 122329
rect 121617 122169 121633 122287
rect 121751 122169 121793 122287
rect 121911 122169 121927 122287
rect 121617 104447 121927 122169
rect 121617 104329 121633 104447
rect 121751 104329 121793 104447
rect 121911 104329 121927 104447
rect 121617 104287 121927 104329
rect 121617 104169 121633 104287
rect 121751 104169 121793 104287
rect 121911 104169 121927 104287
rect 121617 86447 121927 104169
rect 121617 86329 121633 86447
rect 121751 86329 121793 86447
rect 121911 86329 121927 86447
rect 121617 86287 121927 86329
rect 121617 86169 121633 86287
rect 121751 86169 121793 86287
rect 121911 86169 121927 86287
rect 121617 68447 121927 86169
rect 121617 68329 121633 68447
rect 121751 68329 121793 68447
rect 121911 68329 121927 68447
rect 121617 68287 121927 68329
rect 121617 68169 121633 68287
rect 121751 68169 121793 68287
rect 121911 68169 121927 68287
rect 121617 50447 121927 68169
rect 121617 50329 121633 50447
rect 121751 50329 121793 50447
rect 121911 50329 121927 50447
rect 121617 50287 121927 50329
rect 121617 50169 121633 50287
rect 121751 50169 121793 50287
rect 121911 50169 121927 50287
rect 121617 32447 121927 50169
rect 121617 32329 121633 32447
rect 121751 32329 121793 32447
rect 121911 32329 121927 32447
rect 121617 32287 121927 32329
rect 121617 32169 121633 32287
rect 121751 32169 121793 32287
rect 121911 32169 121927 32287
rect 121617 14447 121927 32169
rect 121617 14329 121633 14447
rect 121751 14329 121793 14447
rect 121911 14329 121927 14447
rect 121617 14287 121927 14329
rect 121617 14169 121633 14287
rect 121751 14169 121793 14287
rect 121911 14169 121927 14287
rect 121617 -2573 121927 14169
rect 121617 -2691 121633 -2573
rect 121751 -2691 121793 -2573
rect 121911 -2691 121927 -2573
rect 121617 -2733 121927 -2691
rect 121617 -2851 121633 -2733
rect 121751 -2851 121793 -2733
rect 121911 -2851 121927 -2733
rect 121617 -2867 121927 -2851
rect 123477 340307 123787 355501
rect 132477 355299 132787 355795
rect 132477 355181 132493 355299
rect 132611 355181 132653 355299
rect 132771 355181 132787 355299
rect 132477 355139 132787 355181
rect 132477 355021 132493 355139
rect 132611 355021 132653 355139
rect 132771 355021 132787 355139
rect 130617 354339 130927 354835
rect 130617 354221 130633 354339
rect 130751 354221 130793 354339
rect 130911 354221 130927 354339
rect 130617 354179 130927 354221
rect 130617 354061 130633 354179
rect 130751 354061 130793 354179
rect 130911 354061 130927 354179
rect 128757 353379 129067 353875
rect 128757 353261 128773 353379
rect 128891 353261 128933 353379
rect 129051 353261 129067 353379
rect 128757 353219 129067 353261
rect 128757 353101 128773 353219
rect 128891 353101 128933 353219
rect 129051 353101 129067 353219
rect 123477 340189 123493 340307
rect 123611 340189 123653 340307
rect 123771 340189 123787 340307
rect 123477 340147 123787 340189
rect 123477 340029 123493 340147
rect 123611 340029 123653 340147
rect 123771 340029 123787 340147
rect 123477 322307 123787 340029
rect 123477 322189 123493 322307
rect 123611 322189 123653 322307
rect 123771 322189 123787 322307
rect 123477 322147 123787 322189
rect 123477 322029 123493 322147
rect 123611 322029 123653 322147
rect 123771 322029 123787 322147
rect 123477 304307 123787 322029
rect 123477 304189 123493 304307
rect 123611 304189 123653 304307
rect 123771 304189 123787 304307
rect 123477 304147 123787 304189
rect 123477 304029 123493 304147
rect 123611 304029 123653 304147
rect 123771 304029 123787 304147
rect 123477 286307 123787 304029
rect 123477 286189 123493 286307
rect 123611 286189 123653 286307
rect 123771 286189 123787 286307
rect 123477 286147 123787 286189
rect 123477 286029 123493 286147
rect 123611 286029 123653 286147
rect 123771 286029 123787 286147
rect 123477 268307 123787 286029
rect 123477 268189 123493 268307
rect 123611 268189 123653 268307
rect 123771 268189 123787 268307
rect 123477 268147 123787 268189
rect 123477 268029 123493 268147
rect 123611 268029 123653 268147
rect 123771 268029 123787 268147
rect 123477 250307 123787 268029
rect 123477 250189 123493 250307
rect 123611 250189 123653 250307
rect 123771 250189 123787 250307
rect 123477 250147 123787 250189
rect 123477 250029 123493 250147
rect 123611 250029 123653 250147
rect 123771 250029 123787 250147
rect 123477 232307 123787 250029
rect 123477 232189 123493 232307
rect 123611 232189 123653 232307
rect 123771 232189 123787 232307
rect 123477 232147 123787 232189
rect 123477 232029 123493 232147
rect 123611 232029 123653 232147
rect 123771 232029 123787 232147
rect 123477 214307 123787 232029
rect 123477 214189 123493 214307
rect 123611 214189 123653 214307
rect 123771 214189 123787 214307
rect 123477 214147 123787 214189
rect 123477 214029 123493 214147
rect 123611 214029 123653 214147
rect 123771 214029 123787 214147
rect 123477 196307 123787 214029
rect 123477 196189 123493 196307
rect 123611 196189 123653 196307
rect 123771 196189 123787 196307
rect 123477 196147 123787 196189
rect 123477 196029 123493 196147
rect 123611 196029 123653 196147
rect 123771 196029 123787 196147
rect 123477 178307 123787 196029
rect 123477 178189 123493 178307
rect 123611 178189 123653 178307
rect 123771 178189 123787 178307
rect 123477 178147 123787 178189
rect 123477 178029 123493 178147
rect 123611 178029 123653 178147
rect 123771 178029 123787 178147
rect 123477 160307 123787 178029
rect 123477 160189 123493 160307
rect 123611 160189 123653 160307
rect 123771 160189 123787 160307
rect 123477 160147 123787 160189
rect 123477 160029 123493 160147
rect 123611 160029 123653 160147
rect 123771 160029 123787 160147
rect 123477 142307 123787 160029
rect 123477 142189 123493 142307
rect 123611 142189 123653 142307
rect 123771 142189 123787 142307
rect 123477 142147 123787 142189
rect 123477 142029 123493 142147
rect 123611 142029 123653 142147
rect 123771 142029 123787 142147
rect 123477 124307 123787 142029
rect 123477 124189 123493 124307
rect 123611 124189 123653 124307
rect 123771 124189 123787 124307
rect 123477 124147 123787 124189
rect 123477 124029 123493 124147
rect 123611 124029 123653 124147
rect 123771 124029 123787 124147
rect 123477 106307 123787 124029
rect 123477 106189 123493 106307
rect 123611 106189 123653 106307
rect 123771 106189 123787 106307
rect 123477 106147 123787 106189
rect 123477 106029 123493 106147
rect 123611 106029 123653 106147
rect 123771 106029 123787 106147
rect 123477 88307 123787 106029
rect 123477 88189 123493 88307
rect 123611 88189 123653 88307
rect 123771 88189 123787 88307
rect 123477 88147 123787 88189
rect 123477 88029 123493 88147
rect 123611 88029 123653 88147
rect 123771 88029 123787 88147
rect 123477 70307 123787 88029
rect 123477 70189 123493 70307
rect 123611 70189 123653 70307
rect 123771 70189 123787 70307
rect 123477 70147 123787 70189
rect 123477 70029 123493 70147
rect 123611 70029 123653 70147
rect 123771 70029 123787 70147
rect 123477 52307 123787 70029
rect 123477 52189 123493 52307
rect 123611 52189 123653 52307
rect 123771 52189 123787 52307
rect 123477 52147 123787 52189
rect 123477 52029 123493 52147
rect 123611 52029 123653 52147
rect 123771 52029 123787 52147
rect 123477 34307 123787 52029
rect 123477 34189 123493 34307
rect 123611 34189 123653 34307
rect 123771 34189 123787 34307
rect 123477 34147 123787 34189
rect 123477 34029 123493 34147
rect 123611 34029 123653 34147
rect 123771 34029 123787 34147
rect 123477 16307 123787 34029
rect 123477 16189 123493 16307
rect 123611 16189 123653 16307
rect 123771 16189 123787 16307
rect 123477 16147 123787 16189
rect 123477 16029 123493 16147
rect 123611 16029 123653 16147
rect 123771 16029 123787 16147
rect 114477 -3171 114493 -3053
rect 114611 -3171 114653 -3053
rect 114771 -3171 114787 -3053
rect 114477 -3213 114787 -3171
rect 114477 -3331 114493 -3213
rect 114611 -3331 114653 -3213
rect 114771 -3331 114787 -3213
rect 114477 -3827 114787 -3331
rect 123477 -3533 123787 16029
rect 126897 352419 127207 352915
rect 126897 352301 126913 352419
rect 127031 352301 127073 352419
rect 127191 352301 127207 352419
rect 126897 352259 127207 352301
rect 126897 352141 126913 352259
rect 127031 352141 127073 352259
rect 127191 352141 127207 352259
rect 126897 343727 127207 352141
rect 126897 343609 126913 343727
rect 127031 343609 127073 343727
rect 127191 343609 127207 343727
rect 126897 343567 127207 343609
rect 126897 343449 126913 343567
rect 127031 343449 127073 343567
rect 127191 343449 127207 343567
rect 126897 325727 127207 343449
rect 126897 325609 126913 325727
rect 127031 325609 127073 325727
rect 127191 325609 127207 325727
rect 126897 325567 127207 325609
rect 126897 325449 126913 325567
rect 127031 325449 127073 325567
rect 127191 325449 127207 325567
rect 126897 307727 127207 325449
rect 126897 307609 126913 307727
rect 127031 307609 127073 307727
rect 127191 307609 127207 307727
rect 126897 307567 127207 307609
rect 126897 307449 126913 307567
rect 127031 307449 127073 307567
rect 127191 307449 127207 307567
rect 126897 289727 127207 307449
rect 126897 289609 126913 289727
rect 127031 289609 127073 289727
rect 127191 289609 127207 289727
rect 126897 289567 127207 289609
rect 126897 289449 126913 289567
rect 127031 289449 127073 289567
rect 127191 289449 127207 289567
rect 126897 271727 127207 289449
rect 126897 271609 126913 271727
rect 127031 271609 127073 271727
rect 127191 271609 127207 271727
rect 126897 271567 127207 271609
rect 126897 271449 126913 271567
rect 127031 271449 127073 271567
rect 127191 271449 127207 271567
rect 126897 253727 127207 271449
rect 126897 253609 126913 253727
rect 127031 253609 127073 253727
rect 127191 253609 127207 253727
rect 126897 253567 127207 253609
rect 126897 253449 126913 253567
rect 127031 253449 127073 253567
rect 127191 253449 127207 253567
rect 126897 235727 127207 253449
rect 126897 235609 126913 235727
rect 127031 235609 127073 235727
rect 127191 235609 127207 235727
rect 126897 235567 127207 235609
rect 126897 235449 126913 235567
rect 127031 235449 127073 235567
rect 127191 235449 127207 235567
rect 126897 217727 127207 235449
rect 126897 217609 126913 217727
rect 127031 217609 127073 217727
rect 127191 217609 127207 217727
rect 126897 217567 127207 217609
rect 126897 217449 126913 217567
rect 127031 217449 127073 217567
rect 127191 217449 127207 217567
rect 126897 199727 127207 217449
rect 126897 199609 126913 199727
rect 127031 199609 127073 199727
rect 127191 199609 127207 199727
rect 126897 199567 127207 199609
rect 126897 199449 126913 199567
rect 127031 199449 127073 199567
rect 127191 199449 127207 199567
rect 126897 181727 127207 199449
rect 126897 181609 126913 181727
rect 127031 181609 127073 181727
rect 127191 181609 127207 181727
rect 126897 181567 127207 181609
rect 126897 181449 126913 181567
rect 127031 181449 127073 181567
rect 127191 181449 127207 181567
rect 126897 163727 127207 181449
rect 126897 163609 126913 163727
rect 127031 163609 127073 163727
rect 127191 163609 127207 163727
rect 126897 163567 127207 163609
rect 126897 163449 126913 163567
rect 127031 163449 127073 163567
rect 127191 163449 127207 163567
rect 126897 145727 127207 163449
rect 126897 145609 126913 145727
rect 127031 145609 127073 145727
rect 127191 145609 127207 145727
rect 126897 145567 127207 145609
rect 126897 145449 126913 145567
rect 127031 145449 127073 145567
rect 127191 145449 127207 145567
rect 126897 127727 127207 145449
rect 126897 127609 126913 127727
rect 127031 127609 127073 127727
rect 127191 127609 127207 127727
rect 126897 127567 127207 127609
rect 126897 127449 126913 127567
rect 127031 127449 127073 127567
rect 127191 127449 127207 127567
rect 126897 109727 127207 127449
rect 126897 109609 126913 109727
rect 127031 109609 127073 109727
rect 127191 109609 127207 109727
rect 126897 109567 127207 109609
rect 126897 109449 126913 109567
rect 127031 109449 127073 109567
rect 127191 109449 127207 109567
rect 126897 91727 127207 109449
rect 126897 91609 126913 91727
rect 127031 91609 127073 91727
rect 127191 91609 127207 91727
rect 126897 91567 127207 91609
rect 126897 91449 126913 91567
rect 127031 91449 127073 91567
rect 127191 91449 127207 91567
rect 126897 73727 127207 91449
rect 126897 73609 126913 73727
rect 127031 73609 127073 73727
rect 127191 73609 127207 73727
rect 126897 73567 127207 73609
rect 126897 73449 126913 73567
rect 127031 73449 127073 73567
rect 127191 73449 127207 73567
rect 126897 55727 127207 73449
rect 126897 55609 126913 55727
rect 127031 55609 127073 55727
rect 127191 55609 127207 55727
rect 126897 55567 127207 55609
rect 126897 55449 126913 55567
rect 127031 55449 127073 55567
rect 127191 55449 127207 55567
rect 126897 37727 127207 55449
rect 126897 37609 126913 37727
rect 127031 37609 127073 37727
rect 127191 37609 127207 37727
rect 126897 37567 127207 37609
rect 126897 37449 126913 37567
rect 127031 37449 127073 37567
rect 127191 37449 127207 37567
rect 126897 19727 127207 37449
rect 126897 19609 126913 19727
rect 127031 19609 127073 19727
rect 127191 19609 127207 19727
rect 126897 19567 127207 19609
rect 126897 19449 126913 19567
rect 127031 19449 127073 19567
rect 127191 19449 127207 19567
rect 126897 1727 127207 19449
rect 126897 1609 126913 1727
rect 127031 1609 127073 1727
rect 127191 1609 127207 1727
rect 126897 1567 127207 1609
rect 126897 1449 126913 1567
rect 127031 1449 127073 1567
rect 127191 1449 127207 1567
rect 126897 -173 127207 1449
rect 126897 -291 126913 -173
rect 127031 -291 127073 -173
rect 127191 -291 127207 -173
rect 126897 -333 127207 -291
rect 126897 -451 126913 -333
rect 127031 -451 127073 -333
rect 127191 -451 127207 -333
rect 126897 -947 127207 -451
rect 128757 345587 129067 353101
rect 128757 345469 128773 345587
rect 128891 345469 128933 345587
rect 129051 345469 129067 345587
rect 128757 345427 129067 345469
rect 128757 345309 128773 345427
rect 128891 345309 128933 345427
rect 129051 345309 129067 345427
rect 128757 327587 129067 345309
rect 128757 327469 128773 327587
rect 128891 327469 128933 327587
rect 129051 327469 129067 327587
rect 128757 327427 129067 327469
rect 128757 327309 128773 327427
rect 128891 327309 128933 327427
rect 129051 327309 129067 327427
rect 128757 309587 129067 327309
rect 128757 309469 128773 309587
rect 128891 309469 128933 309587
rect 129051 309469 129067 309587
rect 128757 309427 129067 309469
rect 128757 309309 128773 309427
rect 128891 309309 128933 309427
rect 129051 309309 129067 309427
rect 128757 291587 129067 309309
rect 128757 291469 128773 291587
rect 128891 291469 128933 291587
rect 129051 291469 129067 291587
rect 128757 291427 129067 291469
rect 128757 291309 128773 291427
rect 128891 291309 128933 291427
rect 129051 291309 129067 291427
rect 128757 273587 129067 291309
rect 128757 273469 128773 273587
rect 128891 273469 128933 273587
rect 129051 273469 129067 273587
rect 128757 273427 129067 273469
rect 128757 273309 128773 273427
rect 128891 273309 128933 273427
rect 129051 273309 129067 273427
rect 128757 255587 129067 273309
rect 128757 255469 128773 255587
rect 128891 255469 128933 255587
rect 129051 255469 129067 255587
rect 128757 255427 129067 255469
rect 128757 255309 128773 255427
rect 128891 255309 128933 255427
rect 129051 255309 129067 255427
rect 128757 237587 129067 255309
rect 128757 237469 128773 237587
rect 128891 237469 128933 237587
rect 129051 237469 129067 237587
rect 128757 237427 129067 237469
rect 128757 237309 128773 237427
rect 128891 237309 128933 237427
rect 129051 237309 129067 237427
rect 128757 219587 129067 237309
rect 128757 219469 128773 219587
rect 128891 219469 128933 219587
rect 129051 219469 129067 219587
rect 128757 219427 129067 219469
rect 128757 219309 128773 219427
rect 128891 219309 128933 219427
rect 129051 219309 129067 219427
rect 128757 201587 129067 219309
rect 128757 201469 128773 201587
rect 128891 201469 128933 201587
rect 129051 201469 129067 201587
rect 128757 201427 129067 201469
rect 128757 201309 128773 201427
rect 128891 201309 128933 201427
rect 129051 201309 129067 201427
rect 128757 183587 129067 201309
rect 128757 183469 128773 183587
rect 128891 183469 128933 183587
rect 129051 183469 129067 183587
rect 128757 183427 129067 183469
rect 128757 183309 128773 183427
rect 128891 183309 128933 183427
rect 129051 183309 129067 183427
rect 128757 165587 129067 183309
rect 128757 165469 128773 165587
rect 128891 165469 128933 165587
rect 129051 165469 129067 165587
rect 128757 165427 129067 165469
rect 128757 165309 128773 165427
rect 128891 165309 128933 165427
rect 129051 165309 129067 165427
rect 128757 147587 129067 165309
rect 128757 147469 128773 147587
rect 128891 147469 128933 147587
rect 129051 147469 129067 147587
rect 128757 147427 129067 147469
rect 128757 147309 128773 147427
rect 128891 147309 128933 147427
rect 129051 147309 129067 147427
rect 128757 129587 129067 147309
rect 128757 129469 128773 129587
rect 128891 129469 128933 129587
rect 129051 129469 129067 129587
rect 128757 129427 129067 129469
rect 128757 129309 128773 129427
rect 128891 129309 128933 129427
rect 129051 129309 129067 129427
rect 128757 111587 129067 129309
rect 128757 111469 128773 111587
rect 128891 111469 128933 111587
rect 129051 111469 129067 111587
rect 128757 111427 129067 111469
rect 128757 111309 128773 111427
rect 128891 111309 128933 111427
rect 129051 111309 129067 111427
rect 128757 93587 129067 111309
rect 128757 93469 128773 93587
rect 128891 93469 128933 93587
rect 129051 93469 129067 93587
rect 128757 93427 129067 93469
rect 128757 93309 128773 93427
rect 128891 93309 128933 93427
rect 129051 93309 129067 93427
rect 128757 75587 129067 93309
rect 128757 75469 128773 75587
rect 128891 75469 128933 75587
rect 129051 75469 129067 75587
rect 128757 75427 129067 75469
rect 128757 75309 128773 75427
rect 128891 75309 128933 75427
rect 129051 75309 129067 75427
rect 128757 57587 129067 75309
rect 128757 57469 128773 57587
rect 128891 57469 128933 57587
rect 129051 57469 129067 57587
rect 128757 57427 129067 57469
rect 128757 57309 128773 57427
rect 128891 57309 128933 57427
rect 129051 57309 129067 57427
rect 128757 39587 129067 57309
rect 128757 39469 128773 39587
rect 128891 39469 128933 39587
rect 129051 39469 129067 39587
rect 128757 39427 129067 39469
rect 128757 39309 128773 39427
rect 128891 39309 128933 39427
rect 129051 39309 129067 39427
rect 128757 21587 129067 39309
rect 128757 21469 128773 21587
rect 128891 21469 128933 21587
rect 129051 21469 129067 21587
rect 128757 21427 129067 21469
rect 128757 21309 128773 21427
rect 128891 21309 128933 21427
rect 129051 21309 129067 21427
rect 128757 3587 129067 21309
rect 128757 3469 128773 3587
rect 128891 3469 128933 3587
rect 129051 3469 129067 3587
rect 128757 3427 129067 3469
rect 128757 3309 128773 3427
rect 128891 3309 128933 3427
rect 129051 3309 129067 3427
rect 128757 -1133 129067 3309
rect 128757 -1251 128773 -1133
rect 128891 -1251 128933 -1133
rect 129051 -1251 129067 -1133
rect 128757 -1293 129067 -1251
rect 128757 -1411 128773 -1293
rect 128891 -1411 128933 -1293
rect 129051 -1411 129067 -1293
rect 128757 -1907 129067 -1411
rect 130617 347447 130927 354061
rect 130617 347329 130633 347447
rect 130751 347329 130793 347447
rect 130911 347329 130927 347447
rect 130617 347287 130927 347329
rect 130617 347169 130633 347287
rect 130751 347169 130793 347287
rect 130911 347169 130927 347287
rect 130617 329447 130927 347169
rect 130617 329329 130633 329447
rect 130751 329329 130793 329447
rect 130911 329329 130927 329447
rect 130617 329287 130927 329329
rect 130617 329169 130633 329287
rect 130751 329169 130793 329287
rect 130911 329169 130927 329287
rect 130617 311447 130927 329169
rect 130617 311329 130633 311447
rect 130751 311329 130793 311447
rect 130911 311329 130927 311447
rect 130617 311287 130927 311329
rect 130617 311169 130633 311287
rect 130751 311169 130793 311287
rect 130911 311169 130927 311287
rect 130617 293447 130927 311169
rect 130617 293329 130633 293447
rect 130751 293329 130793 293447
rect 130911 293329 130927 293447
rect 130617 293287 130927 293329
rect 130617 293169 130633 293287
rect 130751 293169 130793 293287
rect 130911 293169 130927 293287
rect 130617 275447 130927 293169
rect 130617 275329 130633 275447
rect 130751 275329 130793 275447
rect 130911 275329 130927 275447
rect 130617 275287 130927 275329
rect 130617 275169 130633 275287
rect 130751 275169 130793 275287
rect 130911 275169 130927 275287
rect 130617 257447 130927 275169
rect 130617 257329 130633 257447
rect 130751 257329 130793 257447
rect 130911 257329 130927 257447
rect 130617 257287 130927 257329
rect 130617 257169 130633 257287
rect 130751 257169 130793 257287
rect 130911 257169 130927 257287
rect 130617 239447 130927 257169
rect 130617 239329 130633 239447
rect 130751 239329 130793 239447
rect 130911 239329 130927 239447
rect 130617 239287 130927 239329
rect 130617 239169 130633 239287
rect 130751 239169 130793 239287
rect 130911 239169 130927 239287
rect 130617 221447 130927 239169
rect 130617 221329 130633 221447
rect 130751 221329 130793 221447
rect 130911 221329 130927 221447
rect 130617 221287 130927 221329
rect 130617 221169 130633 221287
rect 130751 221169 130793 221287
rect 130911 221169 130927 221287
rect 130617 203447 130927 221169
rect 130617 203329 130633 203447
rect 130751 203329 130793 203447
rect 130911 203329 130927 203447
rect 130617 203287 130927 203329
rect 130617 203169 130633 203287
rect 130751 203169 130793 203287
rect 130911 203169 130927 203287
rect 130617 185447 130927 203169
rect 130617 185329 130633 185447
rect 130751 185329 130793 185447
rect 130911 185329 130927 185447
rect 130617 185287 130927 185329
rect 130617 185169 130633 185287
rect 130751 185169 130793 185287
rect 130911 185169 130927 185287
rect 130617 167447 130927 185169
rect 130617 167329 130633 167447
rect 130751 167329 130793 167447
rect 130911 167329 130927 167447
rect 130617 167287 130927 167329
rect 130617 167169 130633 167287
rect 130751 167169 130793 167287
rect 130911 167169 130927 167287
rect 130617 149447 130927 167169
rect 130617 149329 130633 149447
rect 130751 149329 130793 149447
rect 130911 149329 130927 149447
rect 130617 149287 130927 149329
rect 130617 149169 130633 149287
rect 130751 149169 130793 149287
rect 130911 149169 130927 149287
rect 130617 131447 130927 149169
rect 130617 131329 130633 131447
rect 130751 131329 130793 131447
rect 130911 131329 130927 131447
rect 130617 131287 130927 131329
rect 130617 131169 130633 131287
rect 130751 131169 130793 131287
rect 130911 131169 130927 131287
rect 130617 113447 130927 131169
rect 130617 113329 130633 113447
rect 130751 113329 130793 113447
rect 130911 113329 130927 113447
rect 130617 113287 130927 113329
rect 130617 113169 130633 113287
rect 130751 113169 130793 113287
rect 130911 113169 130927 113287
rect 130617 95447 130927 113169
rect 130617 95329 130633 95447
rect 130751 95329 130793 95447
rect 130911 95329 130927 95447
rect 130617 95287 130927 95329
rect 130617 95169 130633 95287
rect 130751 95169 130793 95287
rect 130911 95169 130927 95287
rect 130617 77447 130927 95169
rect 130617 77329 130633 77447
rect 130751 77329 130793 77447
rect 130911 77329 130927 77447
rect 130617 77287 130927 77329
rect 130617 77169 130633 77287
rect 130751 77169 130793 77287
rect 130911 77169 130927 77287
rect 130617 59447 130927 77169
rect 130617 59329 130633 59447
rect 130751 59329 130793 59447
rect 130911 59329 130927 59447
rect 130617 59287 130927 59329
rect 130617 59169 130633 59287
rect 130751 59169 130793 59287
rect 130911 59169 130927 59287
rect 130617 41447 130927 59169
rect 130617 41329 130633 41447
rect 130751 41329 130793 41447
rect 130911 41329 130927 41447
rect 130617 41287 130927 41329
rect 130617 41169 130633 41287
rect 130751 41169 130793 41287
rect 130911 41169 130927 41287
rect 130617 23447 130927 41169
rect 130617 23329 130633 23447
rect 130751 23329 130793 23447
rect 130911 23329 130927 23447
rect 130617 23287 130927 23329
rect 130617 23169 130633 23287
rect 130751 23169 130793 23287
rect 130911 23169 130927 23287
rect 130617 5447 130927 23169
rect 130617 5329 130633 5447
rect 130751 5329 130793 5447
rect 130911 5329 130927 5447
rect 130617 5287 130927 5329
rect 130617 5169 130633 5287
rect 130751 5169 130793 5287
rect 130911 5169 130927 5287
rect 130617 -2093 130927 5169
rect 130617 -2211 130633 -2093
rect 130751 -2211 130793 -2093
rect 130911 -2211 130927 -2093
rect 130617 -2253 130927 -2211
rect 130617 -2371 130633 -2253
rect 130751 -2371 130793 -2253
rect 130911 -2371 130927 -2253
rect 130617 -2867 130927 -2371
rect 132477 349307 132787 355021
rect 141477 355779 141787 355795
rect 141477 355661 141493 355779
rect 141611 355661 141653 355779
rect 141771 355661 141787 355779
rect 141477 355619 141787 355661
rect 141477 355501 141493 355619
rect 141611 355501 141653 355619
rect 141771 355501 141787 355619
rect 139617 354819 139927 354835
rect 139617 354701 139633 354819
rect 139751 354701 139793 354819
rect 139911 354701 139927 354819
rect 139617 354659 139927 354701
rect 139617 354541 139633 354659
rect 139751 354541 139793 354659
rect 139911 354541 139927 354659
rect 137757 353859 138067 353875
rect 137757 353741 137773 353859
rect 137891 353741 137933 353859
rect 138051 353741 138067 353859
rect 137757 353699 138067 353741
rect 137757 353581 137773 353699
rect 137891 353581 137933 353699
rect 138051 353581 138067 353699
rect 132477 349189 132493 349307
rect 132611 349189 132653 349307
rect 132771 349189 132787 349307
rect 132477 349147 132787 349189
rect 132477 349029 132493 349147
rect 132611 349029 132653 349147
rect 132771 349029 132787 349147
rect 132477 331307 132787 349029
rect 132477 331189 132493 331307
rect 132611 331189 132653 331307
rect 132771 331189 132787 331307
rect 132477 331147 132787 331189
rect 132477 331029 132493 331147
rect 132611 331029 132653 331147
rect 132771 331029 132787 331147
rect 132477 313307 132787 331029
rect 132477 313189 132493 313307
rect 132611 313189 132653 313307
rect 132771 313189 132787 313307
rect 132477 313147 132787 313189
rect 132477 313029 132493 313147
rect 132611 313029 132653 313147
rect 132771 313029 132787 313147
rect 132477 295307 132787 313029
rect 132477 295189 132493 295307
rect 132611 295189 132653 295307
rect 132771 295189 132787 295307
rect 132477 295147 132787 295189
rect 132477 295029 132493 295147
rect 132611 295029 132653 295147
rect 132771 295029 132787 295147
rect 132477 277307 132787 295029
rect 132477 277189 132493 277307
rect 132611 277189 132653 277307
rect 132771 277189 132787 277307
rect 132477 277147 132787 277189
rect 132477 277029 132493 277147
rect 132611 277029 132653 277147
rect 132771 277029 132787 277147
rect 132477 259307 132787 277029
rect 132477 259189 132493 259307
rect 132611 259189 132653 259307
rect 132771 259189 132787 259307
rect 132477 259147 132787 259189
rect 132477 259029 132493 259147
rect 132611 259029 132653 259147
rect 132771 259029 132787 259147
rect 132477 241307 132787 259029
rect 132477 241189 132493 241307
rect 132611 241189 132653 241307
rect 132771 241189 132787 241307
rect 132477 241147 132787 241189
rect 132477 241029 132493 241147
rect 132611 241029 132653 241147
rect 132771 241029 132787 241147
rect 132477 223307 132787 241029
rect 132477 223189 132493 223307
rect 132611 223189 132653 223307
rect 132771 223189 132787 223307
rect 132477 223147 132787 223189
rect 132477 223029 132493 223147
rect 132611 223029 132653 223147
rect 132771 223029 132787 223147
rect 132477 205307 132787 223029
rect 132477 205189 132493 205307
rect 132611 205189 132653 205307
rect 132771 205189 132787 205307
rect 132477 205147 132787 205189
rect 132477 205029 132493 205147
rect 132611 205029 132653 205147
rect 132771 205029 132787 205147
rect 132477 187307 132787 205029
rect 132477 187189 132493 187307
rect 132611 187189 132653 187307
rect 132771 187189 132787 187307
rect 132477 187147 132787 187189
rect 132477 187029 132493 187147
rect 132611 187029 132653 187147
rect 132771 187029 132787 187147
rect 132477 169307 132787 187029
rect 132477 169189 132493 169307
rect 132611 169189 132653 169307
rect 132771 169189 132787 169307
rect 132477 169147 132787 169189
rect 132477 169029 132493 169147
rect 132611 169029 132653 169147
rect 132771 169029 132787 169147
rect 132477 151307 132787 169029
rect 132477 151189 132493 151307
rect 132611 151189 132653 151307
rect 132771 151189 132787 151307
rect 132477 151147 132787 151189
rect 132477 151029 132493 151147
rect 132611 151029 132653 151147
rect 132771 151029 132787 151147
rect 132477 133307 132787 151029
rect 132477 133189 132493 133307
rect 132611 133189 132653 133307
rect 132771 133189 132787 133307
rect 132477 133147 132787 133189
rect 132477 133029 132493 133147
rect 132611 133029 132653 133147
rect 132771 133029 132787 133147
rect 132477 115307 132787 133029
rect 132477 115189 132493 115307
rect 132611 115189 132653 115307
rect 132771 115189 132787 115307
rect 132477 115147 132787 115189
rect 132477 115029 132493 115147
rect 132611 115029 132653 115147
rect 132771 115029 132787 115147
rect 132477 97307 132787 115029
rect 132477 97189 132493 97307
rect 132611 97189 132653 97307
rect 132771 97189 132787 97307
rect 132477 97147 132787 97189
rect 132477 97029 132493 97147
rect 132611 97029 132653 97147
rect 132771 97029 132787 97147
rect 132477 79307 132787 97029
rect 132477 79189 132493 79307
rect 132611 79189 132653 79307
rect 132771 79189 132787 79307
rect 132477 79147 132787 79189
rect 132477 79029 132493 79147
rect 132611 79029 132653 79147
rect 132771 79029 132787 79147
rect 132477 61307 132787 79029
rect 132477 61189 132493 61307
rect 132611 61189 132653 61307
rect 132771 61189 132787 61307
rect 132477 61147 132787 61189
rect 132477 61029 132493 61147
rect 132611 61029 132653 61147
rect 132771 61029 132787 61147
rect 132477 43307 132787 61029
rect 132477 43189 132493 43307
rect 132611 43189 132653 43307
rect 132771 43189 132787 43307
rect 132477 43147 132787 43189
rect 132477 43029 132493 43147
rect 132611 43029 132653 43147
rect 132771 43029 132787 43147
rect 132477 25307 132787 43029
rect 132477 25189 132493 25307
rect 132611 25189 132653 25307
rect 132771 25189 132787 25307
rect 132477 25147 132787 25189
rect 132477 25029 132493 25147
rect 132611 25029 132653 25147
rect 132771 25029 132787 25147
rect 132477 7307 132787 25029
rect 132477 7189 132493 7307
rect 132611 7189 132653 7307
rect 132771 7189 132787 7307
rect 132477 7147 132787 7189
rect 132477 7029 132493 7147
rect 132611 7029 132653 7147
rect 132771 7029 132787 7147
rect 123477 -3651 123493 -3533
rect 123611 -3651 123653 -3533
rect 123771 -3651 123787 -3533
rect 123477 -3693 123787 -3651
rect 123477 -3811 123493 -3693
rect 123611 -3811 123653 -3693
rect 123771 -3811 123787 -3693
rect 123477 -3827 123787 -3811
rect 132477 -3053 132787 7029
rect 135897 352899 136207 352915
rect 135897 352781 135913 352899
rect 136031 352781 136073 352899
rect 136191 352781 136207 352899
rect 135897 352739 136207 352781
rect 135897 352621 135913 352739
rect 136031 352621 136073 352739
rect 136191 352621 136207 352739
rect 135897 334727 136207 352621
rect 135897 334609 135913 334727
rect 136031 334609 136073 334727
rect 136191 334609 136207 334727
rect 135897 334567 136207 334609
rect 135897 334449 135913 334567
rect 136031 334449 136073 334567
rect 136191 334449 136207 334567
rect 135897 316727 136207 334449
rect 135897 316609 135913 316727
rect 136031 316609 136073 316727
rect 136191 316609 136207 316727
rect 135897 316567 136207 316609
rect 135897 316449 135913 316567
rect 136031 316449 136073 316567
rect 136191 316449 136207 316567
rect 135897 298727 136207 316449
rect 135897 298609 135913 298727
rect 136031 298609 136073 298727
rect 136191 298609 136207 298727
rect 135897 298567 136207 298609
rect 135897 298449 135913 298567
rect 136031 298449 136073 298567
rect 136191 298449 136207 298567
rect 135897 280727 136207 298449
rect 135897 280609 135913 280727
rect 136031 280609 136073 280727
rect 136191 280609 136207 280727
rect 135897 280567 136207 280609
rect 135897 280449 135913 280567
rect 136031 280449 136073 280567
rect 136191 280449 136207 280567
rect 135897 262727 136207 280449
rect 135897 262609 135913 262727
rect 136031 262609 136073 262727
rect 136191 262609 136207 262727
rect 135897 262567 136207 262609
rect 135897 262449 135913 262567
rect 136031 262449 136073 262567
rect 136191 262449 136207 262567
rect 135897 244727 136207 262449
rect 135897 244609 135913 244727
rect 136031 244609 136073 244727
rect 136191 244609 136207 244727
rect 135897 244567 136207 244609
rect 135897 244449 135913 244567
rect 136031 244449 136073 244567
rect 136191 244449 136207 244567
rect 135897 226727 136207 244449
rect 135897 226609 135913 226727
rect 136031 226609 136073 226727
rect 136191 226609 136207 226727
rect 135897 226567 136207 226609
rect 135897 226449 135913 226567
rect 136031 226449 136073 226567
rect 136191 226449 136207 226567
rect 135897 208727 136207 226449
rect 135897 208609 135913 208727
rect 136031 208609 136073 208727
rect 136191 208609 136207 208727
rect 135897 208567 136207 208609
rect 135897 208449 135913 208567
rect 136031 208449 136073 208567
rect 136191 208449 136207 208567
rect 135897 190727 136207 208449
rect 135897 190609 135913 190727
rect 136031 190609 136073 190727
rect 136191 190609 136207 190727
rect 135897 190567 136207 190609
rect 135897 190449 135913 190567
rect 136031 190449 136073 190567
rect 136191 190449 136207 190567
rect 135897 172727 136207 190449
rect 135897 172609 135913 172727
rect 136031 172609 136073 172727
rect 136191 172609 136207 172727
rect 135897 172567 136207 172609
rect 135897 172449 135913 172567
rect 136031 172449 136073 172567
rect 136191 172449 136207 172567
rect 135897 154727 136207 172449
rect 135897 154609 135913 154727
rect 136031 154609 136073 154727
rect 136191 154609 136207 154727
rect 135897 154567 136207 154609
rect 135897 154449 135913 154567
rect 136031 154449 136073 154567
rect 136191 154449 136207 154567
rect 135897 136727 136207 154449
rect 135897 136609 135913 136727
rect 136031 136609 136073 136727
rect 136191 136609 136207 136727
rect 135897 136567 136207 136609
rect 135897 136449 135913 136567
rect 136031 136449 136073 136567
rect 136191 136449 136207 136567
rect 135897 118727 136207 136449
rect 135897 118609 135913 118727
rect 136031 118609 136073 118727
rect 136191 118609 136207 118727
rect 135897 118567 136207 118609
rect 135897 118449 135913 118567
rect 136031 118449 136073 118567
rect 136191 118449 136207 118567
rect 135897 100727 136207 118449
rect 135897 100609 135913 100727
rect 136031 100609 136073 100727
rect 136191 100609 136207 100727
rect 135897 100567 136207 100609
rect 135897 100449 135913 100567
rect 136031 100449 136073 100567
rect 136191 100449 136207 100567
rect 135897 82727 136207 100449
rect 135897 82609 135913 82727
rect 136031 82609 136073 82727
rect 136191 82609 136207 82727
rect 135897 82567 136207 82609
rect 135897 82449 135913 82567
rect 136031 82449 136073 82567
rect 136191 82449 136207 82567
rect 135897 64727 136207 82449
rect 135897 64609 135913 64727
rect 136031 64609 136073 64727
rect 136191 64609 136207 64727
rect 135897 64567 136207 64609
rect 135897 64449 135913 64567
rect 136031 64449 136073 64567
rect 136191 64449 136207 64567
rect 135897 46727 136207 64449
rect 135897 46609 135913 46727
rect 136031 46609 136073 46727
rect 136191 46609 136207 46727
rect 135897 46567 136207 46609
rect 135897 46449 135913 46567
rect 136031 46449 136073 46567
rect 136191 46449 136207 46567
rect 135897 28727 136207 46449
rect 135897 28609 135913 28727
rect 136031 28609 136073 28727
rect 136191 28609 136207 28727
rect 135897 28567 136207 28609
rect 135897 28449 135913 28567
rect 136031 28449 136073 28567
rect 136191 28449 136207 28567
rect 135897 10727 136207 28449
rect 135897 10609 135913 10727
rect 136031 10609 136073 10727
rect 136191 10609 136207 10727
rect 135897 10567 136207 10609
rect 135897 10449 135913 10567
rect 136031 10449 136073 10567
rect 136191 10449 136207 10567
rect 135897 -653 136207 10449
rect 135897 -771 135913 -653
rect 136031 -771 136073 -653
rect 136191 -771 136207 -653
rect 135897 -813 136207 -771
rect 135897 -931 135913 -813
rect 136031 -931 136073 -813
rect 136191 -931 136207 -813
rect 135897 -947 136207 -931
rect 137757 336587 138067 353581
rect 137757 336469 137773 336587
rect 137891 336469 137933 336587
rect 138051 336469 138067 336587
rect 137757 336427 138067 336469
rect 137757 336309 137773 336427
rect 137891 336309 137933 336427
rect 138051 336309 138067 336427
rect 137757 318587 138067 336309
rect 137757 318469 137773 318587
rect 137891 318469 137933 318587
rect 138051 318469 138067 318587
rect 137757 318427 138067 318469
rect 137757 318309 137773 318427
rect 137891 318309 137933 318427
rect 138051 318309 138067 318427
rect 137757 300587 138067 318309
rect 137757 300469 137773 300587
rect 137891 300469 137933 300587
rect 138051 300469 138067 300587
rect 137757 300427 138067 300469
rect 137757 300309 137773 300427
rect 137891 300309 137933 300427
rect 138051 300309 138067 300427
rect 137757 282587 138067 300309
rect 137757 282469 137773 282587
rect 137891 282469 137933 282587
rect 138051 282469 138067 282587
rect 137757 282427 138067 282469
rect 137757 282309 137773 282427
rect 137891 282309 137933 282427
rect 138051 282309 138067 282427
rect 137757 264587 138067 282309
rect 137757 264469 137773 264587
rect 137891 264469 137933 264587
rect 138051 264469 138067 264587
rect 137757 264427 138067 264469
rect 137757 264309 137773 264427
rect 137891 264309 137933 264427
rect 138051 264309 138067 264427
rect 137757 246587 138067 264309
rect 137757 246469 137773 246587
rect 137891 246469 137933 246587
rect 138051 246469 138067 246587
rect 137757 246427 138067 246469
rect 137757 246309 137773 246427
rect 137891 246309 137933 246427
rect 138051 246309 138067 246427
rect 137757 228587 138067 246309
rect 137757 228469 137773 228587
rect 137891 228469 137933 228587
rect 138051 228469 138067 228587
rect 137757 228427 138067 228469
rect 137757 228309 137773 228427
rect 137891 228309 137933 228427
rect 138051 228309 138067 228427
rect 137757 210587 138067 228309
rect 137757 210469 137773 210587
rect 137891 210469 137933 210587
rect 138051 210469 138067 210587
rect 137757 210427 138067 210469
rect 137757 210309 137773 210427
rect 137891 210309 137933 210427
rect 138051 210309 138067 210427
rect 137757 192587 138067 210309
rect 137757 192469 137773 192587
rect 137891 192469 137933 192587
rect 138051 192469 138067 192587
rect 137757 192427 138067 192469
rect 137757 192309 137773 192427
rect 137891 192309 137933 192427
rect 138051 192309 138067 192427
rect 137757 174587 138067 192309
rect 137757 174469 137773 174587
rect 137891 174469 137933 174587
rect 138051 174469 138067 174587
rect 137757 174427 138067 174469
rect 137757 174309 137773 174427
rect 137891 174309 137933 174427
rect 138051 174309 138067 174427
rect 137757 156587 138067 174309
rect 137757 156469 137773 156587
rect 137891 156469 137933 156587
rect 138051 156469 138067 156587
rect 137757 156427 138067 156469
rect 137757 156309 137773 156427
rect 137891 156309 137933 156427
rect 138051 156309 138067 156427
rect 137757 138587 138067 156309
rect 137757 138469 137773 138587
rect 137891 138469 137933 138587
rect 138051 138469 138067 138587
rect 137757 138427 138067 138469
rect 137757 138309 137773 138427
rect 137891 138309 137933 138427
rect 138051 138309 138067 138427
rect 137757 120587 138067 138309
rect 137757 120469 137773 120587
rect 137891 120469 137933 120587
rect 138051 120469 138067 120587
rect 137757 120427 138067 120469
rect 137757 120309 137773 120427
rect 137891 120309 137933 120427
rect 138051 120309 138067 120427
rect 137757 102587 138067 120309
rect 137757 102469 137773 102587
rect 137891 102469 137933 102587
rect 138051 102469 138067 102587
rect 137757 102427 138067 102469
rect 137757 102309 137773 102427
rect 137891 102309 137933 102427
rect 138051 102309 138067 102427
rect 137757 84587 138067 102309
rect 137757 84469 137773 84587
rect 137891 84469 137933 84587
rect 138051 84469 138067 84587
rect 137757 84427 138067 84469
rect 137757 84309 137773 84427
rect 137891 84309 137933 84427
rect 138051 84309 138067 84427
rect 137757 66587 138067 84309
rect 137757 66469 137773 66587
rect 137891 66469 137933 66587
rect 138051 66469 138067 66587
rect 137757 66427 138067 66469
rect 137757 66309 137773 66427
rect 137891 66309 137933 66427
rect 138051 66309 138067 66427
rect 137757 48587 138067 66309
rect 137757 48469 137773 48587
rect 137891 48469 137933 48587
rect 138051 48469 138067 48587
rect 137757 48427 138067 48469
rect 137757 48309 137773 48427
rect 137891 48309 137933 48427
rect 138051 48309 138067 48427
rect 137757 30587 138067 48309
rect 137757 30469 137773 30587
rect 137891 30469 137933 30587
rect 138051 30469 138067 30587
rect 137757 30427 138067 30469
rect 137757 30309 137773 30427
rect 137891 30309 137933 30427
rect 138051 30309 138067 30427
rect 137757 12587 138067 30309
rect 137757 12469 137773 12587
rect 137891 12469 137933 12587
rect 138051 12469 138067 12587
rect 137757 12427 138067 12469
rect 137757 12309 137773 12427
rect 137891 12309 137933 12427
rect 138051 12309 138067 12427
rect 137757 -1613 138067 12309
rect 137757 -1731 137773 -1613
rect 137891 -1731 137933 -1613
rect 138051 -1731 138067 -1613
rect 137757 -1773 138067 -1731
rect 137757 -1891 137773 -1773
rect 137891 -1891 137933 -1773
rect 138051 -1891 138067 -1773
rect 137757 -1907 138067 -1891
rect 139617 338447 139927 354541
rect 139617 338329 139633 338447
rect 139751 338329 139793 338447
rect 139911 338329 139927 338447
rect 139617 338287 139927 338329
rect 139617 338169 139633 338287
rect 139751 338169 139793 338287
rect 139911 338169 139927 338287
rect 139617 320447 139927 338169
rect 139617 320329 139633 320447
rect 139751 320329 139793 320447
rect 139911 320329 139927 320447
rect 139617 320287 139927 320329
rect 139617 320169 139633 320287
rect 139751 320169 139793 320287
rect 139911 320169 139927 320287
rect 139617 302447 139927 320169
rect 139617 302329 139633 302447
rect 139751 302329 139793 302447
rect 139911 302329 139927 302447
rect 139617 302287 139927 302329
rect 139617 302169 139633 302287
rect 139751 302169 139793 302287
rect 139911 302169 139927 302287
rect 139617 284447 139927 302169
rect 139617 284329 139633 284447
rect 139751 284329 139793 284447
rect 139911 284329 139927 284447
rect 139617 284287 139927 284329
rect 139617 284169 139633 284287
rect 139751 284169 139793 284287
rect 139911 284169 139927 284287
rect 139617 266447 139927 284169
rect 139617 266329 139633 266447
rect 139751 266329 139793 266447
rect 139911 266329 139927 266447
rect 139617 266287 139927 266329
rect 139617 266169 139633 266287
rect 139751 266169 139793 266287
rect 139911 266169 139927 266287
rect 139617 248447 139927 266169
rect 139617 248329 139633 248447
rect 139751 248329 139793 248447
rect 139911 248329 139927 248447
rect 139617 248287 139927 248329
rect 139617 248169 139633 248287
rect 139751 248169 139793 248287
rect 139911 248169 139927 248287
rect 139617 230447 139927 248169
rect 139617 230329 139633 230447
rect 139751 230329 139793 230447
rect 139911 230329 139927 230447
rect 139617 230287 139927 230329
rect 139617 230169 139633 230287
rect 139751 230169 139793 230287
rect 139911 230169 139927 230287
rect 139617 212447 139927 230169
rect 139617 212329 139633 212447
rect 139751 212329 139793 212447
rect 139911 212329 139927 212447
rect 139617 212287 139927 212329
rect 139617 212169 139633 212287
rect 139751 212169 139793 212287
rect 139911 212169 139927 212287
rect 139617 194447 139927 212169
rect 139617 194329 139633 194447
rect 139751 194329 139793 194447
rect 139911 194329 139927 194447
rect 139617 194287 139927 194329
rect 139617 194169 139633 194287
rect 139751 194169 139793 194287
rect 139911 194169 139927 194287
rect 139617 176447 139927 194169
rect 139617 176329 139633 176447
rect 139751 176329 139793 176447
rect 139911 176329 139927 176447
rect 139617 176287 139927 176329
rect 139617 176169 139633 176287
rect 139751 176169 139793 176287
rect 139911 176169 139927 176287
rect 139617 158447 139927 176169
rect 139617 158329 139633 158447
rect 139751 158329 139793 158447
rect 139911 158329 139927 158447
rect 139617 158287 139927 158329
rect 139617 158169 139633 158287
rect 139751 158169 139793 158287
rect 139911 158169 139927 158287
rect 139617 140447 139927 158169
rect 139617 140329 139633 140447
rect 139751 140329 139793 140447
rect 139911 140329 139927 140447
rect 139617 140287 139927 140329
rect 139617 140169 139633 140287
rect 139751 140169 139793 140287
rect 139911 140169 139927 140287
rect 139617 122447 139927 140169
rect 139617 122329 139633 122447
rect 139751 122329 139793 122447
rect 139911 122329 139927 122447
rect 139617 122287 139927 122329
rect 139617 122169 139633 122287
rect 139751 122169 139793 122287
rect 139911 122169 139927 122287
rect 139617 104447 139927 122169
rect 139617 104329 139633 104447
rect 139751 104329 139793 104447
rect 139911 104329 139927 104447
rect 139617 104287 139927 104329
rect 139617 104169 139633 104287
rect 139751 104169 139793 104287
rect 139911 104169 139927 104287
rect 139617 86447 139927 104169
rect 139617 86329 139633 86447
rect 139751 86329 139793 86447
rect 139911 86329 139927 86447
rect 139617 86287 139927 86329
rect 139617 86169 139633 86287
rect 139751 86169 139793 86287
rect 139911 86169 139927 86287
rect 139617 68447 139927 86169
rect 139617 68329 139633 68447
rect 139751 68329 139793 68447
rect 139911 68329 139927 68447
rect 139617 68287 139927 68329
rect 139617 68169 139633 68287
rect 139751 68169 139793 68287
rect 139911 68169 139927 68287
rect 139617 50447 139927 68169
rect 139617 50329 139633 50447
rect 139751 50329 139793 50447
rect 139911 50329 139927 50447
rect 139617 50287 139927 50329
rect 139617 50169 139633 50287
rect 139751 50169 139793 50287
rect 139911 50169 139927 50287
rect 139617 32447 139927 50169
rect 139617 32329 139633 32447
rect 139751 32329 139793 32447
rect 139911 32329 139927 32447
rect 139617 32287 139927 32329
rect 139617 32169 139633 32287
rect 139751 32169 139793 32287
rect 139911 32169 139927 32287
rect 139617 14447 139927 32169
rect 139617 14329 139633 14447
rect 139751 14329 139793 14447
rect 139911 14329 139927 14447
rect 139617 14287 139927 14329
rect 139617 14169 139633 14287
rect 139751 14169 139793 14287
rect 139911 14169 139927 14287
rect 139617 -2573 139927 14169
rect 139617 -2691 139633 -2573
rect 139751 -2691 139793 -2573
rect 139911 -2691 139927 -2573
rect 139617 -2733 139927 -2691
rect 139617 -2851 139633 -2733
rect 139751 -2851 139793 -2733
rect 139911 -2851 139927 -2733
rect 139617 -2867 139927 -2851
rect 141477 340307 141787 355501
rect 150477 355299 150787 355795
rect 150477 355181 150493 355299
rect 150611 355181 150653 355299
rect 150771 355181 150787 355299
rect 150477 355139 150787 355181
rect 150477 355021 150493 355139
rect 150611 355021 150653 355139
rect 150771 355021 150787 355139
rect 148617 354339 148927 354835
rect 148617 354221 148633 354339
rect 148751 354221 148793 354339
rect 148911 354221 148927 354339
rect 148617 354179 148927 354221
rect 148617 354061 148633 354179
rect 148751 354061 148793 354179
rect 148911 354061 148927 354179
rect 146757 353379 147067 353875
rect 146757 353261 146773 353379
rect 146891 353261 146933 353379
rect 147051 353261 147067 353379
rect 146757 353219 147067 353261
rect 146757 353101 146773 353219
rect 146891 353101 146933 353219
rect 147051 353101 147067 353219
rect 141477 340189 141493 340307
rect 141611 340189 141653 340307
rect 141771 340189 141787 340307
rect 141477 340147 141787 340189
rect 141477 340029 141493 340147
rect 141611 340029 141653 340147
rect 141771 340029 141787 340147
rect 141477 322307 141787 340029
rect 141477 322189 141493 322307
rect 141611 322189 141653 322307
rect 141771 322189 141787 322307
rect 141477 322147 141787 322189
rect 141477 322029 141493 322147
rect 141611 322029 141653 322147
rect 141771 322029 141787 322147
rect 141477 304307 141787 322029
rect 141477 304189 141493 304307
rect 141611 304189 141653 304307
rect 141771 304189 141787 304307
rect 141477 304147 141787 304189
rect 141477 304029 141493 304147
rect 141611 304029 141653 304147
rect 141771 304029 141787 304147
rect 141477 286307 141787 304029
rect 141477 286189 141493 286307
rect 141611 286189 141653 286307
rect 141771 286189 141787 286307
rect 141477 286147 141787 286189
rect 141477 286029 141493 286147
rect 141611 286029 141653 286147
rect 141771 286029 141787 286147
rect 141477 268307 141787 286029
rect 141477 268189 141493 268307
rect 141611 268189 141653 268307
rect 141771 268189 141787 268307
rect 141477 268147 141787 268189
rect 141477 268029 141493 268147
rect 141611 268029 141653 268147
rect 141771 268029 141787 268147
rect 141477 250307 141787 268029
rect 141477 250189 141493 250307
rect 141611 250189 141653 250307
rect 141771 250189 141787 250307
rect 141477 250147 141787 250189
rect 141477 250029 141493 250147
rect 141611 250029 141653 250147
rect 141771 250029 141787 250147
rect 141477 232307 141787 250029
rect 141477 232189 141493 232307
rect 141611 232189 141653 232307
rect 141771 232189 141787 232307
rect 141477 232147 141787 232189
rect 141477 232029 141493 232147
rect 141611 232029 141653 232147
rect 141771 232029 141787 232147
rect 141477 214307 141787 232029
rect 141477 214189 141493 214307
rect 141611 214189 141653 214307
rect 141771 214189 141787 214307
rect 141477 214147 141787 214189
rect 141477 214029 141493 214147
rect 141611 214029 141653 214147
rect 141771 214029 141787 214147
rect 141477 196307 141787 214029
rect 141477 196189 141493 196307
rect 141611 196189 141653 196307
rect 141771 196189 141787 196307
rect 141477 196147 141787 196189
rect 141477 196029 141493 196147
rect 141611 196029 141653 196147
rect 141771 196029 141787 196147
rect 141477 178307 141787 196029
rect 141477 178189 141493 178307
rect 141611 178189 141653 178307
rect 141771 178189 141787 178307
rect 141477 178147 141787 178189
rect 141477 178029 141493 178147
rect 141611 178029 141653 178147
rect 141771 178029 141787 178147
rect 141477 160307 141787 178029
rect 141477 160189 141493 160307
rect 141611 160189 141653 160307
rect 141771 160189 141787 160307
rect 141477 160147 141787 160189
rect 141477 160029 141493 160147
rect 141611 160029 141653 160147
rect 141771 160029 141787 160147
rect 141477 142307 141787 160029
rect 141477 142189 141493 142307
rect 141611 142189 141653 142307
rect 141771 142189 141787 142307
rect 141477 142147 141787 142189
rect 141477 142029 141493 142147
rect 141611 142029 141653 142147
rect 141771 142029 141787 142147
rect 141477 124307 141787 142029
rect 141477 124189 141493 124307
rect 141611 124189 141653 124307
rect 141771 124189 141787 124307
rect 141477 124147 141787 124189
rect 141477 124029 141493 124147
rect 141611 124029 141653 124147
rect 141771 124029 141787 124147
rect 141477 106307 141787 124029
rect 141477 106189 141493 106307
rect 141611 106189 141653 106307
rect 141771 106189 141787 106307
rect 141477 106147 141787 106189
rect 141477 106029 141493 106147
rect 141611 106029 141653 106147
rect 141771 106029 141787 106147
rect 141477 88307 141787 106029
rect 141477 88189 141493 88307
rect 141611 88189 141653 88307
rect 141771 88189 141787 88307
rect 141477 88147 141787 88189
rect 141477 88029 141493 88147
rect 141611 88029 141653 88147
rect 141771 88029 141787 88147
rect 141477 70307 141787 88029
rect 141477 70189 141493 70307
rect 141611 70189 141653 70307
rect 141771 70189 141787 70307
rect 141477 70147 141787 70189
rect 141477 70029 141493 70147
rect 141611 70029 141653 70147
rect 141771 70029 141787 70147
rect 141477 52307 141787 70029
rect 141477 52189 141493 52307
rect 141611 52189 141653 52307
rect 141771 52189 141787 52307
rect 141477 52147 141787 52189
rect 141477 52029 141493 52147
rect 141611 52029 141653 52147
rect 141771 52029 141787 52147
rect 141477 34307 141787 52029
rect 141477 34189 141493 34307
rect 141611 34189 141653 34307
rect 141771 34189 141787 34307
rect 141477 34147 141787 34189
rect 141477 34029 141493 34147
rect 141611 34029 141653 34147
rect 141771 34029 141787 34147
rect 141477 16307 141787 34029
rect 141477 16189 141493 16307
rect 141611 16189 141653 16307
rect 141771 16189 141787 16307
rect 141477 16147 141787 16189
rect 141477 16029 141493 16147
rect 141611 16029 141653 16147
rect 141771 16029 141787 16147
rect 132477 -3171 132493 -3053
rect 132611 -3171 132653 -3053
rect 132771 -3171 132787 -3053
rect 132477 -3213 132787 -3171
rect 132477 -3331 132493 -3213
rect 132611 -3331 132653 -3213
rect 132771 -3331 132787 -3213
rect 132477 -3827 132787 -3331
rect 141477 -3533 141787 16029
rect 144897 352419 145207 352915
rect 144897 352301 144913 352419
rect 145031 352301 145073 352419
rect 145191 352301 145207 352419
rect 144897 352259 145207 352301
rect 144897 352141 144913 352259
rect 145031 352141 145073 352259
rect 145191 352141 145207 352259
rect 144897 343727 145207 352141
rect 144897 343609 144913 343727
rect 145031 343609 145073 343727
rect 145191 343609 145207 343727
rect 144897 343567 145207 343609
rect 144897 343449 144913 343567
rect 145031 343449 145073 343567
rect 145191 343449 145207 343567
rect 144897 325727 145207 343449
rect 144897 325609 144913 325727
rect 145031 325609 145073 325727
rect 145191 325609 145207 325727
rect 144897 325567 145207 325609
rect 144897 325449 144913 325567
rect 145031 325449 145073 325567
rect 145191 325449 145207 325567
rect 144897 307727 145207 325449
rect 144897 307609 144913 307727
rect 145031 307609 145073 307727
rect 145191 307609 145207 307727
rect 144897 307567 145207 307609
rect 144897 307449 144913 307567
rect 145031 307449 145073 307567
rect 145191 307449 145207 307567
rect 144897 289727 145207 307449
rect 144897 289609 144913 289727
rect 145031 289609 145073 289727
rect 145191 289609 145207 289727
rect 144897 289567 145207 289609
rect 144897 289449 144913 289567
rect 145031 289449 145073 289567
rect 145191 289449 145207 289567
rect 144897 271727 145207 289449
rect 144897 271609 144913 271727
rect 145031 271609 145073 271727
rect 145191 271609 145207 271727
rect 144897 271567 145207 271609
rect 144897 271449 144913 271567
rect 145031 271449 145073 271567
rect 145191 271449 145207 271567
rect 144897 253727 145207 271449
rect 144897 253609 144913 253727
rect 145031 253609 145073 253727
rect 145191 253609 145207 253727
rect 144897 253567 145207 253609
rect 144897 253449 144913 253567
rect 145031 253449 145073 253567
rect 145191 253449 145207 253567
rect 144897 235727 145207 253449
rect 144897 235609 144913 235727
rect 145031 235609 145073 235727
rect 145191 235609 145207 235727
rect 144897 235567 145207 235609
rect 144897 235449 144913 235567
rect 145031 235449 145073 235567
rect 145191 235449 145207 235567
rect 144897 217727 145207 235449
rect 144897 217609 144913 217727
rect 145031 217609 145073 217727
rect 145191 217609 145207 217727
rect 144897 217567 145207 217609
rect 144897 217449 144913 217567
rect 145031 217449 145073 217567
rect 145191 217449 145207 217567
rect 144897 199727 145207 217449
rect 144897 199609 144913 199727
rect 145031 199609 145073 199727
rect 145191 199609 145207 199727
rect 144897 199567 145207 199609
rect 144897 199449 144913 199567
rect 145031 199449 145073 199567
rect 145191 199449 145207 199567
rect 144897 181727 145207 199449
rect 144897 181609 144913 181727
rect 145031 181609 145073 181727
rect 145191 181609 145207 181727
rect 144897 181567 145207 181609
rect 144897 181449 144913 181567
rect 145031 181449 145073 181567
rect 145191 181449 145207 181567
rect 144897 163727 145207 181449
rect 144897 163609 144913 163727
rect 145031 163609 145073 163727
rect 145191 163609 145207 163727
rect 144897 163567 145207 163609
rect 144897 163449 144913 163567
rect 145031 163449 145073 163567
rect 145191 163449 145207 163567
rect 144897 145727 145207 163449
rect 144897 145609 144913 145727
rect 145031 145609 145073 145727
rect 145191 145609 145207 145727
rect 144897 145567 145207 145609
rect 144897 145449 144913 145567
rect 145031 145449 145073 145567
rect 145191 145449 145207 145567
rect 144897 127727 145207 145449
rect 144897 127609 144913 127727
rect 145031 127609 145073 127727
rect 145191 127609 145207 127727
rect 144897 127567 145207 127609
rect 144897 127449 144913 127567
rect 145031 127449 145073 127567
rect 145191 127449 145207 127567
rect 144897 109727 145207 127449
rect 144897 109609 144913 109727
rect 145031 109609 145073 109727
rect 145191 109609 145207 109727
rect 144897 109567 145207 109609
rect 144897 109449 144913 109567
rect 145031 109449 145073 109567
rect 145191 109449 145207 109567
rect 144897 91727 145207 109449
rect 144897 91609 144913 91727
rect 145031 91609 145073 91727
rect 145191 91609 145207 91727
rect 144897 91567 145207 91609
rect 144897 91449 144913 91567
rect 145031 91449 145073 91567
rect 145191 91449 145207 91567
rect 144897 73727 145207 91449
rect 144897 73609 144913 73727
rect 145031 73609 145073 73727
rect 145191 73609 145207 73727
rect 144897 73567 145207 73609
rect 144897 73449 144913 73567
rect 145031 73449 145073 73567
rect 145191 73449 145207 73567
rect 144897 55727 145207 73449
rect 144897 55609 144913 55727
rect 145031 55609 145073 55727
rect 145191 55609 145207 55727
rect 144897 55567 145207 55609
rect 144897 55449 144913 55567
rect 145031 55449 145073 55567
rect 145191 55449 145207 55567
rect 144897 37727 145207 55449
rect 144897 37609 144913 37727
rect 145031 37609 145073 37727
rect 145191 37609 145207 37727
rect 144897 37567 145207 37609
rect 144897 37449 144913 37567
rect 145031 37449 145073 37567
rect 145191 37449 145207 37567
rect 144897 19727 145207 37449
rect 144897 19609 144913 19727
rect 145031 19609 145073 19727
rect 145191 19609 145207 19727
rect 144897 19567 145207 19609
rect 144897 19449 144913 19567
rect 145031 19449 145073 19567
rect 145191 19449 145207 19567
rect 144897 1727 145207 19449
rect 144897 1609 144913 1727
rect 145031 1609 145073 1727
rect 145191 1609 145207 1727
rect 144897 1567 145207 1609
rect 144897 1449 144913 1567
rect 145031 1449 145073 1567
rect 145191 1449 145207 1567
rect 144897 -173 145207 1449
rect 144897 -291 144913 -173
rect 145031 -291 145073 -173
rect 145191 -291 145207 -173
rect 144897 -333 145207 -291
rect 144897 -451 144913 -333
rect 145031 -451 145073 -333
rect 145191 -451 145207 -333
rect 144897 -947 145207 -451
rect 146757 345587 147067 353101
rect 146757 345469 146773 345587
rect 146891 345469 146933 345587
rect 147051 345469 147067 345587
rect 146757 345427 147067 345469
rect 146757 345309 146773 345427
rect 146891 345309 146933 345427
rect 147051 345309 147067 345427
rect 146757 327587 147067 345309
rect 146757 327469 146773 327587
rect 146891 327469 146933 327587
rect 147051 327469 147067 327587
rect 146757 327427 147067 327469
rect 146757 327309 146773 327427
rect 146891 327309 146933 327427
rect 147051 327309 147067 327427
rect 146757 309587 147067 327309
rect 146757 309469 146773 309587
rect 146891 309469 146933 309587
rect 147051 309469 147067 309587
rect 146757 309427 147067 309469
rect 146757 309309 146773 309427
rect 146891 309309 146933 309427
rect 147051 309309 147067 309427
rect 146757 291587 147067 309309
rect 146757 291469 146773 291587
rect 146891 291469 146933 291587
rect 147051 291469 147067 291587
rect 146757 291427 147067 291469
rect 146757 291309 146773 291427
rect 146891 291309 146933 291427
rect 147051 291309 147067 291427
rect 146757 273587 147067 291309
rect 146757 273469 146773 273587
rect 146891 273469 146933 273587
rect 147051 273469 147067 273587
rect 146757 273427 147067 273469
rect 146757 273309 146773 273427
rect 146891 273309 146933 273427
rect 147051 273309 147067 273427
rect 146757 255587 147067 273309
rect 146757 255469 146773 255587
rect 146891 255469 146933 255587
rect 147051 255469 147067 255587
rect 146757 255427 147067 255469
rect 146757 255309 146773 255427
rect 146891 255309 146933 255427
rect 147051 255309 147067 255427
rect 146757 237587 147067 255309
rect 146757 237469 146773 237587
rect 146891 237469 146933 237587
rect 147051 237469 147067 237587
rect 146757 237427 147067 237469
rect 146757 237309 146773 237427
rect 146891 237309 146933 237427
rect 147051 237309 147067 237427
rect 146757 219587 147067 237309
rect 146757 219469 146773 219587
rect 146891 219469 146933 219587
rect 147051 219469 147067 219587
rect 146757 219427 147067 219469
rect 146757 219309 146773 219427
rect 146891 219309 146933 219427
rect 147051 219309 147067 219427
rect 146757 201587 147067 219309
rect 146757 201469 146773 201587
rect 146891 201469 146933 201587
rect 147051 201469 147067 201587
rect 146757 201427 147067 201469
rect 146757 201309 146773 201427
rect 146891 201309 146933 201427
rect 147051 201309 147067 201427
rect 146757 183587 147067 201309
rect 146757 183469 146773 183587
rect 146891 183469 146933 183587
rect 147051 183469 147067 183587
rect 146757 183427 147067 183469
rect 146757 183309 146773 183427
rect 146891 183309 146933 183427
rect 147051 183309 147067 183427
rect 146757 165587 147067 183309
rect 146757 165469 146773 165587
rect 146891 165469 146933 165587
rect 147051 165469 147067 165587
rect 146757 165427 147067 165469
rect 146757 165309 146773 165427
rect 146891 165309 146933 165427
rect 147051 165309 147067 165427
rect 146757 147587 147067 165309
rect 146757 147469 146773 147587
rect 146891 147469 146933 147587
rect 147051 147469 147067 147587
rect 146757 147427 147067 147469
rect 146757 147309 146773 147427
rect 146891 147309 146933 147427
rect 147051 147309 147067 147427
rect 146757 129587 147067 147309
rect 146757 129469 146773 129587
rect 146891 129469 146933 129587
rect 147051 129469 147067 129587
rect 146757 129427 147067 129469
rect 146757 129309 146773 129427
rect 146891 129309 146933 129427
rect 147051 129309 147067 129427
rect 146757 111587 147067 129309
rect 146757 111469 146773 111587
rect 146891 111469 146933 111587
rect 147051 111469 147067 111587
rect 146757 111427 147067 111469
rect 146757 111309 146773 111427
rect 146891 111309 146933 111427
rect 147051 111309 147067 111427
rect 146757 93587 147067 111309
rect 146757 93469 146773 93587
rect 146891 93469 146933 93587
rect 147051 93469 147067 93587
rect 146757 93427 147067 93469
rect 146757 93309 146773 93427
rect 146891 93309 146933 93427
rect 147051 93309 147067 93427
rect 146757 75587 147067 93309
rect 146757 75469 146773 75587
rect 146891 75469 146933 75587
rect 147051 75469 147067 75587
rect 146757 75427 147067 75469
rect 146757 75309 146773 75427
rect 146891 75309 146933 75427
rect 147051 75309 147067 75427
rect 146757 57587 147067 75309
rect 146757 57469 146773 57587
rect 146891 57469 146933 57587
rect 147051 57469 147067 57587
rect 146757 57427 147067 57469
rect 146757 57309 146773 57427
rect 146891 57309 146933 57427
rect 147051 57309 147067 57427
rect 146757 39587 147067 57309
rect 146757 39469 146773 39587
rect 146891 39469 146933 39587
rect 147051 39469 147067 39587
rect 146757 39427 147067 39469
rect 146757 39309 146773 39427
rect 146891 39309 146933 39427
rect 147051 39309 147067 39427
rect 146757 21587 147067 39309
rect 146757 21469 146773 21587
rect 146891 21469 146933 21587
rect 147051 21469 147067 21587
rect 146757 21427 147067 21469
rect 146757 21309 146773 21427
rect 146891 21309 146933 21427
rect 147051 21309 147067 21427
rect 146757 3587 147067 21309
rect 146757 3469 146773 3587
rect 146891 3469 146933 3587
rect 147051 3469 147067 3587
rect 146757 3427 147067 3469
rect 146757 3309 146773 3427
rect 146891 3309 146933 3427
rect 147051 3309 147067 3427
rect 146757 -1133 147067 3309
rect 146757 -1251 146773 -1133
rect 146891 -1251 146933 -1133
rect 147051 -1251 147067 -1133
rect 146757 -1293 147067 -1251
rect 146757 -1411 146773 -1293
rect 146891 -1411 146933 -1293
rect 147051 -1411 147067 -1293
rect 146757 -1907 147067 -1411
rect 148617 347447 148927 354061
rect 148617 347329 148633 347447
rect 148751 347329 148793 347447
rect 148911 347329 148927 347447
rect 148617 347287 148927 347329
rect 148617 347169 148633 347287
rect 148751 347169 148793 347287
rect 148911 347169 148927 347287
rect 148617 329447 148927 347169
rect 148617 329329 148633 329447
rect 148751 329329 148793 329447
rect 148911 329329 148927 329447
rect 148617 329287 148927 329329
rect 148617 329169 148633 329287
rect 148751 329169 148793 329287
rect 148911 329169 148927 329287
rect 148617 311447 148927 329169
rect 148617 311329 148633 311447
rect 148751 311329 148793 311447
rect 148911 311329 148927 311447
rect 148617 311287 148927 311329
rect 148617 311169 148633 311287
rect 148751 311169 148793 311287
rect 148911 311169 148927 311287
rect 148617 293447 148927 311169
rect 148617 293329 148633 293447
rect 148751 293329 148793 293447
rect 148911 293329 148927 293447
rect 148617 293287 148927 293329
rect 148617 293169 148633 293287
rect 148751 293169 148793 293287
rect 148911 293169 148927 293287
rect 148617 275447 148927 293169
rect 148617 275329 148633 275447
rect 148751 275329 148793 275447
rect 148911 275329 148927 275447
rect 148617 275287 148927 275329
rect 148617 275169 148633 275287
rect 148751 275169 148793 275287
rect 148911 275169 148927 275287
rect 148617 257447 148927 275169
rect 148617 257329 148633 257447
rect 148751 257329 148793 257447
rect 148911 257329 148927 257447
rect 148617 257287 148927 257329
rect 148617 257169 148633 257287
rect 148751 257169 148793 257287
rect 148911 257169 148927 257287
rect 148617 239447 148927 257169
rect 148617 239329 148633 239447
rect 148751 239329 148793 239447
rect 148911 239329 148927 239447
rect 148617 239287 148927 239329
rect 148617 239169 148633 239287
rect 148751 239169 148793 239287
rect 148911 239169 148927 239287
rect 148617 221447 148927 239169
rect 148617 221329 148633 221447
rect 148751 221329 148793 221447
rect 148911 221329 148927 221447
rect 148617 221287 148927 221329
rect 148617 221169 148633 221287
rect 148751 221169 148793 221287
rect 148911 221169 148927 221287
rect 148617 203447 148927 221169
rect 148617 203329 148633 203447
rect 148751 203329 148793 203447
rect 148911 203329 148927 203447
rect 148617 203287 148927 203329
rect 148617 203169 148633 203287
rect 148751 203169 148793 203287
rect 148911 203169 148927 203287
rect 148617 185447 148927 203169
rect 148617 185329 148633 185447
rect 148751 185329 148793 185447
rect 148911 185329 148927 185447
rect 148617 185287 148927 185329
rect 148617 185169 148633 185287
rect 148751 185169 148793 185287
rect 148911 185169 148927 185287
rect 148617 167447 148927 185169
rect 148617 167329 148633 167447
rect 148751 167329 148793 167447
rect 148911 167329 148927 167447
rect 148617 167287 148927 167329
rect 148617 167169 148633 167287
rect 148751 167169 148793 167287
rect 148911 167169 148927 167287
rect 148617 149447 148927 167169
rect 148617 149329 148633 149447
rect 148751 149329 148793 149447
rect 148911 149329 148927 149447
rect 148617 149287 148927 149329
rect 148617 149169 148633 149287
rect 148751 149169 148793 149287
rect 148911 149169 148927 149287
rect 148617 131447 148927 149169
rect 148617 131329 148633 131447
rect 148751 131329 148793 131447
rect 148911 131329 148927 131447
rect 148617 131287 148927 131329
rect 148617 131169 148633 131287
rect 148751 131169 148793 131287
rect 148911 131169 148927 131287
rect 148617 113447 148927 131169
rect 148617 113329 148633 113447
rect 148751 113329 148793 113447
rect 148911 113329 148927 113447
rect 148617 113287 148927 113329
rect 148617 113169 148633 113287
rect 148751 113169 148793 113287
rect 148911 113169 148927 113287
rect 148617 95447 148927 113169
rect 148617 95329 148633 95447
rect 148751 95329 148793 95447
rect 148911 95329 148927 95447
rect 148617 95287 148927 95329
rect 148617 95169 148633 95287
rect 148751 95169 148793 95287
rect 148911 95169 148927 95287
rect 148617 77447 148927 95169
rect 148617 77329 148633 77447
rect 148751 77329 148793 77447
rect 148911 77329 148927 77447
rect 148617 77287 148927 77329
rect 148617 77169 148633 77287
rect 148751 77169 148793 77287
rect 148911 77169 148927 77287
rect 148617 59447 148927 77169
rect 148617 59329 148633 59447
rect 148751 59329 148793 59447
rect 148911 59329 148927 59447
rect 148617 59287 148927 59329
rect 148617 59169 148633 59287
rect 148751 59169 148793 59287
rect 148911 59169 148927 59287
rect 148617 41447 148927 59169
rect 148617 41329 148633 41447
rect 148751 41329 148793 41447
rect 148911 41329 148927 41447
rect 148617 41287 148927 41329
rect 148617 41169 148633 41287
rect 148751 41169 148793 41287
rect 148911 41169 148927 41287
rect 148617 23447 148927 41169
rect 148617 23329 148633 23447
rect 148751 23329 148793 23447
rect 148911 23329 148927 23447
rect 148617 23287 148927 23329
rect 148617 23169 148633 23287
rect 148751 23169 148793 23287
rect 148911 23169 148927 23287
rect 148617 5447 148927 23169
rect 148617 5329 148633 5447
rect 148751 5329 148793 5447
rect 148911 5329 148927 5447
rect 148617 5287 148927 5329
rect 148617 5169 148633 5287
rect 148751 5169 148793 5287
rect 148911 5169 148927 5287
rect 148617 -2093 148927 5169
rect 148617 -2211 148633 -2093
rect 148751 -2211 148793 -2093
rect 148911 -2211 148927 -2093
rect 148617 -2253 148927 -2211
rect 148617 -2371 148633 -2253
rect 148751 -2371 148793 -2253
rect 148911 -2371 148927 -2253
rect 148617 -2867 148927 -2371
rect 150477 349307 150787 355021
rect 159477 355779 159787 355795
rect 159477 355661 159493 355779
rect 159611 355661 159653 355779
rect 159771 355661 159787 355779
rect 159477 355619 159787 355661
rect 159477 355501 159493 355619
rect 159611 355501 159653 355619
rect 159771 355501 159787 355619
rect 157617 354819 157927 354835
rect 157617 354701 157633 354819
rect 157751 354701 157793 354819
rect 157911 354701 157927 354819
rect 157617 354659 157927 354701
rect 157617 354541 157633 354659
rect 157751 354541 157793 354659
rect 157911 354541 157927 354659
rect 155757 353859 156067 353875
rect 155757 353741 155773 353859
rect 155891 353741 155933 353859
rect 156051 353741 156067 353859
rect 155757 353699 156067 353741
rect 155757 353581 155773 353699
rect 155891 353581 155933 353699
rect 156051 353581 156067 353699
rect 150477 349189 150493 349307
rect 150611 349189 150653 349307
rect 150771 349189 150787 349307
rect 150477 349147 150787 349189
rect 150477 349029 150493 349147
rect 150611 349029 150653 349147
rect 150771 349029 150787 349147
rect 150477 331307 150787 349029
rect 150477 331189 150493 331307
rect 150611 331189 150653 331307
rect 150771 331189 150787 331307
rect 150477 331147 150787 331189
rect 150477 331029 150493 331147
rect 150611 331029 150653 331147
rect 150771 331029 150787 331147
rect 150477 313307 150787 331029
rect 150477 313189 150493 313307
rect 150611 313189 150653 313307
rect 150771 313189 150787 313307
rect 150477 313147 150787 313189
rect 150477 313029 150493 313147
rect 150611 313029 150653 313147
rect 150771 313029 150787 313147
rect 150477 295307 150787 313029
rect 150477 295189 150493 295307
rect 150611 295189 150653 295307
rect 150771 295189 150787 295307
rect 150477 295147 150787 295189
rect 150477 295029 150493 295147
rect 150611 295029 150653 295147
rect 150771 295029 150787 295147
rect 150477 277307 150787 295029
rect 150477 277189 150493 277307
rect 150611 277189 150653 277307
rect 150771 277189 150787 277307
rect 150477 277147 150787 277189
rect 150477 277029 150493 277147
rect 150611 277029 150653 277147
rect 150771 277029 150787 277147
rect 150477 259307 150787 277029
rect 150477 259189 150493 259307
rect 150611 259189 150653 259307
rect 150771 259189 150787 259307
rect 150477 259147 150787 259189
rect 150477 259029 150493 259147
rect 150611 259029 150653 259147
rect 150771 259029 150787 259147
rect 150477 241307 150787 259029
rect 150477 241189 150493 241307
rect 150611 241189 150653 241307
rect 150771 241189 150787 241307
rect 150477 241147 150787 241189
rect 150477 241029 150493 241147
rect 150611 241029 150653 241147
rect 150771 241029 150787 241147
rect 150477 223307 150787 241029
rect 150477 223189 150493 223307
rect 150611 223189 150653 223307
rect 150771 223189 150787 223307
rect 150477 223147 150787 223189
rect 150477 223029 150493 223147
rect 150611 223029 150653 223147
rect 150771 223029 150787 223147
rect 150477 205307 150787 223029
rect 150477 205189 150493 205307
rect 150611 205189 150653 205307
rect 150771 205189 150787 205307
rect 150477 205147 150787 205189
rect 150477 205029 150493 205147
rect 150611 205029 150653 205147
rect 150771 205029 150787 205147
rect 150477 187307 150787 205029
rect 150477 187189 150493 187307
rect 150611 187189 150653 187307
rect 150771 187189 150787 187307
rect 150477 187147 150787 187189
rect 150477 187029 150493 187147
rect 150611 187029 150653 187147
rect 150771 187029 150787 187147
rect 150477 169307 150787 187029
rect 150477 169189 150493 169307
rect 150611 169189 150653 169307
rect 150771 169189 150787 169307
rect 150477 169147 150787 169189
rect 150477 169029 150493 169147
rect 150611 169029 150653 169147
rect 150771 169029 150787 169147
rect 150477 151307 150787 169029
rect 150477 151189 150493 151307
rect 150611 151189 150653 151307
rect 150771 151189 150787 151307
rect 150477 151147 150787 151189
rect 150477 151029 150493 151147
rect 150611 151029 150653 151147
rect 150771 151029 150787 151147
rect 150477 133307 150787 151029
rect 150477 133189 150493 133307
rect 150611 133189 150653 133307
rect 150771 133189 150787 133307
rect 150477 133147 150787 133189
rect 150477 133029 150493 133147
rect 150611 133029 150653 133147
rect 150771 133029 150787 133147
rect 150477 115307 150787 133029
rect 150477 115189 150493 115307
rect 150611 115189 150653 115307
rect 150771 115189 150787 115307
rect 150477 115147 150787 115189
rect 150477 115029 150493 115147
rect 150611 115029 150653 115147
rect 150771 115029 150787 115147
rect 150477 97307 150787 115029
rect 150477 97189 150493 97307
rect 150611 97189 150653 97307
rect 150771 97189 150787 97307
rect 150477 97147 150787 97189
rect 150477 97029 150493 97147
rect 150611 97029 150653 97147
rect 150771 97029 150787 97147
rect 150477 79307 150787 97029
rect 150477 79189 150493 79307
rect 150611 79189 150653 79307
rect 150771 79189 150787 79307
rect 150477 79147 150787 79189
rect 150477 79029 150493 79147
rect 150611 79029 150653 79147
rect 150771 79029 150787 79147
rect 150477 61307 150787 79029
rect 150477 61189 150493 61307
rect 150611 61189 150653 61307
rect 150771 61189 150787 61307
rect 150477 61147 150787 61189
rect 150477 61029 150493 61147
rect 150611 61029 150653 61147
rect 150771 61029 150787 61147
rect 150477 43307 150787 61029
rect 150477 43189 150493 43307
rect 150611 43189 150653 43307
rect 150771 43189 150787 43307
rect 150477 43147 150787 43189
rect 150477 43029 150493 43147
rect 150611 43029 150653 43147
rect 150771 43029 150787 43147
rect 150477 25307 150787 43029
rect 150477 25189 150493 25307
rect 150611 25189 150653 25307
rect 150771 25189 150787 25307
rect 150477 25147 150787 25189
rect 150477 25029 150493 25147
rect 150611 25029 150653 25147
rect 150771 25029 150787 25147
rect 150477 7307 150787 25029
rect 150477 7189 150493 7307
rect 150611 7189 150653 7307
rect 150771 7189 150787 7307
rect 150477 7147 150787 7189
rect 150477 7029 150493 7147
rect 150611 7029 150653 7147
rect 150771 7029 150787 7147
rect 141477 -3651 141493 -3533
rect 141611 -3651 141653 -3533
rect 141771 -3651 141787 -3533
rect 141477 -3693 141787 -3651
rect 141477 -3811 141493 -3693
rect 141611 -3811 141653 -3693
rect 141771 -3811 141787 -3693
rect 141477 -3827 141787 -3811
rect 150477 -3053 150787 7029
rect 153897 352899 154207 352915
rect 153897 352781 153913 352899
rect 154031 352781 154073 352899
rect 154191 352781 154207 352899
rect 153897 352739 154207 352781
rect 153897 352621 153913 352739
rect 154031 352621 154073 352739
rect 154191 352621 154207 352739
rect 153897 334727 154207 352621
rect 153897 334609 153913 334727
rect 154031 334609 154073 334727
rect 154191 334609 154207 334727
rect 153897 334567 154207 334609
rect 153897 334449 153913 334567
rect 154031 334449 154073 334567
rect 154191 334449 154207 334567
rect 153897 316727 154207 334449
rect 153897 316609 153913 316727
rect 154031 316609 154073 316727
rect 154191 316609 154207 316727
rect 153897 316567 154207 316609
rect 153897 316449 153913 316567
rect 154031 316449 154073 316567
rect 154191 316449 154207 316567
rect 153897 298727 154207 316449
rect 153897 298609 153913 298727
rect 154031 298609 154073 298727
rect 154191 298609 154207 298727
rect 153897 298567 154207 298609
rect 153897 298449 153913 298567
rect 154031 298449 154073 298567
rect 154191 298449 154207 298567
rect 153897 280727 154207 298449
rect 153897 280609 153913 280727
rect 154031 280609 154073 280727
rect 154191 280609 154207 280727
rect 153897 280567 154207 280609
rect 153897 280449 153913 280567
rect 154031 280449 154073 280567
rect 154191 280449 154207 280567
rect 153897 262727 154207 280449
rect 153897 262609 153913 262727
rect 154031 262609 154073 262727
rect 154191 262609 154207 262727
rect 153897 262567 154207 262609
rect 153897 262449 153913 262567
rect 154031 262449 154073 262567
rect 154191 262449 154207 262567
rect 153897 244727 154207 262449
rect 153897 244609 153913 244727
rect 154031 244609 154073 244727
rect 154191 244609 154207 244727
rect 153897 244567 154207 244609
rect 153897 244449 153913 244567
rect 154031 244449 154073 244567
rect 154191 244449 154207 244567
rect 153897 226727 154207 244449
rect 153897 226609 153913 226727
rect 154031 226609 154073 226727
rect 154191 226609 154207 226727
rect 153897 226567 154207 226609
rect 153897 226449 153913 226567
rect 154031 226449 154073 226567
rect 154191 226449 154207 226567
rect 153897 208727 154207 226449
rect 153897 208609 153913 208727
rect 154031 208609 154073 208727
rect 154191 208609 154207 208727
rect 153897 208567 154207 208609
rect 153897 208449 153913 208567
rect 154031 208449 154073 208567
rect 154191 208449 154207 208567
rect 153897 190727 154207 208449
rect 153897 190609 153913 190727
rect 154031 190609 154073 190727
rect 154191 190609 154207 190727
rect 153897 190567 154207 190609
rect 153897 190449 153913 190567
rect 154031 190449 154073 190567
rect 154191 190449 154207 190567
rect 153897 172727 154207 190449
rect 153897 172609 153913 172727
rect 154031 172609 154073 172727
rect 154191 172609 154207 172727
rect 153897 172567 154207 172609
rect 153897 172449 153913 172567
rect 154031 172449 154073 172567
rect 154191 172449 154207 172567
rect 153897 154727 154207 172449
rect 153897 154609 153913 154727
rect 154031 154609 154073 154727
rect 154191 154609 154207 154727
rect 153897 154567 154207 154609
rect 153897 154449 153913 154567
rect 154031 154449 154073 154567
rect 154191 154449 154207 154567
rect 153897 136727 154207 154449
rect 153897 136609 153913 136727
rect 154031 136609 154073 136727
rect 154191 136609 154207 136727
rect 153897 136567 154207 136609
rect 153897 136449 153913 136567
rect 154031 136449 154073 136567
rect 154191 136449 154207 136567
rect 153897 118727 154207 136449
rect 153897 118609 153913 118727
rect 154031 118609 154073 118727
rect 154191 118609 154207 118727
rect 153897 118567 154207 118609
rect 153897 118449 153913 118567
rect 154031 118449 154073 118567
rect 154191 118449 154207 118567
rect 153897 100727 154207 118449
rect 153897 100609 153913 100727
rect 154031 100609 154073 100727
rect 154191 100609 154207 100727
rect 153897 100567 154207 100609
rect 153897 100449 153913 100567
rect 154031 100449 154073 100567
rect 154191 100449 154207 100567
rect 153897 82727 154207 100449
rect 153897 82609 153913 82727
rect 154031 82609 154073 82727
rect 154191 82609 154207 82727
rect 153897 82567 154207 82609
rect 153897 82449 153913 82567
rect 154031 82449 154073 82567
rect 154191 82449 154207 82567
rect 153897 64727 154207 82449
rect 153897 64609 153913 64727
rect 154031 64609 154073 64727
rect 154191 64609 154207 64727
rect 153897 64567 154207 64609
rect 153897 64449 153913 64567
rect 154031 64449 154073 64567
rect 154191 64449 154207 64567
rect 153897 46727 154207 64449
rect 153897 46609 153913 46727
rect 154031 46609 154073 46727
rect 154191 46609 154207 46727
rect 153897 46567 154207 46609
rect 153897 46449 153913 46567
rect 154031 46449 154073 46567
rect 154191 46449 154207 46567
rect 153897 28727 154207 46449
rect 153897 28609 153913 28727
rect 154031 28609 154073 28727
rect 154191 28609 154207 28727
rect 153897 28567 154207 28609
rect 153897 28449 153913 28567
rect 154031 28449 154073 28567
rect 154191 28449 154207 28567
rect 153897 10727 154207 28449
rect 153897 10609 153913 10727
rect 154031 10609 154073 10727
rect 154191 10609 154207 10727
rect 153897 10567 154207 10609
rect 153897 10449 153913 10567
rect 154031 10449 154073 10567
rect 154191 10449 154207 10567
rect 153897 -653 154207 10449
rect 153897 -771 153913 -653
rect 154031 -771 154073 -653
rect 154191 -771 154207 -653
rect 153897 -813 154207 -771
rect 153897 -931 153913 -813
rect 154031 -931 154073 -813
rect 154191 -931 154207 -813
rect 153897 -947 154207 -931
rect 155757 336587 156067 353581
rect 155757 336469 155773 336587
rect 155891 336469 155933 336587
rect 156051 336469 156067 336587
rect 155757 336427 156067 336469
rect 155757 336309 155773 336427
rect 155891 336309 155933 336427
rect 156051 336309 156067 336427
rect 155757 318587 156067 336309
rect 155757 318469 155773 318587
rect 155891 318469 155933 318587
rect 156051 318469 156067 318587
rect 155757 318427 156067 318469
rect 155757 318309 155773 318427
rect 155891 318309 155933 318427
rect 156051 318309 156067 318427
rect 155757 300587 156067 318309
rect 155757 300469 155773 300587
rect 155891 300469 155933 300587
rect 156051 300469 156067 300587
rect 155757 300427 156067 300469
rect 155757 300309 155773 300427
rect 155891 300309 155933 300427
rect 156051 300309 156067 300427
rect 155757 282587 156067 300309
rect 155757 282469 155773 282587
rect 155891 282469 155933 282587
rect 156051 282469 156067 282587
rect 155757 282427 156067 282469
rect 155757 282309 155773 282427
rect 155891 282309 155933 282427
rect 156051 282309 156067 282427
rect 155757 264587 156067 282309
rect 155757 264469 155773 264587
rect 155891 264469 155933 264587
rect 156051 264469 156067 264587
rect 155757 264427 156067 264469
rect 155757 264309 155773 264427
rect 155891 264309 155933 264427
rect 156051 264309 156067 264427
rect 155757 246587 156067 264309
rect 155757 246469 155773 246587
rect 155891 246469 155933 246587
rect 156051 246469 156067 246587
rect 155757 246427 156067 246469
rect 155757 246309 155773 246427
rect 155891 246309 155933 246427
rect 156051 246309 156067 246427
rect 155757 228587 156067 246309
rect 155757 228469 155773 228587
rect 155891 228469 155933 228587
rect 156051 228469 156067 228587
rect 155757 228427 156067 228469
rect 155757 228309 155773 228427
rect 155891 228309 155933 228427
rect 156051 228309 156067 228427
rect 155757 210587 156067 228309
rect 155757 210469 155773 210587
rect 155891 210469 155933 210587
rect 156051 210469 156067 210587
rect 155757 210427 156067 210469
rect 155757 210309 155773 210427
rect 155891 210309 155933 210427
rect 156051 210309 156067 210427
rect 155757 192587 156067 210309
rect 155757 192469 155773 192587
rect 155891 192469 155933 192587
rect 156051 192469 156067 192587
rect 155757 192427 156067 192469
rect 155757 192309 155773 192427
rect 155891 192309 155933 192427
rect 156051 192309 156067 192427
rect 155757 174587 156067 192309
rect 155757 174469 155773 174587
rect 155891 174469 155933 174587
rect 156051 174469 156067 174587
rect 155757 174427 156067 174469
rect 155757 174309 155773 174427
rect 155891 174309 155933 174427
rect 156051 174309 156067 174427
rect 155757 156587 156067 174309
rect 155757 156469 155773 156587
rect 155891 156469 155933 156587
rect 156051 156469 156067 156587
rect 155757 156427 156067 156469
rect 155757 156309 155773 156427
rect 155891 156309 155933 156427
rect 156051 156309 156067 156427
rect 155757 138587 156067 156309
rect 155757 138469 155773 138587
rect 155891 138469 155933 138587
rect 156051 138469 156067 138587
rect 155757 138427 156067 138469
rect 155757 138309 155773 138427
rect 155891 138309 155933 138427
rect 156051 138309 156067 138427
rect 155757 120587 156067 138309
rect 155757 120469 155773 120587
rect 155891 120469 155933 120587
rect 156051 120469 156067 120587
rect 155757 120427 156067 120469
rect 155757 120309 155773 120427
rect 155891 120309 155933 120427
rect 156051 120309 156067 120427
rect 155757 102587 156067 120309
rect 155757 102469 155773 102587
rect 155891 102469 155933 102587
rect 156051 102469 156067 102587
rect 155757 102427 156067 102469
rect 155757 102309 155773 102427
rect 155891 102309 155933 102427
rect 156051 102309 156067 102427
rect 155757 84587 156067 102309
rect 155757 84469 155773 84587
rect 155891 84469 155933 84587
rect 156051 84469 156067 84587
rect 155757 84427 156067 84469
rect 155757 84309 155773 84427
rect 155891 84309 155933 84427
rect 156051 84309 156067 84427
rect 155757 66587 156067 84309
rect 155757 66469 155773 66587
rect 155891 66469 155933 66587
rect 156051 66469 156067 66587
rect 155757 66427 156067 66469
rect 155757 66309 155773 66427
rect 155891 66309 155933 66427
rect 156051 66309 156067 66427
rect 155757 48587 156067 66309
rect 155757 48469 155773 48587
rect 155891 48469 155933 48587
rect 156051 48469 156067 48587
rect 155757 48427 156067 48469
rect 155757 48309 155773 48427
rect 155891 48309 155933 48427
rect 156051 48309 156067 48427
rect 155757 30587 156067 48309
rect 155757 30469 155773 30587
rect 155891 30469 155933 30587
rect 156051 30469 156067 30587
rect 155757 30427 156067 30469
rect 155757 30309 155773 30427
rect 155891 30309 155933 30427
rect 156051 30309 156067 30427
rect 155757 12587 156067 30309
rect 155757 12469 155773 12587
rect 155891 12469 155933 12587
rect 156051 12469 156067 12587
rect 155757 12427 156067 12469
rect 155757 12309 155773 12427
rect 155891 12309 155933 12427
rect 156051 12309 156067 12427
rect 155757 -1613 156067 12309
rect 155757 -1731 155773 -1613
rect 155891 -1731 155933 -1613
rect 156051 -1731 156067 -1613
rect 155757 -1773 156067 -1731
rect 155757 -1891 155773 -1773
rect 155891 -1891 155933 -1773
rect 156051 -1891 156067 -1773
rect 155757 -1907 156067 -1891
rect 157617 338447 157927 354541
rect 157617 338329 157633 338447
rect 157751 338329 157793 338447
rect 157911 338329 157927 338447
rect 157617 338287 157927 338329
rect 157617 338169 157633 338287
rect 157751 338169 157793 338287
rect 157911 338169 157927 338287
rect 157617 320447 157927 338169
rect 157617 320329 157633 320447
rect 157751 320329 157793 320447
rect 157911 320329 157927 320447
rect 157617 320287 157927 320329
rect 157617 320169 157633 320287
rect 157751 320169 157793 320287
rect 157911 320169 157927 320287
rect 157617 302447 157927 320169
rect 157617 302329 157633 302447
rect 157751 302329 157793 302447
rect 157911 302329 157927 302447
rect 157617 302287 157927 302329
rect 157617 302169 157633 302287
rect 157751 302169 157793 302287
rect 157911 302169 157927 302287
rect 157617 284447 157927 302169
rect 157617 284329 157633 284447
rect 157751 284329 157793 284447
rect 157911 284329 157927 284447
rect 157617 284287 157927 284329
rect 157617 284169 157633 284287
rect 157751 284169 157793 284287
rect 157911 284169 157927 284287
rect 157617 266447 157927 284169
rect 157617 266329 157633 266447
rect 157751 266329 157793 266447
rect 157911 266329 157927 266447
rect 157617 266287 157927 266329
rect 157617 266169 157633 266287
rect 157751 266169 157793 266287
rect 157911 266169 157927 266287
rect 157617 248447 157927 266169
rect 157617 248329 157633 248447
rect 157751 248329 157793 248447
rect 157911 248329 157927 248447
rect 157617 248287 157927 248329
rect 157617 248169 157633 248287
rect 157751 248169 157793 248287
rect 157911 248169 157927 248287
rect 157617 230447 157927 248169
rect 157617 230329 157633 230447
rect 157751 230329 157793 230447
rect 157911 230329 157927 230447
rect 157617 230287 157927 230329
rect 157617 230169 157633 230287
rect 157751 230169 157793 230287
rect 157911 230169 157927 230287
rect 157617 212447 157927 230169
rect 157617 212329 157633 212447
rect 157751 212329 157793 212447
rect 157911 212329 157927 212447
rect 157617 212287 157927 212329
rect 157617 212169 157633 212287
rect 157751 212169 157793 212287
rect 157911 212169 157927 212287
rect 157617 194447 157927 212169
rect 157617 194329 157633 194447
rect 157751 194329 157793 194447
rect 157911 194329 157927 194447
rect 157617 194287 157927 194329
rect 157617 194169 157633 194287
rect 157751 194169 157793 194287
rect 157911 194169 157927 194287
rect 157617 176447 157927 194169
rect 157617 176329 157633 176447
rect 157751 176329 157793 176447
rect 157911 176329 157927 176447
rect 157617 176287 157927 176329
rect 157617 176169 157633 176287
rect 157751 176169 157793 176287
rect 157911 176169 157927 176287
rect 157617 158447 157927 176169
rect 157617 158329 157633 158447
rect 157751 158329 157793 158447
rect 157911 158329 157927 158447
rect 157617 158287 157927 158329
rect 157617 158169 157633 158287
rect 157751 158169 157793 158287
rect 157911 158169 157927 158287
rect 157617 140447 157927 158169
rect 157617 140329 157633 140447
rect 157751 140329 157793 140447
rect 157911 140329 157927 140447
rect 157617 140287 157927 140329
rect 157617 140169 157633 140287
rect 157751 140169 157793 140287
rect 157911 140169 157927 140287
rect 157617 122447 157927 140169
rect 157617 122329 157633 122447
rect 157751 122329 157793 122447
rect 157911 122329 157927 122447
rect 157617 122287 157927 122329
rect 157617 122169 157633 122287
rect 157751 122169 157793 122287
rect 157911 122169 157927 122287
rect 157617 104447 157927 122169
rect 157617 104329 157633 104447
rect 157751 104329 157793 104447
rect 157911 104329 157927 104447
rect 157617 104287 157927 104329
rect 157617 104169 157633 104287
rect 157751 104169 157793 104287
rect 157911 104169 157927 104287
rect 157617 86447 157927 104169
rect 157617 86329 157633 86447
rect 157751 86329 157793 86447
rect 157911 86329 157927 86447
rect 157617 86287 157927 86329
rect 157617 86169 157633 86287
rect 157751 86169 157793 86287
rect 157911 86169 157927 86287
rect 157617 68447 157927 86169
rect 157617 68329 157633 68447
rect 157751 68329 157793 68447
rect 157911 68329 157927 68447
rect 157617 68287 157927 68329
rect 157617 68169 157633 68287
rect 157751 68169 157793 68287
rect 157911 68169 157927 68287
rect 157617 50447 157927 68169
rect 157617 50329 157633 50447
rect 157751 50329 157793 50447
rect 157911 50329 157927 50447
rect 157617 50287 157927 50329
rect 157617 50169 157633 50287
rect 157751 50169 157793 50287
rect 157911 50169 157927 50287
rect 157617 32447 157927 50169
rect 157617 32329 157633 32447
rect 157751 32329 157793 32447
rect 157911 32329 157927 32447
rect 157617 32287 157927 32329
rect 157617 32169 157633 32287
rect 157751 32169 157793 32287
rect 157911 32169 157927 32287
rect 157617 14447 157927 32169
rect 157617 14329 157633 14447
rect 157751 14329 157793 14447
rect 157911 14329 157927 14447
rect 157617 14287 157927 14329
rect 157617 14169 157633 14287
rect 157751 14169 157793 14287
rect 157911 14169 157927 14287
rect 157617 -2573 157927 14169
rect 157617 -2691 157633 -2573
rect 157751 -2691 157793 -2573
rect 157911 -2691 157927 -2573
rect 157617 -2733 157927 -2691
rect 157617 -2851 157633 -2733
rect 157751 -2851 157793 -2733
rect 157911 -2851 157927 -2733
rect 157617 -2867 157927 -2851
rect 159477 340307 159787 355501
rect 168477 355299 168787 355795
rect 168477 355181 168493 355299
rect 168611 355181 168653 355299
rect 168771 355181 168787 355299
rect 168477 355139 168787 355181
rect 168477 355021 168493 355139
rect 168611 355021 168653 355139
rect 168771 355021 168787 355139
rect 166617 354339 166927 354835
rect 166617 354221 166633 354339
rect 166751 354221 166793 354339
rect 166911 354221 166927 354339
rect 166617 354179 166927 354221
rect 166617 354061 166633 354179
rect 166751 354061 166793 354179
rect 166911 354061 166927 354179
rect 164757 353379 165067 353875
rect 164757 353261 164773 353379
rect 164891 353261 164933 353379
rect 165051 353261 165067 353379
rect 164757 353219 165067 353261
rect 164757 353101 164773 353219
rect 164891 353101 164933 353219
rect 165051 353101 165067 353219
rect 159477 340189 159493 340307
rect 159611 340189 159653 340307
rect 159771 340189 159787 340307
rect 159477 340147 159787 340189
rect 159477 340029 159493 340147
rect 159611 340029 159653 340147
rect 159771 340029 159787 340147
rect 159477 322307 159787 340029
rect 159477 322189 159493 322307
rect 159611 322189 159653 322307
rect 159771 322189 159787 322307
rect 159477 322147 159787 322189
rect 159477 322029 159493 322147
rect 159611 322029 159653 322147
rect 159771 322029 159787 322147
rect 159477 304307 159787 322029
rect 159477 304189 159493 304307
rect 159611 304189 159653 304307
rect 159771 304189 159787 304307
rect 159477 304147 159787 304189
rect 159477 304029 159493 304147
rect 159611 304029 159653 304147
rect 159771 304029 159787 304147
rect 159477 286307 159787 304029
rect 159477 286189 159493 286307
rect 159611 286189 159653 286307
rect 159771 286189 159787 286307
rect 159477 286147 159787 286189
rect 159477 286029 159493 286147
rect 159611 286029 159653 286147
rect 159771 286029 159787 286147
rect 159477 268307 159787 286029
rect 159477 268189 159493 268307
rect 159611 268189 159653 268307
rect 159771 268189 159787 268307
rect 159477 268147 159787 268189
rect 159477 268029 159493 268147
rect 159611 268029 159653 268147
rect 159771 268029 159787 268147
rect 159477 250307 159787 268029
rect 159477 250189 159493 250307
rect 159611 250189 159653 250307
rect 159771 250189 159787 250307
rect 159477 250147 159787 250189
rect 159477 250029 159493 250147
rect 159611 250029 159653 250147
rect 159771 250029 159787 250147
rect 159477 232307 159787 250029
rect 159477 232189 159493 232307
rect 159611 232189 159653 232307
rect 159771 232189 159787 232307
rect 159477 232147 159787 232189
rect 159477 232029 159493 232147
rect 159611 232029 159653 232147
rect 159771 232029 159787 232147
rect 159477 214307 159787 232029
rect 159477 214189 159493 214307
rect 159611 214189 159653 214307
rect 159771 214189 159787 214307
rect 159477 214147 159787 214189
rect 159477 214029 159493 214147
rect 159611 214029 159653 214147
rect 159771 214029 159787 214147
rect 159477 196307 159787 214029
rect 159477 196189 159493 196307
rect 159611 196189 159653 196307
rect 159771 196189 159787 196307
rect 159477 196147 159787 196189
rect 159477 196029 159493 196147
rect 159611 196029 159653 196147
rect 159771 196029 159787 196147
rect 159477 178307 159787 196029
rect 159477 178189 159493 178307
rect 159611 178189 159653 178307
rect 159771 178189 159787 178307
rect 159477 178147 159787 178189
rect 159477 178029 159493 178147
rect 159611 178029 159653 178147
rect 159771 178029 159787 178147
rect 159477 160307 159787 178029
rect 159477 160189 159493 160307
rect 159611 160189 159653 160307
rect 159771 160189 159787 160307
rect 159477 160147 159787 160189
rect 159477 160029 159493 160147
rect 159611 160029 159653 160147
rect 159771 160029 159787 160147
rect 159477 142307 159787 160029
rect 159477 142189 159493 142307
rect 159611 142189 159653 142307
rect 159771 142189 159787 142307
rect 159477 142147 159787 142189
rect 159477 142029 159493 142147
rect 159611 142029 159653 142147
rect 159771 142029 159787 142147
rect 159477 124307 159787 142029
rect 159477 124189 159493 124307
rect 159611 124189 159653 124307
rect 159771 124189 159787 124307
rect 159477 124147 159787 124189
rect 159477 124029 159493 124147
rect 159611 124029 159653 124147
rect 159771 124029 159787 124147
rect 159477 106307 159787 124029
rect 159477 106189 159493 106307
rect 159611 106189 159653 106307
rect 159771 106189 159787 106307
rect 159477 106147 159787 106189
rect 159477 106029 159493 106147
rect 159611 106029 159653 106147
rect 159771 106029 159787 106147
rect 159477 88307 159787 106029
rect 159477 88189 159493 88307
rect 159611 88189 159653 88307
rect 159771 88189 159787 88307
rect 159477 88147 159787 88189
rect 159477 88029 159493 88147
rect 159611 88029 159653 88147
rect 159771 88029 159787 88147
rect 159477 70307 159787 88029
rect 159477 70189 159493 70307
rect 159611 70189 159653 70307
rect 159771 70189 159787 70307
rect 159477 70147 159787 70189
rect 159477 70029 159493 70147
rect 159611 70029 159653 70147
rect 159771 70029 159787 70147
rect 159477 52307 159787 70029
rect 159477 52189 159493 52307
rect 159611 52189 159653 52307
rect 159771 52189 159787 52307
rect 159477 52147 159787 52189
rect 159477 52029 159493 52147
rect 159611 52029 159653 52147
rect 159771 52029 159787 52147
rect 159477 34307 159787 52029
rect 159477 34189 159493 34307
rect 159611 34189 159653 34307
rect 159771 34189 159787 34307
rect 159477 34147 159787 34189
rect 159477 34029 159493 34147
rect 159611 34029 159653 34147
rect 159771 34029 159787 34147
rect 159477 16307 159787 34029
rect 159477 16189 159493 16307
rect 159611 16189 159653 16307
rect 159771 16189 159787 16307
rect 159477 16147 159787 16189
rect 159477 16029 159493 16147
rect 159611 16029 159653 16147
rect 159771 16029 159787 16147
rect 150477 -3171 150493 -3053
rect 150611 -3171 150653 -3053
rect 150771 -3171 150787 -3053
rect 150477 -3213 150787 -3171
rect 150477 -3331 150493 -3213
rect 150611 -3331 150653 -3213
rect 150771 -3331 150787 -3213
rect 150477 -3827 150787 -3331
rect 159477 -3533 159787 16029
rect 162897 352419 163207 352915
rect 162897 352301 162913 352419
rect 163031 352301 163073 352419
rect 163191 352301 163207 352419
rect 162897 352259 163207 352301
rect 162897 352141 162913 352259
rect 163031 352141 163073 352259
rect 163191 352141 163207 352259
rect 162897 343727 163207 352141
rect 162897 343609 162913 343727
rect 163031 343609 163073 343727
rect 163191 343609 163207 343727
rect 162897 343567 163207 343609
rect 162897 343449 162913 343567
rect 163031 343449 163073 343567
rect 163191 343449 163207 343567
rect 162897 325727 163207 343449
rect 162897 325609 162913 325727
rect 163031 325609 163073 325727
rect 163191 325609 163207 325727
rect 162897 325567 163207 325609
rect 162897 325449 162913 325567
rect 163031 325449 163073 325567
rect 163191 325449 163207 325567
rect 162897 307727 163207 325449
rect 162897 307609 162913 307727
rect 163031 307609 163073 307727
rect 163191 307609 163207 307727
rect 162897 307567 163207 307609
rect 162897 307449 162913 307567
rect 163031 307449 163073 307567
rect 163191 307449 163207 307567
rect 162897 289727 163207 307449
rect 162897 289609 162913 289727
rect 163031 289609 163073 289727
rect 163191 289609 163207 289727
rect 162897 289567 163207 289609
rect 162897 289449 162913 289567
rect 163031 289449 163073 289567
rect 163191 289449 163207 289567
rect 162897 271727 163207 289449
rect 162897 271609 162913 271727
rect 163031 271609 163073 271727
rect 163191 271609 163207 271727
rect 162897 271567 163207 271609
rect 162897 271449 162913 271567
rect 163031 271449 163073 271567
rect 163191 271449 163207 271567
rect 162897 253727 163207 271449
rect 162897 253609 162913 253727
rect 163031 253609 163073 253727
rect 163191 253609 163207 253727
rect 162897 253567 163207 253609
rect 162897 253449 162913 253567
rect 163031 253449 163073 253567
rect 163191 253449 163207 253567
rect 162897 235727 163207 253449
rect 162897 235609 162913 235727
rect 163031 235609 163073 235727
rect 163191 235609 163207 235727
rect 162897 235567 163207 235609
rect 162897 235449 162913 235567
rect 163031 235449 163073 235567
rect 163191 235449 163207 235567
rect 162897 217727 163207 235449
rect 162897 217609 162913 217727
rect 163031 217609 163073 217727
rect 163191 217609 163207 217727
rect 162897 217567 163207 217609
rect 162897 217449 162913 217567
rect 163031 217449 163073 217567
rect 163191 217449 163207 217567
rect 162897 199727 163207 217449
rect 162897 199609 162913 199727
rect 163031 199609 163073 199727
rect 163191 199609 163207 199727
rect 162897 199567 163207 199609
rect 162897 199449 162913 199567
rect 163031 199449 163073 199567
rect 163191 199449 163207 199567
rect 162897 181727 163207 199449
rect 162897 181609 162913 181727
rect 163031 181609 163073 181727
rect 163191 181609 163207 181727
rect 162897 181567 163207 181609
rect 162897 181449 162913 181567
rect 163031 181449 163073 181567
rect 163191 181449 163207 181567
rect 162897 163727 163207 181449
rect 162897 163609 162913 163727
rect 163031 163609 163073 163727
rect 163191 163609 163207 163727
rect 162897 163567 163207 163609
rect 162897 163449 162913 163567
rect 163031 163449 163073 163567
rect 163191 163449 163207 163567
rect 162897 145727 163207 163449
rect 162897 145609 162913 145727
rect 163031 145609 163073 145727
rect 163191 145609 163207 145727
rect 162897 145567 163207 145609
rect 162897 145449 162913 145567
rect 163031 145449 163073 145567
rect 163191 145449 163207 145567
rect 162897 127727 163207 145449
rect 162897 127609 162913 127727
rect 163031 127609 163073 127727
rect 163191 127609 163207 127727
rect 162897 127567 163207 127609
rect 162897 127449 162913 127567
rect 163031 127449 163073 127567
rect 163191 127449 163207 127567
rect 162897 109727 163207 127449
rect 162897 109609 162913 109727
rect 163031 109609 163073 109727
rect 163191 109609 163207 109727
rect 162897 109567 163207 109609
rect 162897 109449 162913 109567
rect 163031 109449 163073 109567
rect 163191 109449 163207 109567
rect 162897 91727 163207 109449
rect 162897 91609 162913 91727
rect 163031 91609 163073 91727
rect 163191 91609 163207 91727
rect 162897 91567 163207 91609
rect 162897 91449 162913 91567
rect 163031 91449 163073 91567
rect 163191 91449 163207 91567
rect 162897 73727 163207 91449
rect 162897 73609 162913 73727
rect 163031 73609 163073 73727
rect 163191 73609 163207 73727
rect 162897 73567 163207 73609
rect 162897 73449 162913 73567
rect 163031 73449 163073 73567
rect 163191 73449 163207 73567
rect 162897 55727 163207 73449
rect 162897 55609 162913 55727
rect 163031 55609 163073 55727
rect 163191 55609 163207 55727
rect 162897 55567 163207 55609
rect 162897 55449 162913 55567
rect 163031 55449 163073 55567
rect 163191 55449 163207 55567
rect 162897 37727 163207 55449
rect 162897 37609 162913 37727
rect 163031 37609 163073 37727
rect 163191 37609 163207 37727
rect 162897 37567 163207 37609
rect 162897 37449 162913 37567
rect 163031 37449 163073 37567
rect 163191 37449 163207 37567
rect 162897 19727 163207 37449
rect 162897 19609 162913 19727
rect 163031 19609 163073 19727
rect 163191 19609 163207 19727
rect 162897 19567 163207 19609
rect 162897 19449 162913 19567
rect 163031 19449 163073 19567
rect 163191 19449 163207 19567
rect 162897 1727 163207 19449
rect 162897 1609 162913 1727
rect 163031 1609 163073 1727
rect 163191 1609 163207 1727
rect 162897 1567 163207 1609
rect 162897 1449 162913 1567
rect 163031 1449 163073 1567
rect 163191 1449 163207 1567
rect 162897 -173 163207 1449
rect 162897 -291 162913 -173
rect 163031 -291 163073 -173
rect 163191 -291 163207 -173
rect 162897 -333 163207 -291
rect 162897 -451 162913 -333
rect 163031 -451 163073 -333
rect 163191 -451 163207 -333
rect 162897 -947 163207 -451
rect 164757 345587 165067 353101
rect 164757 345469 164773 345587
rect 164891 345469 164933 345587
rect 165051 345469 165067 345587
rect 164757 345427 165067 345469
rect 164757 345309 164773 345427
rect 164891 345309 164933 345427
rect 165051 345309 165067 345427
rect 164757 327587 165067 345309
rect 164757 327469 164773 327587
rect 164891 327469 164933 327587
rect 165051 327469 165067 327587
rect 164757 327427 165067 327469
rect 164757 327309 164773 327427
rect 164891 327309 164933 327427
rect 165051 327309 165067 327427
rect 164757 309587 165067 327309
rect 164757 309469 164773 309587
rect 164891 309469 164933 309587
rect 165051 309469 165067 309587
rect 164757 309427 165067 309469
rect 164757 309309 164773 309427
rect 164891 309309 164933 309427
rect 165051 309309 165067 309427
rect 164757 291587 165067 309309
rect 164757 291469 164773 291587
rect 164891 291469 164933 291587
rect 165051 291469 165067 291587
rect 164757 291427 165067 291469
rect 164757 291309 164773 291427
rect 164891 291309 164933 291427
rect 165051 291309 165067 291427
rect 164757 273587 165067 291309
rect 164757 273469 164773 273587
rect 164891 273469 164933 273587
rect 165051 273469 165067 273587
rect 164757 273427 165067 273469
rect 164757 273309 164773 273427
rect 164891 273309 164933 273427
rect 165051 273309 165067 273427
rect 164757 255587 165067 273309
rect 164757 255469 164773 255587
rect 164891 255469 164933 255587
rect 165051 255469 165067 255587
rect 164757 255427 165067 255469
rect 164757 255309 164773 255427
rect 164891 255309 164933 255427
rect 165051 255309 165067 255427
rect 164757 237587 165067 255309
rect 164757 237469 164773 237587
rect 164891 237469 164933 237587
rect 165051 237469 165067 237587
rect 164757 237427 165067 237469
rect 164757 237309 164773 237427
rect 164891 237309 164933 237427
rect 165051 237309 165067 237427
rect 164757 219587 165067 237309
rect 164757 219469 164773 219587
rect 164891 219469 164933 219587
rect 165051 219469 165067 219587
rect 164757 219427 165067 219469
rect 164757 219309 164773 219427
rect 164891 219309 164933 219427
rect 165051 219309 165067 219427
rect 164757 201587 165067 219309
rect 164757 201469 164773 201587
rect 164891 201469 164933 201587
rect 165051 201469 165067 201587
rect 164757 201427 165067 201469
rect 164757 201309 164773 201427
rect 164891 201309 164933 201427
rect 165051 201309 165067 201427
rect 164757 183587 165067 201309
rect 164757 183469 164773 183587
rect 164891 183469 164933 183587
rect 165051 183469 165067 183587
rect 164757 183427 165067 183469
rect 164757 183309 164773 183427
rect 164891 183309 164933 183427
rect 165051 183309 165067 183427
rect 164757 165587 165067 183309
rect 164757 165469 164773 165587
rect 164891 165469 164933 165587
rect 165051 165469 165067 165587
rect 164757 165427 165067 165469
rect 164757 165309 164773 165427
rect 164891 165309 164933 165427
rect 165051 165309 165067 165427
rect 164757 147587 165067 165309
rect 164757 147469 164773 147587
rect 164891 147469 164933 147587
rect 165051 147469 165067 147587
rect 164757 147427 165067 147469
rect 164757 147309 164773 147427
rect 164891 147309 164933 147427
rect 165051 147309 165067 147427
rect 164757 129587 165067 147309
rect 164757 129469 164773 129587
rect 164891 129469 164933 129587
rect 165051 129469 165067 129587
rect 164757 129427 165067 129469
rect 164757 129309 164773 129427
rect 164891 129309 164933 129427
rect 165051 129309 165067 129427
rect 164757 111587 165067 129309
rect 164757 111469 164773 111587
rect 164891 111469 164933 111587
rect 165051 111469 165067 111587
rect 164757 111427 165067 111469
rect 164757 111309 164773 111427
rect 164891 111309 164933 111427
rect 165051 111309 165067 111427
rect 164757 93587 165067 111309
rect 164757 93469 164773 93587
rect 164891 93469 164933 93587
rect 165051 93469 165067 93587
rect 164757 93427 165067 93469
rect 164757 93309 164773 93427
rect 164891 93309 164933 93427
rect 165051 93309 165067 93427
rect 164757 75587 165067 93309
rect 164757 75469 164773 75587
rect 164891 75469 164933 75587
rect 165051 75469 165067 75587
rect 164757 75427 165067 75469
rect 164757 75309 164773 75427
rect 164891 75309 164933 75427
rect 165051 75309 165067 75427
rect 164757 57587 165067 75309
rect 164757 57469 164773 57587
rect 164891 57469 164933 57587
rect 165051 57469 165067 57587
rect 164757 57427 165067 57469
rect 164757 57309 164773 57427
rect 164891 57309 164933 57427
rect 165051 57309 165067 57427
rect 164757 39587 165067 57309
rect 164757 39469 164773 39587
rect 164891 39469 164933 39587
rect 165051 39469 165067 39587
rect 164757 39427 165067 39469
rect 164757 39309 164773 39427
rect 164891 39309 164933 39427
rect 165051 39309 165067 39427
rect 164757 21587 165067 39309
rect 164757 21469 164773 21587
rect 164891 21469 164933 21587
rect 165051 21469 165067 21587
rect 164757 21427 165067 21469
rect 164757 21309 164773 21427
rect 164891 21309 164933 21427
rect 165051 21309 165067 21427
rect 164757 3587 165067 21309
rect 164757 3469 164773 3587
rect 164891 3469 164933 3587
rect 165051 3469 165067 3587
rect 164757 3427 165067 3469
rect 164757 3309 164773 3427
rect 164891 3309 164933 3427
rect 165051 3309 165067 3427
rect 164757 -1133 165067 3309
rect 164757 -1251 164773 -1133
rect 164891 -1251 164933 -1133
rect 165051 -1251 165067 -1133
rect 164757 -1293 165067 -1251
rect 164757 -1411 164773 -1293
rect 164891 -1411 164933 -1293
rect 165051 -1411 165067 -1293
rect 164757 -1907 165067 -1411
rect 166617 347447 166927 354061
rect 166617 347329 166633 347447
rect 166751 347329 166793 347447
rect 166911 347329 166927 347447
rect 166617 347287 166927 347329
rect 166617 347169 166633 347287
rect 166751 347169 166793 347287
rect 166911 347169 166927 347287
rect 166617 329447 166927 347169
rect 166617 329329 166633 329447
rect 166751 329329 166793 329447
rect 166911 329329 166927 329447
rect 166617 329287 166927 329329
rect 166617 329169 166633 329287
rect 166751 329169 166793 329287
rect 166911 329169 166927 329287
rect 166617 311447 166927 329169
rect 166617 311329 166633 311447
rect 166751 311329 166793 311447
rect 166911 311329 166927 311447
rect 166617 311287 166927 311329
rect 166617 311169 166633 311287
rect 166751 311169 166793 311287
rect 166911 311169 166927 311287
rect 166617 293447 166927 311169
rect 166617 293329 166633 293447
rect 166751 293329 166793 293447
rect 166911 293329 166927 293447
rect 166617 293287 166927 293329
rect 166617 293169 166633 293287
rect 166751 293169 166793 293287
rect 166911 293169 166927 293287
rect 166617 275447 166927 293169
rect 166617 275329 166633 275447
rect 166751 275329 166793 275447
rect 166911 275329 166927 275447
rect 166617 275287 166927 275329
rect 166617 275169 166633 275287
rect 166751 275169 166793 275287
rect 166911 275169 166927 275287
rect 166617 257447 166927 275169
rect 166617 257329 166633 257447
rect 166751 257329 166793 257447
rect 166911 257329 166927 257447
rect 166617 257287 166927 257329
rect 166617 257169 166633 257287
rect 166751 257169 166793 257287
rect 166911 257169 166927 257287
rect 166617 239447 166927 257169
rect 166617 239329 166633 239447
rect 166751 239329 166793 239447
rect 166911 239329 166927 239447
rect 166617 239287 166927 239329
rect 166617 239169 166633 239287
rect 166751 239169 166793 239287
rect 166911 239169 166927 239287
rect 166617 221447 166927 239169
rect 166617 221329 166633 221447
rect 166751 221329 166793 221447
rect 166911 221329 166927 221447
rect 166617 221287 166927 221329
rect 166617 221169 166633 221287
rect 166751 221169 166793 221287
rect 166911 221169 166927 221287
rect 166617 203447 166927 221169
rect 166617 203329 166633 203447
rect 166751 203329 166793 203447
rect 166911 203329 166927 203447
rect 166617 203287 166927 203329
rect 166617 203169 166633 203287
rect 166751 203169 166793 203287
rect 166911 203169 166927 203287
rect 166617 185447 166927 203169
rect 166617 185329 166633 185447
rect 166751 185329 166793 185447
rect 166911 185329 166927 185447
rect 166617 185287 166927 185329
rect 166617 185169 166633 185287
rect 166751 185169 166793 185287
rect 166911 185169 166927 185287
rect 166617 167447 166927 185169
rect 166617 167329 166633 167447
rect 166751 167329 166793 167447
rect 166911 167329 166927 167447
rect 166617 167287 166927 167329
rect 166617 167169 166633 167287
rect 166751 167169 166793 167287
rect 166911 167169 166927 167287
rect 166617 149447 166927 167169
rect 166617 149329 166633 149447
rect 166751 149329 166793 149447
rect 166911 149329 166927 149447
rect 166617 149287 166927 149329
rect 166617 149169 166633 149287
rect 166751 149169 166793 149287
rect 166911 149169 166927 149287
rect 166617 131447 166927 149169
rect 166617 131329 166633 131447
rect 166751 131329 166793 131447
rect 166911 131329 166927 131447
rect 166617 131287 166927 131329
rect 166617 131169 166633 131287
rect 166751 131169 166793 131287
rect 166911 131169 166927 131287
rect 166617 113447 166927 131169
rect 166617 113329 166633 113447
rect 166751 113329 166793 113447
rect 166911 113329 166927 113447
rect 166617 113287 166927 113329
rect 166617 113169 166633 113287
rect 166751 113169 166793 113287
rect 166911 113169 166927 113287
rect 166617 95447 166927 113169
rect 166617 95329 166633 95447
rect 166751 95329 166793 95447
rect 166911 95329 166927 95447
rect 166617 95287 166927 95329
rect 166617 95169 166633 95287
rect 166751 95169 166793 95287
rect 166911 95169 166927 95287
rect 166617 77447 166927 95169
rect 166617 77329 166633 77447
rect 166751 77329 166793 77447
rect 166911 77329 166927 77447
rect 166617 77287 166927 77329
rect 166617 77169 166633 77287
rect 166751 77169 166793 77287
rect 166911 77169 166927 77287
rect 166617 59447 166927 77169
rect 166617 59329 166633 59447
rect 166751 59329 166793 59447
rect 166911 59329 166927 59447
rect 166617 59287 166927 59329
rect 166617 59169 166633 59287
rect 166751 59169 166793 59287
rect 166911 59169 166927 59287
rect 166617 41447 166927 59169
rect 166617 41329 166633 41447
rect 166751 41329 166793 41447
rect 166911 41329 166927 41447
rect 166617 41287 166927 41329
rect 166617 41169 166633 41287
rect 166751 41169 166793 41287
rect 166911 41169 166927 41287
rect 166617 23447 166927 41169
rect 166617 23329 166633 23447
rect 166751 23329 166793 23447
rect 166911 23329 166927 23447
rect 166617 23287 166927 23329
rect 166617 23169 166633 23287
rect 166751 23169 166793 23287
rect 166911 23169 166927 23287
rect 166617 5447 166927 23169
rect 166617 5329 166633 5447
rect 166751 5329 166793 5447
rect 166911 5329 166927 5447
rect 166617 5287 166927 5329
rect 166617 5169 166633 5287
rect 166751 5169 166793 5287
rect 166911 5169 166927 5287
rect 166617 -2093 166927 5169
rect 166617 -2211 166633 -2093
rect 166751 -2211 166793 -2093
rect 166911 -2211 166927 -2093
rect 166617 -2253 166927 -2211
rect 166617 -2371 166633 -2253
rect 166751 -2371 166793 -2253
rect 166911 -2371 166927 -2253
rect 166617 -2867 166927 -2371
rect 168477 349307 168787 355021
rect 177477 355779 177787 355795
rect 177477 355661 177493 355779
rect 177611 355661 177653 355779
rect 177771 355661 177787 355779
rect 177477 355619 177787 355661
rect 177477 355501 177493 355619
rect 177611 355501 177653 355619
rect 177771 355501 177787 355619
rect 175617 354819 175927 354835
rect 175617 354701 175633 354819
rect 175751 354701 175793 354819
rect 175911 354701 175927 354819
rect 175617 354659 175927 354701
rect 175617 354541 175633 354659
rect 175751 354541 175793 354659
rect 175911 354541 175927 354659
rect 173757 353859 174067 353875
rect 173757 353741 173773 353859
rect 173891 353741 173933 353859
rect 174051 353741 174067 353859
rect 173757 353699 174067 353741
rect 173757 353581 173773 353699
rect 173891 353581 173933 353699
rect 174051 353581 174067 353699
rect 168477 349189 168493 349307
rect 168611 349189 168653 349307
rect 168771 349189 168787 349307
rect 168477 349147 168787 349189
rect 168477 349029 168493 349147
rect 168611 349029 168653 349147
rect 168771 349029 168787 349147
rect 168477 331307 168787 349029
rect 168477 331189 168493 331307
rect 168611 331189 168653 331307
rect 168771 331189 168787 331307
rect 168477 331147 168787 331189
rect 168477 331029 168493 331147
rect 168611 331029 168653 331147
rect 168771 331029 168787 331147
rect 168477 313307 168787 331029
rect 168477 313189 168493 313307
rect 168611 313189 168653 313307
rect 168771 313189 168787 313307
rect 168477 313147 168787 313189
rect 168477 313029 168493 313147
rect 168611 313029 168653 313147
rect 168771 313029 168787 313147
rect 168477 295307 168787 313029
rect 168477 295189 168493 295307
rect 168611 295189 168653 295307
rect 168771 295189 168787 295307
rect 168477 295147 168787 295189
rect 168477 295029 168493 295147
rect 168611 295029 168653 295147
rect 168771 295029 168787 295147
rect 168477 277307 168787 295029
rect 168477 277189 168493 277307
rect 168611 277189 168653 277307
rect 168771 277189 168787 277307
rect 168477 277147 168787 277189
rect 168477 277029 168493 277147
rect 168611 277029 168653 277147
rect 168771 277029 168787 277147
rect 168477 259307 168787 277029
rect 168477 259189 168493 259307
rect 168611 259189 168653 259307
rect 168771 259189 168787 259307
rect 168477 259147 168787 259189
rect 168477 259029 168493 259147
rect 168611 259029 168653 259147
rect 168771 259029 168787 259147
rect 168477 241307 168787 259029
rect 168477 241189 168493 241307
rect 168611 241189 168653 241307
rect 168771 241189 168787 241307
rect 168477 241147 168787 241189
rect 168477 241029 168493 241147
rect 168611 241029 168653 241147
rect 168771 241029 168787 241147
rect 168477 223307 168787 241029
rect 168477 223189 168493 223307
rect 168611 223189 168653 223307
rect 168771 223189 168787 223307
rect 168477 223147 168787 223189
rect 168477 223029 168493 223147
rect 168611 223029 168653 223147
rect 168771 223029 168787 223147
rect 168477 205307 168787 223029
rect 168477 205189 168493 205307
rect 168611 205189 168653 205307
rect 168771 205189 168787 205307
rect 168477 205147 168787 205189
rect 168477 205029 168493 205147
rect 168611 205029 168653 205147
rect 168771 205029 168787 205147
rect 168477 187307 168787 205029
rect 168477 187189 168493 187307
rect 168611 187189 168653 187307
rect 168771 187189 168787 187307
rect 168477 187147 168787 187189
rect 168477 187029 168493 187147
rect 168611 187029 168653 187147
rect 168771 187029 168787 187147
rect 168477 169307 168787 187029
rect 168477 169189 168493 169307
rect 168611 169189 168653 169307
rect 168771 169189 168787 169307
rect 168477 169147 168787 169189
rect 168477 169029 168493 169147
rect 168611 169029 168653 169147
rect 168771 169029 168787 169147
rect 168477 151307 168787 169029
rect 168477 151189 168493 151307
rect 168611 151189 168653 151307
rect 168771 151189 168787 151307
rect 168477 151147 168787 151189
rect 168477 151029 168493 151147
rect 168611 151029 168653 151147
rect 168771 151029 168787 151147
rect 168477 133307 168787 151029
rect 168477 133189 168493 133307
rect 168611 133189 168653 133307
rect 168771 133189 168787 133307
rect 168477 133147 168787 133189
rect 168477 133029 168493 133147
rect 168611 133029 168653 133147
rect 168771 133029 168787 133147
rect 168477 115307 168787 133029
rect 168477 115189 168493 115307
rect 168611 115189 168653 115307
rect 168771 115189 168787 115307
rect 168477 115147 168787 115189
rect 168477 115029 168493 115147
rect 168611 115029 168653 115147
rect 168771 115029 168787 115147
rect 168477 97307 168787 115029
rect 168477 97189 168493 97307
rect 168611 97189 168653 97307
rect 168771 97189 168787 97307
rect 168477 97147 168787 97189
rect 168477 97029 168493 97147
rect 168611 97029 168653 97147
rect 168771 97029 168787 97147
rect 168477 79307 168787 97029
rect 168477 79189 168493 79307
rect 168611 79189 168653 79307
rect 168771 79189 168787 79307
rect 168477 79147 168787 79189
rect 168477 79029 168493 79147
rect 168611 79029 168653 79147
rect 168771 79029 168787 79147
rect 168477 61307 168787 79029
rect 168477 61189 168493 61307
rect 168611 61189 168653 61307
rect 168771 61189 168787 61307
rect 168477 61147 168787 61189
rect 168477 61029 168493 61147
rect 168611 61029 168653 61147
rect 168771 61029 168787 61147
rect 168477 43307 168787 61029
rect 168477 43189 168493 43307
rect 168611 43189 168653 43307
rect 168771 43189 168787 43307
rect 168477 43147 168787 43189
rect 168477 43029 168493 43147
rect 168611 43029 168653 43147
rect 168771 43029 168787 43147
rect 168477 25307 168787 43029
rect 168477 25189 168493 25307
rect 168611 25189 168653 25307
rect 168771 25189 168787 25307
rect 168477 25147 168787 25189
rect 168477 25029 168493 25147
rect 168611 25029 168653 25147
rect 168771 25029 168787 25147
rect 168477 7307 168787 25029
rect 168477 7189 168493 7307
rect 168611 7189 168653 7307
rect 168771 7189 168787 7307
rect 168477 7147 168787 7189
rect 168477 7029 168493 7147
rect 168611 7029 168653 7147
rect 168771 7029 168787 7147
rect 159477 -3651 159493 -3533
rect 159611 -3651 159653 -3533
rect 159771 -3651 159787 -3533
rect 159477 -3693 159787 -3651
rect 159477 -3811 159493 -3693
rect 159611 -3811 159653 -3693
rect 159771 -3811 159787 -3693
rect 159477 -3827 159787 -3811
rect 168477 -3053 168787 7029
rect 171897 352899 172207 352915
rect 171897 352781 171913 352899
rect 172031 352781 172073 352899
rect 172191 352781 172207 352899
rect 171897 352739 172207 352781
rect 171897 352621 171913 352739
rect 172031 352621 172073 352739
rect 172191 352621 172207 352739
rect 171897 334727 172207 352621
rect 171897 334609 171913 334727
rect 172031 334609 172073 334727
rect 172191 334609 172207 334727
rect 171897 334567 172207 334609
rect 171897 334449 171913 334567
rect 172031 334449 172073 334567
rect 172191 334449 172207 334567
rect 171897 316727 172207 334449
rect 171897 316609 171913 316727
rect 172031 316609 172073 316727
rect 172191 316609 172207 316727
rect 171897 316567 172207 316609
rect 171897 316449 171913 316567
rect 172031 316449 172073 316567
rect 172191 316449 172207 316567
rect 171897 298727 172207 316449
rect 171897 298609 171913 298727
rect 172031 298609 172073 298727
rect 172191 298609 172207 298727
rect 171897 298567 172207 298609
rect 171897 298449 171913 298567
rect 172031 298449 172073 298567
rect 172191 298449 172207 298567
rect 171897 280727 172207 298449
rect 171897 280609 171913 280727
rect 172031 280609 172073 280727
rect 172191 280609 172207 280727
rect 171897 280567 172207 280609
rect 171897 280449 171913 280567
rect 172031 280449 172073 280567
rect 172191 280449 172207 280567
rect 171897 262727 172207 280449
rect 171897 262609 171913 262727
rect 172031 262609 172073 262727
rect 172191 262609 172207 262727
rect 171897 262567 172207 262609
rect 171897 262449 171913 262567
rect 172031 262449 172073 262567
rect 172191 262449 172207 262567
rect 171897 244727 172207 262449
rect 171897 244609 171913 244727
rect 172031 244609 172073 244727
rect 172191 244609 172207 244727
rect 171897 244567 172207 244609
rect 171897 244449 171913 244567
rect 172031 244449 172073 244567
rect 172191 244449 172207 244567
rect 171897 226727 172207 244449
rect 171897 226609 171913 226727
rect 172031 226609 172073 226727
rect 172191 226609 172207 226727
rect 171897 226567 172207 226609
rect 171897 226449 171913 226567
rect 172031 226449 172073 226567
rect 172191 226449 172207 226567
rect 171897 208727 172207 226449
rect 171897 208609 171913 208727
rect 172031 208609 172073 208727
rect 172191 208609 172207 208727
rect 171897 208567 172207 208609
rect 171897 208449 171913 208567
rect 172031 208449 172073 208567
rect 172191 208449 172207 208567
rect 171897 190727 172207 208449
rect 171897 190609 171913 190727
rect 172031 190609 172073 190727
rect 172191 190609 172207 190727
rect 171897 190567 172207 190609
rect 171897 190449 171913 190567
rect 172031 190449 172073 190567
rect 172191 190449 172207 190567
rect 171897 172727 172207 190449
rect 171897 172609 171913 172727
rect 172031 172609 172073 172727
rect 172191 172609 172207 172727
rect 171897 172567 172207 172609
rect 171897 172449 171913 172567
rect 172031 172449 172073 172567
rect 172191 172449 172207 172567
rect 171897 154727 172207 172449
rect 171897 154609 171913 154727
rect 172031 154609 172073 154727
rect 172191 154609 172207 154727
rect 171897 154567 172207 154609
rect 171897 154449 171913 154567
rect 172031 154449 172073 154567
rect 172191 154449 172207 154567
rect 171897 136727 172207 154449
rect 171897 136609 171913 136727
rect 172031 136609 172073 136727
rect 172191 136609 172207 136727
rect 171897 136567 172207 136609
rect 171897 136449 171913 136567
rect 172031 136449 172073 136567
rect 172191 136449 172207 136567
rect 171897 118727 172207 136449
rect 171897 118609 171913 118727
rect 172031 118609 172073 118727
rect 172191 118609 172207 118727
rect 171897 118567 172207 118609
rect 171897 118449 171913 118567
rect 172031 118449 172073 118567
rect 172191 118449 172207 118567
rect 171897 100727 172207 118449
rect 171897 100609 171913 100727
rect 172031 100609 172073 100727
rect 172191 100609 172207 100727
rect 171897 100567 172207 100609
rect 171897 100449 171913 100567
rect 172031 100449 172073 100567
rect 172191 100449 172207 100567
rect 171897 82727 172207 100449
rect 171897 82609 171913 82727
rect 172031 82609 172073 82727
rect 172191 82609 172207 82727
rect 171897 82567 172207 82609
rect 171897 82449 171913 82567
rect 172031 82449 172073 82567
rect 172191 82449 172207 82567
rect 171897 64727 172207 82449
rect 171897 64609 171913 64727
rect 172031 64609 172073 64727
rect 172191 64609 172207 64727
rect 171897 64567 172207 64609
rect 171897 64449 171913 64567
rect 172031 64449 172073 64567
rect 172191 64449 172207 64567
rect 171897 46727 172207 64449
rect 171897 46609 171913 46727
rect 172031 46609 172073 46727
rect 172191 46609 172207 46727
rect 171897 46567 172207 46609
rect 171897 46449 171913 46567
rect 172031 46449 172073 46567
rect 172191 46449 172207 46567
rect 171897 28727 172207 46449
rect 171897 28609 171913 28727
rect 172031 28609 172073 28727
rect 172191 28609 172207 28727
rect 171897 28567 172207 28609
rect 171897 28449 171913 28567
rect 172031 28449 172073 28567
rect 172191 28449 172207 28567
rect 171897 10727 172207 28449
rect 171897 10609 171913 10727
rect 172031 10609 172073 10727
rect 172191 10609 172207 10727
rect 171897 10567 172207 10609
rect 171897 10449 171913 10567
rect 172031 10449 172073 10567
rect 172191 10449 172207 10567
rect 171897 -653 172207 10449
rect 171897 -771 171913 -653
rect 172031 -771 172073 -653
rect 172191 -771 172207 -653
rect 171897 -813 172207 -771
rect 171897 -931 171913 -813
rect 172031 -931 172073 -813
rect 172191 -931 172207 -813
rect 171897 -947 172207 -931
rect 173757 336587 174067 353581
rect 173757 336469 173773 336587
rect 173891 336469 173933 336587
rect 174051 336469 174067 336587
rect 173757 336427 174067 336469
rect 173757 336309 173773 336427
rect 173891 336309 173933 336427
rect 174051 336309 174067 336427
rect 173757 318587 174067 336309
rect 173757 318469 173773 318587
rect 173891 318469 173933 318587
rect 174051 318469 174067 318587
rect 173757 318427 174067 318469
rect 173757 318309 173773 318427
rect 173891 318309 173933 318427
rect 174051 318309 174067 318427
rect 173757 300587 174067 318309
rect 173757 300469 173773 300587
rect 173891 300469 173933 300587
rect 174051 300469 174067 300587
rect 173757 300427 174067 300469
rect 173757 300309 173773 300427
rect 173891 300309 173933 300427
rect 174051 300309 174067 300427
rect 173757 282587 174067 300309
rect 173757 282469 173773 282587
rect 173891 282469 173933 282587
rect 174051 282469 174067 282587
rect 173757 282427 174067 282469
rect 173757 282309 173773 282427
rect 173891 282309 173933 282427
rect 174051 282309 174067 282427
rect 173757 264587 174067 282309
rect 173757 264469 173773 264587
rect 173891 264469 173933 264587
rect 174051 264469 174067 264587
rect 173757 264427 174067 264469
rect 173757 264309 173773 264427
rect 173891 264309 173933 264427
rect 174051 264309 174067 264427
rect 173757 246587 174067 264309
rect 173757 246469 173773 246587
rect 173891 246469 173933 246587
rect 174051 246469 174067 246587
rect 173757 246427 174067 246469
rect 173757 246309 173773 246427
rect 173891 246309 173933 246427
rect 174051 246309 174067 246427
rect 173757 228587 174067 246309
rect 173757 228469 173773 228587
rect 173891 228469 173933 228587
rect 174051 228469 174067 228587
rect 173757 228427 174067 228469
rect 173757 228309 173773 228427
rect 173891 228309 173933 228427
rect 174051 228309 174067 228427
rect 173757 210587 174067 228309
rect 173757 210469 173773 210587
rect 173891 210469 173933 210587
rect 174051 210469 174067 210587
rect 173757 210427 174067 210469
rect 173757 210309 173773 210427
rect 173891 210309 173933 210427
rect 174051 210309 174067 210427
rect 173757 192587 174067 210309
rect 173757 192469 173773 192587
rect 173891 192469 173933 192587
rect 174051 192469 174067 192587
rect 173757 192427 174067 192469
rect 173757 192309 173773 192427
rect 173891 192309 173933 192427
rect 174051 192309 174067 192427
rect 173757 174587 174067 192309
rect 173757 174469 173773 174587
rect 173891 174469 173933 174587
rect 174051 174469 174067 174587
rect 173757 174427 174067 174469
rect 173757 174309 173773 174427
rect 173891 174309 173933 174427
rect 174051 174309 174067 174427
rect 173757 156587 174067 174309
rect 173757 156469 173773 156587
rect 173891 156469 173933 156587
rect 174051 156469 174067 156587
rect 173757 156427 174067 156469
rect 173757 156309 173773 156427
rect 173891 156309 173933 156427
rect 174051 156309 174067 156427
rect 173757 138587 174067 156309
rect 173757 138469 173773 138587
rect 173891 138469 173933 138587
rect 174051 138469 174067 138587
rect 173757 138427 174067 138469
rect 173757 138309 173773 138427
rect 173891 138309 173933 138427
rect 174051 138309 174067 138427
rect 173757 120587 174067 138309
rect 173757 120469 173773 120587
rect 173891 120469 173933 120587
rect 174051 120469 174067 120587
rect 173757 120427 174067 120469
rect 173757 120309 173773 120427
rect 173891 120309 173933 120427
rect 174051 120309 174067 120427
rect 173757 102587 174067 120309
rect 173757 102469 173773 102587
rect 173891 102469 173933 102587
rect 174051 102469 174067 102587
rect 173757 102427 174067 102469
rect 173757 102309 173773 102427
rect 173891 102309 173933 102427
rect 174051 102309 174067 102427
rect 173757 84587 174067 102309
rect 173757 84469 173773 84587
rect 173891 84469 173933 84587
rect 174051 84469 174067 84587
rect 173757 84427 174067 84469
rect 173757 84309 173773 84427
rect 173891 84309 173933 84427
rect 174051 84309 174067 84427
rect 173757 66587 174067 84309
rect 173757 66469 173773 66587
rect 173891 66469 173933 66587
rect 174051 66469 174067 66587
rect 173757 66427 174067 66469
rect 173757 66309 173773 66427
rect 173891 66309 173933 66427
rect 174051 66309 174067 66427
rect 173757 48587 174067 66309
rect 173757 48469 173773 48587
rect 173891 48469 173933 48587
rect 174051 48469 174067 48587
rect 173757 48427 174067 48469
rect 173757 48309 173773 48427
rect 173891 48309 173933 48427
rect 174051 48309 174067 48427
rect 173757 30587 174067 48309
rect 173757 30469 173773 30587
rect 173891 30469 173933 30587
rect 174051 30469 174067 30587
rect 173757 30427 174067 30469
rect 173757 30309 173773 30427
rect 173891 30309 173933 30427
rect 174051 30309 174067 30427
rect 173757 12587 174067 30309
rect 173757 12469 173773 12587
rect 173891 12469 173933 12587
rect 174051 12469 174067 12587
rect 173757 12427 174067 12469
rect 173757 12309 173773 12427
rect 173891 12309 173933 12427
rect 174051 12309 174067 12427
rect 173757 -1613 174067 12309
rect 173757 -1731 173773 -1613
rect 173891 -1731 173933 -1613
rect 174051 -1731 174067 -1613
rect 173757 -1773 174067 -1731
rect 173757 -1891 173773 -1773
rect 173891 -1891 173933 -1773
rect 174051 -1891 174067 -1773
rect 173757 -1907 174067 -1891
rect 175617 338447 175927 354541
rect 175617 338329 175633 338447
rect 175751 338329 175793 338447
rect 175911 338329 175927 338447
rect 175617 338287 175927 338329
rect 175617 338169 175633 338287
rect 175751 338169 175793 338287
rect 175911 338169 175927 338287
rect 175617 320447 175927 338169
rect 175617 320329 175633 320447
rect 175751 320329 175793 320447
rect 175911 320329 175927 320447
rect 175617 320287 175927 320329
rect 175617 320169 175633 320287
rect 175751 320169 175793 320287
rect 175911 320169 175927 320287
rect 175617 302447 175927 320169
rect 175617 302329 175633 302447
rect 175751 302329 175793 302447
rect 175911 302329 175927 302447
rect 175617 302287 175927 302329
rect 175617 302169 175633 302287
rect 175751 302169 175793 302287
rect 175911 302169 175927 302287
rect 175617 284447 175927 302169
rect 175617 284329 175633 284447
rect 175751 284329 175793 284447
rect 175911 284329 175927 284447
rect 175617 284287 175927 284329
rect 175617 284169 175633 284287
rect 175751 284169 175793 284287
rect 175911 284169 175927 284287
rect 175617 266447 175927 284169
rect 175617 266329 175633 266447
rect 175751 266329 175793 266447
rect 175911 266329 175927 266447
rect 175617 266287 175927 266329
rect 175617 266169 175633 266287
rect 175751 266169 175793 266287
rect 175911 266169 175927 266287
rect 175617 248447 175927 266169
rect 175617 248329 175633 248447
rect 175751 248329 175793 248447
rect 175911 248329 175927 248447
rect 175617 248287 175927 248329
rect 175617 248169 175633 248287
rect 175751 248169 175793 248287
rect 175911 248169 175927 248287
rect 175617 230447 175927 248169
rect 175617 230329 175633 230447
rect 175751 230329 175793 230447
rect 175911 230329 175927 230447
rect 175617 230287 175927 230329
rect 175617 230169 175633 230287
rect 175751 230169 175793 230287
rect 175911 230169 175927 230287
rect 175617 212447 175927 230169
rect 175617 212329 175633 212447
rect 175751 212329 175793 212447
rect 175911 212329 175927 212447
rect 175617 212287 175927 212329
rect 175617 212169 175633 212287
rect 175751 212169 175793 212287
rect 175911 212169 175927 212287
rect 175617 194447 175927 212169
rect 175617 194329 175633 194447
rect 175751 194329 175793 194447
rect 175911 194329 175927 194447
rect 175617 194287 175927 194329
rect 175617 194169 175633 194287
rect 175751 194169 175793 194287
rect 175911 194169 175927 194287
rect 175617 176447 175927 194169
rect 175617 176329 175633 176447
rect 175751 176329 175793 176447
rect 175911 176329 175927 176447
rect 175617 176287 175927 176329
rect 175617 176169 175633 176287
rect 175751 176169 175793 176287
rect 175911 176169 175927 176287
rect 175617 158447 175927 176169
rect 175617 158329 175633 158447
rect 175751 158329 175793 158447
rect 175911 158329 175927 158447
rect 175617 158287 175927 158329
rect 175617 158169 175633 158287
rect 175751 158169 175793 158287
rect 175911 158169 175927 158287
rect 175617 140447 175927 158169
rect 175617 140329 175633 140447
rect 175751 140329 175793 140447
rect 175911 140329 175927 140447
rect 175617 140287 175927 140329
rect 175617 140169 175633 140287
rect 175751 140169 175793 140287
rect 175911 140169 175927 140287
rect 175617 122447 175927 140169
rect 175617 122329 175633 122447
rect 175751 122329 175793 122447
rect 175911 122329 175927 122447
rect 175617 122287 175927 122329
rect 175617 122169 175633 122287
rect 175751 122169 175793 122287
rect 175911 122169 175927 122287
rect 175617 104447 175927 122169
rect 175617 104329 175633 104447
rect 175751 104329 175793 104447
rect 175911 104329 175927 104447
rect 175617 104287 175927 104329
rect 175617 104169 175633 104287
rect 175751 104169 175793 104287
rect 175911 104169 175927 104287
rect 175617 86447 175927 104169
rect 175617 86329 175633 86447
rect 175751 86329 175793 86447
rect 175911 86329 175927 86447
rect 175617 86287 175927 86329
rect 175617 86169 175633 86287
rect 175751 86169 175793 86287
rect 175911 86169 175927 86287
rect 175617 68447 175927 86169
rect 175617 68329 175633 68447
rect 175751 68329 175793 68447
rect 175911 68329 175927 68447
rect 175617 68287 175927 68329
rect 175617 68169 175633 68287
rect 175751 68169 175793 68287
rect 175911 68169 175927 68287
rect 175617 50447 175927 68169
rect 175617 50329 175633 50447
rect 175751 50329 175793 50447
rect 175911 50329 175927 50447
rect 175617 50287 175927 50329
rect 175617 50169 175633 50287
rect 175751 50169 175793 50287
rect 175911 50169 175927 50287
rect 175617 32447 175927 50169
rect 175617 32329 175633 32447
rect 175751 32329 175793 32447
rect 175911 32329 175927 32447
rect 175617 32287 175927 32329
rect 175617 32169 175633 32287
rect 175751 32169 175793 32287
rect 175911 32169 175927 32287
rect 175617 14447 175927 32169
rect 175617 14329 175633 14447
rect 175751 14329 175793 14447
rect 175911 14329 175927 14447
rect 175617 14287 175927 14329
rect 175617 14169 175633 14287
rect 175751 14169 175793 14287
rect 175911 14169 175927 14287
rect 175617 -2573 175927 14169
rect 175617 -2691 175633 -2573
rect 175751 -2691 175793 -2573
rect 175911 -2691 175927 -2573
rect 175617 -2733 175927 -2691
rect 175617 -2851 175633 -2733
rect 175751 -2851 175793 -2733
rect 175911 -2851 175927 -2733
rect 175617 -2867 175927 -2851
rect 177477 340307 177787 355501
rect 186477 355299 186787 355795
rect 186477 355181 186493 355299
rect 186611 355181 186653 355299
rect 186771 355181 186787 355299
rect 186477 355139 186787 355181
rect 186477 355021 186493 355139
rect 186611 355021 186653 355139
rect 186771 355021 186787 355139
rect 184617 354339 184927 354835
rect 184617 354221 184633 354339
rect 184751 354221 184793 354339
rect 184911 354221 184927 354339
rect 184617 354179 184927 354221
rect 184617 354061 184633 354179
rect 184751 354061 184793 354179
rect 184911 354061 184927 354179
rect 182757 353379 183067 353875
rect 182757 353261 182773 353379
rect 182891 353261 182933 353379
rect 183051 353261 183067 353379
rect 182757 353219 183067 353261
rect 182757 353101 182773 353219
rect 182891 353101 182933 353219
rect 183051 353101 183067 353219
rect 177477 340189 177493 340307
rect 177611 340189 177653 340307
rect 177771 340189 177787 340307
rect 177477 340147 177787 340189
rect 177477 340029 177493 340147
rect 177611 340029 177653 340147
rect 177771 340029 177787 340147
rect 177477 322307 177787 340029
rect 177477 322189 177493 322307
rect 177611 322189 177653 322307
rect 177771 322189 177787 322307
rect 177477 322147 177787 322189
rect 177477 322029 177493 322147
rect 177611 322029 177653 322147
rect 177771 322029 177787 322147
rect 177477 304307 177787 322029
rect 177477 304189 177493 304307
rect 177611 304189 177653 304307
rect 177771 304189 177787 304307
rect 177477 304147 177787 304189
rect 177477 304029 177493 304147
rect 177611 304029 177653 304147
rect 177771 304029 177787 304147
rect 177477 286307 177787 304029
rect 177477 286189 177493 286307
rect 177611 286189 177653 286307
rect 177771 286189 177787 286307
rect 177477 286147 177787 286189
rect 177477 286029 177493 286147
rect 177611 286029 177653 286147
rect 177771 286029 177787 286147
rect 177477 268307 177787 286029
rect 177477 268189 177493 268307
rect 177611 268189 177653 268307
rect 177771 268189 177787 268307
rect 177477 268147 177787 268189
rect 177477 268029 177493 268147
rect 177611 268029 177653 268147
rect 177771 268029 177787 268147
rect 177477 250307 177787 268029
rect 177477 250189 177493 250307
rect 177611 250189 177653 250307
rect 177771 250189 177787 250307
rect 177477 250147 177787 250189
rect 177477 250029 177493 250147
rect 177611 250029 177653 250147
rect 177771 250029 177787 250147
rect 177477 232307 177787 250029
rect 177477 232189 177493 232307
rect 177611 232189 177653 232307
rect 177771 232189 177787 232307
rect 177477 232147 177787 232189
rect 177477 232029 177493 232147
rect 177611 232029 177653 232147
rect 177771 232029 177787 232147
rect 177477 214307 177787 232029
rect 177477 214189 177493 214307
rect 177611 214189 177653 214307
rect 177771 214189 177787 214307
rect 177477 214147 177787 214189
rect 177477 214029 177493 214147
rect 177611 214029 177653 214147
rect 177771 214029 177787 214147
rect 177477 196307 177787 214029
rect 177477 196189 177493 196307
rect 177611 196189 177653 196307
rect 177771 196189 177787 196307
rect 177477 196147 177787 196189
rect 177477 196029 177493 196147
rect 177611 196029 177653 196147
rect 177771 196029 177787 196147
rect 177477 178307 177787 196029
rect 177477 178189 177493 178307
rect 177611 178189 177653 178307
rect 177771 178189 177787 178307
rect 177477 178147 177787 178189
rect 177477 178029 177493 178147
rect 177611 178029 177653 178147
rect 177771 178029 177787 178147
rect 177477 160307 177787 178029
rect 177477 160189 177493 160307
rect 177611 160189 177653 160307
rect 177771 160189 177787 160307
rect 177477 160147 177787 160189
rect 177477 160029 177493 160147
rect 177611 160029 177653 160147
rect 177771 160029 177787 160147
rect 177477 142307 177787 160029
rect 177477 142189 177493 142307
rect 177611 142189 177653 142307
rect 177771 142189 177787 142307
rect 177477 142147 177787 142189
rect 177477 142029 177493 142147
rect 177611 142029 177653 142147
rect 177771 142029 177787 142147
rect 177477 124307 177787 142029
rect 177477 124189 177493 124307
rect 177611 124189 177653 124307
rect 177771 124189 177787 124307
rect 177477 124147 177787 124189
rect 177477 124029 177493 124147
rect 177611 124029 177653 124147
rect 177771 124029 177787 124147
rect 177477 106307 177787 124029
rect 177477 106189 177493 106307
rect 177611 106189 177653 106307
rect 177771 106189 177787 106307
rect 177477 106147 177787 106189
rect 177477 106029 177493 106147
rect 177611 106029 177653 106147
rect 177771 106029 177787 106147
rect 177477 88307 177787 106029
rect 177477 88189 177493 88307
rect 177611 88189 177653 88307
rect 177771 88189 177787 88307
rect 177477 88147 177787 88189
rect 177477 88029 177493 88147
rect 177611 88029 177653 88147
rect 177771 88029 177787 88147
rect 177477 70307 177787 88029
rect 177477 70189 177493 70307
rect 177611 70189 177653 70307
rect 177771 70189 177787 70307
rect 177477 70147 177787 70189
rect 177477 70029 177493 70147
rect 177611 70029 177653 70147
rect 177771 70029 177787 70147
rect 177477 52307 177787 70029
rect 177477 52189 177493 52307
rect 177611 52189 177653 52307
rect 177771 52189 177787 52307
rect 177477 52147 177787 52189
rect 177477 52029 177493 52147
rect 177611 52029 177653 52147
rect 177771 52029 177787 52147
rect 177477 34307 177787 52029
rect 177477 34189 177493 34307
rect 177611 34189 177653 34307
rect 177771 34189 177787 34307
rect 177477 34147 177787 34189
rect 177477 34029 177493 34147
rect 177611 34029 177653 34147
rect 177771 34029 177787 34147
rect 177477 16307 177787 34029
rect 177477 16189 177493 16307
rect 177611 16189 177653 16307
rect 177771 16189 177787 16307
rect 177477 16147 177787 16189
rect 177477 16029 177493 16147
rect 177611 16029 177653 16147
rect 177771 16029 177787 16147
rect 168477 -3171 168493 -3053
rect 168611 -3171 168653 -3053
rect 168771 -3171 168787 -3053
rect 168477 -3213 168787 -3171
rect 168477 -3331 168493 -3213
rect 168611 -3331 168653 -3213
rect 168771 -3331 168787 -3213
rect 168477 -3827 168787 -3331
rect 177477 -3533 177787 16029
rect 180897 352419 181207 352915
rect 180897 352301 180913 352419
rect 181031 352301 181073 352419
rect 181191 352301 181207 352419
rect 180897 352259 181207 352301
rect 180897 352141 180913 352259
rect 181031 352141 181073 352259
rect 181191 352141 181207 352259
rect 180897 343727 181207 352141
rect 180897 343609 180913 343727
rect 181031 343609 181073 343727
rect 181191 343609 181207 343727
rect 180897 343567 181207 343609
rect 180897 343449 180913 343567
rect 181031 343449 181073 343567
rect 181191 343449 181207 343567
rect 180897 325727 181207 343449
rect 180897 325609 180913 325727
rect 181031 325609 181073 325727
rect 181191 325609 181207 325727
rect 180897 325567 181207 325609
rect 180897 325449 180913 325567
rect 181031 325449 181073 325567
rect 181191 325449 181207 325567
rect 180897 307727 181207 325449
rect 180897 307609 180913 307727
rect 181031 307609 181073 307727
rect 181191 307609 181207 307727
rect 180897 307567 181207 307609
rect 180897 307449 180913 307567
rect 181031 307449 181073 307567
rect 181191 307449 181207 307567
rect 180897 289727 181207 307449
rect 180897 289609 180913 289727
rect 181031 289609 181073 289727
rect 181191 289609 181207 289727
rect 180897 289567 181207 289609
rect 180897 289449 180913 289567
rect 181031 289449 181073 289567
rect 181191 289449 181207 289567
rect 180897 271727 181207 289449
rect 180897 271609 180913 271727
rect 181031 271609 181073 271727
rect 181191 271609 181207 271727
rect 180897 271567 181207 271609
rect 180897 271449 180913 271567
rect 181031 271449 181073 271567
rect 181191 271449 181207 271567
rect 180897 253727 181207 271449
rect 180897 253609 180913 253727
rect 181031 253609 181073 253727
rect 181191 253609 181207 253727
rect 180897 253567 181207 253609
rect 180897 253449 180913 253567
rect 181031 253449 181073 253567
rect 181191 253449 181207 253567
rect 180897 235727 181207 253449
rect 180897 235609 180913 235727
rect 181031 235609 181073 235727
rect 181191 235609 181207 235727
rect 180897 235567 181207 235609
rect 180897 235449 180913 235567
rect 181031 235449 181073 235567
rect 181191 235449 181207 235567
rect 180897 217727 181207 235449
rect 180897 217609 180913 217727
rect 181031 217609 181073 217727
rect 181191 217609 181207 217727
rect 180897 217567 181207 217609
rect 180897 217449 180913 217567
rect 181031 217449 181073 217567
rect 181191 217449 181207 217567
rect 180897 199727 181207 217449
rect 180897 199609 180913 199727
rect 181031 199609 181073 199727
rect 181191 199609 181207 199727
rect 180897 199567 181207 199609
rect 180897 199449 180913 199567
rect 181031 199449 181073 199567
rect 181191 199449 181207 199567
rect 180897 181727 181207 199449
rect 180897 181609 180913 181727
rect 181031 181609 181073 181727
rect 181191 181609 181207 181727
rect 180897 181567 181207 181609
rect 180897 181449 180913 181567
rect 181031 181449 181073 181567
rect 181191 181449 181207 181567
rect 180897 163727 181207 181449
rect 180897 163609 180913 163727
rect 181031 163609 181073 163727
rect 181191 163609 181207 163727
rect 180897 163567 181207 163609
rect 180897 163449 180913 163567
rect 181031 163449 181073 163567
rect 181191 163449 181207 163567
rect 180897 145727 181207 163449
rect 180897 145609 180913 145727
rect 181031 145609 181073 145727
rect 181191 145609 181207 145727
rect 180897 145567 181207 145609
rect 180897 145449 180913 145567
rect 181031 145449 181073 145567
rect 181191 145449 181207 145567
rect 180897 127727 181207 145449
rect 180897 127609 180913 127727
rect 181031 127609 181073 127727
rect 181191 127609 181207 127727
rect 180897 127567 181207 127609
rect 180897 127449 180913 127567
rect 181031 127449 181073 127567
rect 181191 127449 181207 127567
rect 180897 109727 181207 127449
rect 180897 109609 180913 109727
rect 181031 109609 181073 109727
rect 181191 109609 181207 109727
rect 180897 109567 181207 109609
rect 180897 109449 180913 109567
rect 181031 109449 181073 109567
rect 181191 109449 181207 109567
rect 180897 91727 181207 109449
rect 180897 91609 180913 91727
rect 181031 91609 181073 91727
rect 181191 91609 181207 91727
rect 180897 91567 181207 91609
rect 180897 91449 180913 91567
rect 181031 91449 181073 91567
rect 181191 91449 181207 91567
rect 180897 73727 181207 91449
rect 180897 73609 180913 73727
rect 181031 73609 181073 73727
rect 181191 73609 181207 73727
rect 180897 73567 181207 73609
rect 180897 73449 180913 73567
rect 181031 73449 181073 73567
rect 181191 73449 181207 73567
rect 180897 55727 181207 73449
rect 180897 55609 180913 55727
rect 181031 55609 181073 55727
rect 181191 55609 181207 55727
rect 180897 55567 181207 55609
rect 180897 55449 180913 55567
rect 181031 55449 181073 55567
rect 181191 55449 181207 55567
rect 180897 37727 181207 55449
rect 180897 37609 180913 37727
rect 181031 37609 181073 37727
rect 181191 37609 181207 37727
rect 180897 37567 181207 37609
rect 180897 37449 180913 37567
rect 181031 37449 181073 37567
rect 181191 37449 181207 37567
rect 180897 19727 181207 37449
rect 180897 19609 180913 19727
rect 181031 19609 181073 19727
rect 181191 19609 181207 19727
rect 180897 19567 181207 19609
rect 180897 19449 180913 19567
rect 181031 19449 181073 19567
rect 181191 19449 181207 19567
rect 180897 1727 181207 19449
rect 180897 1609 180913 1727
rect 181031 1609 181073 1727
rect 181191 1609 181207 1727
rect 180897 1567 181207 1609
rect 180897 1449 180913 1567
rect 181031 1449 181073 1567
rect 181191 1449 181207 1567
rect 180897 -173 181207 1449
rect 180897 -291 180913 -173
rect 181031 -291 181073 -173
rect 181191 -291 181207 -173
rect 180897 -333 181207 -291
rect 180897 -451 180913 -333
rect 181031 -451 181073 -333
rect 181191 -451 181207 -333
rect 180897 -947 181207 -451
rect 182757 345587 183067 353101
rect 182757 345469 182773 345587
rect 182891 345469 182933 345587
rect 183051 345469 183067 345587
rect 182757 345427 183067 345469
rect 182757 345309 182773 345427
rect 182891 345309 182933 345427
rect 183051 345309 183067 345427
rect 182757 327587 183067 345309
rect 182757 327469 182773 327587
rect 182891 327469 182933 327587
rect 183051 327469 183067 327587
rect 182757 327427 183067 327469
rect 182757 327309 182773 327427
rect 182891 327309 182933 327427
rect 183051 327309 183067 327427
rect 182757 309587 183067 327309
rect 182757 309469 182773 309587
rect 182891 309469 182933 309587
rect 183051 309469 183067 309587
rect 182757 309427 183067 309469
rect 182757 309309 182773 309427
rect 182891 309309 182933 309427
rect 183051 309309 183067 309427
rect 182757 291587 183067 309309
rect 182757 291469 182773 291587
rect 182891 291469 182933 291587
rect 183051 291469 183067 291587
rect 182757 291427 183067 291469
rect 182757 291309 182773 291427
rect 182891 291309 182933 291427
rect 183051 291309 183067 291427
rect 182757 273587 183067 291309
rect 182757 273469 182773 273587
rect 182891 273469 182933 273587
rect 183051 273469 183067 273587
rect 182757 273427 183067 273469
rect 182757 273309 182773 273427
rect 182891 273309 182933 273427
rect 183051 273309 183067 273427
rect 182757 255587 183067 273309
rect 182757 255469 182773 255587
rect 182891 255469 182933 255587
rect 183051 255469 183067 255587
rect 182757 255427 183067 255469
rect 182757 255309 182773 255427
rect 182891 255309 182933 255427
rect 183051 255309 183067 255427
rect 182757 237587 183067 255309
rect 182757 237469 182773 237587
rect 182891 237469 182933 237587
rect 183051 237469 183067 237587
rect 182757 237427 183067 237469
rect 182757 237309 182773 237427
rect 182891 237309 182933 237427
rect 183051 237309 183067 237427
rect 182757 219587 183067 237309
rect 182757 219469 182773 219587
rect 182891 219469 182933 219587
rect 183051 219469 183067 219587
rect 182757 219427 183067 219469
rect 182757 219309 182773 219427
rect 182891 219309 182933 219427
rect 183051 219309 183067 219427
rect 182757 201587 183067 219309
rect 182757 201469 182773 201587
rect 182891 201469 182933 201587
rect 183051 201469 183067 201587
rect 182757 201427 183067 201469
rect 182757 201309 182773 201427
rect 182891 201309 182933 201427
rect 183051 201309 183067 201427
rect 182757 183587 183067 201309
rect 182757 183469 182773 183587
rect 182891 183469 182933 183587
rect 183051 183469 183067 183587
rect 182757 183427 183067 183469
rect 182757 183309 182773 183427
rect 182891 183309 182933 183427
rect 183051 183309 183067 183427
rect 182757 165587 183067 183309
rect 182757 165469 182773 165587
rect 182891 165469 182933 165587
rect 183051 165469 183067 165587
rect 182757 165427 183067 165469
rect 182757 165309 182773 165427
rect 182891 165309 182933 165427
rect 183051 165309 183067 165427
rect 182757 147587 183067 165309
rect 182757 147469 182773 147587
rect 182891 147469 182933 147587
rect 183051 147469 183067 147587
rect 182757 147427 183067 147469
rect 182757 147309 182773 147427
rect 182891 147309 182933 147427
rect 183051 147309 183067 147427
rect 182757 129587 183067 147309
rect 182757 129469 182773 129587
rect 182891 129469 182933 129587
rect 183051 129469 183067 129587
rect 182757 129427 183067 129469
rect 182757 129309 182773 129427
rect 182891 129309 182933 129427
rect 183051 129309 183067 129427
rect 182757 111587 183067 129309
rect 182757 111469 182773 111587
rect 182891 111469 182933 111587
rect 183051 111469 183067 111587
rect 182757 111427 183067 111469
rect 182757 111309 182773 111427
rect 182891 111309 182933 111427
rect 183051 111309 183067 111427
rect 182757 93587 183067 111309
rect 182757 93469 182773 93587
rect 182891 93469 182933 93587
rect 183051 93469 183067 93587
rect 182757 93427 183067 93469
rect 182757 93309 182773 93427
rect 182891 93309 182933 93427
rect 183051 93309 183067 93427
rect 182757 75587 183067 93309
rect 182757 75469 182773 75587
rect 182891 75469 182933 75587
rect 183051 75469 183067 75587
rect 182757 75427 183067 75469
rect 182757 75309 182773 75427
rect 182891 75309 182933 75427
rect 183051 75309 183067 75427
rect 182757 57587 183067 75309
rect 182757 57469 182773 57587
rect 182891 57469 182933 57587
rect 183051 57469 183067 57587
rect 182757 57427 183067 57469
rect 182757 57309 182773 57427
rect 182891 57309 182933 57427
rect 183051 57309 183067 57427
rect 182757 39587 183067 57309
rect 182757 39469 182773 39587
rect 182891 39469 182933 39587
rect 183051 39469 183067 39587
rect 182757 39427 183067 39469
rect 182757 39309 182773 39427
rect 182891 39309 182933 39427
rect 183051 39309 183067 39427
rect 182757 21587 183067 39309
rect 182757 21469 182773 21587
rect 182891 21469 182933 21587
rect 183051 21469 183067 21587
rect 182757 21427 183067 21469
rect 182757 21309 182773 21427
rect 182891 21309 182933 21427
rect 183051 21309 183067 21427
rect 182757 3587 183067 21309
rect 182757 3469 182773 3587
rect 182891 3469 182933 3587
rect 183051 3469 183067 3587
rect 182757 3427 183067 3469
rect 182757 3309 182773 3427
rect 182891 3309 182933 3427
rect 183051 3309 183067 3427
rect 182757 -1133 183067 3309
rect 182757 -1251 182773 -1133
rect 182891 -1251 182933 -1133
rect 183051 -1251 183067 -1133
rect 182757 -1293 183067 -1251
rect 182757 -1411 182773 -1293
rect 182891 -1411 182933 -1293
rect 183051 -1411 183067 -1293
rect 182757 -1907 183067 -1411
rect 184617 347447 184927 354061
rect 184617 347329 184633 347447
rect 184751 347329 184793 347447
rect 184911 347329 184927 347447
rect 184617 347287 184927 347329
rect 184617 347169 184633 347287
rect 184751 347169 184793 347287
rect 184911 347169 184927 347287
rect 184617 329447 184927 347169
rect 184617 329329 184633 329447
rect 184751 329329 184793 329447
rect 184911 329329 184927 329447
rect 184617 329287 184927 329329
rect 184617 329169 184633 329287
rect 184751 329169 184793 329287
rect 184911 329169 184927 329287
rect 184617 311447 184927 329169
rect 184617 311329 184633 311447
rect 184751 311329 184793 311447
rect 184911 311329 184927 311447
rect 184617 311287 184927 311329
rect 184617 311169 184633 311287
rect 184751 311169 184793 311287
rect 184911 311169 184927 311287
rect 184617 293447 184927 311169
rect 184617 293329 184633 293447
rect 184751 293329 184793 293447
rect 184911 293329 184927 293447
rect 184617 293287 184927 293329
rect 184617 293169 184633 293287
rect 184751 293169 184793 293287
rect 184911 293169 184927 293287
rect 184617 275447 184927 293169
rect 184617 275329 184633 275447
rect 184751 275329 184793 275447
rect 184911 275329 184927 275447
rect 184617 275287 184927 275329
rect 184617 275169 184633 275287
rect 184751 275169 184793 275287
rect 184911 275169 184927 275287
rect 184617 257447 184927 275169
rect 184617 257329 184633 257447
rect 184751 257329 184793 257447
rect 184911 257329 184927 257447
rect 184617 257287 184927 257329
rect 184617 257169 184633 257287
rect 184751 257169 184793 257287
rect 184911 257169 184927 257287
rect 184617 239447 184927 257169
rect 184617 239329 184633 239447
rect 184751 239329 184793 239447
rect 184911 239329 184927 239447
rect 184617 239287 184927 239329
rect 184617 239169 184633 239287
rect 184751 239169 184793 239287
rect 184911 239169 184927 239287
rect 184617 221447 184927 239169
rect 184617 221329 184633 221447
rect 184751 221329 184793 221447
rect 184911 221329 184927 221447
rect 184617 221287 184927 221329
rect 184617 221169 184633 221287
rect 184751 221169 184793 221287
rect 184911 221169 184927 221287
rect 184617 203447 184927 221169
rect 184617 203329 184633 203447
rect 184751 203329 184793 203447
rect 184911 203329 184927 203447
rect 184617 203287 184927 203329
rect 184617 203169 184633 203287
rect 184751 203169 184793 203287
rect 184911 203169 184927 203287
rect 184617 185447 184927 203169
rect 184617 185329 184633 185447
rect 184751 185329 184793 185447
rect 184911 185329 184927 185447
rect 184617 185287 184927 185329
rect 184617 185169 184633 185287
rect 184751 185169 184793 185287
rect 184911 185169 184927 185287
rect 184617 167447 184927 185169
rect 184617 167329 184633 167447
rect 184751 167329 184793 167447
rect 184911 167329 184927 167447
rect 184617 167287 184927 167329
rect 184617 167169 184633 167287
rect 184751 167169 184793 167287
rect 184911 167169 184927 167287
rect 184617 149447 184927 167169
rect 184617 149329 184633 149447
rect 184751 149329 184793 149447
rect 184911 149329 184927 149447
rect 184617 149287 184927 149329
rect 184617 149169 184633 149287
rect 184751 149169 184793 149287
rect 184911 149169 184927 149287
rect 184617 131447 184927 149169
rect 184617 131329 184633 131447
rect 184751 131329 184793 131447
rect 184911 131329 184927 131447
rect 184617 131287 184927 131329
rect 184617 131169 184633 131287
rect 184751 131169 184793 131287
rect 184911 131169 184927 131287
rect 184617 113447 184927 131169
rect 184617 113329 184633 113447
rect 184751 113329 184793 113447
rect 184911 113329 184927 113447
rect 184617 113287 184927 113329
rect 184617 113169 184633 113287
rect 184751 113169 184793 113287
rect 184911 113169 184927 113287
rect 184617 95447 184927 113169
rect 184617 95329 184633 95447
rect 184751 95329 184793 95447
rect 184911 95329 184927 95447
rect 184617 95287 184927 95329
rect 184617 95169 184633 95287
rect 184751 95169 184793 95287
rect 184911 95169 184927 95287
rect 184617 77447 184927 95169
rect 184617 77329 184633 77447
rect 184751 77329 184793 77447
rect 184911 77329 184927 77447
rect 184617 77287 184927 77329
rect 184617 77169 184633 77287
rect 184751 77169 184793 77287
rect 184911 77169 184927 77287
rect 184617 59447 184927 77169
rect 184617 59329 184633 59447
rect 184751 59329 184793 59447
rect 184911 59329 184927 59447
rect 184617 59287 184927 59329
rect 184617 59169 184633 59287
rect 184751 59169 184793 59287
rect 184911 59169 184927 59287
rect 184617 41447 184927 59169
rect 184617 41329 184633 41447
rect 184751 41329 184793 41447
rect 184911 41329 184927 41447
rect 184617 41287 184927 41329
rect 184617 41169 184633 41287
rect 184751 41169 184793 41287
rect 184911 41169 184927 41287
rect 184617 23447 184927 41169
rect 184617 23329 184633 23447
rect 184751 23329 184793 23447
rect 184911 23329 184927 23447
rect 184617 23287 184927 23329
rect 184617 23169 184633 23287
rect 184751 23169 184793 23287
rect 184911 23169 184927 23287
rect 184617 5447 184927 23169
rect 184617 5329 184633 5447
rect 184751 5329 184793 5447
rect 184911 5329 184927 5447
rect 184617 5287 184927 5329
rect 184617 5169 184633 5287
rect 184751 5169 184793 5287
rect 184911 5169 184927 5287
rect 184617 -2093 184927 5169
rect 184617 -2211 184633 -2093
rect 184751 -2211 184793 -2093
rect 184911 -2211 184927 -2093
rect 184617 -2253 184927 -2211
rect 184617 -2371 184633 -2253
rect 184751 -2371 184793 -2253
rect 184911 -2371 184927 -2253
rect 184617 -2867 184927 -2371
rect 186477 349307 186787 355021
rect 195477 355779 195787 355795
rect 195477 355661 195493 355779
rect 195611 355661 195653 355779
rect 195771 355661 195787 355779
rect 195477 355619 195787 355661
rect 195477 355501 195493 355619
rect 195611 355501 195653 355619
rect 195771 355501 195787 355619
rect 193617 354819 193927 354835
rect 193617 354701 193633 354819
rect 193751 354701 193793 354819
rect 193911 354701 193927 354819
rect 193617 354659 193927 354701
rect 193617 354541 193633 354659
rect 193751 354541 193793 354659
rect 193911 354541 193927 354659
rect 191757 353859 192067 353875
rect 191757 353741 191773 353859
rect 191891 353741 191933 353859
rect 192051 353741 192067 353859
rect 191757 353699 192067 353741
rect 191757 353581 191773 353699
rect 191891 353581 191933 353699
rect 192051 353581 192067 353699
rect 186477 349189 186493 349307
rect 186611 349189 186653 349307
rect 186771 349189 186787 349307
rect 186477 349147 186787 349189
rect 186477 349029 186493 349147
rect 186611 349029 186653 349147
rect 186771 349029 186787 349147
rect 186477 331307 186787 349029
rect 186477 331189 186493 331307
rect 186611 331189 186653 331307
rect 186771 331189 186787 331307
rect 186477 331147 186787 331189
rect 186477 331029 186493 331147
rect 186611 331029 186653 331147
rect 186771 331029 186787 331147
rect 186477 313307 186787 331029
rect 186477 313189 186493 313307
rect 186611 313189 186653 313307
rect 186771 313189 186787 313307
rect 186477 313147 186787 313189
rect 186477 313029 186493 313147
rect 186611 313029 186653 313147
rect 186771 313029 186787 313147
rect 186477 295307 186787 313029
rect 186477 295189 186493 295307
rect 186611 295189 186653 295307
rect 186771 295189 186787 295307
rect 186477 295147 186787 295189
rect 186477 295029 186493 295147
rect 186611 295029 186653 295147
rect 186771 295029 186787 295147
rect 186477 277307 186787 295029
rect 186477 277189 186493 277307
rect 186611 277189 186653 277307
rect 186771 277189 186787 277307
rect 186477 277147 186787 277189
rect 186477 277029 186493 277147
rect 186611 277029 186653 277147
rect 186771 277029 186787 277147
rect 186477 259307 186787 277029
rect 186477 259189 186493 259307
rect 186611 259189 186653 259307
rect 186771 259189 186787 259307
rect 186477 259147 186787 259189
rect 186477 259029 186493 259147
rect 186611 259029 186653 259147
rect 186771 259029 186787 259147
rect 186477 241307 186787 259029
rect 186477 241189 186493 241307
rect 186611 241189 186653 241307
rect 186771 241189 186787 241307
rect 186477 241147 186787 241189
rect 186477 241029 186493 241147
rect 186611 241029 186653 241147
rect 186771 241029 186787 241147
rect 186477 223307 186787 241029
rect 186477 223189 186493 223307
rect 186611 223189 186653 223307
rect 186771 223189 186787 223307
rect 186477 223147 186787 223189
rect 186477 223029 186493 223147
rect 186611 223029 186653 223147
rect 186771 223029 186787 223147
rect 186477 205307 186787 223029
rect 186477 205189 186493 205307
rect 186611 205189 186653 205307
rect 186771 205189 186787 205307
rect 186477 205147 186787 205189
rect 186477 205029 186493 205147
rect 186611 205029 186653 205147
rect 186771 205029 186787 205147
rect 186477 187307 186787 205029
rect 186477 187189 186493 187307
rect 186611 187189 186653 187307
rect 186771 187189 186787 187307
rect 186477 187147 186787 187189
rect 186477 187029 186493 187147
rect 186611 187029 186653 187147
rect 186771 187029 186787 187147
rect 186477 169307 186787 187029
rect 186477 169189 186493 169307
rect 186611 169189 186653 169307
rect 186771 169189 186787 169307
rect 186477 169147 186787 169189
rect 186477 169029 186493 169147
rect 186611 169029 186653 169147
rect 186771 169029 186787 169147
rect 186477 151307 186787 169029
rect 186477 151189 186493 151307
rect 186611 151189 186653 151307
rect 186771 151189 186787 151307
rect 186477 151147 186787 151189
rect 186477 151029 186493 151147
rect 186611 151029 186653 151147
rect 186771 151029 186787 151147
rect 186477 133307 186787 151029
rect 186477 133189 186493 133307
rect 186611 133189 186653 133307
rect 186771 133189 186787 133307
rect 186477 133147 186787 133189
rect 186477 133029 186493 133147
rect 186611 133029 186653 133147
rect 186771 133029 186787 133147
rect 186477 115307 186787 133029
rect 186477 115189 186493 115307
rect 186611 115189 186653 115307
rect 186771 115189 186787 115307
rect 186477 115147 186787 115189
rect 186477 115029 186493 115147
rect 186611 115029 186653 115147
rect 186771 115029 186787 115147
rect 186477 97307 186787 115029
rect 186477 97189 186493 97307
rect 186611 97189 186653 97307
rect 186771 97189 186787 97307
rect 186477 97147 186787 97189
rect 186477 97029 186493 97147
rect 186611 97029 186653 97147
rect 186771 97029 186787 97147
rect 186477 79307 186787 97029
rect 186477 79189 186493 79307
rect 186611 79189 186653 79307
rect 186771 79189 186787 79307
rect 186477 79147 186787 79189
rect 186477 79029 186493 79147
rect 186611 79029 186653 79147
rect 186771 79029 186787 79147
rect 186477 61307 186787 79029
rect 186477 61189 186493 61307
rect 186611 61189 186653 61307
rect 186771 61189 186787 61307
rect 186477 61147 186787 61189
rect 186477 61029 186493 61147
rect 186611 61029 186653 61147
rect 186771 61029 186787 61147
rect 186477 43307 186787 61029
rect 186477 43189 186493 43307
rect 186611 43189 186653 43307
rect 186771 43189 186787 43307
rect 186477 43147 186787 43189
rect 186477 43029 186493 43147
rect 186611 43029 186653 43147
rect 186771 43029 186787 43147
rect 186477 25307 186787 43029
rect 186477 25189 186493 25307
rect 186611 25189 186653 25307
rect 186771 25189 186787 25307
rect 186477 25147 186787 25189
rect 186477 25029 186493 25147
rect 186611 25029 186653 25147
rect 186771 25029 186787 25147
rect 186477 7307 186787 25029
rect 186477 7189 186493 7307
rect 186611 7189 186653 7307
rect 186771 7189 186787 7307
rect 186477 7147 186787 7189
rect 186477 7029 186493 7147
rect 186611 7029 186653 7147
rect 186771 7029 186787 7147
rect 177477 -3651 177493 -3533
rect 177611 -3651 177653 -3533
rect 177771 -3651 177787 -3533
rect 177477 -3693 177787 -3651
rect 177477 -3811 177493 -3693
rect 177611 -3811 177653 -3693
rect 177771 -3811 177787 -3693
rect 177477 -3827 177787 -3811
rect 186477 -3053 186787 7029
rect 189897 352899 190207 352915
rect 189897 352781 189913 352899
rect 190031 352781 190073 352899
rect 190191 352781 190207 352899
rect 189897 352739 190207 352781
rect 189897 352621 189913 352739
rect 190031 352621 190073 352739
rect 190191 352621 190207 352739
rect 189897 334727 190207 352621
rect 189897 334609 189913 334727
rect 190031 334609 190073 334727
rect 190191 334609 190207 334727
rect 189897 334567 190207 334609
rect 189897 334449 189913 334567
rect 190031 334449 190073 334567
rect 190191 334449 190207 334567
rect 189897 316727 190207 334449
rect 189897 316609 189913 316727
rect 190031 316609 190073 316727
rect 190191 316609 190207 316727
rect 189897 316567 190207 316609
rect 189897 316449 189913 316567
rect 190031 316449 190073 316567
rect 190191 316449 190207 316567
rect 189897 298727 190207 316449
rect 189897 298609 189913 298727
rect 190031 298609 190073 298727
rect 190191 298609 190207 298727
rect 189897 298567 190207 298609
rect 189897 298449 189913 298567
rect 190031 298449 190073 298567
rect 190191 298449 190207 298567
rect 189897 280727 190207 298449
rect 189897 280609 189913 280727
rect 190031 280609 190073 280727
rect 190191 280609 190207 280727
rect 189897 280567 190207 280609
rect 189897 280449 189913 280567
rect 190031 280449 190073 280567
rect 190191 280449 190207 280567
rect 189897 262727 190207 280449
rect 189897 262609 189913 262727
rect 190031 262609 190073 262727
rect 190191 262609 190207 262727
rect 189897 262567 190207 262609
rect 189897 262449 189913 262567
rect 190031 262449 190073 262567
rect 190191 262449 190207 262567
rect 189897 244727 190207 262449
rect 189897 244609 189913 244727
rect 190031 244609 190073 244727
rect 190191 244609 190207 244727
rect 189897 244567 190207 244609
rect 189897 244449 189913 244567
rect 190031 244449 190073 244567
rect 190191 244449 190207 244567
rect 189897 226727 190207 244449
rect 189897 226609 189913 226727
rect 190031 226609 190073 226727
rect 190191 226609 190207 226727
rect 189897 226567 190207 226609
rect 189897 226449 189913 226567
rect 190031 226449 190073 226567
rect 190191 226449 190207 226567
rect 189897 208727 190207 226449
rect 189897 208609 189913 208727
rect 190031 208609 190073 208727
rect 190191 208609 190207 208727
rect 189897 208567 190207 208609
rect 189897 208449 189913 208567
rect 190031 208449 190073 208567
rect 190191 208449 190207 208567
rect 189897 190727 190207 208449
rect 189897 190609 189913 190727
rect 190031 190609 190073 190727
rect 190191 190609 190207 190727
rect 189897 190567 190207 190609
rect 189897 190449 189913 190567
rect 190031 190449 190073 190567
rect 190191 190449 190207 190567
rect 189897 172727 190207 190449
rect 189897 172609 189913 172727
rect 190031 172609 190073 172727
rect 190191 172609 190207 172727
rect 189897 172567 190207 172609
rect 189897 172449 189913 172567
rect 190031 172449 190073 172567
rect 190191 172449 190207 172567
rect 189897 154727 190207 172449
rect 189897 154609 189913 154727
rect 190031 154609 190073 154727
rect 190191 154609 190207 154727
rect 189897 154567 190207 154609
rect 189897 154449 189913 154567
rect 190031 154449 190073 154567
rect 190191 154449 190207 154567
rect 189897 136727 190207 154449
rect 189897 136609 189913 136727
rect 190031 136609 190073 136727
rect 190191 136609 190207 136727
rect 189897 136567 190207 136609
rect 189897 136449 189913 136567
rect 190031 136449 190073 136567
rect 190191 136449 190207 136567
rect 189897 118727 190207 136449
rect 189897 118609 189913 118727
rect 190031 118609 190073 118727
rect 190191 118609 190207 118727
rect 189897 118567 190207 118609
rect 189897 118449 189913 118567
rect 190031 118449 190073 118567
rect 190191 118449 190207 118567
rect 189897 100727 190207 118449
rect 189897 100609 189913 100727
rect 190031 100609 190073 100727
rect 190191 100609 190207 100727
rect 189897 100567 190207 100609
rect 189897 100449 189913 100567
rect 190031 100449 190073 100567
rect 190191 100449 190207 100567
rect 189897 82727 190207 100449
rect 189897 82609 189913 82727
rect 190031 82609 190073 82727
rect 190191 82609 190207 82727
rect 189897 82567 190207 82609
rect 189897 82449 189913 82567
rect 190031 82449 190073 82567
rect 190191 82449 190207 82567
rect 189897 64727 190207 82449
rect 189897 64609 189913 64727
rect 190031 64609 190073 64727
rect 190191 64609 190207 64727
rect 189897 64567 190207 64609
rect 189897 64449 189913 64567
rect 190031 64449 190073 64567
rect 190191 64449 190207 64567
rect 189897 46727 190207 64449
rect 189897 46609 189913 46727
rect 190031 46609 190073 46727
rect 190191 46609 190207 46727
rect 189897 46567 190207 46609
rect 189897 46449 189913 46567
rect 190031 46449 190073 46567
rect 190191 46449 190207 46567
rect 189897 28727 190207 46449
rect 189897 28609 189913 28727
rect 190031 28609 190073 28727
rect 190191 28609 190207 28727
rect 189897 28567 190207 28609
rect 189897 28449 189913 28567
rect 190031 28449 190073 28567
rect 190191 28449 190207 28567
rect 189897 10727 190207 28449
rect 189897 10609 189913 10727
rect 190031 10609 190073 10727
rect 190191 10609 190207 10727
rect 189897 10567 190207 10609
rect 189897 10449 189913 10567
rect 190031 10449 190073 10567
rect 190191 10449 190207 10567
rect 189897 -653 190207 10449
rect 189897 -771 189913 -653
rect 190031 -771 190073 -653
rect 190191 -771 190207 -653
rect 189897 -813 190207 -771
rect 189897 -931 189913 -813
rect 190031 -931 190073 -813
rect 190191 -931 190207 -813
rect 189897 -947 190207 -931
rect 191757 336587 192067 353581
rect 191757 336469 191773 336587
rect 191891 336469 191933 336587
rect 192051 336469 192067 336587
rect 191757 336427 192067 336469
rect 191757 336309 191773 336427
rect 191891 336309 191933 336427
rect 192051 336309 192067 336427
rect 191757 318587 192067 336309
rect 191757 318469 191773 318587
rect 191891 318469 191933 318587
rect 192051 318469 192067 318587
rect 191757 318427 192067 318469
rect 191757 318309 191773 318427
rect 191891 318309 191933 318427
rect 192051 318309 192067 318427
rect 191757 300587 192067 318309
rect 191757 300469 191773 300587
rect 191891 300469 191933 300587
rect 192051 300469 192067 300587
rect 191757 300427 192067 300469
rect 191757 300309 191773 300427
rect 191891 300309 191933 300427
rect 192051 300309 192067 300427
rect 191757 282587 192067 300309
rect 191757 282469 191773 282587
rect 191891 282469 191933 282587
rect 192051 282469 192067 282587
rect 191757 282427 192067 282469
rect 191757 282309 191773 282427
rect 191891 282309 191933 282427
rect 192051 282309 192067 282427
rect 191757 264587 192067 282309
rect 191757 264469 191773 264587
rect 191891 264469 191933 264587
rect 192051 264469 192067 264587
rect 191757 264427 192067 264469
rect 191757 264309 191773 264427
rect 191891 264309 191933 264427
rect 192051 264309 192067 264427
rect 191757 246587 192067 264309
rect 191757 246469 191773 246587
rect 191891 246469 191933 246587
rect 192051 246469 192067 246587
rect 191757 246427 192067 246469
rect 191757 246309 191773 246427
rect 191891 246309 191933 246427
rect 192051 246309 192067 246427
rect 191757 228587 192067 246309
rect 191757 228469 191773 228587
rect 191891 228469 191933 228587
rect 192051 228469 192067 228587
rect 191757 228427 192067 228469
rect 191757 228309 191773 228427
rect 191891 228309 191933 228427
rect 192051 228309 192067 228427
rect 191757 210587 192067 228309
rect 191757 210469 191773 210587
rect 191891 210469 191933 210587
rect 192051 210469 192067 210587
rect 191757 210427 192067 210469
rect 191757 210309 191773 210427
rect 191891 210309 191933 210427
rect 192051 210309 192067 210427
rect 191757 192587 192067 210309
rect 191757 192469 191773 192587
rect 191891 192469 191933 192587
rect 192051 192469 192067 192587
rect 191757 192427 192067 192469
rect 191757 192309 191773 192427
rect 191891 192309 191933 192427
rect 192051 192309 192067 192427
rect 191757 174587 192067 192309
rect 191757 174469 191773 174587
rect 191891 174469 191933 174587
rect 192051 174469 192067 174587
rect 191757 174427 192067 174469
rect 191757 174309 191773 174427
rect 191891 174309 191933 174427
rect 192051 174309 192067 174427
rect 191757 156587 192067 174309
rect 191757 156469 191773 156587
rect 191891 156469 191933 156587
rect 192051 156469 192067 156587
rect 191757 156427 192067 156469
rect 191757 156309 191773 156427
rect 191891 156309 191933 156427
rect 192051 156309 192067 156427
rect 191757 138587 192067 156309
rect 191757 138469 191773 138587
rect 191891 138469 191933 138587
rect 192051 138469 192067 138587
rect 191757 138427 192067 138469
rect 191757 138309 191773 138427
rect 191891 138309 191933 138427
rect 192051 138309 192067 138427
rect 191757 120587 192067 138309
rect 191757 120469 191773 120587
rect 191891 120469 191933 120587
rect 192051 120469 192067 120587
rect 191757 120427 192067 120469
rect 191757 120309 191773 120427
rect 191891 120309 191933 120427
rect 192051 120309 192067 120427
rect 191757 102587 192067 120309
rect 191757 102469 191773 102587
rect 191891 102469 191933 102587
rect 192051 102469 192067 102587
rect 191757 102427 192067 102469
rect 191757 102309 191773 102427
rect 191891 102309 191933 102427
rect 192051 102309 192067 102427
rect 191757 84587 192067 102309
rect 191757 84469 191773 84587
rect 191891 84469 191933 84587
rect 192051 84469 192067 84587
rect 191757 84427 192067 84469
rect 191757 84309 191773 84427
rect 191891 84309 191933 84427
rect 192051 84309 192067 84427
rect 191757 66587 192067 84309
rect 191757 66469 191773 66587
rect 191891 66469 191933 66587
rect 192051 66469 192067 66587
rect 191757 66427 192067 66469
rect 191757 66309 191773 66427
rect 191891 66309 191933 66427
rect 192051 66309 192067 66427
rect 191757 48587 192067 66309
rect 191757 48469 191773 48587
rect 191891 48469 191933 48587
rect 192051 48469 192067 48587
rect 191757 48427 192067 48469
rect 191757 48309 191773 48427
rect 191891 48309 191933 48427
rect 192051 48309 192067 48427
rect 191757 30587 192067 48309
rect 191757 30469 191773 30587
rect 191891 30469 191933 30587
rect 192051 30469 192067 30587
rect 191757 30427 192067 30469
rect 191757 30309 191773 30427
rect 191891 30309 191933 30427
rect 192051 30309 192067 30427
rect 191757 12587 192067 30309
rect 191757 12469 191773 12587
rect 191891 12469 191933 12587
rect 192051 12469 192067 12587
rect 191757 12427 192067 12469
rect 191757 12309 191773 12427
rect 191891 12309 191933 12427
rect 192051 12309 192067 12427
rect 191757 -1613 192067 12309
rect 191757 -1731 191773 -1613
rect 191891 -1731 191933 -1613
rect 192051 -1731 192067 -1613
rect 191757 -1773 192067 -1731
rect 191757 -1891 191773 -1773
rect 191891 -1891 191933 -1773
rect 192051 -1891 192067 -1773
rect 191757 -1907 192067 -1891
rect 193617 338447 193927 354541
rect 193617 338329 193633 338447
rect 193751 338329 193793 338447
rect 193911 338329 193927 338447
rect 193617 338287 193927 338329
rect 193617 338169 193633 338287
rect 193751 338169 193793 338287
rect 193911 338169 193927 338287
rect 193617 320447 193927 338169
rect 193617 320329 193633 320447
rect 193751 320329 193793 320447
rect 193911 320329 193927 320447
rect 193617 320287 193927 320329
rect 193617 320169 193633 320287
rect 193751 320169 193793 320287
rect 193911 320169 193927 320287
rect 193617 302447 193927 320169
rect 193617 302329 193633 302447
rect 193751 302329 193793 302447
rect 193911 302329 193927 302447
rect 193617 302287 193927 302329
rect 193617 302169 193633 302287
rect 193751 302169 193793 302287
rect 193911 302169 193927 302287
rect 193617 284447 193927 302169
rect 193617 284329 193633 284447
rect 193751 284329 193793 284447
rect 193911 284329 193927 284447
rect 193617 284287 193927 284329
rect 193617 284169 193633 284287
rect 193751 284169 193793 284287
rect 193911 284169 193927 284287
rect 193617 266447 193927 284169
rect 193617 266329 193633 266447
rect 193751 266329 193793 266447
rect 193911 266329 193927 266447
rect 193617 266287 193927 266329
rect 193617 266169 193633 266287
rect 193751 266169 193793 266287
rect 193911 266169 193927 266287
rect 193617 248447 193927 266169
rect 193617 248329 193633 248447
rect 193751 248329 193793 248447
rect 193911 248329 193927 248447
rect 193617 248287 193927 248329
rect 193617 248169 193633 248287
rect 193751 248169 193793 248287
rect 193911 248169 193927 248287
rect 193617 230447 193927 248169
rect 193617 230329 193633 230447
rect 193751 230329 193793 230447
rect 193911 230329 193927 230447
rect 193617 230287 193927 230329
rect 193617 230169 193633 230287
rect 193751 230169 193793 230287
rect 193911 230169 193927 230287
rect 193617 212447 193927 230169
rect 193617 212329 193633 212447
rect 193751 212329 193793 212447
rect 193911 212329 193927 212447
rect 193617 212287 193927 212329
rect 193617 212169 193633 212287
rect 193751 212169 193793 212287
rect 193911 212169 193927 212287
rect 193617 194447 193927 212169
rect 193617 194329 193633 194447
rect 193751 194329 193793 194447
rect 193911 194329 193927 194447
rect 193617 194287 193927 194329
rect 193617 194169 193633 194287
rect 193751 194169 193793 194287
rect 193911 194169 193927 194287
rect 193617 176447 193927 194169
rect 193617 176329 193633 176447
rect 193751 176329 193793 176447
rect 193911 176329 193927 176447
rect 193617 176287 193927 176329
rect 193617 176169 193633 176287
rect 193751 176169 193793 176287
rect 193911 176169 193927 176287
rect 193617 158447 193927 176169
rect 193617 158329 193633 158447
rect 193751 158329 193793 158447
rect 193911 158329 193927 158447
rect 193617 158287 193927 158329
rect 193617 158169 193633 158287
rect 193751 158169 193793 158287
rect 193911 158169 193927 158287
rect 193617 140447 193927 158169
rect 193617 140329 193633 140447
rect 193751 140329 193793 140447
rect 193911 140329 193927 140447
rect 193617 140287 193927 140329
rect 193617 140169 193633 140287
rect 193751 140169 193793 140287
rect 193911 140169 193927 140287
rect 193617 122447 193927 140169
rect 193617 122329 193633 122447
rect 193751 122329 193793 122447
rect 193911 122329 193927 122447
rect 193617 122287 193927 122329
rect 193617 122169 193633 122287
rect 193751 122169 193793 122287
rect 193911 122169 193927 122287
rect 193617 104447 193927 122169
rect 193617 104329 193633 104447
rect 193751 104329 193793 104447
rect 193911 104329 193927 104447
rect 193617 104287 193927 104329
rect 193617 104169 193633 104287
rect 193751 104169 193793 104287
rect 193911 104169 193927 104287
rect 193617 86447 193927 104169
rect 193617 86329 193633 86447
rect 193751 86329 193793 86447
rect 193911 86329 193927 86447
rect 193617 86287 193927 86329
rect 193617 86169 193633 86287
rect 193751 86169 193793 86287
rect 193911 86169 193927 86287
rect 193617 68447 193927 86169
rect 193617 68329 193633 68447
rect 193751 68329 193793 68447
rect 193911 68329 193927 68447
rect 193617 68287 193927 68329
rect 193617 68169 193633 68287
rect 193751 68169 193793 68287
rect 193911 68169 193927 68287
rect 193617 50447 193927 68169
rect 193617 50329 193633 50447
rect 193751 50329 193793 50447
rect 193911 50329 193927 50447
rect 193617 50287 193927 50329
rect 193617 50169 193633 50287
rect 193751 50169 193793 50287
rect 193911 50169 193927 50287
rect 193617 32447 193927 50169
rect 193617 32329 193633 32447
rect 193751 32329 193793 32447
rect 193911 32329 193927 32447
rect 193617 32287 193927 32329
rect 193617 32169 193633 32287
rect 193751 32169 193793 32287
rect 193911 32169 193927 32287
rect 193617 14447 193927 32169
rect 193617 14329 193633 14447
rect 193751 14329 193793 14447
rect 193911 14329 193927 14447
rect 193617 14287 193927 14329
rect 193617 14169 193633 14287
rect 193751 14169 193793 14287
rect 193911 14169 193927 14287
rect 193617 -2573 193927 14169
rect 193617 -2691 193633 -2573
rect 193751 -2691 193793 -2573
rect 193911 -2691 193927 -2573
rect 193617 -2733 193927 -2691
rect 193617 -2851 193633 -2733
rect 193751 -2851 193793 -2733
rect 193911 -2851 193927 -2733
rect 193617 -2867 193927 -2851
rect 195477 340307 195787 355501
rect 204477 355299 204787 355795
rect 204477 355181 204493 355299
rect 204611 355181 204653 355299
rect 204771 355181 204787 355299
rect 204477 355139 204787 355181
rect 204477 355021 204493 355139
rect 204611 355021 204653 355139
rect 204771 355021 204787 355139
rect 202617 354339 202927 354835
rect 202617 354221 202633 354339
rect 202751 354221 202793 354339
rect 202911 354221 202927 354339
rect 202617 354179 202927 354221
rect 202617 354061 202633 354179
rect 202751 354061 202793 354179
rect 202911 354061 202927 354179
rect 200757 353379 201067 353875
rect 200757 353261 200773 353379
rect 200891 353261 200933 353379
rect 201051 353261 201067 353379
rect 200757 353219 201067 353261
rect 200757 353101 200773 353219
rect 200891 353101 200933 353219
rect 201051 353101 201067 353219
rect 195477 340189 195493 340307
rect 195611 340189 195653 340307
rect 195771 340189 195787 340307
rect 195477 340147 195787 340189
rect 195477 340029 195493 340147
rect 195611 340029 195653 340147
rect 195771 340029 195787 340147
rect 195477 322307 195787 340029
rect 195477 322189 195493 322307
rect 195611 322189 195653 322307
rect 195771 322189 195787 322307
rect 195477 322147 195787 322189
rect 195477 322029 195493 322147
rect 195611 322029 195653 322147
rect 195771 322029 195787 322147
rect 195477 304307 195787 322029
rect 195477 304189 195493 304307
rect 195611 304189 195653 304307
rect 195771 304189 195787 304307
rect 195477 304147 195787 304189
rect 195477 304029 195493 304147
rect 195611 304029 195653 304147
rect 195771 304029 195787 304147
rect 195477 286307 195787 304029
rect 195477 286189 195493 286307
rect 195611 286189 195653 286307
rect 195771 286189 195787 286307
rect 195477 286147 195787 286189
rect 195477 286029 195493 286147
rect 195611 286029 195653 286147
rect 195771 286029 195787 286147
rect 195477 268307 195787 286029
rect 195477 268189 195493 268307
rect 195611 268189 195653 268307
rect 195771 268189 195787 268307
rect 195477 268147 195787 268189
rect 195477 268029 195493 268147
rect 195611 268029 195653 268147
rect 195771 268029 195787 268147
rect 195477 250307 195787 268029
rect 195477 250189 195493 250307
rect 195611 250189 195653 250307
rect 195771 250189 195787 250307
rect 195477 250147 195787 250189
rect 195477 250029 195493 250147
rect 195611 250029 195653 250147
rect 195771 250029 195787 250147
rect 195477 232307 195787 250029
rect 195477 232189 195493 232307
rect 195611 232189 195653 232307
rect 195771 232189 195787 232307
rect 195477 232147 195787 232189
rect 195477 232029 195493 232147
rect 195611 232029 195653 232147
rect 195771 232029 195787 232147
rect 195477 214307 195787 232029
rect 195477 214189 195493 214307
rect 195611 214189 195653 214307
rect 195771 214189 195787 214307
rect 195477 214147 195787 214189
rect 195477 214029 195493 214147
rect 195611 214029 195653 214147
rect 195771 214029 195787 214147
rect 195477 196307 195787 214029
rect 195477 196189 195493 196307
rect 195611 196189 195653 196307
rect 195771 196189 195787 196307
rect 195477 196147 195787 196189
rect 195477 196029 195493 196147
rect 195611 196029 195653 196147
rect 195771 196029 195787 196147
rect 195477 178307 195787 196029
rect 195477 178189 195493 178307
rect 195611 178189 195653 178307
rect 195771 178189 195787 178307
rect 195477 178147 195787 178189
rect 195477 178029 195493 178147
rect 195611 178029 195653 178147
rect 195771 178029 195787 178147
rect 195477 160307 195787 178029
rect 195477 160189 195493 160307
rect 195611 160189 195653 160307
rect 195771 160189 195787 160307
rect 195477 160147 195787 160189
rect 195477 160029 195493 160147
rect 195611 160029 195653 160147
rect 195771 160029 195787 160147
rect 195477 142307 195787 160029
rect 195477 142189 195493 142307
rect 195611 142189 195653 142307
rect 195771 142189 195787 142307
rect 195477 142147 195787 142189
rect 195477 142029 195493 142147
rect 195611 142029 195653 142147
rect 195771 142029 195787 142147
rect 195477 124307 195787 142029
rect 195477 124189 195493 124307
rect 195611 124189 195653 124307
rect 195771 124189 195787 124307
rect 195477 124147 195787 124189
rect 195477 124029 195493 124147
rect 195611 124029 195653 124147
rect 195771 124029 195787 124147
rect 195477 106307 195787 124029
rect 195477 106189 195493 106307
rect 195611 106189 195653 106307
rect 195771 106189 195787 106307
rect 195477 106147 195787 106189
rect 195477 106029 195493 106147
rect 195611 106029 195653 106147
rect 195771 106029 195787 106147
rect 195477 88307 195787 106029
rect 195477 88189 195493 88307
rect 195611 88189 195653 88307
rect 195771 88189 195787 88307
rect 195477 88147 195787 88189
rect 195477 88029 195493 88147
rect 195611 88029 195653 88147
rect 195771 88029 195787 88147
rect 195477 70307 195787 88029
rect 195477 70189 195493 70307
rect 195611 70189 195653 70307
rect 195771 70189 195787 70307
rect 195477 70147 195787 70189
rect 195477 70029 195493 70147
rect 195611 70029 195653 70147
rect 195771 70029 195787 70147
rect 195477 52307 195787 70029
rect 195477 52189 195493 52307
rect 195611 52189 195653 52307
rect 195771 52189 195787 52307
rect 195477 52147 195787 52189
rect 195477 52029 195493 52147
rect 195611 52029 195653 52147
rect 195771 52029 195787 52147
rect 195477 34307 195787 52029
rect 195477 34189 195493 34307
rect 195611 34189 195653 34307
rect 195771 34189 195787 34307
rect 195477 34147 195787 34189
rect 195477 34029 195493 34147
rect 195611 34029 195653 34147
rect 195771 34029 195787 34147
rect 195477 16307 195787 34029
rect 195477 16189 195493 16307
rect 195611 16189 195653 16307
rect 195771 16189 195787 16307
rect 195477 16147 195787 16189
rect 195477 16029 195493 16147
rect 195611 16029 195653 16147
rect 195771 16029 195787 16147
rect 186477 -3171 186493 -3053
rect 186611 -3171 186653 -3053
rect 186771 -3171 186787 -3053
rect 186477 -3213 186787 -3171
rect 186477 -3331 186493 -3213
rect 186611 -3331 186653 -3213
rect 186771 -3331 186787 -3213
rect 186477 -3827 186787 -3331
rect 195477 -3533 195787 16029
rect 198897 352419 199207 352915
rect 198897 352301 198913 352419
rect 199031 352301 199073 352419
rect 199191 352301 199207 352419
rect 198897 352259 199207 352301
rect 198897 352141 198913 352259
rect 199031 352141 199073 352259
rect 199191 352141 199207 352259
rect 198897 343727 199207 352141
rect 198897 343609 198913 343727
rect 199031 343609 199073 343727
rect 199191 343609 199207 343727
rect 198897 343567 199207 343609
rect 198897 343449 198913 343567
rect 199031 343449 199073 343567
rect 199191 343449 199207 343567
rect 198897 325727 199207 343449
rect 198897 325609 198913 325727
rect 199031 325609 199073 325727
rect 199191 325609 199207 325727
rect 198897 325567 199207 325609
rect 198897 325449 198913 325567
rect 199031 325449 199073 325567
rect 199191 325449 199207 325567
rect 198897 307727 199207 325449
rect 198897 307609 198913 307727
rect 199031 307609 199073 307727
rect 199191 307609 199207 307727
rect 198897 307567 199207 307609
rect 198897 307449 198913 307567
rect 199031 307449 199073 307567
rect 199191 307449 199207 307567
rect 198897 289727 199207 307449
rect 198897 289609 198913 289727
rect 199031 289609 199073 289727
rect 199191 289609 199207 289727
rect 198897 289567 199207 289609
rect 198897 289449 198913 289567
rect 199031 289449 199073 289567
rect 199191 289449 199207 289567
rect 198897 271727 199207 289449
rect 198897 271609 198913 271727
rect 199031 271609 199073 271727
rect 199191 271609 199207 271727
rect 198897 271567 199207 271609
rect 198897 271449 198913 271567
rect 199031 271449 199073 271567
rect 199191 271449 199207 271567
rect 198897 253727 199207 271449
rect 198897 253609 198913 253727
rect 199031 253609 199073 253727
rect 199191 253609 199207 253727
rect 198897 253567 199207 253609
rect 198897 253449 198913 253567
rect 199031 253449 199073 253567
rect 199191 253449 199207 253567
rect 198897 235727 199207 253449
rect 198897 235609 198913 235727
rect 199031 235609 199073 235727
rect 199191 235609 199207 235727
rect 198897 235567 199207 235609
rect 198897 235449 198913 235567
rect 199031 235449 199073 235567
rect 199191 235449 199207 235567
rect 198897 217727 199207 235449
rect 198897 217609 198913 217727
rect 199031 217609 199073 217727
rect 199191 217609 199207 217727
rect 198897 217567 199207 217609
rect 198897 217449 198913 217567
rect 199031 217449 199073 217567
rect 199191 217449 199207 217567
rect 198897 199727 199207 217449
rect 198897 199609 198913 199727
rect 199031 199609 199073 199727
rect 199191 199609 199207 199727
rect 198897 199567 199207 199609
rect 198897 199449 198913 199567
rect 199031 199449 199073 199567
rect 199191 199449 199207 199567
rect 198897 181727 199207 199449
rect 198897 181609 198913 181727
rect 199031 181609 199073 181727
rect 199191 181609 199207 181727
rect 198897 181567 199207 181609
rect 198897 181449 198913 181567
rect 199031 181449 199073 181567
rect 199191 181449 199207 181567
rect 198897 163727 199207 181449
rect 198897 163609 198913 163727
rect 199031 163609 199073 163727
rect 199191 163609 199207 163727
rect 198897 163567 199207 163609
rect 198897 163449 198913 163567
rect 199031 163449 199073 163567
rect 199191 163449 199207 163567
rect 198897 145727 199207 163449
rect 198897 145609 198913 145727
rect 199031 145609 199073 145727
rect 199191 145609 199207 145727
rect 198897 145567 199207 145609
rect 198897 145449 198913 145567
rect 199031 145449 199073 145567
rect 199191 145449 199207 145567
rect 198897 127727 199207 145449
rect 198897 127609 198913 127727
rect 199031 127609 199073 127727
rect 199191 127609 199207 127727
rect 198897 127567 199207 127609
rect 198897 127449 198913 127567
rect 199031 127449 199073 127567
rect 199191 127449 199207 127567
rect 198897 109727 199207 127449
rect 198897 109609 198913 109727
rect 199031 109609 199073 109727
rect 199191 109609 199207 109727
rect 198897 109567 199207 109609
rect 198897 109449 198913 109567
rect 199031 109449 199073 109567
rect 199191 109449 199207 109567
rect 198897 91727 199207 109449
rect 198897 91609 198913 91727
rect 199031 91609 199073 91727
rect 199191 91609 199207 91727
rect 198897 91567 199207 91609
rect 198897 91449 198913 91567
rect 199031 91449 199073 91567
rect 199191 91449 199207 91567
rect 198897 73727 199207 91449
rect 198897 73609 198913 73727
rect 199031 73609 199073 73727
rect 199191 73609 199207 73727
rect 198897 73567 199207 73609
rect 198897 73449 198913 73567
rect 199031 73449 199073 73567
rect 199191 73449 199207 73567
rect 198897 55727 199207 73449
rect 198897 55609 198913 55727
rect 199031 55609 199073 55727
rect 199191 55609 199207 55727
rect 198897 55567 199207 55609
rect 198897 55449 198913 55567
rect 199031 55449 199073 55567
rect 199191 55449 199207 55567
rect 198897 37727 199207 55449
rect 198897 37609 198913 37727
rect 199031 37609 199073 37727
rect 199191 37609 199207 37727
rect 198897 37567 199207 37609
rect 198897 37449 198913 37567
rect 199031 37449 199073 37567
rect 199191 37449 199207 37567
rect 198897 19727 199207 37449
rect 198897 19609 198913 19727
rect 199031 19609 199073 19727
rect 199191 19609 199207 19727
rect 198897 19567 199207 19609
rect 198897 19449 198913 19567
rect 199031 19449 199073 19567
rect 199191 19449 199207 19567
rect 198897 1727 199207 19449
rect 198897 1609 198913 1727
rect 199031 1609 199073 1727
rect 199191 1609 199207 1727
rect 198897 1567 199207 1609
rect 198897 1449 198913 1567
rect 199031 1449 199073 1567
rect 199191 1449 199207 1567
rect 198897 -173 199207 1449
rect 198897 -291 198913 -173
rect 199031 -291 199073 -173
rect 199191 -291 199207 -173
rect 198897 -333 199207 -291
rect 198897 -451 198913 -333
rect 199031 -451 199073 -333
rect 199191 -451 199207 -333
rect 198897 -947 199207 -451
rect 200757 345587 201067 353101
rect 200757 345469 200773 345587
rect 200891 345469 200933 345587
rect 201051 345469 201067 345587
rect 200757 345427 201067 345469
rect 200757 345309 200773 345427
rect 200891 345309 200933 345427
rect 201051 345309 201067 345427
rect 200757 327587 201067 345309
rect 200757 327469 200773 327587
rect 200891 327469 200933 327587
rect 201051 327469 201067 327587
rect 200757 327427 201067 327469
rect 200757 327309 200773 327427
rect 200891 327309 200933 327427
rect 201051 327309 201067 327427
rect 200757 309587 201067 327309
rect 200757 309469 200773 309587
rect 200891 309469 200933 309587
rect 201051 309469 201067 309587
rect 200757 309427 201067 309469
rect 200757 309309 200773 309427
rect 200891 309309 200933 309427
rect 201051 309309 201067 309427
rect 200757 291587 201067 309309
rect 200757 291469 200773 291587
rect 200891 291469 200933 291587
rect 201051 291469 201067 291587
rect 200757 291427 201067 291469
rect 200757 291309 200773 291427
rect 200891 291309 200933 291427
rect 201051 291309 201067 291427
rect 200757 273587 201067 291309
rect 200757 273469 200773 273587
rect 200891 273469 200933 273587
rect 201051 273469 201067 273587
rect 200757 273427 201067 273469
rect 200757 273309 200773 273427
rect 200891 273309 200933 273427
rect 201051 273309 201067 273427
rect 200757 255587 201067 273309
rect 200757 255469 200773 255587
rect 200891 255469 200933 255587
rect 201051 255469 201067 255587
rect 200757 255427 201067 255469
rect 200757 255309 200773 255427
rect 200891 255309 200933 255427
rect 201051 255309 201067 255427
rect 200757 237587 201067 255309
rect 200757 237469 200773 237587
rect 200891 237469 200933 237587
rect 201051 237469 201067 237587
rect 200757 237427 201067 237469
rect 200757 237309 200773 237427
rect 200891 237309 200933 237427
rect 201051 237309 201067 237427
rect 200757 219587 201067 237309
rect 200757 219469 200773 219587
rect 200891 219469 200933 219587
rect 201051 219469 201067 219587
rect 200757 219427 201067 219469
rect 200757 219309 200773 219427
rect 200891 219309 200933 219427
rect 201051 219309 201067 219427
rect 200757 201587 201067 219309
rect 200757 201469 200773 201587
rect 200891 201469 200933 201587
rect 201051 201469 201067 201587
rect 200757 201427 201067 201469
rect 200757 201309 200773 201427
rect 200891 201309 200933 201427
rect 201051 201309 201067 201427
rect 200757 183587 201067 201309
rect 200757 183469 200773 183587
rect 200891 183469 200933 183587
rect 201051 183469 201067 183587
rect 200757 183427 201067 183469
rect 200757 183309 200773 183427
rect 200891 183309 200933 183427
rect 201051 183309 201067 183427
rect 200757 165587 201067 183309
rect 200757 165469 200773 165587
rect 200891 165469 200933 165587
rect 201051 165469 201067 165587
rect 200757 165427 201067 165469
rect 200757 165309 200773 165427
rect 200891 165309 200933 165427
rect 201051 165309 201067 165427
rect 200757 147587 201067 165309
rect 200757 147469 200773 147587
rect 200891 147469 200933 147587
rect 201051 147469 201067 147587
rect 200757 147427 201067 147469
rect 200757 147309 200773 147427
rect 200891 147309 200933 147427
rect 201051 147309 201067 147427
rect 200757 129587 201067 147309
rect 200757 129469 200773 129587
rect 200891 129469 200933 129587
rect 201051 129469 201067 129587
rect 200757 129427 201067 129469
rect 200757 129309 200773 129427
rect 200891 129309 200933 129427
rect 201051 129309 201067 129427
rect 200757 111587 201067 129309
rect 200757 111469 200773 111587
rect 200891 111469 200933 111587
rect 201051 111469 201067 111587
rect 200757 111427 201067 111469
rect 200757 111309 200773 111427
rect 200891 111309 200933 111427
rect 201051 111309 201067 111427
rect 200757 93587 201067 111309
rect 200757 93469 200773 93587
rect 200891 93469 200933 93587
rect 201051 93469 201067 93587
rect 200757 93427 201067 93469
rect 200757 93309 200773 93427
rect 200891 93309 200933 93427
rect 201051 93309 201067 93427
rect 200757 75587 201067 93309
rect 200757 75469 200773 75587
rect 200891 75469 200933 75587
rect 201051 75469 201067 75587
rect 200757 75427 201067 75469
rect 200757 75309 200773 75427
rect 200891 75309 200933 75427
rect 201051 75309 201067 75427
rect 200757 57587 201067 75309
rect 200757 57469 200773 57587
rect 200891 57469 200933 57587
rect 201051 57469 201067 57587
rect 200757 57427 201067 57469
rect 200757 57309 200773 57427
rect 200891 57309 200933 57427
rect 201051 57309 201067 57427
rect 200757 39587 201067 57309
rect 200757 39469 200773 39587
rect 200891 39469 200933 39587
rect 201051 39469 201067 39587
rect 200757 39427 201067 39469
rect 200757 39309 200773 39427
rect 200891 39309 200933 39427
rect 201051 39309 201067 39427
rect 200757 21587 201067 39309
rect 200757 21469 200773 21587
rect 200891 21469 200933 21587
rect 201051 21469 201067 21587
rect 200757 21427 201067 21469
rect 200757 21309 200773 21427
rect 200891 21309 200933 21427
rect 201051 21309 201067 21427
rect 200757 3587 201067 21309
rect 200757 3469 200773 3587
rect 200891 3469 200933 3587
rect 201051 3469 201067 3587
rect 200757 3427 201067 3469
rect 200757 3309 200773 3427
rect 200891 3309 200933 3427
rect 201051 3309 201067 3427
rect 200757 -1133 201067 3309
rect 200757 -1251 200773 -1133
rect 200891 -1251 200933 -1133
rect 201051 -1251 201067 -1133
rect 200757 -1293 201067 -1251
rect 200757 -1411 200773 -1293
rect 200891 -1411 200933 -1293
rect 201051 -1411 201067 -1293
rect 200757 -1907 201067 -1411
rect 202617 347447 202927 354061
rect 202617 347329 202633 347447
rect 202751 347329 202793 347447
rect 202911 347329 202927 347447
rect 202617 347287 202927 347329
rect 202617 347169 202633 347287
rect 202751 347169 202793 347287
rect 202911 347169 202927 347287
rect 202617 329447 202927 347169
rect 202617 329329 202633 329447
rect 202751 329329 202793 329447
rect 202911 329329 202927 329447
rect 202617 329287 202927 329329
rect 202617 329169 202633 329287
rect 202751 329169 202793 329287
rect 202911 329169 202927 329287
rect 202617 311447 202927 329169
rect 202617 311329 202633 311447
rect 202751 311329 202793 311447
rect 202911 311329 202927 311447
rect 202617 311287 202927 311329
rect 202617 311169 202633 311287
rect 202751 311169 202793 311287
rect 202911 311169 202927 311287
rect 202617 293447 202927 311169
rect 202617 293329 202633 293447
rect 202751 293329 202793 293447
rect 202911 293329 202927 293447
rect 202617 293287 202927 293329
rect 202617 293169 202633 293287
rect 202751 293169 202793 293287
rect 202911 293169 202927 293287
rect 202617 275447 202927 293169
rect 202617 275329 202633 275447
rect 202751 275329 202793 275447
rect 202911 275329 202927 275447
rect 202617 275287 202927 275329
rect 202617 275169 202633 275287
rect 202751 275169 202793 275287
rect 202911 275169 202927 275287
rect 202617 257447 202927 275169
rect 202617 257329 202633 257447
rect 202751 257329 202793 257447
rect 202911 257329 202927 257447
rect 202617 257287 202927 257329
rect 202617 257169 202633 257287
rect 202751 257169 202793 257287
rect 202911 257169 202927 257287
rect 202617 239447 202927 257169
rect 202617 239329 202633 239447
rect 202751 239329 202793 239447
rect 202911 239329 202927 239447
rect 202617 239287 202927 239329
rect 202617 239169 202633 239287
rect 202751 239169 202793 239287
rect 202911 239169 202927 239287
rect 202617 221447 202927 239169
rect 202617 221329 202633 221447
rect 202751 221329 202793 221447
rect 202911 221329 202927 221447
rect 202617 221287 202927 221329
rect 202617 221169 202633 221287
rect 202751 221169 202793 221287
rect 202911 221169 202927 221287
rect 202617 203447 202927 221169
rect 202617 203329 202633 203447
rect 202751 203329 202793 203447
rect 202911 203329 202927 203447
rect 202617 203287 202927 203329
rect 202617 203169 202633 203287
rect 202751 203169 202793 203287
rect 202911 203169 202927 203287
rect 202617 185447 202927 203169
rect 202617 185329 202633 185447
rect 202751 185329 202793 185447
rect 202911 185329 202927 185447
rect 202617 185287 202927 185329
rect 202617 185169 202633 185287
rect 202751 185169 202793 185287
rect 202911 185169 202927 185287
rect 202617 167447 202927 185169
rect 202617 167329 202633 167447
rect 202751 167329 202793 167447
rect 202911 167329 202927 167447
rect 202617 167287 202927 167329
rect 202617 167169 202633 167287
rect 202751 167169 202793 167287
rect 202911 167169 202927 167287
rect 202617 149447 202927 167169
rect 202617 149329 202633 149447
rect 202751 149329 202793 149447
rect 202911 149329 202927 149447
rect 202617 149287 202927 149329
rect 202617 149169 202633 149287
rect 202751 149169 202793 149287
rect 202911 149169 202927 149287
rect 202617 131447 202927 149169
rect 202617 131329 202633 131447
rect 202751 131329 202793 131447
rect 202911 131329 202927 131447
rect 202617 131287 202927 131329
rect 202617 131169 202633 131287
rect 202751 131169 202793 131287
rect 202911 131169 202927 131287
rect 202617 113447 202927 131169
rect 202617 113329 202633 113447
rect 202751 113329 202793 113447
rect 202911 113329 202927 113447
rect 202617 113287 202927 113329
rect 202617 113169 202633 113287
rect 202751 113169 202793 113287
rect 202911 113169 202927 113287
rect 202617 95447 202927 113169
rect 202617 95329 202633 95447
rect 202751 95329 202793 95447
rect 202911 95329 202927 95447
rect 202617 95287 202927 95329
rect 202617 95169 202633 95287
rect 202751 95169 202793 95287
rect 202911 95169 202927 95287
rect 202617 77447 202927 95169
rect 202617 77329 202633 77447
rect 202751 77329 202793 77447
rect 202911 77329 202927 77447
rect 202617 77287 202927 77329
rect 202617 77169 202633 77287
rect 202751 77169 202793 77287
rect 202911 77169 202927 77287
rect 202617 59447 202927 77169
rect 202617 59329 202633 59447
rect 202751 59329 202793 59447
rect 202911 59329 202927 59447
rect 202617 59287 202927 59329
rect 202617 59169 202633 59287
rect 202751 59169 202793 59287
rect 202911 59169 202927 59287
rect 202617 41447 202927 59169
rect 202617 41329 202633 41447
rect 202751 41329 202793 41447
rect 202911 41329 202927 41447
rect 202617 41287 202927 41329
rect 202617 41169 202633 41287
rect 202751 41169 202793 41287
rect 202911 41169 202927 41287
rect 202617 23447 202927 41169
rect 202617 23329 202633 23447
rect 202751 23329 202793 23447
rect 202911 23329 202927 23447
rect 202617 23287 202927 23329
rect 202617 23169 202633 23287
rect 202751 23169 202793 23287
rect 202911 23169 202927 23287
rect 202617 5447 202927 23169
rect 202617 5329 202633 5447
rect 202751 5329 202793 5447
rect 202911 5329 202927 5447
rect 202617 5287 202927 5329
rect 202617 5169 202633 5287
rect 202751 5169 202793 5287
rect 202911 5169 202927 5287
rect 202617 -2093 202927 5169
rect 202617 -2211 202633 -2093
rect 202751 -2211 202793 -2093
rect 202911 -2211 202927 -2093
rect 202617 -2253 202927 -2211
rect 202617 -2371 202633 -2253
rect 202751 -2371 202793 -2253
rect 202911 -2371 202927 -2253
rect 202617 -2867 202927 -2371
rect 204477 349307 204787 355021
rect 213477 355779 213787 355795
rect 213477 355661 213493 355779
rect 213611 355661 213653 355779
rect 213771 355661 213787 355779
rect 213477 355619 213787 355661
rect 213477 355501 213493 355619
rect 213611 355501 213653 355619
rect 213771 355501 213787 355619
rect 211617 354819 211927 354835
rect 211617 354701 211633 354819
rect 211751 354701 211793 354819
rect 211911 354701 211927 354819
rect 211617 354659 211927 354701
rect 211617 354541 211633 354659
rect 211751 354541 211793 354659
rect 211911 354541 211927 354659
rect 209757 353859 210067 353875
rect 209757 353741 209773 353859
rect 209891 353741 209933 353859
rect 210051 353741 210067 353859
rect 209757 353699 210067 353741
rect 209757 353581 209773 353699
rect 209891 353581 209933 353699
rect 210051 353581 210067 353699
rect 204477 349189 204493 349307
rect 204611 349189 204653 349307
rect 204771 349189 204787 349307
rect 204477 349147 204787 349189
rect 204477 349029 204493 349147
rect 204611 349029 204653 349147
rect 204771 349029 204787 349147
rect 204477 331307 204787 349029
rect 204477 331189 204493 331307
rect 204611 331189 204653 331307
rect 204771 331189 204787 331307
rect 204477 331147 204787 331189
rect 204477 331029 204493 331147
rect 204611 331029 204653 331147
rect 204771 331029 204787 331147
rect 204477 313307 204787 331029
rect 204477 313189 204493 313307
rect 204611 313189 204653 313307
rect 204771 313189 204787 313307
rect 204477 313147 204787 313189
rect 204477 313029 204493 313147
rect 204611 313029 204653 313147
rect 204771 313029 204787 313147
rect 204477 295307 204787 313029
rect 204477 295189 204493 295307
rect 204611 295189 204653 295307
rect 204771 295189 204787 295307
rect 204477 295147 204787 295189
rect 204477 295029 204493 295147
rect 204611 295029 204653 295147
rect 204771 295029 204787 295147
rect 204477 277307 204787 295029
rect 204477 277189 204493 277307
rect 204611 277189 204653 277307
rect 204771 277189 204787 277307
rect 204477 277147 204787 277189
rect 204477 277029 204493 277147
rect 204611 277029 204653 277147
rect 204771 277029 204787 277147
rect 204477 259307 204787 277029
rect 204477 259189 204493 259307
rect 204611 259189 204653 259307
rect 204771 259189 204787 259307
rect 204477 259147 204787 259189
rect 204477 259029 204493 259147
rect 204611 259029 204653 259147
rect 204771 259029 204787 259147
rect 204477 241307 204787 259029
rect 204477 241189 204493 241307
rect 204611 241189 204653 241307
rect 204771 241189 204787 241307
rect 204477 241147 204787 241189
rect 204477 241029 204493 241147
rect 204611 241029 204653 241147
rect 204771 241029 204787 241147
rect 204477 223307 204787 241029
rect 204477 223189 204493 223307
rect 204611 223189 204653 223307
rect 204771 223189 204787 223307
rect 204477 223147 204787 223189
rect 204477 223029 204493 223147
rect 204611 223029 204653 223147
rect 204771 223029 204787 223147
rect 204477 205307 204787 223029
rect 204477 205189 204493 205307
rect 204611 205189 204653 205307
rect 204771 205189 204787 205307
rect 204477 205147 204787 205189
rect 204477 205029 204493 205147
rect 204611 205029 204653 205147
rect 204771 205029 204787 205147
rect 204477 187307 204787 205029
rect 204477 187189 204493 187307
rect 204611 187189 204653 187307
rect 204771 187189 204787 187307
rect 204477 187147 204787 187189
rect 204477 187029 204493 187147
rect 204611 187029 204653 187147
rect 204771 187029 204787 187147
rect 204477 169307 204787 187029
rect 204477 169189 204493 169307
rect 204611 169189 204653 169307
rect 204771 169189 204787 169307
rect 204477 169147 204787 169189
rect 204477 169029 204493 169147
rect 204611 169029 204653 169147
rect 204771 169029 204787 169147
rect 204477 151307 204787 169029
rect 204477 151189 204493 151307
rect 204611 151189 204653 151307
rect 204771 151189 204787 151307
rect 204477 151147 204787 151189
rect 204477 151029 204493 151147
rect 204611 151029 204653 151147
rect 204771 151029 204787 151147
rect 204477 133307 204787 151029
rect 204477 133189 204493 133307
rect 204611 133189 204653 133307
rect 204771 133189 204787 133307
rect 204477 133147 204787 133189
rect 204477 133029 204493 133147
rect 204611 133029 204653 133147
rect 204771 133029 204787 133147
rect 204477 115307 204787 133029
rect 204477 115189 204493 115307
rect 204611 115189 204653 115307
rect 204771 115189 204787 115307
rect 204477 115147 204787 115189
rect 204477 115029 204493 115147
rect 204611 115029 204653 115147
rect 204771 115029 204787 115147
rect 204477 97307 204787 115029
rect 204477 97189 204493 97307
rect 204611 97189 204653 97307
rect 204771 97189 204787 97307
rect 204477 97147 204787 97189
rect 204477 97029 204493 97147
rect 204611 97029 204653 97147
rect 204771 97029 204787 97147
rect 204477 79307 204787 97029
rect 204477 79189 204493 79307
rect 204611 79189 204653 79307
rect 204771 79189 204787 79307
rect 204477 79147 204787 79189
rect 204477 79029 204493 79147
rect 204611 79029 204653 79147
rect 204771 79029 204787 79147
rect 204477 61307 204787 79029
rect 204477 61189 204493 61307
rect 204611 61189 204653 61307
rect 204771 61189 204787 61307
rect 204477 61147 204787 61189
rect 204477 61029 204493 61147
rect 204611 61029 204653 61147
rect 204771 61029 204787 61147
rect 204477 43307 204787 61029
rect 204477 43189 204493 43307
rect 204611 43189 204653 43307
rect 204771 43189 204787 43307
rect 204477 43147 204787 43189
rect 204477 43029 204493 43147
rect 204611 43029 204653 43147
rect 204771 43029 204787 43147
rect 204477 25307 204787 43029
rect 204477 25189 204493 25307
rect 204611 25189 204653 25307
rect 204771 25189 204787 25307
rect 204477 25147 204787 25189
rect 204477 25029 204493 25147
rect 204611 25029 204653 25147
rect 204771 25029 204787 25147
rect 204477 7307 204787 25029
rect 204477 7189 204493 7307
rect 204611 7189 204653 7307
rect 204771 7189 204787 7307
rect 204477 7147 204787 7189
rect 204477 7029 204493 7147
rect 204611 7029 204653 7147
rect 204771 7029 204787 7147
rect 195477 -3651 195493 -3533
rect 195611 -3651 195653 -3533
rect 195771 -3651 195787 -3533
rect 195477 -3693 195787 -3651
rect 195477 -3811 195493 -3693
rect 195611 -3811 195653 -3693
rect 195771 -3811 195787 -3693
rect 195477 -3827 195787 -3811
rect 204477 -3053 204787 7029
rect 207897 352899 208207 352915
rect 207897 352781 207913 352899
rect 208031 352781 208073 352899
rect 208191 352781 208207 352899
rect 207897 352739 208207 352781
rect 207897 352621 207913 352739
rect 208031 352621 208073 352739
rect 208191 352621 208207 352739
rect 207897 334727 208207 352621
rect 207897 334609 207913 334727
rect 208031 334609 208073 334727
rect 208191 334609 208207 334727
rect 207897 334567 208207 334609
rect 207897 334449 207913 334567
rect 208031 334449 208073 334567
rect 208191 334449 208207 334567
rect 207897 316727 208207 334449
rect 207897 316609 207913 316727
rect 208031 316609 208073 316727
rect 208191 316609 208207 316727
rect 207897 316567 208207 316609
rect 207897 316449 207913 316567
rect 208031 316449 208073 316567
rect 208191 316449 208207 316567
rect 207897 298727 208207 316449
rect 207897 298609 207913 298727
rect 208031 298609 208073 298727
rect 208191 298609 208207 298727
rect 207897 298567 208207 298609
rect 207897 298449 207913 298567
rect 208031 298449 208073 298567
rect 208191 298449 208207 298567
rect 207897 280727 208207 298449
rect 207897 280609 207913 280727
rect 208031 280609 208073 280727
rect 208191 280609 208207 280727
rect 207897 280567 208207 280609
rect 207897 280449 207913 280567
rect 208031 280449 208073 280567
rect 208191 280449 208207 280567
rect 207897 262727 208207 280449
rect 207897 262609 207913 262727
rect 208031 262609 208073 262727
rect 208191 262609 208207 262727
rect 207897 262567 208207 262609
rect 207897 262449 207913 262567
rect 208031 262449 208073 262567
rect 208191 262449 208207 262567
rect 207897 244727 208207 262449
rect 207897 244609 207913 244727
rect 208031 244609 208073 244727
rect 208191 244609 208207 244727
rect 207897 244567 208207 244609
rect 207897 244449 207913 244567
rect 208031 244449 208073 244567
rect 208191 244449 208207 244567
rect 207897 226727 208207 244449
rect 207897 226609 207913 226727
rect 208031 226609 208073 226727
rect 208191 226609 208207 226727
rect 207897 226567 208207 226609
rect 207897 226449 207913 226567
rect 208031 226449 208073 226567
rect 208191 226449 208207 226567
rect 207897 208727 208207 226449
rect 207897 208609 207913 208727
rect 208031 208609 208073 208727
rect 208191 208609 208207 208727
rect 207897 208567 208207 208609
rect 207897 208449 207913 208567
rect 208031 208449 208073 208567
rect 208191 208449 208207 208567
rect 207897 190727 208207 208449
rect 207897 190609 207913 190727
rect 208031 190609 208073 190727
rect 208191 190609 208207 190727
rect 207897 190567 208207 190609
rect 207897 190449 207913 190567
rect 208031 190449 208073 190567
rect 208191 190449 208207 190567
rect 207897 172727 208207 190449
rect 207897 172609 207913 172727
rect 208031 172609 208073 172727
rect 208191 172609 208207 172727
rect 207897 172567 208207 172609
rect 207897 172449 207913 172567
rect 208031 172449 208073 172567
rect 208191 172449 208207 172567
rect 207897 154727 208207 172449
rect 207897 154609 207913 154727
rect 208031 154609 208073 154727
rect 208191 154609 208207 154727
rect 207897 154567 208207 154609
rect 207897 154449 207913 154567
rect 208031 154449 208073 154567
rect 208191 154449 208207 154567
rect 207897 136727 208207 154449
rect 207897 136609 207913 136727
rect 208031 136609 208073 136727
rect 208191 136609 208207 136727
rect 207897 136567 208207 136609
rect 207897 136449 207913 136567
rect 208031 136449 208073 136567
rect 208191 136449 208207 136567
rect 207897 118727 208207 136449
rect 207897 118609 207913 118727
rect 208031 118609 208073 118727
rect 208191 118609 208207 118727
rect 207897 118567 208207 118609
rect 207897 118449 207913 118567
rect 208031 118449 208073 118567
rect 208191 118449 208207 118567
rect 207897 100727 208207 118449
rect 207897 100609 207913 100727
rect 208031 100609 208073 100727
rect 208191 100609 208207 100727
rect 207897 100567 208207 100609
rect 207897 100449 207913 100567
rect 208031 100449 208073 100567
rect 208191 100449 208207 100567
rect 207897 82727 208207 100449
rect 207897 82609 207913 82727
rect 208031 82609 208073 82727
rect 208191 82609 208207 82727
rect 207897 82567 208207 82609
rect 207897 82449 207913 82567
rect 208031 82449 208073 82567
rect 208191 82449 208207 82567
rect 207897 64727 208207 82449
rect 207897 64609 207913 64727
rect 208031 64609 208073 64727
rect 208191 64609 208207 64727
rect 207897 64567 208207 64609
rect 207897 64449 207913 64567
rect 208031 64449 208073 64567
rect 208191 64449 208207 64567
rect 207897 46727 208207 64449
rect 207897 46609 207913 46727
rect 208031 46609 208073 46727
rect 208191 46609 208207 46727
rect 207897 46567 208207 46609
rect 207897 46449 207913 46567
rect 208031 46449 208073 46567
rect 208191 46449 208207 46567
rect 207897 28727 208207 46449
rect 207897 28609 207913 28727
rect 208031 28609 208073 28727
rect 208191 28609 208207 28727
rect 207897 28567 208207 28609
rect 207897 28449 207913 28567
rect 208031 28449 208073 28567
rect 208191 28449 208207 28567
rect 207897 10727 208207 28449
rect 207897 10609 207913 10727
rect 208031 10609 208073 10727
rect 208191 10609 208207 10727
rect 207897 10567 208207 10609
rect 207897 10449 207913 10567
rect 208031 10449 208073 10567
rect 208191 10449 208207 10567
rect 207897 -653 208207 10449
rect 207897 -771 207913 -653
rect 208031 -771 208073 -653
rect 208191 -771 208207 -653
rect 207897 -813 208207 -771
rect 207897 -931 207913 -813
rect 208031 -931 208073 -813
rect 208191 -931 208207 -813
rect 207897 -947 208207 -931
rect 209757 336587 210067 353581
rect 209757 336469 209773 336587
rect 209891 336469 209933 336587
rect 210051 336469 210067 336587
rect 209757 336427 210067 336469
rect 209757 336309 209773 336427
rect 209891 336309 209933 336427
rect 210051 336309 210067 336427
rect 209757 318587 210067 336309
rect 209757 318469 209773 318587
rect 209891 318469 209933 318587
rect 210051 318469 210067 318587
rect 209757 318427 210067 318469
rect 209757 318309 209773 318427
rect 209891 318309 209933 318427
rect 210051 318309 210067 318427
rect 209757 300587 210067 318309
rect 209757 300469 209773 300587
rect 209891 300469 209933 300587
rect 210051 300469 210067 300587
rect 209757 300427 210067 300469
rect 209757 300309 209773 300427
rect 209891 300309 209933 300427
rect 210051 300309 210067 300427
rect 209757 282587 210067 300309
rect 209757 282469 209773 282587
rect 209891 282469 209933 282587
rect 210051 282469 210067 282587
rect 209757 282427 210067 282469
rect 209757 282309 209773 282427
rect 209891 282309 209933 282427
rect 210051 282309 210067 282427
rect 209757 264587 210067 282309
rect 209757 264469 209773 264587
rect 209891 264469 209933 264587
rect 210051 264469 210067 264587
rect 209757 264427 210067 264469
rect 209757 264309 209773 264427
rect 209891 264309 209933 264427
rect 210051 264309 210067 264427
rect 209757 246587 210067 264309
rect 209757 246469 209773 246587
rect 209891 246469 209933 246587
rect 210051 246469 210067 246587
rect 209757 246427 210067 246469
rect 209757 246309 209773 246427
rect 209891 246309 209933 246427
rect 210051 246309 210067 246427
rect 209757 228587 210067 246309
rect 209757 228469 209773 228587
rect 209891 228469 209933 228587
rect 210051 228469 210067 228587
rect 209757 228427 210067 228469
rect 209757 228309 209773 228427
rect 209891 228309 209933 228427
rect 210051 228309 210067 228427
rect 209757 210587 210067 228309
rect 209757 210469 209773 210587
rect 209891 210469 209933 210587
rect 210051 210469 210067 210587
rect 209757 210427 210067 210469
rect 209757 210309 209773 210427
rect 209891 210309 209933 210427
rect 210051 210309 210067 210427
rect 209757 192587 210067 210309
rect 209757 192469 209773 192587
rect 209891 192469 209933 192587
rect 210051 192469 210067 192587
rect 209757 192427 210067 192469
rect 209757 192309 209773 192427
rect 209891 192309 209933 192427
rect 210051 192309 210067 192427
rect 209757 174587 210067 192309
rect 209757 174469 209773 174587
rect 209891 174469 209933 174587
rect 210051 174469 210067 174587
rect 209757 174427 210067 174469
rect 209757 174309 209773 174427
rect 209891 174309 209933 174427
rect 210051 174309 210067 174427
rect 209757 156587 210067 174309
rect 209757 156469 209773 156587
rect 209891 156469 209933 156587
rect 210051 156469 210067 156587
rect 209757 156427 210067 156469
rect 209757 156309 209773 156427
rect 209891 156309 209933 156427
rect 210051 156309 210067 156427
rect 209757 138587 210067 156309
rect 209757 138469 209773 138587
rect 209891 138469 209933 138587
rect 210051 138469 210067 138587
rect 209757 138427 210067 138469
rect 209757 138309 209773 138427
rect 209891 138309 209933 138427
rect 210051 138309 210067 138427
rect 209757 120587 210067 138309
rect 209757 120469 209773 120587
rect 209891 120469 209933 120587
rect 210051 120469 210067 120587
rect 209757 120427 210067 120469
rect 209757 120309 209773 120427
rect 209891 120309 209933 120427
rect 210051 120309 210067 120427
rect 209757 102587 210067 120309
rect 209757 102469 209773 102587
rect 209891 102469 209933 102587
rect 210051 102469 210067 102587
rect 209757 102427 210067 102469
rect 209757 102309 209773 102427
rect 209891 102309 209933 102427
rect 210051 102309 210067 102427
rect 209757 84587 210067 102309
rect 209757 84469 209773 84587
rect 209891 84469 209933 84587
rect 210051 84469 210067 84587
rect 209757 84427 210067 84469
rect 209757 84309 209773 84427
rect 209891 84309 209933 84427
rect 210051 84309 210067 84427
rect 209757 66587 210067 84309
rect 209757 66469 209773 66587
rect 209891 66469 209933 66587
rect 210051 66469 210067 66587
rect 209757 66427 210067 66469
rect 209757 66309 209773 66427
rect 209891 66309 209933 66427
rect 210051 66309 210067 66427
rect 209757 48587 210067 66309
rect 209757 48469 209773 48587
rect 209891 48469 209933 48587
rect 210051 48469 210067 48587
rect 209757 48427 210067 48469
rect 209757 48309 209773 48427
rect 209891 48309 209933 48427
rect 210051 48309 210067 48427
rect 209757 30587 210067 48309
rect 209757 30469 209773 30587
rect 209891 30469 209933 30587
rect 210051 30469 210067 30587
rect 209757 30427 210067 30469
rect 209757 30309 209773 30427
rect 209891 30309 209933 30427
rect 210051 30309 210067 30427
rect 209757 12587 210067 30309
rect 209757 12469 209773 12587
rect 209891 12469 209933 12587
rect 210051 12469 210067 12587
rect 209757 12427 210067 12469
rect 209757 12309 209773 12427
rect 209891 12309 209933 12427
rect 210051 12309 210067 12427
rect 209757 -1613 210067 12309
rect 209757 -1731 209773 -1613
rect 209891 -1731 209933 -1613
rect 210051 -1731 210067 -1613
rect 209757 -1773 210067 -1731
rect 209757 -1891 209773 -1773
rect 209891 -1891 209933 -1773
rect 210051 -1891 210067 -1773
rect 209757 -1907 210067 -1891
rect 211617 338447 211927 354541
rect 211617 338329 211633 338447
rect 211751 338329 211793 338447
rect 211911 338329 211927 338447
rect 211617 338287 211927 338329
rect 211617 338169 211633 338287
rect 211751 338169 211793 338287
rect 211911 338169 211927 338287
rect 211617 320447 211927 338169
rect 211617 320329 211633 320447
rect 211751 320329 211793 320447
rect 211911 320329 211927 320447
rect 211617 320287 211927 320329
rect 211617 320169 211633 320287
rect 211751 320169 211793 320287
rect 211911 320169 211927 320287
rect 211617 302447 211927 320169
rect 211617 302329 211633 302447
rect 211751 302329 211793 302447
rect 211911 302329 211927 302447
rect 211617 302287 211927 302329
rect 211617 302169 211633 302287
rect 211751 302169 211793 302287
rect 211911 302169 211927 302287
rect 211617 284447 211927 302169
rect 211617 284329 211633 284447
rect 211751 284329 211793 284447
rect 211911 284329 211927 284447
rect 211617 284287 211927 284329
rect 211617 284169 211633 284287
rect 211751 284169 211793 284287
rect 211911 284169 211927 284287
rect 211617 266447 211927 284169
rect 211617 266329 211633 266447
rect 211751 266329 211793 266447
rect 211911 266329 211927 266447
rect 211617 266287 211927 266329
rect 211617 266169 211633 266287
rect 211751 266169 211793 266287
rect 211911 266169 211927 266287
rect 211617 248447 211927 266169
rect 211617 248329 211633 248447
rect 211751 248329 211793 248447
rect 211911 248329 211927 248447
rect 211617 248287 211927 248329
rect 211617 248169 211633 248287
rect 211751 248169 211793 248287
rect 211911 248169 211927 248287
rect 211617 230447 211927 248169
rect 211617 230329 211633 230447
rect 211751 230329 211793 230447
rect 211911 230329 211927 230447
rect 211617 230287 211927 230329
rect 211617 230169 211633 230287
rect 211751 230169 211793 230287
rect 211911 230169 211927 230287
rect 211617 212447 211927 230169
rect 211617 212329 211633 212447
rect 211751 212329 211793 212447
rect 211911 212329 211927 212447
rect 211617 212287 211927 212329
rect 211617 212169 211633 212287
rect 211751 212169 211793 212287
rect 211911 212169 211927 212287
rect 211617 194447 211927 212169
rect 211617 194329 211633 194447
rect 211751 194329 211793 194447
rect 211911 194329 211927 194447
rect 211617 194287 211927 194329
rect 211617 194169 211633 194287
rect 211751 194169 211793 194287
rect 211911 194169 211927 194287
rect 211617 176447 211927 194169
rect 211617 176329 211633 176447
rect 211751 176329 211793 176447
rect 211911 176329 211927 176447
rect 211617 176287 211927 176329
rect 211617 176169 211633 176287
rect 211751 176169 211793 176287
rect 211911 176169 211927 176287
rect 211617 158447 211927 176169
rect 211617 158329 211633 158447
rect 211751 158329 211793 158447
rect 211911 158329 211927 158447
rect 211617 158287 211927 158329
rect 211617 158169 211633 158287
rect 211751 158169 211793 158287
rect 211911 158169 211927 158287
rect 211617 140447 211927 158169
rect 211617 140329 211633 140447
rect 211751 140329 211793 140447
rect 211911 140329 211927 140447
rect 211617 140287 211927 140329
rect 211617 140169 211633 140287
rect 211751 140169 211793 140287
rect 211911 140169 211927 140287
rect 211617 122447 211927 140169
rect 211617 122329 211633 122447
rect 211751 122329 211793 122447
rect 211911 122329 211927 122447
rect 211617 122287 211927 122329
rect 211617 122169 211633 122287
rect 211751 122169 211793 122287
rect 211911 122169 211927 122287
rect 211617 104447 211927 122169
rect 211617 104329 211633 104447
rect 211751 104329 211793 104447
rect 211911 104329 211927 104447
rect 211617 104287 211927 104329
rect 211617 104169 211633 104287
rect 211751 104169 211793 104287
rect 211911 104169 211927 104287
rect 211617 86447 211927 104169
rect 211617 86329 211633 86447
rect 211751 86329 211793 86447
rect 211911 86329 211927 86447
rect 211617 86287 211927 86329
rect 211617 86169 211633 86287
rect 211751 86169 211793 86287
rect 211911 86169 211927 86287
rect 211617 68447 211927 86169
rect 211617 68329 211633 68447
rect 211751 68329 211793 68447
rect 211911 68329 211927 68447
rect 211617 68287 211927 68329
rect 211617 68169 211633 68287
rect 211751 68169 211793 68287
rect 211911 68169 211927 68287
rect 211617 50447 211927 68169
rect 211617 50329 211633 50447
rect 211751 50329 211793 50447
rect 211911 50329 211927 50447
rect 211617 50287 211927 50329
rect 211617 50169 211633 50287
rect 211751 50169 211793 50287
rect 211911 50169 211927 50287
rect 211617 32447 211927 50169
rect 211617 32329 211633 32447
rect 211751 32329 211793 32447
rect 211911 32329 211927 32447
rect 211617 32287 211927 32329
rect 211617 32169 211633 32287
rect 211751 32169 211793 32287
rect 211911 32169 211927 32287
rect 211617 14447 211927 32169
rect 211617 14329 211633 14447
rect 211751 14329 211793 14447
rect 211911 14329 211927 14447
rect 211617 14287 211927 14329
rect 211617 14169 211633 14287
rect 211751 14169 211793 14287
rect 211911 14169 211927 14287
rect 211617 -2573 211927 14169
rect 211617 -2691 211633 -2573
rect 211751 -2691 211793 -2573
rect 211911 -2691 211927 -2573
rect 211617 -2733 211927 -2691
rect 211617 -2851 211633 -2733
rect 211751 -2851 211793 -2733
rect 211911 -2851 211927 -2733
rect 211617 -2867 211927 -2851
rect 213477 340307 213787 355501
rect 222477 355299 222787 355795
rect 222477 355181 222493 355299
rect 222611 355181 222653 355299
rect 222771 355181 222787 355299
rect 222477 355139 222787 355181
rect 222477 355021 222493 355139
rect 222611 355021 222653 355139
rect 222771 355021 222787 355139
rect 220617 354339 220927 354835
rect 220617 354221 220633 354339
rect 220751 354221 220793 354339
rect 220911 354221 220927 354339
rect 220617 354179 220927 354221
rect 220617 354061 220633 354179
rect 220751 354061 220793 354179
rect 220911 354061 220927 354179
rect 218757 353379 219067 353875
rect 218757 353261 218773 353379
rect 218891 353261 218933 353379
rect 219051 353261 219067 353379
rect 218757 353219 219067 353261
rect 218757 353101 218773 353219
rect 218891 353101 218933 353219
rect 219051 353101 219067 353219
rect 213477 340189 213493 340307
rect 213611 340189 213653 340307
rect 213771 340189 213787 340307
rect 213477 340147 213787 340189
rect 213477 340029 213493 340147
rect 213611 340029 213653 340147
rect 213771 340029 213787 340147
rect 213477 322307 213787 340029
rect 213477 322189 213493 322307
rect 213611 322189 213653 322307
rect 213771 322189 213787 322307
rect 213477 322147 213787 322189
rect 213477 322029 213493 322147
rect 213611 322029 213653 322147
rect 213771 322029 213787 322147
rect 213477 304307 213787 322029
rect 213477 304189 213493 304307
rect 213611 304189 213653 304307
rect 213771 304189 213787 304307
rect 213477 304147 213787 304189
rect 213477 304029 213493 304147
rect 213611 304029 213653 304147
rect 213771 304029 213787 304147
rect 213477 286307 213787 304029
rect 213477 286189 213493 286307
rect 213611 286189 213653 286307
rect 213771 286189 213787 286307
rect 213477 286147 213787 286189
rect 213477 286029 213493 286147
rect 213611 286029 213653 286147
rect 213771 286029 213787 286147
rect 213477 268307 213787 286029
rect 213477 268189 213493 268307
rect 213611 268189 213653 268307
rect 213771 268189 213787 268307
rect 213477 268147 213787 268189
rect 213477 268029 213493 268147
rect 213611 268029 213653 268147
rect 213771 268029 213787 268147
rect 213477 250307 213787 268029
rect 213477 250189 213493 250307
rect 213611 250189 213653 250307
rect 213771 250189 213787 250307
rect 213477 250147 213787 250189
rect 213477 250029 213493 250147
rect 213611 250029 213653 250147
rect 213771 250029 213787 250147
rect 213477 232307 213787 250029
rect 213477 232189 213493 232307
rect 213611 232189 213653 232307
rect 213771 232189 213787 232307
rect 213477 232147 213787 232189
rect 213477 232029 213493 232147
rect 213611 232029 213653 232147
rect 213771 232029 213787 232147
rect 213477 214307 213787 232029
rect 213477 214189 213493 214307
rect 213611 214189 213653 214307
rect 213771 214189 213787 214307
rect 213477 214147 213787 214189
rect 213477 214029 213493 214147
rect 213611 214029 213653 214147
rect 213771 214029 213787 214147
rect 213477 196307 213787 214029
rect 213477 196189 213493 196307
rect 213611 196189 213653 196307
rect 213771 196189 213787 196307
rect 213477 196147 213787 196189
rect 213477 196029 213493 196147
rect 213611 196029 213653 196147
rect 213771 196029 213787 196147
rect 213477 178307 213787 196029
rect 213477 178189 213493 178307
rect 213611 178189 213653 178307
rect 213771 178189 213787 178307
rect 213477 178147 213787 178189
rect 213477 178029 213493 178147
rect 213611 178029 213653 178147
rect 213771 178029 213787 178147
rect 213477 160307 213787 178029
rect 213477 160189 213493 160307
rect 213611 160189 213653 160307
rect 213771 160189 213787 160307
rect 213477 160147 213787 160189
rect 213477 160029 213493 160147
rect 213611 160029 213653 160147
rect 213771 160029 213787 160147
rect 213477 142307 213787 160029
rect 213477 142189 213493 142307
rect 213611 142189 213653 142307
rect 213771 142189 213787 142307
rect 213477 142147 213787 142189
rect 213477 142029 213493 142147
rect 213611 142029 213653 142147
rect 213771 142029 213787 142147
rect 213477 124307 213787 142029
rect 213477 124189 213493 124307
rect 213611 124189 213653 124307
rect 213771 124189 213787 124307
rect 213477 124147 213787 124189
rect 213477 124029 213493 124147
rect 213611 124029 213653 124147
rect 213771 124029 213787 124147
rect 213477 106307 213787 124029
rect 213477 106189 213493 106307
rect 213611 106189 213653 106307
rect 213771 106189 213787 106307
rect 213477 106147 213787 106189
rect 213477 106029 213493 106147
rect 213611 106029 213653 106147
rect 213771 106029 213787 106147
rect 213477 88307 213787 106029
rect 213477 88189 213493 88307
rect 213611 88189 213653 88307
rect 213771 88189 213787 88307
rect 213477 88147 213787 88189
rect 213477 88029 213493 88147
rect 213611 88029 213653 88147
rect 213771 88029 213787 88147
rect 213477 70307 213787 88029
rect 213477 70189 213493 70307
rect 213611 70189 213653 70307
rect 213771 70189 213787 70307
rect 213477 70147 213787 70189
rect 213477 70029 213493 70147
rect 213611 70029 213653 70147
rect 213771 70029 213787 70147
rect 213477 52307 213787 70029
rect 213477 52189 213493 52307
rect 213611 52189 213653 52307
rect 213771 52189 213787 52307
rect 213477 52147 213787 52189
rect 213477 52029 213493 52147
rect 213611 52029 213653 52147
rect 213771 52029 213787 52147
rect 213477 34307 213787 52029
rect 213477 34189 213493 34307
rect 213611 34189 213653 34307
rect 213771 34189 213787 34307
rect 213477 34147 213787 34189
rect 213477 34029 213493 34147
rect 213611 34029 213653 34147
rect 213771 34029 213787 34147
rect 213477 16307 213787 34029
rect 213477 16189 213493 16307
rect 213611 16189 213653 16307
rect 213771 16189 213787 16307
rect 213477 16147 213787 16189
rect 213477 16029 213493 16147
rect 213611 16029 213653 16147
rect 213771 16029 213787 16147
rect 204477 -3171 204493 -3053
rect 204611 -3171 204653 -3053
rect 204771 -3171 204787 -3053
rect 204477 -3213 204787 -3171
rect 204477 -3331 204493 -3213
rect 204611 -3331 204653 -3213
rect 204771 -3331 204787 -3213
rect 204477 -3827 204787 -3331
rect 213477 -3533 213787 16029
rect 216897 352419 217207 352915
rect 216897 352301 216913 352419
rect 217031 352301 217073 352419
rect 217191 352301 217207 352419
rect 216897 352259 217207 352301
rect 216897 352141 216913 352259
rect 217031 352141 217073 352259
rect 217191 352141 217207 352259
rect 216897 343727 217207 352141
rect 216897 343609 216913 343727
rect 217031 343609 217073 343727
rect 217191 343609 217207 343727
rect 216897 343567 217207 343609
rect 216897 343449 216913 343567
rect 217031 343449 217073 343567
rect 217191 343449 217207 343567
rect 216897 325727 217207 343449
rect 216897 325609 216913 325727
rect 217031 325609 217073 325727
rect 217191 325609 217207 325727
rect 216897 325567 217207 325609
rect 216897 325449 216913 325567
rect 217031 325449 217073 325567
rect 217191 325449 217207 325567
rect 216897 307727 217207 325449
rect 216897 307609 216913 307727
rect 217031 307609 217073 307727
rect 217191 307609 217207 307727
rect 216897 307567 217207 307609
rect 216897 307449 216913 307567
rect 217031 307449 217073 307567
rect 217191 307449 217207 307567
rect 216897 289727 217207 307449
rect 216897 289609 216913 289727
rect 217031 289609 217073 289727
rect 217191 289609 217207 289727
rect 216897 289567 217207 289609
rect 216897 289449 216913 289567
rect 217031 289449 217073 289567
rect 217191 289449 217207 289567
rect 216897 271727 217207 289449
rect 216897 271609 216913 271727
rect 217031 271609 217073 271727
rect 217191 271609 217207 271727
rect 216897 271567 217207 271609
rect 216897 271449 216913 271567
rect 217031 271449 217073 271567
rect 217191 271449 217207 271567
rect 216897 253727 217207 271449
rect 216897 253609 216913 253727
rect 217031 253609 217073 253727
rect 217191 253609 217207 253727
rect 216897 253567 217207 253609
rect 216897 253449 216913 253567
rect 217031 253449 217073 253567
rect 217191 253449 217207 253567
rect 216897 235727 217207 253449
rect 216897 235609 216913 235727
rect 217031 235609 217073 235727
rect 217191 235609 217207 235727
rect 216897 235567 217207 235609
rect 216897 235449 216913 235567
rect 217031 235449 217073 235567
rect 217191 235449 217207 235567
rect 216897 217727 217207 235449
rect 216897 217609 216913 217727
rect 217031 217609 217073 217727
rect 217191 217609 217207 217727
rect 216897 217567 217207 217609
rect 216897 217449 216913 217567
rect 217031 217449 217073 217567
rect 217191 217449 217207 217567
rect 216897 199727 217207 217449
rect 216897 199609 216913 199727
rect 217031 199609 217073 199727
rect 217191 199609 217207 199727
rect 216897 199567 217207 199609
rect 216897 199449 216913 199567
rect 217031 199449 217073 199567
rect 217191 199449 217207 199567
rect 216897 181727 217207 199449
rect 216897 181609 216913 181727
rect 217031 181609 217073 181727
rect 217191 181609 217207 181727
rect 216897 181567 217207 181609
rect 216897 181449 216913 181567
rect 217031 181449 217073 181567
rect 217191 181449 217207 181567
rect 216897 163727 217207 181449
rect 216897 163609 216913 163727
rect 217031 163609 217073 163727
rect 217191 163609 217207 163727
rect 216897 163567 217207 163609
rect 216897 163449 216913 163567
rect 217031 163449 217073 163567
rect 217191 163449 217207 163567
rect 216897 145727 217207 163449
rect 216897 145609 216913 145727
rect 217031 145609 217073 145727
rect 217191 145609 217207 145727
rect 216897 145567 217207 145609
rect 216897 145449 216913 145567
rect 217031 145449 217073 145567
rect 217191 145449 217207 145567
rect 216897 127727 217207 145449
rect 216897 127609 216913 127727
rect 217031 127609 217073 127727
rect 217191 127609 217207 127727
rect 216897 127567 217207 127609
rect 216897 127449 216913 127567
rect 217031 127449 217073 127567
rect 217191 127449 217207 127567
rect 216897 109727 217207 127449
rect 216897 109609 216913 109727
rect 217031 109609 217073 109727
rect 217191 109609 217207 109727
rect 216897 109567 217207 109609
rect 216897 109449 216913 109567
rect 217031 109449 217073 109567
rect 217191 109449 217207 109567
rect 216897 91727 217207 109449
rect 216897 91609 216913 91727
rect 217031 91609 217073 91727
rect 217191 91609 217207 91727
rect 216897 91567 217207 91609
rect 216897 91449 216913 91567
rect 217031 91449 217073 91567
rect 217191 91449 217207 91567
rect 216897 73727 217207 91449
rect 216897 73609 216913 73727
rect 217031 73609 217073 73727
rect 217191 73609 217207 73727
rect 216897 73567 217207 73609
rect 216897 73449 216913 73567
rect 217031 73449 217073 73567
rect 217191 73449 217207 73567
rect 216897 55727 217207 73449
rect 216897 55609 216913 55727
rect 217031 55609 217073 55727
rect 217191 55609 217207 55727
rect 216897 55567 217207 55609
rect 216897 55449 216913 55567
rect 217031 55449 217073 55567
rect 217191 55449 217207 55567
rect 216897 37727 217207 55449
rect 216897 37609 216913 37727
rect 217031 37609 217073 37727
rect 217191 37609 217207 37727
rect 216897 37567 217207 37609
rect 216897 37449 216913 37567
rect 217031 37449 217073 37567
rect 217191 37449 217207 37567
rect 216897 19727 217207 37449
rect 216897 19609 216913 19727
rect 217031 19609 217073 19727
rect 217191 19609 217207 19727
rect 216897 19567 217207 19609
rect 216897 19449 216913 19567
rect 217031 19449 217073 19567
rect 217191 19449 217207 19567
rect 216897 1727 217207 19449
rect 216897 1609 216913 1727
rect 217031 1609 217073 1727
rect 217191 1609 217207 1727
rect 216897 1567 217207 1609
rect 216897 1449 216913 1567
rect 217031 1449 217073 1567
rect 217191 1449 217207 1567
rect 216897 -173 217207 1449
rect 216897 -291 216913 -173
rect 217031 -291 217073 -173
rect 217191 -291 217207 -173
rect 216897 -333 217207 -291
rect 216897 -451 216913 -333
rect 217031 -451 217073 -333
rect 217191 -451 217207 -333
rect 216897 -947 217207 -451
rect 218757 345587 219067 353101
rect 218757 345469 218773 345587
rect 218891 345469 218933 345587
rect 219051 345469 219067 345587
rect 218757 345427 219067 345469
rect 218757 345309 218773 345427
rect 218891 345309 218933 345427
rect 219051 345309 219067 345427
rect 218757 327587 219067 345309
rect 218757 327469 218773 327587
rect 218891 327469 218933 327587
rect 219051 327469 219067 327587
rect 218757 327427 219067 327469
rect 218757 327309 218773 327427
rect 218891 327309 218933 327427
rect 219051 327309 219067 327427
rect 218757 309587 219067 327309
rect 218757 309469 218773 309587
rect 218891 309469 218933 309587
rect 219051 309469 219067 309587
rect 218757 309427 219067 309469
rect 218757 309309 218773 309427
rect 218891 309309 218933 309427
rect 219051 309309 219067 309427
rect 218757 291587 219067 309309
rect 218757 291469 218773 291587
rect 218891 291469 218933 291587
rect 219051 291469 219067 291587
rect 218757 291427 219067 291469
rect 218757 291309 218773 291427
rect 218891 291309 218933 291427
rect 219051 291309 219067 291427
rect 218757 273587 219067 291309
rect 218757 273469 218773 273587
rect 218891 273469 218933 273587
rect 219051 273469 219067 273587
rect 218757 273427 219067 273469
rect 218757 273309 218773 273427
rect 218891 273309 218933 273427
rect 219051 273309 219067 273427
rect 218757 255587 219067 273309
rect 218757 255469 218773 255587
rect 218891 255469 218933 255587
rect 219051 255469 219067 255587
rect 218757 255427 219067 255469
rect 218757 255309 218773 255427
rect 218891 255309 218933 255427
rect 219051 255309 219067 255427
rect 218757 237587 219067 255309
rect 218757 237469 218773 237587
rect 218891 237469 218933 237587
rect 219051 237469 219067 237587
rect 218757 237427 219067 237469
rect 218757 237309 218773 237427
rect 218891 237309 218933 237427
rect 219051 237309 219067 237427
rect 218757 219587 219067 237309
rect 218757 219469 218773 219587
rect 218891 219469 218933 219587
rect 219051 219469 219067 219587
rect 218757 219427 219067 219469
rect 218757 219309 218773 219427
rect 218891 219309 218933 219427
rect 219051 219309 219067 219427
rect 218757 201587 219067 219309
rect 218757 201469 218773 201587
rect 218891 201469 218933 201587
rect 219051 201469 219067 201587
rect 218757 201427 219067 201469
rect 218757 201309 218773 201427
rect 218891 201309 218933 201427
rect 219051 201309 219067 201427
rect 218757 183587 219067 201309
rect 218757 183469 218773 183587
rect 218891 183469 218933 183587
rect 219051 183469 219067 183587
rect 218757 183427 219067 183469
rect 218757 183309 218773 183427
rect 218891 183309 218933 183427
rect 219051 183309 219067 183427
rect 218757 165587 219067 183309
rect 218757 165469 218773 165587
rect 218891 165469 218933 165587
rect 219051 165469 219067 165587
rect 218757 165427 219067 165469
rect 218757 165309 218773 165427
rect 218891 165309 218933 165427
rect 219051 165309 219067 165427
rect 218757 147587 219067 165309
rect 218757 147469 218773 147587
rect 218891 147469 218933 147587
rect 219051 147469 219067 147587
rect 218757 147427 219067 147469
rect 218757 147309 218773 147427
rect 218891 147309 218933 147427
rect 219051 147309 219067 147427
rect 218757 129587 219067 147309
rect 218757 129469 218773 129587
rect 218891 129469 218933 129587
rect 219051 129469 219067 129587
rect 218757 129427 219067 129469
rect 218757 129309 218773 129427
rect 218891 129309 218933 129427
rect 219051 129309 219067 129427
rect 218757 111587 219067 129309
rect 218757 111469 218773 111587
rect 218891 111469 218933 111587
rect 219051 111469 219067 111587
rect 218757 111427 219067 111469
rect 218757 111309 218773 111427
rect 218891 111309 218933 111427
rect 219051 111309 219067 111427
rect 218757 93587 219067 111309
rect 218757 93469 218773 93587
rect 218891 93469 218933 93587
rect 219051 93469 219067 93587
rect 218757 93427 219067 93469
rect 218757 93309 218773 93427
rect 218891 93309 218933 93427
rect 219051 93309 219067 93427
rect 218757 75587 219067 93309
rect 218757 75469 218773 75587
rect 218891 75469 218933 75587
rect 219051 75469 219067 75587
rect 218757 75427 219067 75469
rect 218757 75309 218773 75427
rect 218891 75309 218933 75427
rect 219051 75309 219067 75427
rect 218757 57587 219067 75309
rect 218757 57469 218773 57587
rect 218891 57469 218933 57587
rect 219051 57469 219067 57587
rect 218757 57427 219067 57469
rect 218757 57309 218773 57427
rect 218891 57309 218933 57427
rect 219051 57309 219067 57427
rect 218757 39587 219067 57309
rect 218757 39469 218773 39587
rect 218891 39469 218933 39587
rect 219051 39469 219067 39587
rect 218757 39427 219067 39469
rect 218757 39309 218773 39427
rect 218891 39309 218933 39427
rect 219051 39309 219067 39427
rect 218757 21587 219067 39309
rect 218757 21469 218773 21587
rect 218891 21469 218933 21587
rect 219051 21469 219067 21587
rect 218757 21427 219067 21469
rect 218757 21309 218773 21427
rect 218891 21309 218933 21427
rect 219051 21309 219067 21427
rect 218757 3587 219067 21309
rect 218757 3469 218773 3587
rect 218891 3469 218933 3587
rect 219051 3469 219067 3587
rect 218757 3427 219067 3469
rect 218757 3309 218773 3427
rect 218891 3309 218933 3427
rect 219051 3309 219067 3427
rect 218757 -1133 219067 3309
rect 218757 -1251 218773 -1133
rect 218891 -1251 218933 -1133
rect 219051 -1251 219067 -1133
rect 218757 -1293 219067 -1251
rect 218757 -1411 218773 -1293
rect 218891 -1411 218933 -1293
rect 219051 -1411 219067 -1293
rect 218757 -1907 219067 -1411
rect 220617 347447 220927 354061
rect 220617 347329 220633 347447
rect 220751 347329 220793 347447
rect 220911 347329 220927 347447
rect 220617 347287 220927 347329
rect 220617 347169 220633 347287
rect 220751 347169 220793 347287
rect 220911 347169 220927 347287
rect 220617 329447 220927 347169
rect 220617 329329 220633 329447
rect 220751 329329 220793 329447
rect 220911 329329 220927 329447
rect 220617 329287 220927 329329
rect 220617 329169 220633 329287
rect 220751 329169 220793 329287
rect 220911 329169 220927 329287
rect 220617 311447 220927 329169
rect 220617 311329 220633 311447
rect 220751 311329 220793 311447
rect 220911 311329 220927 311447
rect 220617 311287 220927 311329
rect 220617 311169 220633 311287
rect 220751 311169 220793 311287
rect 220911 311169 220927 311287
rect 220617 293447 220927 311169
rect 220617 293329 220633 293447
rect 220751 293329 220793 293447
rect 220911 293329 220927 293447
rect 220617 293287 220927 293329
rect 220617 293169 220633 293287
rect 220751 293169 220793 293287
rect 220911 293169 220927 293287
rect 220617 275447 220927 293169
rect 220617 275329 220633 275447
rect 220751 275329 220793 275447
rect 220911 275329 220927 275447
rect 220617 275287 220927 275329
rect 220617 275169 220633 275287
rect 220751 275169 220793 275287
rect 220911 275169 220927 275287
rect 220617 257447 220927 275169
rect 220617 257329 220633 257447
rect 220751 257329 220793 257447
rect 220911 257329 220927 257447
rect 220617 257287 220927 257329
rect 220617 257169 220633 257287
rect 220751 257169 220793 257287
rect 220911 257169 220927 257287
rect 220617 239447 220927 257169
rect 220617 239329 220633 239447
rect 220751 239329 220793 239447
rect 220911 239329 220927 239447
rect 220617 239287 220927 239329
rect 220617 239169 220633 239287
rect 220751 239169 220793 239287
rect 220911 239169 220927 239287
rect 220617 221447 220927 239169
rect 220617 221329 220633 221447
rect 220751 221329 220793 221447
rect 220911 221329 220927 221447
rect 220617 221287 220927 221329
rect 220617 221169 220633 221287
rect 220751 221169 220793 221287
rect 220911 221169 220927 221287
rect 220617 203447 220927 221169
rect 220617 203329 220633 203447
rect 220751 203329 220793 203447
rect 220911 203329 220927 203447
rect 220617 203287 220927 203329
rect 220617 203169 220633 203287
rect 220751 203169 220793 203287
rect 220911 203169 220927 203287
rect 220617 185447 220927 203169
rect 220617 185329 220633 185447
rect 220751 185329 220793 185447
rect 220911 185329 220927 185447
rect 220617 185287 220927 185329
rect 220617 185169 220633 185287
rect 220751 185169 220793 185287
rect 220911 185169 220927 185287
rect 220617 167447 220927 185169
rect 220617 167329 220633 167447
rect 220751 167329 220793 167447
rect 220911 167329 220927 167447
rect 220617 167287 220927 167329
rect 220617 167169 220633 167287
rect 220751 167169 220793 167287
rect 220911 167169 220927 167287
rect 220617 149447 220927 167169
rect 220617 149329 220633 149447
rect 220751 149329 220793 149447
rect 220911 149329 220927 149447
rect 220617 149287 220927 149329
rect 220617 149169 220633 149287
rect 220751 149169 220793 149287
rect 220911 149169 220927 149287
rect 220617 131447 220927 149169
rect 220617 131329 220633 131447
rect 220751 131329 220793 131447
rect 220911 131329 220927 131447
rect 220617 131287 220927 131329
rect 220617 131169 220633 131287
rect 220751 131169 220793 131287
rect 220911 131169 220927 131287
rect 220617 113447 220927 131169
rect 220617 113329 220633 113447
rect 220751 113329 220793 113447
rect 220911 113329 220927 113447
rect 220617 113287 220927 113329
rect 220617 113169 220633 113287
rect 220751 113169 220793 113287
rect 220911 113169 220927 113287
rect 220617 95447 220927 113169
rect 220617 95329 220633 95447
rect 220751 95329 220793 95447
rect 220911 95329 220927 95447
rect 220617 95287 220927 95329
rect 220617 95169 220633 95287
rect 220751 95169 220793 95287
rect 220911 95169 220927 95287
rect 220617 77447 220927 95169
rect 220617 77329 220633 77447
rect 220751 77329 220793 77447
rect 220911 77329 220927 77447
rect 220617 77287 220927 77329
rect 220617 77169 220633 77287
rect 220751 77169 220793 77287
rect 220911 77169 220927 77287
rect 220617 59447 220927 77169
rect 220617 59329 220633 59447
rect 220751 59329 220793 59447
rect 220911 59329 220927 59447
rect 220617 59287 220927 59329
rect 220617 59169 220633 59287
rect 220751 59169 220793 59287
rect 220911 59169 220927 59287
rect 220617 41447 220927 59169
rect 220617 41329 220633 41447
rect 220751 41329 220793 41447
rect 220911 41329 220927 41447
rect 220617 41287 220927 41329
rect 220617 41169 220633 41287
rect 220751 41169 220793 41287
rect 220911 41169 220927 41287
rect 220617 23447 220927 41169
rect 220617 23329 220633 23447
rect 220751 23329 220793 23447
rect 220911 23329 220927 23447
rect 220617 23287 220927 23329
rect 220617 23169 220633 23287
rect 220751 23169 220793 23287
rect 220911 23169 220927 23287
rect 220617 5447 220927 23169
rect 220617 5329 220633 5447
rect 220751 5329 220793 5447
rect 220911 5329 220927 5447
rect 220617 5287 220927 5329
rect 220617 5169 220633 5287
rect 220751 5169 220793 5287
rect 220911 5169 220927 5287
rect 220617 -2093 220927 5169
rect 220617 -2211 220633 -2093
rect 220751 -2211 220793 -2093
rect 220911 -2211 220927 -2093
rect 220617 -2253 220927 -2211
rect 220617 -2371 220633 -2253
rect 220751 -2371 220793 -2253
rect 220911 -2371 220927 -2253
rect 220617 -2867 220927 -2371
rect 222477 349307 222787 355021
rect 231477 355779 231787 355795
rect 231477 355661 231493 355779
rect 231611 355661 231653 355779
rect 231771 355661 231787 355779
rect 231477 355619 231787 355661
rect 231477 355501 231493 355619
rect 231611 355501 231653 355619
rect 231771 355501 231787 355619
rect 229617 354819 229927 354835
rect 229617 354701 229633 354819
rect 229751 354701 229793 354819
rect 229911 354701 229927 354819
rect 229617 354659 229927 354701
rect 229617 354541 229633 354659
rect 229751 354541 229793 354659
rect 229911 354541 229927 354659
rect 227757 353859 228067 353875
rect 227757 353741 227773 353859
rect 227891 353741 227933 353859
rect 228051 353741 228067 353859
rect 227757 353699 228067 353741
rect 227757 353581 227773 353699
rect 227891 353581 227933 353699
rect 228051 353581 228067 353699
rect 222477 349189 222493 349307
rect 222611 349189 222653 349307
rect 222771 349189 222787 349307
rect 222477 349147 222787 349189
rect 222477 349029 222493 349147
rect 222611 349029 222653 349147
rect 222771 349029 222787 349147
rect 222477 331307 222787 349029
rect 222477 331189 222493 331307
rect 222611 331189 222653 331307
rect 222771 331189 222787 331307
rect 222477 331147 222787 331189
rect 222477 331029 222493 331147
rect 222611 331029 222653 331147
rect 222771 331029 222787 331147
rect 222477 313307 222787 331029
rect 222477 313189 222493 313307
rect 222611 313189 222653 313307
rect 222771 313189 222787 313307
rect 222477 313147 222787 313189
rect 222477 313029 222493 313147
rect 222611 313029 222653 313147
rect 222771 313029 222787 313147
rect 222477 295307 222787 313029
rect 222477 295189 222493 295307
rect 222611 295189 222653 295307
rect 222771 295189 222787 295307
rect 222477 295147 222787 295189
rect 222477 295029 222493 295147
rect 222611 295029 222653 295147
rect 222771 295029 222787 295147
rect 222477 277307 222787 295029
rect 222477 277189 222493 277307
rect 222611 277189 222653 277307
rect 222771 277189 222787 277307
rect 222477 277147 222787 277189
rect 222477 277029 222493 277147
rect 222611 277029 222653 277147
rect 222771 277029 222787 277147
rect 222477 259307 222787 277029
rect 222477 259189 222493 259307
rect 222611 259189 222653 259307
rect 222771 259189 222787 259307
rect 222477 259147 222787 259189
rect 222477 259029 222493 259147
rect 222611 259029 222653 259147
rect 222771 259029 222787 259147
rect 222477 241307 222787 259029
rect 222477 241189 222493 241307
rect 222611 241189 222653 241307
rect 222771 241189 222787 241307
rect 222477 241147 222787 241189
rect 222477 241029 222493 241147
rect 222611 241029 222653 241147
rect 222771 241029 222787 241147
rect 222477 223307 222787 241029
rect 222477 223189 222493 223307
rect 222611 223189 222653 223307
rect 222771 223189 222787 223307
rect 222477 223147 222787 223189
rect 222477 223029 222493 223147
rect 222611 223029 222653 223147
rect 222771 223029 222787 223147
rect 222477 205307 222787 223029
rect 222477 205189 222493 205307
rect 222611 205189 222653 205307
rect 222771 205189 222787 205307
rect 222477 205147 222787 205189
rect 222477 205029 222493 205147
rect 222611 205029 222653 205147
rect 222771 205029 222787 205147
rect 222477 187307 222787 205029
rect 222477 187189 222493 187307
rect 222611 187189 222653 187307
rect 222771 187189 222787 187307
rect 222477 187147 222787 187189
rect 222477 187029 222493 187147
rect 222611 187029 222653 187147
rect 222771 187029 222787 187147
rect 222477 169307 222787 187029
rect 222477 169189 222493 169307
rect 222611 169189 222653 169307
rect 222771 169189 222787 169307
rect 222477 169147 222787 169189
rect 222477 169029 222493 169147
rect 222611 169029 222653 169147
rect 222771 169029 222787 169147
rect 222477 151307 222787 169029
rect 222477 151189 222493 151307
rect 222611 151189 222653 151307
rect 222771 151189 222787 151307
rect 222477 151147 222787 151189
rect 222477 151029 222493 151147
rect 222611 151029 222653 151147
rect 222771 151029 222787 151147
rect 222477 133307 222787 151029
rect 222477 133189 222493 133307
rect 222611 133189 222653 133307
rect 222771 133189 222787 133307
rect 222477 133147 222787 133189
rect 222477 133029 222493 133147
rect 222611 133029 222653 133147
rect 222771 133029 222787 133147
rect 222477 115307 222787 133029
rect 222477 115189 222493 115307
rect 222611 115189 222653 115307
rect 222771 115189 222787 115307
rect 222477 115147 222787 115189
rect 222477 115029 222493 115147
rect 222611 115029 222653 115147
rect 222771 115029 222787 115147
rect 222477 97307 222787 115029
rect 222477 97189 222493 97307
rect 222611 97189 222653 97307
rect 222771 97189 222787 97307
rect 222477 97147 222787 97189
rect 222477 97029 222493 97147
rect 222611 97029 222653 97147
rect 222771 97029 222787 97147
rect 222477 79307 222787 97029
rect 222477 79189 222493 79307
rect 222611 79189 222653 79307
rect 222771 79189 222787 79307
rect 222477 79147 222787 79189
rect 222477 79029 222493 79147
rect 222611 79029 222653 79147
rect 222771 79029 222787 79147
rect 222477 61307 222787 79029
rect 222477 61189 222493 61307
rect 222611 61189 222653 61307
rect 222771 61189 222787 61307
rect 222477 61147 222787 61189
rect 222477 61029 222493 61147
rect 222611 61029 222653 61147
rect 222771 61029 222787 61147
rect 222477 43307 222787 61029
rect 222477 43189 222493 43307
rect 222611 43189 222653 43307
rect 222771 43189 222787 43307
rect 222477 43147 222787 43189
rect 222477 43029 222493 43147
rect 222611 43029 222653 43147
rect 222771 43029 222787 43147
rect 222477 25307 222787 43029
rect 222477 25189 222493 25307
rect 222611 25189 222653 25307
rect 222771 25189 222787 25307
rect 222477 25147 222787 25189
rect 222477 25029 222493 25147
rect 222611 25029 222653 25147
rect 222771 25029 222787 25147
rect 222477 7307 222787 25029
rect 222477 7189 222493 7307
rect 222611 7189 222653 7307
rect 222771 7189 222787 7307
rect 222477 7147 222787 7189
rect 222477 7029 222493 7147
rect 222611 7029 222653 7147
rect 222771 7029 222787 7147
rect 213477 -3651 213493 -3533
rect 213611 -3651 213653 -3533
rect 213771 -3651 213787 -3533
rect 213477 -3693 213787 -3651
rect 213477 -3811 213493 -3693
rect 213611 -3811 213653 -3693
rect 213771 -3811 213787 -3693
rect 213477 -3827 213787 -3811
rect 222477 -3053 222787 7029
rect 225897 352899 226207 352915
rect 225897 352781 225913 352899
rect 226031 352781 226073 352899
rect 226191 352781 226207 352899
rect 225897 352739 226207 352781
rect 225897 352621 225913 352739
rect 226031 352621 226073 352739
rect 226191 352621 226207 352739
rect 225897 334727 226207 352621
rect 225897 334609 225913 334727
rect 226031 334609 226073 334727
rect 226191 334609 226207 334727
rect 225897 334567 226207 334609
rect 225897 334449 225913 334567
rect 226031 334449 226073 334567
rect 226191 334449 226207 334567
rect 225897 316727 226207 334449
rect 225897 316609 225913 316727
rect 226031 316609 226073 316727
rect 226191 316609 226207 316727
rect 225897 316567 226207 316609
rect 225897 316449 225913 316567
rect 226031 316449 226073 316567
rect 226191 316449 226207 316567
rect 225897 298727 226207 316449
rect 225897 298609 225913 298727
rect 226031 298609 226073 298727
rect 226191 298609 226207 298727
rect 225897 298567 226207 298609
rect 225897 298449 225913 298567
rect 226031 298449 226073 298567
rect 226191 298449 226207 298567
rect 225897 280727 226207 298449
rect 225897 280609 225913 280727
rect 226031 280609 226073 280727
rect 226191 280609 226207 280727
rect 225897 280567 226207 280609
rect 225897 280449 225913 280567
rect 226031 280449 226073 280567
rect 226191 280449 226207 280567
rect 225897 262727 226207 280449
rect 225897 262609 225913 262727
rect 226031 262609 226073 262727
rect 226191 262609 226207 262727
rect 225897 262567 226207 262609
rect 225897 262449 225913 262567
rect 226031 262449 226073 262567
rect 226191 262449 226207 262567
rect 225897 244727 226207 262449
rect 225897 244609 225913 244727
rect 226031 244609 226073 244727
rect 226191 244609 226207 244727
rect 225897 244567 226207 244609
rect 225897 244449 225913 244567
rect 226031 244449 226073 244567
rect 226191 244449 226207 244567
rect 225897 226727 226207 244449
rect 225897 226609 225913 226727
rect 226031 226609 226073 226727
rect 226191 226609 226207 226727
rect 225897 226567 226207 226609
rect 225897 226449 225913 226567
rect 226031 226449 226073 226567
rect 226191 226449 226207 226567
rect 225897 208727 226207 226449
rect 225897 208609 225913 208727
rect 226031 208609 226073 208727
rect 226191 208609 226207 208727
rect 225897 208567 226207 208609
rect 225897 208449 225913 208567
rect 226031 208449 226073 208567
rect 226191 208449 226207 208567
rect 225897 190727 226207 208449
rect 225897 190609 225913 190727
rect 226031 190609 226073 190727
rect 226191 190609 226207 190727
rect 225897 190567 226207 190609
rect 225897 190449 225913 190567
rect 226031 190449 226073 190567
rect 226191 190449 226207 190567
rect 225897 172727 226207 190449
rect 225897 172609 225913 172727
rect 226031 172609 226073 172727
rect 226191 172609 226207 172727
rect 225897 172567 226207 172609
rect 225897 172449 225913 172567
rect 226031 172449 226073 172567
rect 226191 172449 226207 172567
rect 225897 154727 226207 172449
rect 225897 154609 225913 154727
rect 226031 154609 226073 154727
rect 226191 154609 226207 154727
rect 225897 154567 226207 154609
rect 225897 154449 225913 154567
rect 226031 154449 226073 154567
rect 226191 154449 226207 154567
rect 225897 136727 226207 154449
rect 225897 136609 225913 136727
rect 226031 136609 226073 136727
rect 226191 136609 226207 136727
rect 225897 136567 226207 136609
rect 225897 136449 225913 136567
rect 226031 136449 226073 136567
rect 226191 136449 226207 136567
rect 225897 118727 226207 136449
rect 225897 118609 225913 118727
rect 226031 118609 226073 118727
rect 226191 118609 226207 118727
rect 225897 118567 226207 118609
rect 225897 118449 225913 118567
rect 226031 118449 226073 118567
rect 226191 118449 226207 118567
rect 225897 100727 226207 118449
rect 225897 100609 225913 100727
rect 226031 100609 226073 100727
rect 226191 100609 226207 100727
rect 225897 100567 226207 100609
rect 225897 100449 225913 100567
rect 226031 100449 226073 100567
rect 226191 100449 226207 100567
rect 225897 82727 226207 100449
rect 225897 82609 225913 82727
rect 226031 82609 226073 82727
rect 226191 82609 226207 82727
rect 225897 82567 226207 82609
rect 225897 82449 225913 82567
rect 226031 82449 226073 82567
rect 226191 82449 226207 82567
rect 225897 64727 226207 82449
rect 225897 64609 225913 64727
rect 226031 64609 226073 64727
rect 226191 64609 226207 64727
rect 225897 64567 226207 64609
rect 225897 64449 225913 64567
rect 226031 64449 226073 64567
rect 226191 64449 226207 64567
rect 225897 46727 226207 64449
rect 225897 46609 225913 46727
rect 226031 46609 226073 46727
rect 226191 46609 226207 46727
rect 225897 46567 226207 46609
rect 225897 46449 225913 46567
rect 226031 46449 226073 46567
rect 226191 46449 226207 46567
rect 225897 28727 226207 46449
rect 225897 28609 225913 28727
rect 226031 28609 226073 28727
rect 226191 28609 226207 28727
rect 225897 28567 226207 28609
rect 225897 28449 225913 28567
rect 226031 28449 226073 28567
rect 226191 28449 226207 28567
rect 225897 10727 226207 28449
rect 225897 10609 225913 10727
rect 226031 10609 226073 10727
rect 226191 10609 226207 10727
rect 225897 10567 226207 10609
rect 225897 10449 225913 10567
rect 226031 10449 226073 10567
rect 226191 10449 226207 10567
rect 225897 -653 226207 10449
rect 225897 -771 225913 -653
rect 226031 -771 226073 -653
rect 226191 -771 226207 -653
rect 225897 -813 226207 -771
rect 225897 -931 225913 -813
rect 226031 -931 226073 -813
rect 226191 -931 226207 -813
rect 225897 -947 226207 -931
rect 227757 336587 228067 353581
rect 227757 336469 227773 336587
rect 227891 336469 227933 336587
rect 228051 336469 228067 336587
rect 227757 336427 228067 336469
rect 227757 336309 227773 336427
rect 227891 336309 227933 336427
rect 228051 336309 228067 336427
rect 227757 318587 228067 336309
rect 227757 318469 227773 318587
rect 227891 318469 227933 318587
rect 228051 318469 228067 318587
rect 227757 318427 228067 318469
rect 227757 318309 227773 318427
rect 227891 318309 227933 318427
rect 228051 318309 228067 318427
rect 227757 300587 228067 318309
rect 227757 300469 227773 300587
rect 227891 300469 227933 300587
rect 228051 300469 228067 300587
rect 227757 300427 228067 300469
rect 227757 300309 227773 300427
rect 227891 300309 227933 300427
rect 228051 300309 228067 300427
rect 227757 282587 228067 300309
rect 227757 282469 227773 282587
rect 227891 282469 227933 282587
rect 228051 282469 228067 282587
rect 227757 282427 228067 282469
rect 227757 282309 227773 282427
rect 227891 282309 227933 282427
rect 228051 282309 228067 282427
rect 227757 264587 228067 282309
rect 227757 264469 227773 264587
rect 227891 264469 227933 264587
rect 228051 264469 228067 264587
rect 227757 264427 228067 264469
rect 227757 264309 227773 264427
rect 227891 264309 227933 264427
rect 228051 264309 228067 264427
rect 227757 246587 228067 264309
rect 227757 246469 227773 246587
rect 227891 246469 227933 246587
rect 228051 246469 228067 246587
rect 227757 246427 228067 246469
rect 227757 246309 227773 246427
rect 227891 246309 227933 246427
rect 228051 246309 228067 246427
rect 227757 228587 228067 246309
rect 227757 228469 227773 228587
rect 227891 228469 227933 228587
rect 228051 228469 228067 228587
rect 227757 228427 228067 228469
rect 227757 228309 227773 228427
rect 227891 228309 227933 228427
rect 228051 228309 228067 228427
rect 227757 210587 228067 228309
rect 227757 210469 227773 210587
rect 227891 210469 227933 210587
rect 228051 210469 228067 210587
rect 227757 210427 228067 210469
rect 227757 210309 227773 210427
rect 227891 210309 227933 210427
rect 228051 210309 228067 210427
rect 227757 192587 228067 210309
rect 227757 192469 227773 192587
rect 227891 192469 227933 192587
rect 228051 192469 228067 192587
rect 227757 192427 228067 192469
rect 227757 192309 227773 192427
rect 227891 192309 227933 192427
rect 228051 192309 228067 192427
rect 227757 174587 228067 192309
rect 227757 174469 227773 174587
rect 227891 174469 227933 174587
rect 228051 174469 228067 174587
rect 227757 174427 228067 174469
rect 227757 174309 227773 174427
rect 227891 174309 227933 174427
rect 228051 174309 228067 174427
rect 227757 156587 228067 174309
rect 227757 156469 227773 156587
rect 227891 156469 227933 156587
rect 228051 156469 228067 156587
rect 227757 156427 228067 156469
rect 227757 156309 227773 156427
rect 227891 156309 227933 156427
rect 228051 156309 228067 156427
rect 227757 138587 228067 156309
rect 227757 138469 227773 138587
rect 227891 138469 227933 138587
rect 228051 138469 228067 138587
rect 227757 138427 228067 138469
rect 227757 138309 227773 138427
rect 227891 138309 227933 138427
rect 228051 138309 228067 138427
rect 227757 120587 228067 138309
rect 227757 120469 227773 120587
rect 227891 120469 227933 120587
rect 228051 120469 228067 120587
rect 227757 120427 228067 120469
rect 227757 120309 227773 120427
rect 227891 120309 227933 120427
rect 228051 120309 228067 120427
rect 227757 102587 228067 120309
rect 227757 102469 227773 102587
rect 227891 102469 227933 102587
rect 228051 102469 228067 102587
rect 227757 102427 228067 102469
rect 227757 102309 227773 102427
rect 227891 102309 227933 102427
rect 228051 102309 228067 102427
rect 227757 84587 228067 102309
rect 227757 84469 227773 84587
rect 227891 84469 227933 84587
rect 228051 84469 228067 84587
rect 227757 84427 228067 84469
rect 227757 84309 227773 84427
rect 227891 84309 227933 84427
rect 228051 84309 228067 84427
rect 227757 66587 228067 84309
rect 227757 66469 227773 66587
rect 227891 66469 227933 66587
rect 228051 66469 228067 66587
rect 227757 66427 228067 66469
rect 227757 66309 227773 66427
rect 227891 66309 227933 66427
rect 228051 66309 228067 66427
rect 227757 48587 228067 66309
rect 227757 48469 227773 48587
rect 227891 48469 227933 48587
rect 228051 48469 228067 48587
rect 227757 48427 228067 48469
rect 227757 48309 227773 48427
rect 227891 48309 227933 48427
rect 228051 48309 228067 48427
rect 227757 30587 228067 48309
rect 227757 30469 227773 30587
rect 227891 30469 227933 30587
rect 228051 30469 228067 30587
rect 227757 30427 228067 30469
rect 227757 30309 227773 30427
rect 227891 30309 227933 30427
rect 228051 30309 228067 30427
rect 227757 12587 228067 30309
rect 227757 12469 227773 12587
rect 227891 12469 227933 12587
rect 228051 12469 228067 12587
rect 227757 12427 228067 12469
rect 227757 12309 227773 12427
rect 227891 12309 227933 12427
rect 228051 12309 228067 12427
rect 227757 -1613 228067 12309
rect 227757 -1731 227773 -1613
rect 227891 -1731 227933 -1613
rect 228051 -1731 228067 -1613
rect 227757 -1773 228067 -1731
rect 227757 -1891 227773 -1773
rect 227891 -1891 227933 -1773
rect 228051 -1891 228067 -1773
rect 227757 -1907 228067 -1891
rect 229617 338447 229927 354541
rect 229617 338329 229633 338447
rect 229751 338329 229793 338447
rect 229911 338329 229927 338447
rect 229617 338287 229927 338329
rect 229617 338169 229633 338287
rect 229751 338169 229793 338287
rect 229911 338169 229927 338287
rect 229617 320447 229927 338169
rect 229617 320329 229633 320447
rect 229751 320329 229793 320447
rect 229911 320329 229927 320447
rect 229617 320287 229927 320329
rect 229617 320169 229633 320287
rect 229751 320169 229793 320287
rect 229911 320169 229927 320287
rect 229617 302447 229927 320169
rect 229617 302329 229633 302447
rect 229751 302329 229793 302447
rect 229911 302329 229927 302447
rect 229617 302287 229927 302329
rect 229617 302169 229633 302287
rect 229751 302169 229793 302287
rect 229911 302169 229927 302287
rect 229617 284447 229927 302169
rect 229617 284329 229633 284447
rect 229751 284329 229793 284447
rect 229911 284329 229927 284447
rect 229617 284287 229927 284329
rect 229617 284169 229633 284287
rect 229751 284169 229793 284287
rect 229911 284169 229927 284287
rect 229617 266447 229927 284169
rect 229617 266329 229633 266447
rect 229751 266329 229793 266447
rect 229911 266329 229927 266447
rect 229617 266287 229927 266329
rect 229617 266169 229633 266287
rect 229751 266169 229793 266287
rect 229911 266169 229927 266287
rect 229617 248447 229927 266169
rect 229617 248329 229633 248447
rect 229751 248329 229793 248447
rect 229911 248329 229927 248447
rect 229617 248287 229927 248329
rect 229617 248169 229633 248287
rect 229751 248169 229793 248287
rect 229911 248169 229927 248287
rect 229617 230447 229927 248169
rect 229617 230329 229633 230447
rect 229751 230329 229793 230447
rect 229911 230329 229927 230447
rect 229617 230287 229927 230329
rect 229617 230169 229633 230287
rect 229751 230169 229793 230287
rect 229911 230169 229927 230287
rect 229617 212447 229927 230169
rect 229617 212329 229633 212447
rect 229751 212329 229793 212447
rect 229911 212329 229927 212447
rect 229617 212287 229927 212329
rect 229617 212169 229633 212287
rect 229751 212169 229793 212287
rect 229911 212169 229927 212287
rect 229617 194447 229927 212169
rect 229617 194329 229633 194447
rect 229751 194329 229793 194447
rect 229911 194329 229927 194447
rect 229617 194287 229927 194329
rect 229617 194169 229633 194287
rect 229751 194169 229793 194287
rect 229911 194169 229927 194287
rect 229617 176447 229927 194169
rect 229617 176329 229633 176447
rect 229751 176329 229793 176447
rect 229911 176329 229927 176447
rect 229617 176287 229927 176329
rect 229617 176169 229633 176287
rect 229751 176169 229793 176287
rect 229911 176169 229927 176287
rect 229617 158447 229927 176169
rect 229617 158329 229633 158447
rect 229751 158329 229793 158447
rect 229911 158329 229927 158447
rect 229617 158287 229927 158329
rect 229617 158169 229633 158287
rect 229751 158169 229793 158287
rect 229911 158169 229927 158287
rect 229617 140447 229927 158169
rect 229617 140329 229633 140447
rect 229751 140329 229793 140447
rect 229911 140329 229927 140447
rect 229617 140287 229927 140329
rect 229617 140169 229633 140287
rect 229751 140169 229793 140287
rect 229911 140169 229927 140287
rect 229617 122447 229927 140169
rect 229617 122329 229633 122447
rect 229751 122329 229793 122447
rect 229911 122329 229927 122447
rect 229617 122287 229927 122329
rect 229617 122169 229633 122287
rect 229751 122169 229793 122287
rect 229911 122169 229927 122287
rect 229617 104447 229927 122169
rect 229617 104329 229633 104447
rect 229751 104329 229793 104447
rect 229911 104329 229927 104447
rect 229617 104287 229927 104329
rect 229617 104169 229633 104287
rect 229751 104169 229793 104287
rect 229911 104169 229927 104287
rect 229617 86447 229927 104169
rect 229617 86329 229633 86447
rect 229751 86329 229793 86447
rect 229911 86329 229927 86447
rect 229617 86287 229927 86329
rect 229617 86169 229633 86287
rect 229751 86169 229793 86287
rect 229911 86169 229927 86287
rect 229617 68447 229927 86169
rect 229617 68329 229633 68447
rect 229751 68329 229793 68447
rect 229911 68329 229927 68447
rect 229617 68287 229927 68329
rect 229617 68169 229633 68287
rect 229751 68169 229793 68287
rect 229911 68169 229927 68287
rect 229617 50447 229927 68169
rect 229617 50329 229633 50447
rect 229751 50329 229793 50447
rect 229911 50329 229927 50447
rect 229617 50287 229927 50329
rect 229617 50169 229633 50287
rect 229751 50169 229793 50287
rect 229911 50169 229927 50287
rect 229617 32447 229927 50169
rect 229617 32329 229633 32447
rect 229751 32329 229793 32447
rect 229911 32329 229927 32447
rect 229617 32287 229927 32329
rect 229617 32169 229633 32287
rect 229751 32169 229793 32287
rect 229911 32169 229927 32287
rect 229617 14447 229927 32169
rect 229617 14329 229633 14447
rect 229751 14329 229793 14447
rect 229911 14329 229927 14447
rect 229617 14287 229927 14329
rect 229617 14169 229633 14287
rect 229751 14169 229793 14287
rect 229911 14169 229927 14287
rect 229617 -2573 229927 14169
rect 229617 -2691 229633 -2573
rect 229751 -2691 229793 -2573
rect 229911 -2691 229927 -2573
rect 229617 -2733 229927 -2691
rect 229617 -2851 229633 -2733
rect 229751 -2851 229793 -2733
rect 229911 -2851 229927 -2733
rect 229617 -2867 229927 -2851
rect 231477 340307 231787 355501
rect 240477 355299 240787 355795
rect 240477 355181 240493 355299
rect 240611 355181 240653 355299
rect 240771 355181 240787 355299
rect 240477 355139 240787 355181
rect 240477 355021 240493 355139
rect 240611 355021 240653 355139
rect 240771 355021 240787 355139
rect 238617 354339 238927 354835
rect 238617 354221 238633 354339
rect 238751 354221 238793 354339
rect 238911 354221 238927 354339
rect 238617 354179 238927 354221
rect 238617 354061 238633 354179
rect 238751 354061 238793 354179
rect 238911 354061 238927 354179
rect 236757 353379 237067 353875
rect 236757 353261 236773 353379
rect 236891 353261 236933 353379
rect 237051 353261 237067 353379
rect 236757 353219 237067 353261
rect 236757 353101 236773 353219
rect 236891 353101 236933 353219
rect 237051 353101 237067 353219
rect 231477 340189 231493 340307
rect 231611 340189 231653 340307
rect 231771 340189 231787 340307
rect 231477 340147 231787 340189
rect 231477 340029 231493 340147
rect 231611 340029 231653 340147
rect 231771 340029 231787 340147
rect 231477 322307 231787 340029
rect 231477 322189 231493 322307
rect 231611 322189 231653 322307
rect 231771 322189 231787 322307
rect 231477 322147 231787 322189
rect 231477 322029 231493 322147
rect 231611 322029 231653 322147
rect 231771 322029 231787 322147
rect 231477 304307 231787 322029
rect 231477 304189 231493 304307
rect 231611 304189 231653 304307
rect 231771 304189 231787 304307
rect 231477 304147 231787 304189
rect 231477 304029 231493 304147
rect 231611 304029 231653 304147
rect 231771 304029 231787 304147
rect 231477 286307 231787 304029
rect 231477 286189 231493 286307
rect 231611 286189 231653 286307
rect 231771 286189 231787 286307
rect 231477 286147 231787 286189
rect 231477 286029 231493 286147
rect 231611 286029 231653 286147
rect 231771 286029 231787 286147
rect 231477 268307 231787 286029
rect 231477 268189 231493 268307
rect 231611 268189 231653 268307
rect 231771 268189 231787 268307
rect 231477 268147 231787 268189
rect 231477 268029 231493 268147
rect 231611 268029 231653 268147
rect 231771 268029 231787 268147
rect 231477 250307 231787 268029
rect 231477 250189 231493 250307
rect 231611 250189 231653 250307
rect 231771 250189 231787 250307
rect 231477 250147 231787 250189
rect 231477 250029 231493 250147
rect 231611 250029 231653 250147
rect 231771 250029 231787 250147
rect 231477 232307 231787 250029
rect 231477 232189 231493 232307
rect 231611 232189 231653 232307
rect 231771 232189 231787 232307
rect 231477 232147 231787 232189
rect 231477 232029 231493 232147
rect 231611 232029 231653 232147
rect 231771 232029 231787 232147
rect 231477 214307 231787 232029
rect 231477 214189 231493 214307
rect 231611 214189 231653 214307
rect 231771 214189 231787 214307
rect 231477 214147 231787 214189
rect 231477 214029 231493 214147
rect 231611 214029 231653 214147
rect 231771 214029 231787 214147
rect 231477 196307 231787 214029
rect 231477 196189 231493 196307
rect 231611 196189 231653 196307
rect 231771 196189 231787 196307
rect 231477 196147 231787 196189
rect 231477 196029 231493 196147
rect 231611 196029 231653 196147
rect 231771 196029 231787 196147
rect 231477 178307 231787 196029
rect 231477 178189 231493 178307
rect 231611 178189 231653 178307
rect 231771 178189 231787 178307
rect 231477 178147 231787 178189
rect 231477 178029 231493 178147
rect 231611 178029 231653 178147
rect 231771 178029 231787 178147
rect 231477 160307 231787 178029
rect 231477 160189 231493 160307
rect 231611 160189 231653 160307
rect 231771 160189 231787 160307
rect 231477 160147 231787 160189
rect 231477 160029 231493 160147
rect 231611 160029 231653 160147
rect 231771 160029 231787 160147
rect 231477 142307 231787 160029
rect 231477 142189 231493 142307
rect 231611 142189 231653 142307
rect 231771 142189 231787 142307
rect 231477 142147 231787 142189
rect 231477 142029 231493 142147
rect 231611 142029 231653 142147
rect 231771 142029 231787 142147
rect 231477 124307 231787 142029
rect 231477 124189 231493 124307
rect 231611 124189 231653 124307
rect 231771 124189 231787 124307
rect 231477 124147 231787 124189
rect 231477 124029 231493 124147
rect 231611 124029 231653 124147
rect 231771 124029 231787 124147
rect 231477 106307 231787 124029
rect 231477 106189 231493 106307
rect 231611 106189 231653 106307
rect 231771 106189 231787 106307
rect 231477 106147 231787 106189
rect 231477 106029 231493 106147
rect 231611 106029 231653 106147
rect 231771 106029 231787 106147
rect 231477 88307 231787 106029
rect 231477 88189 231493 88307
rect 231611 88189 231653 88307
rect 231771 88189 231787 88307
rect 231477 88147 231787 88189
rect 231477 88029 231493 88147
rect 231611 88029 231653 88147
rect 231771 88029 231787 88147
rect 231477 70307 231787 88029
rect 231477 70189 231493 70307
rect 231611 70189 231653 70307
rect 231771 70189 231787 70307
rect 231477 70147 231787 70189
rect 231477 70029 231493 70147
rect 231611 70029 231653 70147
rect 231771 70029 231787 70147
rect 231477 52307 231787 70029
rect 231477 52189 231493 52307
rect 231611 52189 231653 52307
rect 231771 52189 231787 52307
rect 231477 52147 231787 52189
rect 231477 52029 231493 52147
rect 231611 52029 231653 52147
rect 231771 52029 231787 52147
rect 231477 34307 231787 52029
rect 231477 34189 231493 34307
rect 231611 34189 231653 34307
rect 231771 34189 231787 34307
rect 231477 34147 231787 34189
rect 231477 34029 231493 34147
rect 231611 34029 231653 34147
rect 231771 34029 231787 34147
rect 231477 16307 231787 34029
rect 231477 16189 231493 16307
rect 231611 16189 231653 16307
rect 231771 16189 231787 16307
rect 231477 16147 231787 16189
rect 231477 16029 231493 16147
rect 231611 16029 231653 16147
rect 231771 16029 231787 16147
rect 222477 -3171 222493 -3053
rect 222611 -3171 222653 -3053
rect 222771 -3171 222787 -3053
rect 222477 -3213 222787 -3171
rect 222477 -3331 222493 -3213
rect 222611 -3331 222653 -3213
rect 222771 -3331 222787 -3213
rect 222477 -3827 222787 -3331
rect 231477 -3533 231787 16029
rect 234897 352419 235207 352915
rect 234897 352301 234913 352419
rect 235031 352301 235073 352419
rect 235191 352301 235207 352419
rect 234897 352259 235207 352301
rect 234897 352141 234913 352259
rect 235031 352141 235073 352259
rect 235191 352141 235207 352259
rect 234897 343727 235207 352141
rect 234897 343609 234913 343727
rect 235031 343609 235073 343727
rect 235191 343609 235207 343727
rect 234897 343567 235207 343609
rect 234897 343449 234913 343567
rect 235031 343449 235073 343567
rect 235191 343449 235207 343567
rect 234897 325727 235207 343449
rect 234897 325609 234913 325727
rect 235031 325609 235073 325727
rect 235191 325609 235207 325727
rect 234897 325567 235207 325609
rect 234897 325449 234913 325567
rect 235031 325449 235073 325567
rect 235191 325449 235207 325567
rect 234897 307727 235207 325449
rect 234897 307609 234913 307727
rect 235031 307609 235073 307727
rect 235191 307609 235207 307727
rect 234897 307567 235207 307609
rect 234897 307449 234913 307567
rect 235031 307449 235073 307567
rect 235191 307449 235207 307567
rect 234897 289727 235207 307449
rect 234897 289609 234913 289727
rect 235031 289609 235073 289727
rect 235191 289609 235207 289727
rect 234897 289567 235207 289609
rect 234897 289449 234913 289567
rect 235031 289449 235073 289567
rect 235191 289449 235207 289567
rect 234897 271727 235207 289449
rect 234897 271609 234913 271727
rect 235031 271609 235073 271727
rect 235191 271609 235207 271727
rect 234897 271567 235207 271609
rect 234897 271449 234913 271567
rect 235031 271449 235073 271567
rect 235191 271449 235207 271567
rect 234897 253727 235207 271449
rect 234897 253609 234913 253727
rect 235031 253609 235073 253727
rect 235191 253609 235207 253727
rect 234897 253567 235207 253609
rect 234897 253449 234913 253567
rect 235031 253449 235073 253567
rect 235191 253449 235207 253567
rect 234897 235727 235207 253449
rect 234897 235609 234913 235727
rect 235031 235609 235073 235727
rect 235191 235609 235207 235727
rect 234897 235567 235207 235609
rect 234897 235449 234913 235567
rect 235031 235449 235073 235567
rect 235191 235449 235207 235567
rect 234897 217727 235207 235449
rect 234897 217609 234913 217727
rect 235031 217609 235073 217727
rect 235191 217609 235207 217727
rect 234897 217567 235207 217609
rect 234897 217449 234913 217567
rect 235031 217449 235073 217567
rect 235191 217449 235207 217567
rect 234897 199727 235207 217449
rect 234897 199609 234913 199727
rect 235031 199609 235073 199727
rect 235191 199609 235207 199727
rect 234897 199567 235207 199609
rect 234897 199449 234913 199567
rect 235031 199449 235073 199567
rect 235191 199449 235207 199567
rect 234897 181727 235207 199449
rect 234897 181609 234913 181727
rect 235031 181609 235073 181727
rect 235191 181609 235207 181727
rect 234897 181567 235207 181609
rect 234897 181449 234913 181567
rect 235031 181449 235073 181567
rect 235191 181449 235207 181567
rect 234897 163727 235207 181449
rect 234897 163609 234913 163727
rect 235031 163609 235073 163727
rect 235191 163609 235207 163727
rect 234897 163567 235207 163609
rect 234897 163449 234913 163567
rect 235031 163449 235073 163567
rect 235191 163449 235207 163567
rect 234897 145727 235207 163449
rect 234897 145609 234913 145727
rect 235031 145609 235073 145727
rect 235191 145609 235207 145727
rect 234897 145567 235207 145609
rect 234897 145449 234913 145567
rect 235031 145449 235073 145567
rect 235191 145449 235207 145567
rect 234897 127727 235207 145449
rect 234897 127609 234913 127727
rect 235031 127609 235073 127727
rect 235191 127609 235207 127727
rect 234897 127567 235207 127609
rect 234897 127449 234913 127567
rect 235031 127449 235073 127567
rect 235191 127449 235207 127567
rect 234897 109727 235207 127449
rect 234897 109609 234913 109727
rect 235031 109609 235073 109727
rect 235191 109609 235207 109727
rect 234897 109567 235207 109609
rect 234897 109449 234913 109567
rect 235031 109449 235073 109567
rect 235191 109449 235207 109567
rect 234897 91727 235207 109449
rect 234897 91609 234913 91727
rect 235031 91609 235073 91727
rect 235191 91609 235207 91727
rect 234897 91567 235207 91609
rect 234897 91449 234913 91567
rect 235031 91449 235073 91567
rect 235191 91449 235207 91567
rect 234897 73727 235207 91449
rect 234897 73609 234913 73727
rect 235031 73609 235073 73727
rect 235191 73609 235207 73727
rect 234897 73567 235207 73609
rect 234897 73449 234913 73567
rect 235031 73449 235073 73567
rect 235191 73449 235207 73567
rect 234897 55727 235207 73449
rect 234897 55609 234913 55727
rect 235031 55609 235073 55727
rect 235191 55609 235207 55727
rect 234897 55567 235207 55609
rect 234897 55449 234913 55567
rect 235031 55449 235073 55567
rect 235191 55449 235207 55567
rect 234897 37727 235207 55449
rect 234897 37609 234913 37727
rect 235031 37609 235073 37727
rect 235191 37609 235207 37727
rect 234897 37567 235207 37609
rect 234897 37449 234913 37567
rect 235031 37449 235073 37567
rect 235191 37449 235207 37567
rect 234897 19727 235207 37449
rect 234897 19609 234913 19727
rect 235031 19609 235073 19727
rect 235191 19609 235207 19727
rect 234897 19567 235207 19609
rect 234897 19449 234913 19567
rect 235031 19449 235073 19567
rect 235191 19449 235207 19567
rect 234897 1727 235207 19449
rect 234897 1609 234913 1727
rect 235031 1609 235073 1727
rect 235191 1609 235207 1727
rect 234897 1567 235207 1609
rect 234897 1449 234913 1567
rect 235031 1449 235073 1567
rect 235191 1449 235207 1567
rect 234897 -173 235207 1449
rect 234897 -291 234913 -173
rect 235031 -291 235073 -173
rect 235191 -291 235207 -173
rect 234897 -333 235207 -291
rect 234897 -451 234913 -333
rect 235031 -451 235073 -333
rect 235191 -451 235207 -333
rect 234897 -947 235207 -451
rect 236757 345587 237067 353101
rect 236757 345469 236773 345587
rect 236891 345469 236933 345587
rect 237051 345469 237067 345587
rect 236757 345427 237067 345469
rect 236757 345309 236773 345427
rect 236891 345309 236933 345427
rect 237051 345309 237067 345427
rect 236757 327587 237067 345309
rect 236757 327469 236773 327587
rect 236891 327469 236933 327587
rect 237051 327469 237067 327587
rect 236757 327427 237067 327469
rect 236757 327309 236773 327427
rect 236891 327309 236933 327427
rect 237051 327309 237067 327427
rect 236757 309587 237067 327309
rect 236757 309469 236773 309587
rect 236891 309469 236933 309587
rect 237051 309469 237067 309587
rect 236757 309427 237067 309469
rect 236757 309309 236773 309427
rect 236891 309309 236933 309427
rect 237051 309309 237067 309427
rect 236757 291587 237067 309309
rect 236757 291469 236773 291587
rect 236891 291469 236933 291587
rect 237051 291469 237067 291587
rect 236757 291427 237067 291469
rect 236757 291309 236773 291427
rect 236891 291309 236933 291427
rect 237051 291309 237067 291427
rect 236757 273587 237067 291309
rect 236757 273469 236773 273587
rect 236891 273469 236933 273587
rect 237051 273469 237067 273587
rect 236757 273427 237067 273469
rect 236757 273309 236773 273427
rect 236891 273309 236933 273427
rect 237051 273309 237067 273427
rect 236757 255587 237067 273309
rect 236757 255469 236773 255587
rect 236891 255469 236933 255587
rect 237051 255469 237067 255587
rect 236757 255427 237067 255469
rect 236757 255309 236773 255427
rect 236891 255309 236933 255427
rect 237051 255309 237067 255427
rect 236757 237587 237067 255309
rect 236757 237469 236773 237587
rect 236891 237469 236933 237587
rect 237051 237469 237067 237587
rect 236757 237427 237067 237469
rect 236757 237309 236773 237427
rect 236891 237309 236933 237427
rect 237051 237309 237067 237427
rect 236757 219587 237067 237309
rect 236757 219469 236773 219587
rect 236891 219469 236933 219587
rect 237051 219469 237067 219587
rect 236757 219427 237067 219469
rect 236757 219309 236773 219427
rect 236891 219309 236933 219427
rect 237051 219309 237067 219427
rect 236757 201587 237067 219309
rect 236757 201469 236773 201587
rect 236891 201469 236933 201587
rect 237051 201469 237067 201587
rect 236757 201427 237067 201469
rect 236757 201309 236773 201427
rect 236891 201309 236933 201427
rect 237051 201309 237067 201427
rect 236757 183587 237067 201309
rect 236757 183469 236773 183587
rect 236891 183469 236933 183587
rect 237051 183469 237067 183587
rect 236757 183427 237067 183469
rect 236757 183309 236773 183427
rect 236891 183309 236933 183427
rect 237051 183309 237067 183427
rect 236757 165587 237067 183309
rect 236757 165469 236773 165587
rect 236891 165469 236933 165587
rect 237051 165469 237067 165587
rect 236757 165427 237067 165469
rect 236757 165309 236773 165427
rect 236891 165309 236933 165427
rect 237051 165309 237067 165427
rect 236757 147587 237067 165309
rect 236757 147469 236773 147587
rect 236891 147469 236933 147587
rect 237051 147469 237067 147587
rect 236757 147427 237067 147469
rect 236757 147309 236773 147427
rect 236891 147309 236933 147427
rect 237051 147309 237067 147427
rect 236757 129587 237067 147309
rect 236757 129469 236773 129587
rect 236891 129469 236933 129587
rect 237051 129469 237067 129587
rect 236757 129427 237067 129469
rect 236757 129309 236773 129427
rect 236891 129309 236933 129427
rect 237051 129309 237067 129427
rect 236757 111587 237067 129309
rect 236757 111469 236773 111587
rect 236891 111469 236933 111587
rect 237051 111469 237067 111587
rect 236757 111427 237067 111469
rect 236757 111309 236773 111427
rect 236891 111309 236933 111427
rect 237051 111309 237067 111427
rect 236757 93587 237067 111309
rect 236757 93469 236773 93587
rect 236891 93469 236933 93587
rect 237051 93469 237067 93587
rect 236757 93427 237067 93469
rect 236757 93309 236773 93427
rect 236891 93309 236933 93427
rect 237051 93309 237067 93427
rect 236757 75587 237067 93309
rect 236757 75469 236773 75587
rect 236891 75469 236933 75587
rect 237051 75469 237067 75587
rect 236757 75427 237067 75469
rect 236757 75309 236773 75427
rect 236891 75309 236933 75427
rect 237051 75309 237067 75427
rect 236757 57587 237067 75309
rect 236757 57469 236773 57587
rect 236891 57469 236933 57587
rect 237051 57469 237067 57587
rect 236757 57427 237067 57469
rect 236757 57309 236773 57427
rect 236891 57309 236933 57427
rect 237051 57309 237067 57427
rect 236757 39587 237067 57309
rect 236757 39469 236773 39587
rect 236891 39469 236933 39587
rect 237051 39469 237067 39587
rect 236757 39427 237067 39469
rect 236757 39309 236773 39427
rect 236891 39309 236933 39427
rect 237051 39309 237067 39427
rect 236757 21587 237067 39309
rect 236757 21469 236773 21587
rect 236891 21469 236933 21587
rect 237051 21469 237067 21587
rect 236757 21427 237067 21469
rect 236757 21309 236773 21427
rect 236891 21309 236933 21427
rect 237051 21309 237067 21427
rect 236757 3587 237067 21309
rect 236757 3469 236773 3587
rect 236891 3469 236933 3587
rect 237051 3469 237067 3587
rect 236757 3427 237067 3469
rect 236757 3309 236773 3427
rect 236891 3309 236933 3427
rect 237051 3309 237067 3427
rect 236757 -1133 237067 3309
rect 236757 -1251 236773 -1133
rect 236891 -1251 236933 -1133
rect 237051 -1251 237067 -1133
rect 236757 -1293 237067 -1251
rect 236757 -1411 236773 -1293
rect 236891 -1411 236933 -1293
rect 237051 -1411 237067 -1293
rect 236757 -1907 237067 -1411
rect 238617 347447 238927 354061
rect 238617 347329 238633 347447
rect 238751 347329 238793 347447
rect 238911 347329 238927 347447
rect 238617 347287 238927 347329
rect 238617 347169 238633 347287
rect 238751 347169 238793 347287
rect 238911 347169 238927 347287
rect 238617 329447 238927 347169
rect 238617 329329 238633 329447
rect 238751 329329 238793 329447
rect 238911 329329 238927 329447
rect 238617 329287 238927 329329
rect 238617 329169 238633 329287
rect 238751 329169 238793 329287
rect 238911 329169 238927 329287
rect 238617 311447 238927 329169
rect 238617 311329 238633 311447
rect 238751 311329 238793 311447
rect 238911 311329 238927 311447
rect 238617 311287 238927 311329
rect 238617 311169 238633 311287
rect 238751 311169 238793 311287
rect 238911 311169 238927 311287
rect 238617 293447 238927 311169
rect 238617 293329 238633 293447
rect 238751 293329 238793 293447
rect 238911 293329 238927 293447
rect 238617 293287 238927 293329
rect 238617 293169 238633 293287
rect 238751 293169 238793 293287
rect 238911 293169 238927 293287
rect 238617 275447 238927 293169
rect 238617 275329 238633 275447
rect 238751 275329 238793 275447
rect 238911 275329 238927 275447
rect 238617 275287 238927 275329
rect 238617 275169 238633 275287
rect 238751 275169 238793 275287
rect 238911 275169 238927 275287
rect 238617 257447 238927 275169
rect 238617 257329 238633 257447
rect 238751 257329 238793 257447
rect 238911 257329 238927 257447
rect 238617 257287 238927 257329
rect 238617 257169 238633 257287
rect 238751 257169 238793 257287
rect 238911 257169 238927 257287
rect 238617 239447 238927 257169
rect 238617 239329 238633 239447
rect 238751 239329 238793 239447
rect 238911 239329 238927 239447
rect 238617 239287 238927 239329
rect 238617 239169 238633 239287
rect 238751 239169 238793 239287
rect 238911 239169 238927 239287
rect 238617 221447 238927 239169
rect 238617 221329 238633 221447
rect 238751 221329 238793 221447
rect 238911 221329 238927 221447
rect 238617 221287 238927 221329
rect 238617 221169 238633 221287
rect 238751 221169 238793 221287
rect 238911 221169 238927 221287
rect 238617 203447 238927 221169
rect 238617 203329 238633 203447
rect 238751 203329 238793 203447
rect 238911 203329 238927 203447
rect 238617 203287 238927 203329
rect 238617 203169 238633 203287
rect 238751 203169 238793 203287
rect 238911 203169 238927 203287
rect 238617 185447 238927 203169
rect 238617 185329 238633 185447
rect 238751 185329 238793 185447
rect 238911 185329 238927 185447
rect 238617 185287 238927 185329
rect 238617 185169 238633 185287
rect 238751 185169 238793 185287
rect 238911 185169 238927 185287
rect 238617 167447 238927 185169
rect 238617 167329 238633 167447
rect 238751 167329 238793 167447
rect 238911 167329 238927 167447
rect 238617 167287 238927 167329
rect 238617 167169 238633 167287
rect 238751 167169 238793 167287
rect 238911 167169 238927 167287
rect 238617 149447 238927 167169
rect 238617 149329 238633 149447
rect 238751 149329 238793 149447
rect 238911 149329 238927 149447
rect 238617 149287 238927 149329
rect 238617 149169 238633 149287
rect 238751 149169 238793 149287
rect 238911 149169 238927 149287
rect 238617 131447 238927 149169
rect 238617 131329 238633 131447
rect 238751 131329 238793 131447
rect 238911 131329 238927 131447
rect 238617 131287 238927 131329
rect 238617 131169 238633 131287
rect 238751 131169 238793 131287
rect 238911 131169 238927 131287
rect 238617 113447 238927 131169
rect 238617 113329 238633 113447
rect 238751 113329 238793 113447
rect 238911 113329 238927 113447
rect 238617 113287 238927 113329
rect 238617 113169 238633 113287
rect 238751 113169 238793 113287
rect 238911 113169 238927 113287
rect 238617 95447 238927 113169
rect 238617 95329 238633 95447
rect 238751 95329 238793 95447
rect 238911 95329 238927 95447
rect 238617 95287 238927 95329
rect 238617 95169 238633 95287
rect 238751 95169 238793 95287
rect 238911 95169 238927 95287
rect 238617 77447 238927 95169
rect 238617 77329 238633 77447
rect 238751 77329 238793 77447
rect 238911 77329 238927 77447
rect 238617 77287 238927 77329
rect 238617 77169 238633 77287
rect 238751 77169 238793 77287
rect 238911 77169 238927 77287
rect 238617 59447 238927 77169
rect 238617 59329 238633 59447
rect 238751 59329 238793 59447
rect 238911 59329 238927 59447
rect 238617 59287 238927 59329
rect 238617 59169 238633 59287
rect 238751 59169 238793 59287
rect 238911 59169 238927 59287
rect 238617 41447 238927 59169
rect 238617 41329 238633 41447
rect 238751 41329 238793 41447
rect 238911 41329 238927 41447
rect 238617 41287 238927 41329
rect 238617 41169 238633 41287
rect 238751 41169 238793 41287
rect 238911 41169 238927 41287
rect 238617 23447 238927 41169
rect 238617 23329 238633 23447
rect 238751 23329 238793 23447
rect 238911 23329 238927 23447
rect 238617 23287 238927 23329
rect 238617 23169 238633 23287
rect 238751 23169 238793 23287
rect 238911 23169 238927 23287
rect 238617 5447 238927 23169
rect 238617 5329 238633 5447
rect 238751 5329 238793 5447
rect 238911 5329 238927 5447
rect 238617 5287 238927 5329
rect 238617 5169 238633 5287
rect 238751 5169 238793 5287
rect 238911 5169 238927 5287
rect 238617 -2093 238927 5169
rect 238617 -2211 238633 -2093
rect 238751 -2211 238793 -2093
rect 238911 -2211 238927 -2093
rect 238617 -2253 238927 -2211
rect 238617 -2371 238633 -2253
rect 238751 -2371 238793 -2253
rect 238911 -2371 238927 -2253
rect 238617 -2867 238927 -2371
rect 240477 349307 240787 355021
rect 249477 355779 249787 355795
rect 249477 355661 249493 355779
rect 249611 355661 249653 355779
rect 249771 355661 249787 355779
rect 249477 355619 249787 355661
rect 249477 355501 249493 355619
rect 249611 355501 249653 355619
rect 249771 355501 249787 355619
rect 247617 354819 247927 354835
rect 247617 354701 247633 354819
rect 247751 354701 247793 354819
rect 247911 354701 247927 354819
rect 247617 354659 247927 354701
rect 247617 354541 247633 354659
rect 247751 354541 247793 354659
rect 247911 354541 247927 354659
rect 245757 353859 246067 353875
rect 245757 353741 245773 353859
rect 245891 353741 245933 353859
rect 246051 353741 246067 353859
rect 245757 353699 246067 353741
rect 245757 353581 245773 353699
rect 245891 353581 245933 353699
rect 246051 353581 246067 353699
rect 240477 349189 240493 349307
rect 240611 349189 240653 349307
rect 240771 349189 240787 349307
rect 240477 349147 240787 349189
rect 240477 349029 240493 349147
rect 240611 349029 240653 349147
rect 240771 349029 240787 349147
rect 240477 331307 240787 349029
rect 240477 331189 240493 331307
rect 240611 331189 240653 331307
rect 240771 331189 240787 331307
rect 240477 331147 240787 331189
rect 240477 331029 240493 331147
rect 240611 331029 240653 331147
rect 240771 331029 240787 331147
rect 240477 313307 240787 331029
rect 240477 313189 240493 313307
rect 240611 313189 240653 313307
rect 240771 313189 240787 313307
rect 240477 313147 240787 313189
rect 240477 313029 240493 313147
rect 240611 313029 240653 313147
rect 240771 313029 240787 313147
rect 240477 295307 240787 313029
rect 240477 295189 240493 295307
rect 240611 295189 240653 295307
rect 240771 295189 240787 295307
rect 240477 295147 240787 295189
rect 240477 295029 240493 295147
rect 240611 295029 240653 295147
rect 240771 295029 240787 295147
rect 240477 277307 240787 295029
rect 240477 277189 240493 277307
rect 240611 277189 240653 277307
rect 240771 277189 240787 277307
rect 240477 277147 240787 277189
rect 240477 277029 240493 277147
rect 240611 277029 240653 277147
rect 240771 277029 240787 277147
rect 240477 259307 240787 277029
rect 240477 259189 240493 259307
rect 240611 259189 240653 259307
rect 240771 259189 240787 259307
rect 240477 259147 240787 259189
rect 240477 259029 240493 259147
rect 240611 259029 240653 259147
rect 240771 259029 240787 259147
rect 240477 241307 240787 259029
rect 240477 241189 240493 241307
rect 240611 241189 240653 241307
rect 240771 241189 240787 241307
rect 240477 241147 240787 241189
rect 240477 241029 240493 241147
rect 240611 241029 240653 241147
rect 240771 241029 240787 241147
rect 240477 223307 240787 241029
rect 240477 223189 240493 223307
rect 240611 223189 240653 223307
rect 240771 223189 240787 223307
rect 240477 223147 240787 223189
rect 240477 223029 240493 223147
rect 240611 223029 240653 223147
rect 240771 223029 240787 223147
rect 240477 205307 240787 223029
rect 240477 205189 240493 205307
rect 240611 205189 240653 205307
rect 240771 205189 240787 205307
rect 240477 205147 240787 205189
rect 240477 205029 240493 205147
rect 240611 205029 240653 205147
rect 240771 205029 240787 205147
rect 240477 187307 240787 205029
rect 240477 187189 240493 187307
rect 240611 187189 240653 187307
rect 240771 187189 240787 187307
rect 240477 187147 240787 187189
rect 240477 187029 240493 187147
rect 240611 187029 240653 187147
rect 240771 187029 240787 187147
rect 240477 169307 240787 187029
rect 240477 169189 240493 169307
rect 240611 169189 240653 169307
rect 240771 169189 240787 169307
rect 240477 169147 240787 169189
rect 240477 169029 240493 169147
rect 240611 169029 240653 169147
rect 240771 169029 240787 169147
rect 240477 151307 240787 169029
rect 240477 151189 240493 151307
rect 240611 151189 240653 151307
rect 240771 151189 240787 151307
rect 240477 151147 240787 151189
rect 240477 151029 240493 151147
rect 240611 151029 240653 151147
rect 240771 151029 240787 151147
rect 240477 133307 240787 151029
rect 240477 133189 240493 133307
rect 240611 133189 240653 133307
rect 240771 133189 240787 133307
rect 240477 133147 240787 133189
rect 240477 133029 240493 133147
rect 240611 133029 240653 133147
rect 240771 133029 240787 133147
rect 240477 115307 240787 133029
rect 240477 115189 240493 115307
rect 240611 115189 240653 115307
rect 240771 115189 240787 115307
rect 240477 115147 240787 115189
rect 240477 115029 240493 115147
rect 240611 115029 240653 115147
rect 240771 115029 240787 115147
rect 240477 97307 240787 115029
rect 240477 97189 240493 97307
rect 240611 97189 240653 97307
rect 240771 97189 240787 97307
rect 240477 97147 240787 97189
rect 240477 97029 240493 97147
rect 240611 97029 240653 97147
rect 240771 97029 240787 97147
rect 240477 79307 240787 97029
rect 240477 79189 240493 79307
rect 240611 79189 240653 79307
rect 240771 79189 240787 79307
rect 240477 79147 240787 79189
rect 240477 79029 240493 79147
rect 240611 79029 240653 79147
rect 240771 79029 240787 79147
rect 240477 61307 240787 79029
rect 240477 61189 240493 61307
rect 240611 61189 240653 61307
rect 240771 61189 240787 61307
rect 240477 61147 240787 61189
rect 240477 61029 240493 61147
rect 240611 61029 240653 61147
rect 240771 61029 240787 61147
rect 240477 43307 240787 61029
rect 240477 43189 240493 43307
rect 240611 43189 240653 43307
rect 240771 43189 240787 43307
rect 240477 43147 240787 43189
rect 240477 43029 240493 43147
rect 240611 43029 240653 43147
rect 240771 43029 240787 43147
rect 240477 25307 240787 43029
rect 240477 25189 240493 25307
rect 240611 25189 240653 25307
rect 240771 25189 240787 25307
rect 240477 25147 240787 25189
rect 240477 25029 240493 25147
rect 240611 25029 240653 25147
rect 240771 25029 240787 25147
rect 240477 7307 240787 25029
rect 240477 7189 240493 7307
rect 240611 7189 240653 7307
rect 240771 7189 240787 7307
rect 240477 7147 240787 7189
rect 240477 7029 240493 7147
rect 240611 7029 240653 7147
rect 240771 7029 240787 7147
rect 231477 -3651 231493 -3533
rect 231611 -3651 231653 -3533
rect 231771 -3651 231787 -3533
rect 231477 -3693 231787 -3651
rect 231477 -3811 231493 -3693
rect 231611 -3811 231653 -3693
rect 231771 -3811 231787 -3693
rect 231477 -3827 231787 -3811
rect 240477 -3053 240787 7029
rect 243897 352899 244207 352915
rect 243897 352781 243913 352899
rect 244031 352781 244073 352899
rect 244191 352781 244207 352899
rect 243897 352739 244207 352781
rect 243897 352621 243913 352739
rect 244031 352621 244073 352739
rect 244191 352621 244207 352739
rect 243897 334727 244207 352621
rect 243897 334609 243913 334727
rect 244031 334609 244073 334727
rect 244191 334609 244207 334727
rect 243897 334567 244207 334609
rect 243897 334449 243913 334567
rect 244031 334449 244073 334567
rect 244191 334449 244207 334567
rect 243897 316727 244207 334449
rect 243897 316609 243913 316727
rect 244031 316609 244073 316727
rect 244191 316609 244207 316727
rect 243897 316567 244207 316609
rect 243897 316449 243913 316567
rect 244031 316449 244073 316567
rect 244191 316449 244207 316567
rect 243897 298727 244207 316449
rect 243897 298609 243913 298727
rect 244031 298609 244073 298727
rect 244191 298609 244207 298727
rect 243897 298567 244207 298609
rect 243897 298449 243913 298567
rect 244031 298449 244073 298567
rect 244191 298449 244207 298567
rect 243897 280727 244207 298449
rect 243897 280609 243913 280727
rect 244031 280609 244073 280727
rect 244191 280609 244207 280727
rect 243897 280567 244207 280609
rect 243897 280449 243913 280567
rect 244031 280449 244073 280567
rect 244191 280449 244207 280567
rect 243897 262727 244207 280449
rect 243897 262609 243913 262727
rect 244031 262609 244073 262727
rect 244191 262609 244207 262727
rect 243897 262567 244207 262609
rect 243897 262449 243913 262567
rect 244031 262449 244073 262567
rect 244191 262449 244207 262567
rect 243897 244727 244207 262449
rect 243897 244609 243913 244727
rect 244031 244609 244073 244727
rect 244191 244609 244207 244727
rect 243897 244567 244207 244609
rect 243897 244449 243913 244567
rect 244031 244449 244073 244567
rect 244191 244449 244207 244567
rect 243897 226727 244207 244449
rect 243897 226609 243913 226727
rect 244031 226609 244073 226727
rect 244191 226609 244207 226727
rect 243897 226567 244207 226609
rect 243897 226449 243913 226567
rect 244031 226449 244073 226567
rect 244191 226449 244207 226567
rect 243897 208727 244207 226449
rect 243897 208609 243913 208727
rect 244031 208609 244073 208727
rect 244191 208609 244207 208727
rect 243897 208567 244207 208609
rect 243897 208449 243913 208567
rect 244031 208449 244073 208567
rect 244191 208449 244207 208567
rect 243897 190727 244207 208449
rect 243897 190609 243913 190727
rect 244031 190609 244073 190727
rect 244191 190609 244207 190727
rect 243897 190567 244207 190609
rect 243897 190449 243913 190567
rect 244031 190449 244073 190567
rect 244191 190449 244207 190567
rect 243897 172727 244207 190449
rect 243897 172609 243913 172727
rect 244031 172609 244073 172727
rect 244191 172609 244207 172727
rect 243897 172567 244207 172609
rect 243897 172449 243913 172567
rect 244031 172449 244073 172567
rect 244191 172449 244207 172567
rect 243897 154727 244207 172449
rect 243897 154609 243913 154727
rect 244031 154609 244073 154727
rect 244191 154609 244207 154727
rect 243897 154567 244207 154609
rect 243897 154449 243913 154567
rect 244031 154449 244073 154567
rect 244191 154449 244207 154567
rect 243897 136727 244207 154449
rect 243897 136609 243913 136727
rect 244031 136609 244073 136727
rect 244191 136609 244207 136727
rect 243897 136567 244207 136609
rect 243897 136449 243913 136567
rect 244031 136449 244073 136567
rect 244191 136449 244207 136567
rect 243897 118727 244207 136449
rect 243897 118609 243913 118727
rect 244031 118609 244073 118727
rect 244191 118609 244207 118727
rect 243897 118567 244207 118609
rect 243897 118449 243913 118567
rect 244031 118449 244073 118567
rect 244191 118449 244207 118567
rect 243897 100727 244207 118449
rect 243897 100609 243913 100727
rect 244031 100609 244073 100727
rect 244191 100609 244207 100727
rect 243897 100567 244207 100609
rect 243897 100449 243913 100567
rect 244031 100449 244073 100567
rect 244191 100449 244207 100567
rect 243897 82727 244207 100449
rect 243897 82609 243913 82727
rect 244031 82609 244073 82727
rect 244191 82609 244207 82727
rect 243897 82567 244207 82609
rect 243897 82449 243913 82567
rect 244031 82449 244073 82567
rect 244191 82449 244207 82567
rect 243897 64727 244207 82449
rect 243897 64609 243913 64727
rect 244031 64609 244073 64727
rect 244191 64609 244207 64727
rect 243897 64567 244207 64609
rect 243897 64449 243913 64567
rect 244031 64449 244073 64567
rect 244191 64449 244207 64567
rect 243897 46727 244207 64449
rect 243897 46609 243913 46727
rect 244031 46609 244073 46727
rect 244191 46609 244207 46727
rect 243897 46567 244207 46609
rect 243897 46449 243913 46567
rect 244031 46449 244073 46567
rect 244191 46449 244207 46567
rect 243897 28727 244207 46449
rect 243897 28609 243913 28727
rect 244031 28609 244073 28727
rect 244191 28609 244207 28727
rect 243897 28567 244207 28609
rect 243897 28449 243913 28567
rect 244031 28449 244073 28567
rect 244191 28449 244207 28567
rect 243897 10727 244207 28449
rect 243897 10609 243913 10727
rect 244031 10609 244073 10727
rect 244191 10609 244207 10727
rect 243897 10567 244207 10609
rect 243897 10449 243913 10567
rect 244031 10449 244073 10567
rect 244191 10449 244207 10567
rect 243897 -653 244207 10449
rect 243897 -771 243913 -653
rect 244031 -771 244073 -653
rect 244191 -771 244207 -653
rect 243897 -813 244207 -771
rect 243897 -931 243913 -813
rect 244031 -931 244073 -813
rect 244191 -931 244207 -813
rect 243897 -947 244207 -931
rect 245757 336587 246067 353581
rect 245757 336469 245773 336587
rect 245891 336469 245933 336587
rect 246051 336469 246067 336587
rect 245757 336427 246067 336469
rect 245757 336309 245773 336427
rect 245891 336309 245933 336427
rect 246051 336309 246067 336427
rect 245757 318587 246067 336309
rect 245757 318469 245773 318587
rect 245891 318469 245933 318587
rect 246051 318469 246067 318587
rect 245757 318427 246067 318469
rect 245757 318309 245773 318427
rect 245891 318309 245933 318427
rect 246051 318309 246067 318427
rect 245757 300587 246067 318309
rect 245757 300469 245773 300587
rect 245891 300469 245933 300587
rect 246051 300469 246067 300587
rect 245757 300427 246067 300469
rect 245757 300309 245773 300427
rect 245891 300309 245933 300427
rect 246051 300309 246067 300427
rect 245757 282587 246067 300309
rect 245757 282469 245773 282587
rect 245891 282469 245933 282587
rect 246051 282469 246067 282587
rect 245757 282427 246067 282469
rect 245757 282309 245773 282427
rect 245891 282309 245933 282427
rect 246051 282309 246067 282427
rect 245757 264587 246067 282309
rect 245757 264469 245773 264587
rect 245891 264469 245933 264587
rect 246051 264469 246067 264587
rect 245757 264427 246067 264469
rect 245757 264309 245773 264427
rect 245891 264309 245933 264427
rect 246051 264309 246067 264427
rect 245757 246587 246067 264309
rect 245757 246469 245773 246587
rect 245891 246469 245933 246587
rect 246051 246469 246067 246587
rect 245757 246427 246067 246469
rect 245757 246309 245773 246427
rect 245891 246309 245933 246427
rect 246051 246309 246067 246427
rect 245757 228587 246067 246309
rect 245757 228469 245773 228587
rect 245891 228469 245933 228587
rect 246051 228469 246067 228587
rect 245757 228427 246067 228469
rect 245757 228309 245773 228427
rect 245891 228309 245933 228427
rect 246051 228309 246067 228427
rect 245757 210587 246067 228309
rect 245757 210469 245773 210587
rect 245891 210469 245933 210587
rect 246051 210469 246067 210587
rect 245757 210427 246067 210469
rect 245757 210309 245773 210427
rect 245891 210309 245933 210427
rect 246051 210309 246067 210427
rect 245757 192587 246067 210309
rect 245757 192469 245773 192587
rect 245891 192469 245933 192587
rect 246051 192469 246067 192587
rect 245757 192427 246067 192469
rect 245757 192309 245773 192427
rect 245891 192309 245933 192427
rect 246051 192309 246067 192427
rect 245757 174587 246067 192309
rect 245757 174469 245773 174587
rect 245891 174469 245933 174587
rect 246051 174469 246067 174587
rect 245757 174427 246067 174469
rect 245757 174309 245773 174427
rect 245891 174309 245933 174427
rect 246051 174309 246067 174427
rect 245757 156587 246067 174309
rect 245757 156469 245773 156587
rect 245891 156469 245933 156587
rect 246051 156469 246067 156587
rect 245757 156427 246067 156469
rect 245757 156309 245773 156427
rect 245891 156309 245933 156427
rect 246051 156309 246067 156427
rect 245757 138587 246067 156309
rect 245757 138469 245773 138587
rect 245891 138469 245933 138587
rect 246051 138469 246067 138587
rect 245757 138427 246067 138469
rect 245757 138309 245773 138427
rect 245891 138309 245933 138427
rect 246051 138309 246067 138427
rect 245757 120587 246067 138309
rect 245757 120469 245773 120587
rect 245891 120469 245933 120587
rect 246051 120469 246067 120587
rect 245757 120427 246067 120469
rect 245757 120309 245773 120427
rect 245891 120309 245933 120427
rect 246051 120309 246067 120427
rect 245757 102587 246067 120309
rect 245757 102469 245773 102587
rect 245891 102469 245933 102587
rect 246051 102469 246067 102587
rect 245757 102427 246067 102469
rect 245757 102309 245773 102427
rect 245891 102309 245933 102427
rect 246051 102309 246067 102427
rect 245757 84587 246067 102309
rect 245757 84469 245773 84587
rect 245891 84469 245933 84587
rect 246051 84469 246067 84587
rect 245757 84427 246067 84469
rect 245757 84309 245773 84427
rect 245891 84309 245933 84427
rect 246051 84309 246067 84427
rect 245757 66587 246067 84309
rect 245757 66469 245773 66587
rect 245891 66469 245933 66587
rect 246051 66469 246067 66587
rect 245757 66427 246067 66469
rect 245757 66309 245773 66427
rect 245891 66309 245933 66427
rect 246051 66309 246067 66427
rect 245757 48587 246067 66309
rect 245757 48469 245773 48587
rect 245891 48469 245933 48587
rect 246051 48469 246067 48587
rect 245757 48427 246067 48469
rect 245757 48309 245773 48427
rect 245891 48309 245933 48427
rect 246051 48309 246067 48427
rect 245757 30587 246067 48309
rect 245757 30469 245773 30587
rect 245891 30469 245933 30587
rect 246051 30469 246067 30587
rect 245757 30427 246067 30469
rect 245757 30309 245773 30427
rect 245891 30309 245933 30427
rect 246051 30309 246067 30427
rect 245757 12587 246067 30309
rect 245757 12469 245773 12587
rect 245891 12469 245933 12587
rect 246051 12469 246067 12587
rect 245757 12427 246067 12469
rect 245757 12309 245773 12427
rect 245891 12309 245933 12427
rect 246051 12309 246067 12427
rect 245757 -1613 246067 12309
rect 245757 -1731 245773 -1613
rect 245891 -1731 245933 -1613
rect 246051 -1731 246067 -1613
rect 245757 -1773 246067 -1731
rect 245757 -1891 245773 -1773
rect 245891 -1891 245933 -1773
rect 246051 -1891 246067 -1773
rect 245757 -1907 246067 -1891
rect 247617 338447 247927 354541
rect 247617 338329 247633 338447
rect 247751 338329 247793 338447
rect 247911 338329 247927 338447
rect 247617 338287 247927 338329
rect 247617 338169 247633 338287
rect 247751 338169 247793 338287
rect 247911 338169 247927 338287
rect 247617 320447 247927 338169
rect 247617 320329 247633 320447
rect 247751 320329 247793 320447
rect 247911 320329 247927 320447
rect 247617 320287 247927 320329
rect 247617 320169 247633 320287
rect 247751 320169 247793 320287
rect 247911 320169 247927 320287
rect 247617 302447 247927 320169
rect 247617 302329 247633 302447
rect 247751 302329 247793 302447
rect 247911 302329 247927 302447
rect 247617 302287 247927 302329
rect 247617 302169 247633 302287
rect 247751 302169 247793 302287
rect 247911 302169 247927 302287
rect 247617 284447 247927 302169
rect 247617 284329 247633 284447
rect 247751 284329 247793 284447
rect 247911 284329 247927 284447
rect 247617 284287 247927 284329
rect 247617 284169 247633 284287
rect 247751 284169 247793 284287
rect 247911 284169 247927 284287
rect 247617 266447 247927 284169
rect 247617 266329 247633 266447
rect 247751 266329 247793 266447
rect 247911 266329 247927 266447
rect 247617 266287 247927 266329
rect 247617 266169 247633 266287
rect 247751 266169 247793 266287
rect 247911 266169 247927 266287
rect 247617 248447 247927 266169
rect 247617 248329 247633 248447
rect 247751 248329 247793 248447
rect 247911 248329 247927 248447
rect 247617 248287 247927 248329
rect 247617 248169 247633 248287
rect 247751 248169 247793 248287
rect 247911 248169 247927 248287
rect 247617 230447 247927 248169
rect 247617 230329 247633 230447
rect 247751 230329 247793 230447
rect 247911 230329 247927 230447
rect 247617 230287 247927 230329
rect 247617 230169 247633 230287
rect 247751 230169 247793 230287
rect 247911 230169 247927 230287
rect 247617 212447 247927 230169
rect 247617 212329 247633 212447
rect 247751 212329 247793 212447
rect 247911 212329 247927 212447
rect 247617 212287 247927 212329
rect 247617 212169 247633 212287
rect 247751 212169 247793 212287
rect 247911 212169 247927 212287
rect 247617 194447 247927 212169
rect 247617 194329 247633 194447
rect 247751 194329 247793 194447
rect 247911 194329 247927 194447
rect 247617 194287 247927 194329
rect 247617 194169 247633 194287
rect 247751 194169 247793 194287
rect 247911 194169 247927 194287
rect 247617 176447 247927 194169
rect 247617 176329 247633 176447
rect 247751 176329 247793 176447
rect 247911 176329 247927 176447
rect 247617 176287 247927 176329
rect 247617 176169 247633 176287
rect 247751 176169 247793 176287
rect 247911 176169 247927 176287
rect 247617 158447 247927 176169
rect 247617 158329 247633 158447
rect 247751 158329 247793 158447
rect 247911 158329 247927 158447
rect 247617 158287 247927 158329
rect 247617 158169 247633 158287
rect 247751 158169 247793 158287
rect 247911 158169 247927 158287
rect 247617 140447 247927 158169
rect 247617 140329 247633 140447
rect 247751 140329 247793 140447
rect 247911 140329 247927 140447
rect 247617 140287 247927 140329
rect 247617 140169 247633 140287
rect 247751 140169 247793 140287
rect 247911 140169 247927 140287
rect 247617 122447 247927 140169
rect 247617 122329 247633 122447
rect 247751 122329 247793 122447
rect 247911 122329 247927 122447
rect 247617 122287 247927 122329
rect 247617 122169 247633 122287
rect 247751 122169 247793 122287
rect 247911 122169 247927 122287
rect 247617 104447 247927 122169
rect 247617 104329 247633 104447
rect 247751 104329 247793 104447
rect 247911 104329 247927 104447
rect 247617 104287 247927 104329
rect 247617 104169 247633 104287
rect 247751 104169 247793 104287
rect 247911 104169 247927 104287
rect 247617 86447 247927 104169
rect 247617 86329 247633 86447
rect 247751 86329 247793 86447
rect 247911 86329 247927 86447
rect 247617 86287 247927 86329
rect 247617 86169 247633 86287
rect 247751 86169 247793 86287
rect 247911 86169 247927 86287
rect 247617 68447 247927 86169
rect 247617 68329 247633 68447
rect 247751 68329 247793 68447
rect 247911 68329 247927 68447
rect 247617 68287 247927 68329
rect 247617 68169 247633 68287
rect 247751 68169 247793 68287
rect 247911 68169 247927 68287
rect 247617 50447 247927 68169
rect 247617 50329 247633 50447
rect 247751 50329 247793 50447
rect 247911 50329 247927 50447
rect 247617 50287 247927 50329
rect 247617 50169 247633 50287
rect 247751 50169 247793 50287
rect 247911 50169 247927 50287
rect 247617 32447 247927 50169
rect 247617 32329 247633 32447
rect 247751 32329 247793 32447
rect 247911 32329 247927 32447
rect 247617 32287 247927 32329
rect 247617 32169 247633 32287
rect 247751 32169 247793 32287
rect 247911 32169 247927 32287
rect 247617 14447 247927 32169
rect 247617 14329 247633 14447
rect 247751 14329 247793 14447
rect 247911 14329 247927 14447
rect 247617 14287 247927 14329
rect 247617 14169 247633 14287
rect 247751 14169 247793 14287
rect 247911 14169 247927 14287
rect 247617 -2573 247927 14169
rect 247617 -2691 247633 -2573
rect 247751 -2691 247793 -2573
rect 247911 -2691 247927 -2573
rect 247617 -2733 247927 -2691
rect 247617 -2851 247633 -2733
rect 247751 -2851 247793 -2733
rect 247911 -2851 247927 -2733
rect 247617 -2867 247927 -2851
rect 249477 340307 249787 355501
rect 258477 355299 258787 355795
rect 258477 355181 258493 355299
rect 258611 355181 258653 355299
rect 258771 355181 258787 355299
rect 258477 355139 258787 355181
rect 258477 355021 258493 355139
rect 258611 355021 258653 355139
rect 258771 355021 258787 355139
rect 256617 354339 256927 354835
rect 256617 354221 256633 354339
rect 256751 354221 256793 354339
rect 256911 354221 256927 354339
rect 256617 354179 256927 354221
rect 256617 354061 256633 354179
rect 256751 354061 256793 354179
rect 256911 354061 256927 354179
rect 254757 353379 255067 353875
rect 254757 353261 254773 353379
rect 254891 353261 254933 353379
rect 255051 353261 255067 353379
rect 254757 353219 255067 353261
rect 254757 353101 254773 353219
rect 254891 353101 254933 353219
rect 255051 353101 255067 353219
rect 249477 340189 249493 340307
rect 249611 340189 249653 340307
rect 249771 340189 249787 340307
rect 249477 340147 249787 340189
rect 249477 340029 249493 340147
rect 249611 340029 249653 340147
rect 249771 340029 249787 340147
rect 249477 322307 249787 340029
rect 249477 322189 249493 322307
rect 249611 322189 249653 322307
rect 249771 322189 249787 322307
rect 249477 322147 249787 322189
rect 249477 322029 249493 322147
rect 249611 322029 249653 322147
rect 249771 322029 249787 322147
rect 249477 304307 249787 322029
rect 249477 304189 249493 304307
rect 249611 304189 249653 304307
rect 249771 304189 249787 304307
rect 249477 304147 249787 304189
rect 249477 304029 249493 304147
rect 249611 304029 249653 304147
rect 249771 304029 249787 304147
rect 249477 286307 249787 304029
rect 249477 286189 249493 286307
rect 249611 286189 249653 286307
rect 249771 286189 249787 286307
rect 249477 286147 249787 286189
rect 249477 286029 249493 286147
rect 249611 286029 249653 286147
rect 249771 286029 249787 286147
rect 249477 268307 249787 286029
rect 249477 268189 249493 268307
rect 249611 268189 249653 268307
rect 249771 268189 249787 268307
rect 249477 268147 249787 268189
rect 249477 268029 249493 268147
rect 249611 268029 249653 268147
rect 249771 268029 249787 268147
rect 249477 250307 249787 268029
rect 249477 250189 249493 250307
rect 249611 250189 249653 250307
rect 249771 250189 249787 250307
rect 249477 250147 249787 250189
rect 249477 250029 249493 250147
rect 249611 250029 249653 250147
rect 249771 250029 249787 250147
rect 249477 232307 249787 250029
rect 249477 232189 249493 232307
rect 249611 232189 249653 232307
rect 249771 232189 249787 232307
rect 249477 232147 249787 232189
rect 249477 232029 249493 232147
rect 249611 232029 249653 232147
rect 249771 232029 249787 232147
rect 249477 214307 249787 232029
rect 249477 214189 249493 214307
rect 249611 214189 249653 214307
rect 249771 214189 249787 214307
rect 249477 214147 249787 214189
rect 249477 214029 249493 214147
rect 249611 214029 249653 214147
rect 249771 214029 249787 214147
rect 249477 196307 249787 214029
rect 249477 196189 249493 196307
rect 249611 196189 249653 196307
rect 249771 196189 249787 196307
rect 249477 196147 249787 196189
rect 249477 196029 249493 196147
rect 249611 196029 249653 196147
rect 249771 196029 249787 196147
rect 249477 178307 249787 196029
rect 249477 178189 249493 178307
rect 249611 178189 249653 178307
rect 249771 178189 249787 178307
rect 249477 178147 249787 178189
rect 249477 178029 249493 178147
rect 249611 178029 249653 178147
rect 249771 178029 249787 178147
rect 249477 160307 249787 178029
rect 249477 160189 249493 160307
rect 249611 160189 249653 160307
rect 249771 160189 249787 160307
rect 249477 160147 249787 160189
rect 249477 160029 249493 160147
rect 249611 160029 249653 160147
rect 249771 160029 249787 160147
rect 249477 142307 249787 160029
rect 249477 142189 249493 142307
rect 249611 142189 249653 142307
rect 249771 142189 249787 142307
rect 249477 142147 249787 142189
rect 249477 142029 249493 142147
rect 249611 142029 249653 142147
rect 249771 142029 249787 142147
rect 249477 124307 249787 142029
rect 249477 124189 249493 124307
rect 249611 124189 249653 124307
rect 249771 124189 249787 124307
rect 249477 124147 249787 124189
rect 249477 124029 249493 124147
rect 249611 124029 249653 124147
rect 249771 124029 249787 124147
rect 249477 106307 249787 124029
rect 249477 106189 249493 106307
rect 249611 106189 249653 106307
rect 249771 106189 249787 106307
rect 249477 106147 249787 106189
rect 249477 106029 249493 106147
rect 249611 106029 249653 106147
rect 249771 106029 249787 106147
rect 249477 88307 249787 106029
rect 249477 88189 249493 88307
rect 249611 88189 249653 88307
rect 249771 88189 249787 88307
rect 249477 88147 249787 88189
rect 249477 88029 249493 88147
rect 249611 88029 249653 88147
rect 249771 88029 249787 88147
rect 249477 70307 249787 88029
rect 249477 70189 249493 70307
rect 249611 70189 249653 70307
rect 249771 70189 249787 70307
rect 249477 70147 249787 70189
rect 249477 70029 249493 70147
rect 249611 70029 249653 70147
rect 249771 70029 249787 70147
rect 249477 52307 249787 70029
rect 249477 52189 249493 52307
rect 249611 52189 249653 52307
rect 249771 52189 249787 52307
rect 249477 52147 249787 52189
rect 249477 52029 249493 52147
rect 249611 52029 249653 52147
rect 249771 52029 249787 52147
rect 249477 34307 249787 52029
rect 249477 34189 249493 34307
rect 249611 34189 249653 34307
rect 249771 34189 249787 34307
rect 249477 34147 249787 34189
rect 249477 34029 249493 34147
rect 249611 34029 249653 34147
rect 249771 34029 249787 34147
rect 249477 16307 249787 34029
rect 249477 16189 249493 16307
rect 249611 16189 249653 16307
rect 249771 16189 249787 16307
rect 249477 16147 249787 16189
rect 249477 16029 249493 16147
rect 249611 16029 249653 16147
rect 249771 16029 249787 16147
rect 240477 -3171 240493 -3053
rect 240611 -3171 240653 -3053
rect 240771 -3171 240787 -3053
rect 240477 -3213 240787 -3171
rect 240477 -3331 240493 -3213
rect 240611 -3331 240653 -3213
rect 240771 -3331 240787 -3213
rect 240477 -3827 240787 -3331
rect 249477 -3533 249787 16029
rect 252897 352419 253207 352915
rect 252897 352301 252913 352419
rect 253031 352301 253073 352419
rect 253191 352301 253207 352419
rect 252897 352259 253207 352301
rect 252897 352141 252913 352259
rect 253031 352141 253073 352259
rect 253191 352141 253207 352259
rect 252897 343727 253207 352141
rect 252897 343609 252913 343727
rect 253031 343609 253073 343727
rect 253191 343609 253207 343727
rect 252897 343567 253207 343609
rect 252897 343449 252913 343567
rect 253031 343449 253073 343567
rect 253191 343449 253207 343567
rect 252897 325727 253207 343449
rect 252897 325609 252913 325727
rect 253031 325609 253073 325727
rect 253191 325609 253207 325727
rect 252897 325567 253207 325609
rect 252897 325449 252913 325567
rect 253031 325449 253073 325567
rect 253191 325449 253207 325567
rect 252897 307727 253207 325449
rect 252897 307609 252913 307727
rect 253031 307609 253073 307727
rect 253191 307609 253207 307727
rect 252897 307567 253207 307609
rect 252897 307449 252913 307567
rect 253031 307449 253073 307567
rect 253191 307449 253207 307567
rect 252897 289727 253207 307449
rect 252897 289609 252913 289727
rect 253031 289609 253073 289727
rect 253191 289609 253207 289727
rect 252897 289567 253207 289609
rect 252897 289449 252913 289567
rect 253031 289449 253073 289567
rect 253191 289449 253207 289567
rect 252897 271727 253207 289449
rect 252897 271609 252913 271727
rect 253031 271609 253073 271727
rect 253191 271609 253207 271727
rect 252897 271567 253207 271609
rect 252897 271449 252913 271567
rect 253031 271449 253073 271567
rect 253191 271449 253207 271567
rect 252897 253727 253207 271449
rect 252897 253609 252913 253727
rect 253031 253609 253073 253727
rect 253191 253609 253207 253727
rect 252897 253567 253207 253609
rect 252897 253449 252913 253567
rect 253031 253449 253073 253567
rect 253191 253449 253207 253567
rect 252897 235727 253207 253449
rect 252897 235609 252913 235727
rect 253031 235609 253073 235727
rect 253191 235609 253207 235727
rect 252897 235567 253207 235609
rect 252897 235449 252913 235567
rect 253031 235449 253073 235567
rect 253191 235449 253207 235567
rect 252897 217727 253207 235449
rect 252897 217609 252913 217727
rect 253031 217609 253073 217727
rect 253191 217609 253207 217727
rect 252897 217567 253207 217609
rect 252897 217449 252913 217567
rect 253031 217449 253073 217567
rect 253191 217449 253207 217567
rect 252897 199727 253207 217449
rect 252897 199609 252913 199727
rect 253031 199609 253073 199727
rect 253191 199609 253207 199727
rect 252897 199567 253207 199609
rect 252897 199449 252913 199567
rect 253031 199449 253073 199567
rect 253191 199449 253207 199567
rect 252897 181727 253207 199449
rect 252897 181609 252913 181727
rect 253031 181609 253073 181727
rect 253191 181609 253207 181727
rect 252897 181567 253207 181609
rect 252897 181449 252913 181567
rect 253031 181449 253073 181567
rect 253191 181449 253207 181567
rect 252897 163727 253207 181449
rect 252897 163609 252913 163727
rect 253031 163609 253073 163727
rect 253191 163609 253207 163727
rect 252897 163567 253207 163609
rect 252897 163449 252913 163567
rect 253031 163449 253073 163567
rect 253191 163449 253207 163567
rect 252897 145727 253207 163449
rect 252897 145609 252913 145727
rect 253031 145609 253073 145727
rect 253191 145609 253207 145727
rect 252897 145567 253207 145609
rect 252897 145449 252913 145567
rect 253031 145449 253073 145567
rect 253191 145449 253207 145567
rect 252897 127727 253207 145449
rect 252897 127609 252913 127727
rect 253031 127609 253073 127727
rect 253191 127609 253207 127727
rect 252897 127567 253207 127609
rect 252897 127449 252913 127567
rect 253031 127449 253073 127567
rect 253191 127449 253207 127567
rect 252897 109727 253207 127449
rect 252897 109609 252913 109727
rect 253031 109609 253073 109727
rect 253191 109609 253207 109727
rect 252897 109567 253207 109609
rect 252897 109449 252913 109567
rect 253031 109449 253073 109567
rect 253191 109449 253207 109567
rect 252897 91727 253207 109449
rect 252897 91609 252913 91727
rect 253031 91609 253073 91727
rect 253191 91609 253207 91727
rect 252897 91567 253207 91609
rect 252897 91449 252913 91567
rect 253031 91449 253073 91567
rect 253191 91449 253207 91567
rect 252897 73727 253207 91449
rect 252897 73609 252913 73727
rect 253031 73609 253073 73727
rect 253191 73609 253207 73727
rect 252897 73567 253207 73609
rect 252897 73449 252913 73567
rect 253031 73449 253073 73567
rect 253191 73449 253207 73567
rect 252897 55727 253207 73449
rect 252897 55609 252913 55727
rect 253031 55609 253073 55727
rect 253191 55609 253207 55727
rect 252897 55567 253207 55609
rect 252897 55449 252913 55567
rect 253031 55449 253073 55567
rect 253191 55449 253207 55567
rect 252897 37727 253207 55449
rect 252897 37609 252913 37727
rect 253031 37609 253073 37727
rect 253191 37609 253207 37727
rect 252897 37567 253207 37609
rect 252897 37449 252913 37567
rect 253031 37449 253073 37567
rect 253191 37449 253207 37567
rect 252897 19727 253207 37449
rect 252897 19609 252913 19727
rect 253031 19609 253073 19727
rect 253191 19609 253207 19727
rect 252897 19567 253207 19609
rect 252897 19449 252913 19567
rect 253031 19449 253073 19567
rect 253191 19449 253207 19567
rect 252897 1727 253207 19449
rect 252897 1609 252913 1727
rect 253031 1609 253073 1727
rect 253191 1609 253207 1727
rect 252897 1567 253207 1609
rect 252897 1449 252913 1567
rect 253031 1449 253073 1567
rect 253191 1449 253207 1567
rect 252897 -173 253207 1449
rect 252897 -291 252913 -173
rect 253031 -291 253073 -173
rect 253191 -291 253207 -173
rect 252897 -333 253207 -291
rect 252897 -451 252913 -333
rect 253031 -451 253073 -333
rect 253191 -451 253207 -333
rect 252897 -947 253207 -451
rect 254757 345587 255067 353101
rect 254757 345469 254773 345587
rect 254891 345469 254933 345587
rect 255051 345469 255067 345587
rect 254757 345427 255067 345469
rect 254757 345309 254773 345427
rect 254891 345309 254933 345427
rect 255051 345309 255067 345427
rect 254757 327587 255067 345309
rect 254757 327469 254773 327587
rect 254891 327469 254933 327587
rect 255051 327469 255067 327587
rect 254757 327427 255067 327469
rect 254757 327309 254773 327427
rect 254891 327309 254933 327427
rect 255051 327309 255067 327427
rect 254757 309587 255067 327309
rect 254757 309469 254773 309587
rect 254891 309469 254933 309587
rect 255051 309469 255067 309587
rect 254757 309427 255067 309469
rect 254757 309309 254773 309427
rect 254891 309309 254933 309427
rect 255051 309309 255067 309427
rect 254757 291587 255067 309309
rect 254757 291469 254773 291587
rect 254891 291469 254933 291587
rect 255051 291469 255067 291587
rect 254757 291427 255067 291469
rect 254757 291309 254773 291427
rect 254891 291309 254933 291427
rect 255051 291309 255067 291427
rect 254757 273587 255067 291309
rect 254757 273469 254773 273587
rect 254891 273469 254933 273587
rect 255051 273469 255067 273587
rect 254757 273427 255067 273469
rect 254757 273309 254773 273427
rect 254891 273309 254933 273427
rect 255051 273309 255067 273427
rect 254757 255587 255067 273309
rect 254757 255469 254773 255587
rect 254891 255469 254933 255587
rect 255051 255469 255067 255587
rect 254757 255427 255067 255469
rect 254757 255309 254773 255427
rect 254891 255309 254933 255427
rect 255051 255309 255067 255427
rect 254757 237587 255067 255309
rect 254757 237469 254773 237587
rect 254891 237469 254933 237587
rect 255051 237469 255067 237587
rect 254757 237427 255067 237469
rect 254757 237309 254773 237427
rect 254891 237309 254933 237427
rect 255051 237309 255067 237427
rect 254757 219587 255067 237309
rect 254757 219469 254773 219587
rect 254891 219469 254933 219587
rect 255051 219469 255067 219587
rect 254757 219427 255067 219469
rect 254757 219309 254773 219427
rect 254891 219309 254933 219427
rect 255051 219309 255067 219427
rect 254757 201587 255067 219309
rect 254757 201469 254773 201587
rect 254891 201469 254933 201587
rect 255051 201469 255067 201587
rect 254757 201427 255067 201469
rect 254757 201309 254773 201427
rect 254891 201309 254933 201427
rect 255051 201309 255067 201427
rect 254757 183587 255067 201309
rect 254757 183469 254773 183587
rect 254891 183469 254933 183587
rect 255051 183469 255067 183587
rect 254757 183427 255067 183469
rect 254757 183309 254773 183427
rect 254891 183309 254933 183427
rect 255051 183309 255067 183427
rect 254757 165587 255067 183309
rect 254757 165469 254773 165587
rect 254891 165469 254933 165587
rect 255051 165469 255067 165587
rect 254757 165427 255067 165469
rect 254757 165309 254773 165427
rect 254891 165309 254933 165427
rect 255051 165309 255067 165427
rect 254757 147587 255067 165309
rect 254757 147469 254773 147587
rect 254891 147469 254933 147587
rect 255051 147469 255067 147587
rect 254757 147427 255067 147469
rect 254757 147309 254773 147427
rect 254891 147309 254933 147427
rect 255051 147309 255067 147427
rect 254757 129587 255067 147309
rect 254757 129469 254773 129587
rect 254891 129469 254933 129587
rect 255051 129469 255067 129587
rect 254757 129427 255067 129469
rect 254757 129309 254773 129427
rect 254891 129309 254933 129427
rect 255051 129309 255067 129427
rect 254757 111587 255067 129309
rect 254757 111469 254773 111587
rect 254891 111469 254933 111587
rect 255051 111469 255067 111587
rect 254757 111427 255067 111469
rect 254757 111309 254773 111427
rect 254891 111309 254933 111427
rect 255051 111309 255067 111427
rect 254757 93587 255067 111309
rect 254757 93469 254773 93587
rect 254891 93469 254933 93587
rect 255051 93469 255067 93587
rect 254757 93427 255067 93469
rect 254757 93309 254773 93427
rect 254891 93309 254933 93427
rect 255051 93309 255067 93427
rect 254757 75587 255067 93309
rect 254757 75469 254773 75587
rect 254891 75469 254933 75587
rect 255051 75469 255067 75587
rect 254757 75427 255067 75469
rect 254757 75309 254773 75427
rect 254891 75309 254933 75427
rect 255051 75309 255067 75427
rect 254757 57587 255067 75309
rect 254757 57469 254773 57587
rect 254891 57469 254933 57587
rect 255051 57469 255067 57587
rect 254757 57427 255067 57469
rect 254757 57309 254773 57427
rect 254891 57309 254933 57427
rect 255051 57309 255067 57427
rect 254757 39587 255067 57309
rect 254757 39469 254773 39587
rect 254891 39469 254933 39587
rect 255051 39469 255067 39587
rect 254757 39427 255067 39469
rect 254757 39309 254773 39427
rect 254891 39309 254933 39427
rect 255051 39309 255067 39427
rect 254757 21587 255067 39309
rect 254757 21469 254773 21587
rect 254891 21469 254933 21587
rect 255051 21469 255067 21587
rect 254757 21427 255067 21469
rect 254757 21309 254773 21427
rect 254891 21309 254933 21427
rect 255051 21309 255067 21427
rect 254757 3587 255067 21309
rect 254757 3469 254773 3587
rect 254891 3469 254933 3587
rect 255051 3469 255067 3587
rect 254757 3427 255067 3469
rect 254757 3309 254773 3427
rect 254891 3309 254933 3427
rect 255051 3309 255067 3427
rect 254757 -1133 255067 3309
rect 254757 -1251 254773 -1133
rect 254891 -1251 254933 -1133
rect 255051 -1251 255067 -1133
rect 254757 -1293 255067 -1251
rect 254757 -1411 254773 -1293
rect 254891 -1411 254933 -1293
rect 255051 -1411 255067 -1293
rect 254757 -1907 255067 -1411
rect 256617 347447 256927 354061
rect 256617 347329 256633 347447
rect 256751 347329 256793 347447
rect 256911 347329 256927 347447
rect 256617 347287 256927 347329
rect 256617 347169 256633 347287
rect 256751 347169 256793 347287
rect 256911 347169 256927 347287
rect 256617 329447 256927 347169
rect 256617 329329 256633 329447
rect 256751 329329 256793 329447
rect 256911 329329 256927 329447
rect 256617 329287 256927 329329
rect 256617 329169 256633 329287
rect 256751 329169 256793 329287
rect 256911 329169 256927 329287
rect 256617 311447 256927 329169
rect 256617 311329 256633 311447
rect 256751 311329 256793 311447
rect 256911 311329 256927 311447
rect 256617 311287 256927 311329
rect 256617 311169 256633 311287
rect 256751 311169 256793 311287
rect 256911 311169 256927 311287
rect 256617 293447 256927 311169
rect 256617 293329 256633 293447
rect 256751 293329 256793 293447
rect 256911 293329 256927 293447
rect 256617 293287 256927 293329
rect 256617 293169 256633 293287
rect 256751 293169 256793 293287
rect 256911 293169 256927 293287
rect 256617 275447 256927 293169
rect 256617 275329 256633 275447
rect 256751 275329 256793 275447
rect 256911 275329 256927 275447
rect 256617 275287 256927 275329
rect 256617 275169 256633 275287
rect 256751 275169 256793 275287
rect 256911 275169 256927 275287
rect 256617 257447 256927 275169
rect 256617 257329 256633 257447
rect 256751 257329 256793 257447
rect 256911 257329 256927 257447
rect 256617 257287 256927 257329
rect 256617 257169 256633 257287
rect 256751 257169 256793 257287
rect 256911 257169 256927 257287
rect 256617 239447 256927 257169
rect 256617 239329 256633 239447
rect 256751 239329 256793 239447
rect 256911 239329 256927 239447
rect 256617 239287 256927 239329
rect 256617 239169 256633 239287
rect 256751 239169 256793 239287
rect 256911 239169 256927 239287
rect 256617 221447 256927 239169
rect 256617 221329 256633 221447
rect 256751 221329 256793 221447
rect 256911 221329 256927 221447
rect 256617 221287 256927 221329
rect 256617 221169 256633 221287
rect 256751 221169 256793 221287
rect 256911 221169 256927 221287
rect 256617 203447 256927 221169
rect 256617 203329 256633 203447
rect 256751 203329 256793 203447
rect 256911 203329 256927 203447
rect 256617 203287 256927 203329
rect 256617 203169 256633 203287
rect 256751 203169 256793 203287
rect 256911 203169 256927 203287
rect 256617 185447 256927 203169
rect 256617 185329 256633 185447
rect 256751 185329 256793 185447
rect 256911 185329 256927 185447
rect 256617 185287 256927 185329
rect 256617 185169 256633 185287
rect 256751 185169 256793 185287
rect 256911 185169 256927 185287
rect 256617 167447 256927 185169
rect 256617 167329 256633 167447
rect 256751 167329 256793 167447
rect 256911 167329 256927 167447
rect 256617 167287 256927 167329
rect 256617 167169 256633 167287
rect 256751 167169 256793 167287
rect 256911 167169 256927 167287
rect 256617 149447 256927 167169
rect 256617 149329 256633 149447
rect 256751 149329 256793 149447
rect 256911 149329 256927 149447
rect 256617 149287 256927 149329
rect 256617 149169 256633 149287
rect 256751 149169 256793 149287
rect 256911 149169 256927 149287
rect 256617 131447 256927 149169
rect 256617 131329 256633 131447
rect 256751 131329 256793 131447
rect 256911 131329 256927 131447
rect 256617 131287 256927 131329
rect 256617 131169 256633 131287
rect 256751 131169 256793 131287
rect 256911 131169 256927 131287
rect 256617 113447 256927 131169
rect 256617 113329 256633 113447
rect 256751 113329 256793 113447
rect 256911 113329 256927 113447
rect 256617 113287 256927 113329
rect 256617 113169 256633 113287
rect 256751 113169 256793 113287
rect 256911 113169 256927 113287
rect 256617 95447 256927 113169
rect 256617 95329 256633 95447
rect 256751 95329 256793 95447
rect 256911 95329 256927 95447
rect 256617 95287 256927 95329
rect 256617 95169 256633 95287
rect 256751 95169 256793 95287
rect 256911 95169 256927 95287
rect 256617 77447 256927 95169
rect 256617 77329 256633 77447
rect 256751 77329 256793 77447
rect 256911 77329 256927 77447
rect 256617 77287 256927 77329
rect 256617 77169 256633 77287
rect 256751 77169 256793 77287
rect 256911 77169 256927 77287
rect 256617 59447 256927 77169
rect 256617 59329 256633 59447
rect 256751 59329 256793 59447
rect 256911 59329 256927 59447
rect 256617 59287 256927 59329
rect 256617 59169 256633 59287
rect 256751 59169 256793 59287
rect 256911 59169 256927 59287
rect 256617 41447 256927 59169
rect 256617 41329 256633 41447
rect 256751 41329 256793 41447
rect 256911 41329 256927 41447
rect 256617 41287 256927 41329
rect 256617 41169 256633 41287
rect 256751 41169 256793 41287
rect 256911 41169 256927 41287
rect 256617 23447 256927 41169
rect 256617 23329 256633 23447
rect 256751 23329 256793 23447
rect 256911 23329 256927 23447
rect 256617 23287 256927 23329
rect 256617 23169 256633 23287
rect 256751 23169 256793 23287
rect 256911 23169 256927 23287
rect 256617 5447 256927 23169
rect 256617 5329 256633 5447
rect 256751 5329 256793 5447
rect 256911 5329 256927 5447
rect 256617 5287 256927 5329
rect 256617 5169 256633 5287
rect 256751 5169 256793 5287
rect 256911 5169 256927 5287
rect 256617 -2093 256927 5169
rect 256617 -2211 256633 -2093
rect 256751 -2211 256793 -2093
rect 256911 -2211 256927 -2093
rect 256617 -2253 256927 -2211
rect 256617 -2371 256633 -2253
rect 256751 -2371 256793 -2253
rect 256911 -2371 256927 -2253
rect 256617 -2867 256927 -2371
rect 258477 349307 258787 355021
rect 267477 355779 267787 355795
rect 267477 355661 267493 355779
rect 267611 355661 267653 355779
rect 267771 355661 267787 355779
rect 267477 355619 267787 355661
rect 267477 355501 267493 355619
rect 267611 355501 267653 355619
rect 267771 355501 267787 355619
rect 265617 354819 265927 354835
rect 265617 354701 265633 354819
rect 265751 354701 265793 354819
rect 265911 354701 265927 354819
rect 265617 354659 265927 354701
rect 265617 354541 265633 354659
rect 265751 354541 265793 354659
rect 265911 354541 265927 354659
rect 263757 353859 264067 353875
rect 263757 353741 263773 353859
rect 263891 353741 263933 353859
rect 264051 353741 264067 353859
rect 263757 353699 264067 353741
rect 263757 353581 263773 353699
rect 263891 353581 263933 353699
rect 264051 353581 264067 353699
rect 258477 349189 258493 349307
rect 258611 349189 258653 349307
rect 258771 349189 258787 349307
rect 258477 349147 258787 349189
rect 258477 349029 258493 349147
rect 258611 349029 258653 349147
rect 258771 349029 258787 349147
rect 258477 331307 258787 349029
rect 258477 331189 258493 331307
rect 258611 331189 258653 331307
rect 258771 331189 258787 331307
rect 258477 331147 258787 331189
rect 258477 331029 258493 331147
rect 258611 331029 258653 331147
rect 258771 331029 258787 331147
rect 258477 313307 258787 331029
rect 258477 313189 258493 313307
rect 258611 313189 258653 313307
rect 258771 313189 258787 313307
rect 258477 313147 258787 313189
rect 258477 313029 258493 313147
rect 258611 313029 258653 313147
rect 258771 313029 258787 313147
rect 258477 295307 258787 313029
rect 258477 295189 258493 295307
rect 258611 295189 258653 295307
rect 258771 295189 258787 295307
rect 258477 295147 258787 295189
rect 258477 295029 258493 295147
rect 258611 295029 258653 295147
rect 258771 295029 258787 295147
rect 258477 277307 258787 295029
rect 258477 277189 258493 277307
rect 258611 277189 258653 277307
rect 258771 277189 258787 277307
rect 258477 277147 258787 277189
rect 258477 277029 258493 277147
rect 258611 277029 258653 277147
rect 258771 277029 258787 277147
rect 258477 259307 258787 277029
rect 258477 259189 258493 259307
rect 258611 259189 258653 259307
rect 258771 259189 258787 259307
rect 258477 259147 258787 259189
rect 258477 259029 258493 259147
rect 258611 259029 258653 259147
rect 258771 259029 258787 259147
rect 258477 241307 258787 259029
rect 258477 241189 258493 241307
rect 258611 241189 258653 241307
rect 258771 241189 258787 241307
rect 258477 241147 258787 241189
rect 258477 241029 258493 241147
rect 258611 241029 258653 241147
rect 258771 241029 258787 241147
rect 258477 223307 258787 241029
rect 258477 223189 258493 223307
rect 258611 223189 258653 223307
rect 258771 223189 258787 223307
rect 258477 223147 258787 223189
rect 258477 223029 258493 223147
rect 258611 223029 258653 223147
rect 258771 223029 258787 223147
rect 258477 205307 258787 223029
rect 258477 205189 258493 205307
rect 258611 205189 258653 205307
rect 258771 205189 258787 205307
rect 258477 205147 258787 205189
rect 258477 205029 258493 205147
rect 258611 205029 258653 205147
rect 258771 205029 258787 205147
rect 258477 187307 258787 205029
rect 258477 187189 258493 187307
rect 258611 187189 258653 187307
rect 258771 187189 258787 187307
rect 258477 187147 258787 187189
rect 258477 187029 258493 187147
rect 258611 187029 258653 187147
rect 258771 187029 258787 187147
rect 258477 169307 258787 187029
rect 258477 169189 258493 169307
rect 258611 169189 258653 169307
rect 258771 169189 258787 169307
rect 258477 169147 258787 169189
rect 258477 169029 258493 169147
rect 258611 169029 258653 169147
rect 258771 169029 258787 169147
rect 258477 151307 258787 169029
rect 258477 151189 258493 151307
rect 258611 151189 258653 151307
rect 258771 151189 258787 151307
rect 258477 151147 258787 151189
rect 258477 151029 258493 151147
rect 258611 151029 258653 151147
rect 258771 151029 258787 151147
rect 258477 133307 258787 151029
rect 258477 133189 258493 133307
rect 258611 133189 258653 133307
rect 258771 133189 258787 133307
rect 258477 133147 258787 133189
rect 258477 133029 258493 133147
rect 258611 133029 258653 133147
rect 258771 133029 258787 133147
rect 258477 115307 258787 133029
rect 258477 115189 258493 115307
rect 258611 115189 258653 115307
rect 258771 115189 258787 115307
rect 258477 115147 258787 115189
rect 258477 115029 258493 115147
rect 258611 115029 258653 115147
rect 258771 115029 258787 115147
rect 258477 97307 258787 115029
rect 258477 97189 258493 97307
rect 258611 97189 258653 97307
rect 258771 97189 258787 97307
rect 258477 97147 258787 97189
rect 258477 97029 258493 97147
rect 258611 97029 258653 97147
rect 258771 97029 258787 97147
rect 258477 79307 258787 97029
rect 258477 79189 258493 79307
rect 258611 79189 258653 79307
rect 258771 79189 258787 79307
rect 258477 79147 258787 79189
rect 258477 79029 258493 79147
rect 258611 79029 258653 79147
rect 258771 79029 258787 79147
rect 258477 61307 258787 79029
rect 258477 61189 258493 61307
rect 258611 61189 258653 61307
rect 258771 61189 258787 61307
rect 258477 61147 258787 61189
rect 258477 61029 258493 61147
rect 258611 61029 258653 61147
rect 258771 61029 258787 61147
rect 258477 43307 258787 61029
rect 258477 43189 258493 43307
rect 258611 43189 258653 43307
rect 258771 43189 258787 43307
rect 258477 43147 258787 43189
rect 258477 43029 258493 43147
rect 258611 43029 258653 43147
rect 258771 43029 258787 43147
rect 258477 25307 258787 43029
rect 258477 25189 258493 25307
rect 258611 25189 258653 25307
rect 258771 25189 258787 25307
rect 258477 25147 258787 25189
rect 258477 25029 258493 25147
rect 258611 25029 258653 25147
rect 258771 25029 258787 25147
rect 258477 7307 258787 25029
rect 258477 7189 258493 7307
rect 258611 7189 258653 7307
rect 258771 7189 258787 7307
rect 258477 7147 258787 7189
rect 258477 7029 258493 7147
rect 258611 7029 258653 7147
rect 258771 7029 258787 7147
rect 249477 -3651 249493 -3533
rect 249611 -3651 249653 -3533
rect 249771 -3651 249787 -3533
rect 249477 -3693 249787 -3651
rect 249477 -3811 249493 -3693
rect 249611 -3811 249653 -3693
rect 249771 -3811 249787 -3693
rect 249477 -3827 249787 -3811
rect 258477 -3053 258787 7029
rect 261897 352899 262207 352915
rect 261897 352781 261913 352899
rect 262031 352781 262073 352899
rect 262191 352781 262207 352899
rect 261897 352739 262207 352781
rect 261897 352621 261913 352739
rect 262031 352621 262073 352739
rect 262191 352621 262207 352739
rect 261897 334727 262207 352621
rect 261897 334609 261913 334727
rect 262031 334609 262073 334727
rect 262191 334609 262207 334727
rect 261897 334567 262207 334609
rect 261897 334449 261913 334567
rect 262031 334449 262073 334567
rect 262191 334449 262207 334567
rect 261897 316727 262207 334449
rect 261897 316609 261913 316727
rect 262031 316609 262073 316727
rect 262191 316609 262207 316727
rect 261897 316567 262207 316609
rect 261897 316449 261913 316567
rect 262031 316449 262073 316567
rect 262191 316449 262207 316567
rect 261897 298727 262207 316449
rect 261897 298609 261913 298727
rect 262031 298609 262073 298727
rect 262191 298609 262207 298727
rect 261897 298567 262207 298609
rect 261897 298449 261913 298567
rect 262031 298449 262073 298567
rect 262191 298449 262207 298567
rect 261897 280727 262207 298449
rect 261897 280609 261913 280727
rect 262031 280609 262073 280727
rect 262191 280609 262207 280727
rect 261897 280567 262207 280609
rect 261897 280449 261913 280567
rect 262031 280449 262073 280567
rect 262191 280449 262207 280567
rect 261897 262727 262207 280449
rect 261897 262609 261913 262727
rect 262031 262609 262073 262727
rect 262191 262609 262207 262727
rect 261897 262567 262207 262609
rect 261897 262449 261913 262567
rect 262031 262449 262073 262567
rect 262191 262449 262207 262567
rect 261897 244727 262207 262449
rect 261897 244609 261913 244727
rect 262031 244609 262073 244727
rect 262191 244609 262207 244727
rect 261897 244567 262207 244609
rect 261897 244449 261913 244567
rect 262031 244449 262073 244567
rect 262191 244449 262207 244567
rect 261897 226727 262207 244449
rect 261897 226609 261913 226727
rect 262031 226609 262073 226727
rect 262191 226609 262207 226727
rect 261897 226567 262207 226609
rect 261897 226449 261913 226567
rect 262031 226449 262073 226567
rect 262191 226449 262207 226567
rect 261897 208727 262207 226449
rect 261897 208609 261913 208727
rect 262031 208609 262073 208727
rect 262191 208609 262207 208727
rect 261897 208567 262207 208609
rect 261897 208449 261913 208567
rect 262031 208449 262073 208567
rect 262191 208449 262207 208567
rect 261897 190727 262207 208449
rect 261897 190609 261913 190727
rect 262031 190609 262073 190727
rect 262191 190609 262207 190727
rect 261897 190567 262207 190609
rect 261897 190449 261913 190567
rect 262031 190449 262073 190567
rect 262191 190449 262207 190567
rect 261897 172727 262207 190449
rect 261897 172609 261913 172727
rect 262031 172609 262073 172727
rect 262191 172609 262207 172727
rect 261897 172567 262207 172609
rect 261897 172449 261913 172567
rect 262031 172449 262073 172567
rect 262191 172449 262207 172567
rect 261897 154727 262207 172449
rect 261897 154609 261913 154727
rect 262031 154609 262073 154727
rect 262191 154609 262207 154727
rect 261897 154567 262207 154609
rect 261897 154449 261913 154567
rect 262031 154449 262073 154567
rect 262191 154449 262207 154567
rect 261897 136727 262207 154449
rect 261897 136609 261913 136727
rect 262031 136609 262073 136727
rect 262191 136609 262207 136727
rect 261897 136567 262207 136609
rect 261897 136449 261913 136567
rect 262031 136449 262073 136567
rect 262191 136449 262207 136567
rect 261897 118727 262207 136449
rect 261897 118609 261913 118727
rect 262031 118609 262073 118727
rect 262191 118609 262207 118727
rect 261897 118567 262207 118609
rect 261897 118449 261913 118567
rect 262031 118449 262073 118567
rect 262191 118449 262207 118567
rect 261897 100727 262207 118449
rect 261897 100609 261913 100727
rect 262031 100609 262073 100727
rect 262191 100609 262207 100727
rect 261897 100567 262207 100609
rect 261897 100449 261913 100567
rect 262031 100449 262073 100567
rect 262191 100449 262207 100567
rect 261897 82727 262207 100449
rect 261897 82609 261913 82727
rect 262031 82609 262073 82727
rect 262191 82609 262207 82727
rect 261897 82567 262207 82609
rect 261897 82449 261913 82567
rect 262031 82449 262073 82567
rect 262191 82449 262207 82567
rect 261897 64727 262207 82449
rect 261897 64609 261913 64727
rect 262031 64609 262073 64727
rect 262191 64609 262207 64727
rect 261897 64567 262207 64609
rect 261897 64449 261913 64567
rect 262031 64449 262073 64567
rect 262191 64449 262207 64567
rect 261897 46727 262207 64449
rect 261897 46609 261913 46727
rect 262031 46609 262073 46727
rect 262191 46609 262207 46727
rect 261897 46567 262207 46609
rect 261897 46449 261913 46567
rect 262031 46449 262073 46567
rect 262191 46449 262207 46567
rect 261897 28727 262207 46449
rect 261897 28609 261913 28727
rect 262031 28609 262073 28727
rect 262191 28609 262207 28727
rect 261897 28567 262207 28609
rect 261897 28449 261913 28567
rect 262031 28449 262073 28567
rect 262191 28449 262207 28567
rect 261897 10727 262207 28449
rect 261897 10609 261913 10727
rect 262031 10609 262073 10727
rect 262191 10609 262207 10727
rect 261897 10567 262207 10609
rect 261897 10449 261913 10567
rect 262031 10449 262073 10567
rect 262191 10449 262207 10567
rect 261897 -653 262207 10449
rect 261897 -771 261913 -653
rect 262031 -771 262073 -653
rect 262191 -771 262207 -653
rect 261897 -813 262207 -771
rect 261897 -931 261913 -813
rect 262031 -931 262073 -813
rect 262191 -931 262207 -813
rect 261897 -947 262207 -931
rect 263757 336587 264067 353581
rect 263757 336469 263773 336587
rect 263891 336469 263933 336587
rect 264051 336469 264067 336587
rect 263757 336427 264067 336469
rect 263757 336309 263773 336427
rect 263891 336309 263933 336427
rect 264051 336309 264067 336427
rect 263757 318587 264067 336309
rect 263757 318469 263773 318587
rect 263891 318469 263933 318587
rect 264051 318469 264067 318587
rect 263757 318427 264067 318469
rect 263757 318309 263773 318427
rect 263891 318309 263933 318427
rect 264051 318309 264067 318427
rect 263757 300587 264067 318309
rect 263757 300469 263773 300587
rect 263891 300469 263933 300587
rect 264051 300469 264067 300587
rect 263757 300427 264067 300469
rect 263757 300309 263773 300427
rect 263891 300309 263933 300427
rect 264051 300309 264067 300427
rect 263757 282587 264067 300309
rect 263757 282469 263773 282587
rect 263891 282469 263933 282587
rect 264051 282469 264067 282587
rect 263757 282427 264067 282469
rect 263757 282309 263773 282427
rect 263891 282309 263933 282427
rect 264051 282309 264067 282427
rect 263757 264587 264067 282309
rect 263757 264469 263773 264587
rect 263891 264469 263933 264587
rect 264051 264469 264067 264587
rect 263757 264427 264067 264469
rect 263757 264309 263773 264427
rect 263891 264309 263933 264427
rect 264051 264309 264067 264427
rect 263757 246587 264067 264309
rect 263757 246469 263773 246587
rect 263891 246469 263933 246587
rect 264051 246469 264067 246587
rect 263757 246427 264067 246469
rect 263757 246309 263773 246427
rect 263891 246309 263933 246427
rect 264051 246309 264067 246427
rect 263757 228587 264067 246309
rect 263757 228469 263773 228587
rect 263891 228469 263933 228587
rect 264051 228469 264067 228587
rect 263757 228427 264067 228469
rect 263757 228309 263773 228427
rect 263891 228309 263933 228427
rect 264051 228309 264067 228427
rect 263757 210587 264067 228309
rect 263757 210469 263773 210587
rect 263891 210469 263933 210587
rect 264051 210469 264067 210587
rect 263757 210427 264067 210469
rect 263757 210309 263773 210427
rect 263891 210309 263933 210427
rect 264051 210309 264067 210427
rect 263757 192587 264067 210309
rect 263757 192469 263773 192587
rect 263891 192469 263933 192587
rect 264051 192469 264067 192587
rect 263757 192427 264067 192469
rect 263757 192309 263773 192427
rect 263891 192309 263933 192427
rect 264051 192309 264067 192427
rect 263757 174587 264067 192309
rect 263757 174469 263773 174587
rect 263891 174469 263933 174587
rect 264051 174469 264067 174587
rect 263757 174427 264067 174469
rect 263757 174309 263773 174427
rect 263891 174309 263933 174427
rect 264051 174309 264067 174427
rect 263757 156587 264067 174309
rect 263757 156469 263773 156587
rect 263891 156469 263933 156587
rect 264051 156469 264067 156587
rect 263757 156427 264067 156469
rect 263757 156309 263773 156427
rect 263891 156309 263933 156427
rect 264051 156309 264067 156427
rect 263757 138587 264067 156309
rect 263757 138469 263773 138587
rect 263891 138469 263933 138587
rect 264051 138469 264067 138587
rect 263757 138427 264067 138469
rect 263757 138309 263773 138427
rect 263891 138309 263933 138427
rect 264051 138309 264067 138427
rect 263757 120587 264067 138309
rect 263757 120469 263773 120587
rect 263891 120469 263933 120587
rect 264051 120469 264067 120587
rect 263757 120427 264067 120469
rect 263757 120309 263773 120427
rect 263891 120309 263933 120427
rect 264051 120309 264067 120427
rect 263757 102587 264067 120309
rect 263757 102469 263773 102587
rect 263891 102469 263933 102587
rect 264051 102469 264067 102587
rect 263757 102427 264067 102469
rect 263757 102309 263773 102427
rect 263891 102309 263933 102427
rect 264051 102309 264067 102427
rect 263757 84587 264067 102309
rect 263757 84469 263773 84587
rect 263891 84469 263933 84587
rect 264051 84469 264067 84587
rect 263757 84427 264067 84469
rect 263757 84309 263773 84427
rect 263891 84309 263933 84427
rect 264051 84309 264067 84427
rect 263757 66587 264067 84309
rect 263757 66469 263773 66587
rect 263891 66469 263933 66587
rect 264051 66469 264067 66587
rect 263757 66427 264067 66469
rect 263757 66309 263773 66427
rect 263891 66309 263933 66427
rect 264051 66309 264067 66427
rect 263757 48587 264067 66309
rect 263757 48469 263773 48587
rect 263891 48469 263933 48587
rect 264051 48469 264067 48587
rect 263757 48427 264067 48469
rect 263757 48309 263773 48427
rect 263891 48309 263933 48427
rect 264051 48309 264067 48427
rect 263757 30587 264067 48309
rect 263757 30469 263773 30587
rect 263891 30469 263933 30587
rect 264051 30469 264067 30587
rect 263757 30427 264067 30469
rect 263757 30309 263773 30427
rect 263891 30309 263933 30427
rect 264051 30309 264067 30427
rect 263757 12587 264067 30309
rect 263757 12469 263773 12587
rect 263891 12469 263933 12587
rect 264051 12469 264067 12587
rect 263757 12427 264067 12469
rect 263757 12309 263773 12427
rect 263891 12309 263933 12427
rect 264051 12309 264067 12427
rect 263757 -1613 264067 12309
rect 263757 -1731 263773 -1613
rect 263891 -1731 263933 -1613
rect 264051 -1731 264067 -1613
rect 263757 -1773 264067 -1731
rect 263757 -1891 263773 -1773
rect 263891 -1891 263933 -1773
rect 264051 -1891 264067 -1773
rect 263757 -1907 264067 -1891
rect 265617 338447 265927 354541
rect 265617 338329 265633 338447
rect 265751 338329 265793 338447
rect 265911 338329 265927 338447
rect 265617 338287 265927 338329
rect 265617 338169 265633 338287
rect 265751 338169 265793 338287
rect 265911 338169 265927 338287
rect 265617 320447 265927 338169
rect 265617 320329 265633 320447
rect 265751 320329 265793 320447
rect 265911 320329 265927 320447
rect 265617 320287 265927 320329
rect 265617 320169 265633 320287
rect 265751 320169 265793 320287
rect 265911 320169 265927 320287
rect 265617 302447 265927 320169
rect 265617 302329 265633 302447
rect 265751 302329 265793 302447
rect 265911 302329 265927 302447
rect 265617 302287 265927 302329
rect 265617 302169 265633 302287
rect 265751 302169 265793 302287
rect 265911 302169 265927 302287
rect 265617 284447 265927 302169
rect 265617 284329 265633 284447
rect 265751 284329 265793 284447
rect 265911 284329 265927 284447
rect 265617 284287 265927 284329
rect 265617 284169 265633 284287
rect 265751 284169 265793 284287
rect 265911 284169 265927 284287
rect 265617 266447 265927 284169
rect 265617 266329 265633 266447
rect 265751 266329 265793 266447
rect 265911 266329 265927 266447
rect 265617 266287 265927 266329
rect 265617 266169 265633 266287
rect 265751 266169 265793 266287
rect 265911 266169 265927 266287
rect 265617 248447 265927 266169
rect 265617 248329 265633 248447
rect 265751 248329 265793 248447
rect 265911 248329 265927 248447
rect 265617 248287 265927 248329
rect 265617 248169 265633 248287
rect 265751 248169 265793 248287
rect 265911 248169 265927 248287
rect 265617 230447 265927 248169
rect 265617 230329 265633 230447
rect 265751 230329 265793 230447
rect 265911 230329 265927 230447
rect 265617 230287 265927 230329
rect 265617 230169 265633 230287
rect 265751 230169 265793 230287
rect 265911 230169 265927 230287
rect 265617 212447 265927 230169
rect 265617 212329 265633 212447
rect 265751 212329 265793 212447
rect 265911 212329 265927 212447
rect 265617 212287 265927 212329
rect 265617 212169 265633 212287
rect 265751 212169 265793 212287
rect 265911 212169 265927 212287
rect 265617 194447 265927 212169
rect 265617 194329 265633 194447
rect 265751 194329 265793 194447
rect 265911 194329 265927 194447
rect 265617 194287 265927 194329
rect 265617 194169 265633 194287
rect 265751 194169 265793 194287
rect 265911 194169 265927 194287
rect 265617 176447 265927 194169
rect 265617 176329 265633 176447
rect 265751 176329 265793 176447
rect 265911 176329 265927 176447
rect 265617 176287 265927 176329
rect 265617 176169 265633 176287
rect 265751 176169 265793 176287
rect 265911 176169 265927 176287
rect 265617 158447 265927 176169
rect 265617 158329 265633 158447
rect 265751 158329 265793 158447
rect 265911 158329 265927 158447
rect 265617 158287 265927 158329
rect 265617 158169 265633 158287
rect 265751 158169 265793 158287
rect 265911 158169 265927 158287
rect 265617 140447 265927 158169
rect 265617 140329 265633 140447
rect 265751 140329 265793 140447
rect 265911 140329 265927 140447
rect 265617 140287 265927 140329
rect 265617 140169 265633 140287
rect 265751 140169 265793 140287
rect 265911 140169 265927 140287
rect 265617 122447 265927 140169
rect 265617 122329 265633 122447
rect 265751 122329 265793 122447
rect 265911 122329 265927 122447
rect 265617 122287 265927 122329
rect 265617 122169 265633 122287
rect 265751 122169 265793 122287
rect 265911 122169 265927 122287
rect 265617 104447 265927 122169
rect 265617 104329 265633 104447
rect 265751 104329 265793 104447
rect 265911 104329 265927 104447
rect 265617 104287 265927 104329
rect 265617 104169 265633 104287
rect 265751 104169 265793 104287
rect 265911 104169 265927 104287
rect 265617 86447 265927 104169
rect 265617 86329 265633 86447
rect 265751 86329 265793 86447
rect 265911 86329 265927 86447
rect 265617 86287 265927 86329
rect 265617 86169 265633 86287
rect 265751 86169 265793 86287
rect 265911 86169 265927 86287
rect 265617 68447 265927 86169
rect 265617 68329 265633 68447
rect 265751 68329 265793 68447
rect 265911 68329 265927 68447
rect 265617 68287 265927 68329
rect 265617 68169 265633 68287
rect 265751 68169 265793 68287
rect 265911 68169 265927 68287
rect 265617 50447 265927 68169
rect 265617 50329 265633 50447
rect 265751 50329 265793 50447
rect 265911 50329 265927 50447
rect 265617 50287 265927 50329
rect 265617 50169 265633 50287
rect 265751 50169 265793 50287
rect 265911 50169 265927 50287
rect 265617 32447 265927 50169
rect 265617 32329 265633 32447
rect 265751 32329 265793 32447
rect 265911 32329 265927 32447
rect 265617 32287 265927 32329
rect 265617 32169 265633 32287
rect 265751 32169 265793 32287
rect 265911 32169 265927 32287
rect 265617 14447 265927 32169
rect 265617 14329 265633 14447
rect 265751 14329 265793 14447
rect 265911 14329 265927 14447
rect 265617 14287 265927 14329
rect 265617 14169 265633 14287
rect 265751 14169 265793 14287
rect 265911 14169 265927 14287
rect 265617 -2573 265927 14169
rect 265617 -2691 265633 -2573
rect 265751 -2691 265793 -2573
rect 265911 -2691 265927 -2573
rect 265617 -2733 265927 -2691
rect 265617 -2851 265633 -2733
rect 265751 -2851 265793 -2733
rect 265911 -2851 265927 -2733
rect 265617 -2867 265927 -2851
rect 267477 340307 267787 355501
rect 276477 355299 276787 355795
rect 276477 355181 276493 355299
rect 276611 355181 276653 355299
rect 276771 355181 276787 355299
rect 276477 355139 276787 355181
rect 276477 355021 276493 355139
rect 276611 355021 276653 355139
rect 276771 355021 276787 355139
rect 274617 354339 274927 354835
rect 274617 354221 274633 354339
rect 274751 354221 274793 354339
rect 274911 354221 274927 354339
rect 274617 354179 274927 354221
rect 274617 354061 274633 354179
rect 274751 354061 274793 354179
rect 274911 354061 274927 354179
rect 272757 353379 273067 353875
rect 272757 353261 272773 353379
rect 272891 353261 272933 353379
rect 273051 353261 273067 353379
rect 272757 353219 273067 353261
rect 272757 353101 272773 353219
rect 272891 353101 272933 353219
rect 273051 353101 273067 353219
rect 267477 340189 267493 340307
rect 267611 340189 267653 340307
rect 267771 340189 267787 340307
rect 267477 340147 267787 340189
rect 267477 340029 267493 340147
rect 267611 340029 267653 340147
rect 267771 340029 267787 340147
rect 267477 322307 267787 340029
rect 267477 322189 267493 322307
rect 267611 322189 267653 322307
rect 267771 322189 267787 322307
rect 267477 322147 267787 322189
rect 267477 322029 267493 322147
rect 267611 322029 267653 322147
rect 267771 322029 267787 322147
rect 267477 304307 267787 322029
rect 267477 304189 267493 304307
rect 267611 304189 267653 304307
rect 267771 304189 267787 304307
rect 267477 304147 267787 304189
rect 267477 304029 267493 304147
rect 267611 304029 267653 304147
rect 267771 304029 267787 304147
rect 267477 286307 267787 304029
rect 267477 286189 267493 286307
rect 267611 286189 267653 286307
rect 267771 286189 267787 286307
rect 267477 286147 267787 286189
rect 267477 286029 267493 286147
rect 267611 286029 267653 286147
rect 267771 286029 267787 286147
rect 267477 268307 267787 286029
rect 267477 268189 267493 268307
rect 267611 268189 267653 268307
rect 267771 268189 267787 268307
rect 267477 268147 267787 268189
rect 267477 268029 267493 268147
rect 267611 268029 267653 268147
rect 267771 268029 267787 268147
rect 267477 250307 267787 268029
rect 267477 250189 267493 250307
rect 267611 250189 267653 250307
rect 267771 250189 267787 250307
rect 267477 250147 267787 250189
rect 267477 250029 267493 250147
rect 267611 250029 267653 250147
rect 267771 250029 267787 250147
rect 267477 232307 267787 250029
rect 267477 232189 267493 232307
rect 267611 232189 267653 232307
rect 267771 232189 267787 232307
rect 267477 232147 267787 232189
rect 267477 232029 267493 232147
rect 267611 232029 267653 232147
rect 267771 232029 267787 232147
rect 267477 214307 267787 232029
rect 267477 214189 267493 214307
rect 267611 214189 267653 214307
rect 267771 214189 267787 214307
rect 267477 214147 267787 214189
rect 267477 214029 267493 214147
rect 267611 214029 267653 214147
rect 267771 214029 267787 214147
rect 267477 196307 267787 214029
rect 267477 196189 267493 196307
rect 267611 196189 267653 196307
rect 267771 196189 267787 196307
rect 267477 196147 267787 196189
rect 267477 196029 267493 196147
rect 267611 196029 267653 196147
rect 267771 196029 267787 196147
rect 267477 178307 267787 196029
rect 267477 178189 267493 178307
rect 267611 178189 267653 178307
rect 267771 178189 267787 178307
rect 267477 178147 267787 178189
rect 267477 178029 267493 178147
rect 267611 178029 267653 178147
rect 267771 178029 267787 178147
rect 267477 160307 267787 178029
rect 267477 160189 267493 160307
rect 267611 160189 267653 160307
rect 267771 160189 267787 160307
rect 267477 160147 267787 160189
rect 267477 160029 267493 160147
rect 267611 160029 267653 160147
rect 267771 160029 267787 160147
rect 267477 142307 267787 160029
rect 267477 142189 267493 142307
rect 267611 142189 267653 142307
rect 267771 142189 267787 142307
rect 267477 142147 267787 142189
rect 267477 142029 267493 142147
rect 267611 142029 267653 142147
rect 267771 142029 267787 142147
rect 267477 124307 267787 142029
rect 267477 124189 267493 124307
rect 267611 124189 267653 124307
rect 267771 124189 267787 124307
rect 267477 124147 267787 124189
rect 267477 124029 267493 124147
rect 267611 124029 267653 124147
rect 267771 124029 267787 124147
rect 267477 106307 267787 124029
rect 267477 106189 267493 106307
rect 267611 106189 267653 106307
rect 267771 106189 267787 106307
rect 267477 106147 267787 106189
rect 267477 106029 267493 106147
rect 267611 106029 267653 106147
rect 267771 106029 267787 106147
rect 267477 88307 267787 106029
rect 267477 88189 267493 88307
rect 267611 88189 267653 88307
rect 267771 88189 267787 88307
rect 267477 88147 267787 88189
rect 267477 88029 267493 88147
rect 267611 88029 267653 88147
rect 267771 88029 267787 88147
rect 267477 70307 267787 88029
rect 267477 70189 267493 70307
rect 267611 70189 267653 70307
rect 267771 70189 267787 70307
rect 267477 70147 267787 70189
rect 267477 70029 267493 70147
rect 267611 70029 267653 70147
rect 267771 70029 267787 70147
rect 267477 52307 267787 70029
rect 267477 52189 267493 52307
rect 267611 52189 267653 52307
rect 267771 52189 267787 52307
rect 267477 52147 267787 52189
rect 267477 52029 267493 52147
rect 267611 52029 267653 52147
rect 267771 52029 267787 52147
rect 267477 34307 267787 52029
rect 267477 34189 267493 34307
rect 267611 34189 267653 34307
rect 267771 34189 267787 34307
rect 267477 34147 267787 34189
rect 267477 34029 267493 34147
rect 267611 34029 267653 34147
rect 267771 34029 267787 34147
rect 267477 16307 267787 34029
rect 267477 16189 267493 16307
rect 267611 16189 267653 16307
rect 267771 16189 267787 16307
rect 267477 16147 267787 16189
rect 267477 16029 267493 16147
rect 267611 16029 267653 16147
rect 267771 16029 267787 16147
rect 258477 -3171 258493 -3053
rect 258611 -3171 258653 -3053
rect 258771 -3171 258787 -3053
rect 258477 -3213 258787 -3171
rect 258477 -3331 258493 -3213
rect 258611 -3331 258653 -3213
rect 258771 -3331 258787 -3213
rect 258477 -3827 258787 -3331
rect 267477 -3533 267787 16029
rect 270897 352419 271207 352915
rect 270897 352301 270913 352419
rect 271031 352301 271073 352419
rect 271191 352301 271207 352419
rect 270897 352259 271207 352301
rect 270897 352141 270913 352259
rect 271031 352141 271073 352259
rect 271191 352141 271207 352259
rect 270897 343727 271207 352141
rect 270897 343609 270913 343727
rect 271031 343609 271073 343727
rect 271191 343609 271207 343727
rect 270897 343567 271207 343609
rect 270897 343449 270913 343567
rect 271031 343449 271073 343567
rect 271191 343449 271207 343567
rect 270897 325727 271207 343449
rect 270897 325609 270913 325727
rect 271031 325609 271073 325727
rect 271191 325609 271207 325727
rect 270897 325567 271207 325609
rect 270897 325449 270913 325567
rect 271031 325449 271073 325567
rect 271191 325449 271207 325567
rect 270897 307727 271207 325449
rect 270897 307609 270913 307727
rect 271031 307609 271073 307727
rect 271191 307609 271207 307727
rect 270897 307567 271207 307609
rect 270897 307449 270913 307567
rect 271031 307449 271073 307567
rect 271191 307449 271207 307567
rect 270897 289727 271207 307449
rect 270897 289609 270913 289727
rect 271031 289609 271073 289727
rect 271191 289609 271207 289727
rect 270897 289567 271207 289609
rect 270897 289449 270913 289567
rect 271031 289449 271073 289567
rect 271191 289449 271207 289567
rect 270897 271727 271207 289449
rect 270897 271609 270913 271727
rect 271031 271609 271073 271727
rect 271191 271609 271207 271727
rect 270897 271567 271207 271609
rect 270897 271449 270913 271567
rect 271031 271449 271073 271567
rect 271191 271449 271207 271567
rect 270897 253727 271207 271449
rect 270897 253609 270913 253727
rect 271031 253609 271073 253727
rect 271191 253609 271207 253727
rect 270897 253567 271207 253609
rect 270897 253449 270913 253567
rect 271031 253449 271073 253567
rect 271191 253449 271207 253567
rect 270897 235727 271207 253449
rect 270897 235609 270913 235727
rect 271031 235609 271073 235727
rect 271191 235609 271207 235727
rect 270897 235567 271207 235609
rect 270897 235449 270913 235567
rect 271031 235449 271073 235567
rect 271191 235449 271207 235567
rect 270897 217727 271207 235449
rect 270897 217609 270913 217727
rect 271031 217609 271073 217727
rect 271191 217609 271207 217727
rect 270897 217567 271207 217609
rect 270897 217449 270913 217567
rect 271031 217449 271073 217567
rect 271191 217449 271207 217567
rect 270897 199727 271207 217449
rect 270897 199609 270913 199727
rect 271031 199609 271073 199727
rect 271191 199609 271207 199727
rect 270897 199567 271207 199609
rect 270897 199449 270913 199567
rect 271031 199449 271073 199567
rect 271191 199449 271207 199567
rect 270897 181727 271207 199449
rect 270897 181609 270913 181727
rect 271031 181609 271073 181727
rect 271191 181609 271207 181727
rect 270897 181567 271207 181609
rect 270897 181449 270913 181567
rect 271031 181449 271073 181567
rect 271191 181449 271207 181567
rect 270897 163727 271207 181449
rect 270897 163609 270913 163727
rect 271031 163609 271073 163727
rect 271191 163609 271207 163727
rect 270897 163567 271207 163609
rect 270897 163449 270913 163567
rect 271031 163449 271073 163567
rect 271191 163449 271207 163567
rect 270897 145727 271207 163449
rect 270897 145609 270913 145727
rect 271031 145609 271073 145727
rect 271191 145609 271207 145727
rect 270897 145567 271207 145609
rect 270897 145449 270913 145567
rect 271031 145449 271073 145567
rect 271191 145449 271207 145567
rect 270897 127727 271207 145449
rect 270897 127609 270913 127727
rect 271031 127609 271073 127727
rect 271191 127609 271207 127727
rect 270897 127567 271207 127609
rect 270897 127449 270913 127567
rect 271031 127449 271073 127567
rect 271191 127449 271207 127567
rect 270897 109727 271207 127449
rect 270897 109609 270913 109727
rect 271031 109609 271073 109727
rect 271191 109609 271207 109727
rect 270897 109567 271207 109609
rect 270897 109449 270913 109567
rect 271031 109449 271073 109567
rect 271191 109449 271207 109567
rect 270897 91727 271207 109449
rect 270897 91609 270913 91727
rect 271031 91609 271073 91727
rect 271191 91609 271207 91727
rect 270897 91567 271207 91609
rect 270897 91449 270913 91567
rect 271031 91449 271073 91567
rect 271191 91449 271207 91567
rect 270897 73727 271207 91449
rect 270897 73609 270913 73727
rect 271031 73609 271073 73727
rect 271191 73609 271207 73727
rect 270897 73567 271207 73609
rect 270897 73449 270913 73567
rect 271031 73449 271073 73567
rect 271191 73449 271207 73567
rect 270897 55727 271207 73449
rect 270897 55609 270913 55727
rect 271031 55609 271073 55727
rect 271191 55609 271207 55727
rect 270897 55567 271207 55609
rect 270897 55449 270913 55567
rect 271031 55449 271073 55567
rect 271191 55449 271207 55567
rect 270897 37727 271207 55449
rect 270897 37609 270913 37727
rect 271031 37609 271073 37727
rect 271191 37609 271207 37727
rect 270897 37567 271207 37609
rect 270897 37449 270913 37567
rect 271031 37449 271073 37567
rect 271191 37449 271207 37567
rect 270897 19727 271207 37449
rect 270897 19609 270913 19727
rect 271031 19609 271073 19727
rect 271191 19609 271207 19727
rect 270897 19567 271207 19609
rect 270897 19449 270913 19567
rect 271031 19449 271073 19567
rect 271191 19449 271207 19567
rect 270897 1727 271207 19449
rect 270897 1609 270913 1727
rect 271031 1609 271073 1727
rect 271191 1609 271207 1727
rect 270897 1567 271207 1609
rect 270897 1449 270913 1567
rect 271031 1449 271073 1567
rect 271191 1449 271207 1567
rect 270897 -173 271207 1449
rect 270897 -291 270913 -173
rect 271031 -291 271073 -173
rect 271191 -291 271207 -173
rect 270897 -333 271207 -291
rect 270897 -451 270913 -333
rect 271031 -451 271073 -333
rect 271191 -451 271207 -333
rect 270897 -947 271207 -451
rect 272757 345587 273067 353101
rect 272757 345469 272773 345587
rect 272891 345469 272933 345587
rect 273051 345469 273067 345587
rect 272757 345427 273067 345469
rect 272757 345309 272773 345427
rect 272891 345309 272933 345427
rect 273051 345309 273067 345427
rect 272757 327587 273067 345309
rect 272757 327469 272773 327587
rect 272891 327469 272933 327587
rect 273051 327469 273067 327587
rect 272757 327427 273067 327469
rect 272757 327309 272773 327427
rect 272891 327309 272933 327427
rect 273051 327309 273067 327427
rect 272757 309587 273067 327309
rect 272757 309469 272773 309587
rect 272891 309469 272933 309587
rect 273051 309469 273067 309587
rect 272757 309427 273067 309469
rect 272757 309309 272773 309427
rect 272891 309309 272933 309427
rect 273051 309309 273067 309427
rect 272757 291587 273067 309309
rect 272757 291469 272773 291587
rect 272891 291469 272933 291587
rect 273051 291469 273067 291587
rect 272757 291427 273067 291469
rect 272757 291309 272773 291427
rect 272891 291309 272933 291427
rect 273051 291309 273067 291427
rect 272757 273587 273067 291309
rect 272757 273469 272773 273587
rect 272891 273469 272933 273587
rect 273051 273469 273067 273587
rect 272757 273427 273067 273469
rect 272757 273309 272773 273427
rect 272891 273309 272933 273427
rect 273051 273309 273067 273427
rect 272757 255587 273067 273309
rect 272757 255469 272773 255587
rect 272891 255469 272933 255587
rect 273051 255469 273067 255587
rect 272757 255427 273067 255469
rect 272757 255309 272773 255427
rect 272891 255309 272933 255427
rect 273051 255309 273067 255427
rect 272757 237587 273067 255309
rect 272757 237469 272773 237587
rect 272891 237469 272933 237587
rect 273051 237469 273067 237587
rect 272757 237427 273067 237469
rect 272757 237309 272773 237427
rect 272891 237309 272933 237427
rect 273051 237309 273067 237427
rect 272757 219587 273067 237309
rect 272757 219469 272773 219587
rect 272891 219469 272933 219587
rect 273051 219469 273067 219587
rect 272757 219427 273067 219469
rect 272757 219309 272773 219427
rect 272891 219309 272933 219427
rect 273051 219309 273067 219427
rect 272757 201587 273067 219309
rect 272757 201469 272773 201587
rect 272891 201469 272933 201587
rect 273051 201469 273067 201587
rect 272757 201427 273067 201469
rect 272757 201309 272773 201427
rect 272891 201309 272933 201427
rect 273051 201309 273067 201427
rect 272757 183587 273067 201309
rect 272757 183469 272773 183587
rect 272891 183469 272933 183587
rect 273051 183469 273067 183587
rect 272757 183427 273067 183469
rect 272757 183309 272773 183427
rect 272891 183309 272933 183427
rect 273051 183309 273067 183427
rect 272757 165587 273067 183309
rect 272757 165469 272773 165587
rect 272891 165469 272933 165587
rect 273051 165469 273067 165587
rect 272757 165427 273067 165469
rect 272757 165309 272773 165427
rect 272891 165309 272933 165427
rect 273051 165309 273067 165427
rect 272757 147587 273067 165309
rect 272757 147469 272773 147587
rect 272891 147469 272933 147587
rect 273051 147469 273067 147587
rect 272757 147427 273067 147469
rect 272757 147309 272773 147427
rect 272891 147309 272933 147427
rect 273051 147309 273067 147427
rect 272757 129587 273067 147309
rect 272757 129469 272773 129587
rect 272891 129469 272933 129587
rect 273051 129469 273067 129587
rect 272757 129427 273067 129469
rect 272757 129309 272773 129427
rect 272891 129309 272933 129427
rect 273051 129309 273067 129427
rect 272757 111587 273067 129309
rect 272757 111469 272773 111587
rect 272891 111469 272933 111587
rect 273051 111469 273067 111587
rect 272757 111427 273067 111469
rect 272757 111309 272773 111427
rect 272891 111309 272933 111427
rect 273051 111309 273067 111427
rect 272757 93587 273067 111309
rect 272757 93469 272773 93587
rect 272891 93469 272933 93587
rect 273051 93469 273067 93587
rect 272757 93427 273067 93469
rect 272757 93309 272773 93427
rect 272891 93309 272933 93427
rect 273051 93309 273067 93427
rect 272757 75587 273067 93309
rect 272757 75469 272773 75587
rect 272891 75469 272933 75587
rect 273051 75469 273067 75587
rect 272757 75427 273067 75469
rect 272757 75309 272773 75427
rect 272891 75309 272933 75427
rect 273051 75309 273067 75427
rect 272757 57587 273067 75309
rect 272757 57469 272773 57587
rect 272891 57469 272933 57587
rect 273051 57469 273067 57587
rect 272757 57427 273067 57469
rect 272757 57309 272773 57427
rect 272891 57309 272933 57427
rect 273051 57309 273067 57427
rect 272757 39587 273067 57309
rect 272757 39469 272773 39587
rect 272891 39469 272933 39587
rect 273051 39469 273067 39587
rect 272757 39427 273067 39469
rect 272757 39309 272773 39427
rect 272891 39309 272933 39427
rect 273051 39309 273067 39427
rect 272757 21587 273067 39309
rect 272757 21469 272773 21587
rect 272891 21469 272933 21587
rect 273051 21469 273067 21587
rect 272757 21427 273067 21469
rect 272757 21309 272773 21427
rect 272891 21309 272933 21427
rect 273051 21309 273067 21427
rect 272757 3587 273067 21309
rect 272757 3469 272773 3587
rect 272891 3469 272933 3587
rect 273051 3469 273067 3587
rect 272757 3427 273067 3469
rect 272757 3309 272773 3427
rect 272891 3309 272933 3427
rect 273051 3309 273067 3427
rect 272757 -1133 273067 3309
rect 272757 -1251 272773 -1133
rect 272891 -1251 272933 -1133
rect 273051 -1251 273067 -1133
rect 272757 -1293 273067 -1251
rect 272757 -1411 272773 -1293
rect 272891 -1411 272933 -1293
rect 273051 -1411 273067 -1293
rect 272757 -1907 273067 -1411
rect 274617 347447 274927 354061
rect 274617 347329 274633 347447
rect 274751 347329 274793 347447
rect 274911 347329 274927 347447
rect 274617 347287 274927 347329
rect 274617 347169 274633 347287
rect 274751 347169 274793 347287
rect 274911 347169 274927 347287
rect 274617 329447 274927 347169
rect 274617 329329 274633 329447
rect 274751 329329 274793 329447
rect 274911 329329 274927 329447
rect 274617 329287 274927 329329
rect 274617 329169 274633 329287
rect 274751 329169 274793 329287
rect 274911 329169 274927 329287
rect 274617 311447 274927 329169
rect 274617 311329 274633 311447
rect 274751 311329 274793 311447
rect 274911 311329 274927 311447
rect 274617 311287 274927 311329
rect 274617 311169 274633 311287
rect 274751 311169 274793 311287
rect 274911 311169 274927 311287
rect 274617 293447 274927 311169
rect 274617 293329 274633 293447
rect 274751 293329 274793 293447
rect 274911 293329 274927 293447
rect 274617 293287 274927 293329
rect 274617 293169 274633 293287
rect 274751 293169 274793 293287
rect 274911 293169 274927 293287
rect 274617 275447 274927 293169
rect 274617 275329 274633 275447
rect 274751 275329 274793 275447
rect 274911 275329 274927 275447
rect 274617 275287 274927 275329
rect 274617 275169 274633 275287
rect 274751 275169 274793 275287
rect 274911 275169 274927 275287
rect 274617 257447 274927 275169
rect 274617 257329 274633 257447
rect 274751 257329 274793 257447
rect 274911 257329 274927 257447
rect 274617 257287 274927 257329
rect 274617 257169 274633 257287
rect 274751 257169 274793 257287
rect 274911 257169 274927 257287
rect 274617 239447 274927 257169
rect 274617 239329 274633 239447
rect 274751 239329 274793 239447
rect 274911 239329 274927 239447
rect 274617 239287 274927 239329
rect 274617 239169 274633 239287
rect 274751 239169 274793 239287
rect 274911 239169 274927 239287
rect 274617 221447 274927 239169
rect 274617 221329 274633 221447
rect 274751 221329 274793 221447
rect 274911 221329 274927 221447
rect 274617 221287 274927 221329
rect 274617 221169 274633 221287
rect 274751 221169 274793 221287
rect 274911 221169 274927 221287
rect 274617 203447 274927 221169
rect 274617 203329 274633 203447
rect 274751 203329 274793 203447
rect 274911 203329 274927 203447
rect 274617 203287 274927 203329
rect 274617 203169 274633 203287
rect 274751 203169 274793 203287
rect 274911 203169 274927 203287
rect 274617 185447 274927 203169
rect 274617 185329 274633 185447
rect 274751 185329 274793 185447
rect 274911 185329 274927 185447
rect 274617 185287 274927 185329
rect 274617 185169 274633 185287
rect 274751 185169 274793 185287
rect 274911 185169 274927 185287
rect 274617 167447 274927 185169
rect 274617 167329 274633 167447
rect 274751 167329 274793 167447
rect 274911 167329 274927 167447
rect 274617 167287 274927 167329
rect 274617 167169 274633 167287
rect 274751 167169 274793 167287
rect 274911 167169 274927 167287
rect 274617 149447 274927 167169
rect 274617 149329 274633 149447
rect 274751 149329 274793 149447
rect 274911 149329 274927 149447
rect 274617 149287 274927 149329
rect 274617 149169 274633 149287
rect 274751 149169 274793 149287
rect 274911 149169 274927 149287
rect 274617 131447 274927 149169
rect 274617 131329 274633 131447
rect 274751 131329 274793 131447
rect 274911 131329 274927 131447
rect 274617 131287 274927 131329
rect 274617 131169 274633 131287
rect 274751 131169 274793 131287
rect 274911 131169 274927 131287
rect 274617 113447 274927 131169
rect 274617 113329 274633 113447
rect 274751 113329 274793 113447
rect 274911 113329 274927 113447
rect 274617 113287 274927 113329
rect 274617 113169 274633 113287
rect 274751 113169 274793 113287
rect 274911 113169 274927 113287
rect 274617 95447 274927 113169
rect 274617 95329 274633 95447
rect 274751 95329 274793 95447
rect 274911 95329 274927 95447
rect 274617 95287 274927 95329
rect 274617 95169 274633 95287
rect 274751 95169 274793 95287
rect 274911 95169 274927 95287
rect 274617 77447 274927 95169
rect 274617 77329 274633 77447
rect 274751 77329 274793 77447
rect 274911 77329 274927 77447
rect 274617 77287 274927 77329
rect 274617 77169 274633 77287
rect 274751 77169 274793 77287
rect 274911 77169 274927 77287
rect 274617 59447 274927 77169
rect 274617 59329 274633 59447
rect 274751 59329 274793 59447
rect 274911 59329 274927 59447
rect 274617 59287 274927 59329
rect 274617 59169 274633 59287
rect 274751 59169 274793 59287
rect 274911 59169 274927 59287
rect 274617 41447 274927 59169
rect 274617 41329 274633 41447
rect 274751 41329 274793 41447
rect 274911 41329 274927 41447
rect 274617 41287 274927 41329
rect 274617 41169 274633 41287
rect 274751 41169 274793 41287
rect 274911 41169 274927 41287
rect 274617 23447 274927 41169
rect 274617 23329 274633 23447
rect 274751 23329 274793 23447
rect 274911 23329 274927 23447
rect 274617 23287 274927 23329
rect 274617 23169 274633 23287
rect 274751 23169 274793 23287
rect 274911 23169 274927 23287
rect 274617 5447 274927 23169
rect 274617 5329 274633 5447
rect 274751 5329 274793 5447
rect 274911 5329 274927 5447
rect 274617 5287 274927 5329
rect 274617 5169 274633 5287
rect 274751 5169 274793 5287
rect 274911 5169 274927 5287
rect 274617 -2093 274927 5169
rect 274617 -2211 274633 -2093
rect 274751 -2211 274793 -2093
rect 274911 -2211 274927 -2093
rect 274617 -2253 274927 -2211
rect 274617 -2371 274633 -2253
rect 274751 -2371 274793 -2253
rect 274911 -2371 274927 -2253
rect 274617 -2867 274927 -2371
rect 276477 349307 276787 355021
rect 285477 355779 285787 355795
rect 285477 355661 285493 355779
rect 285611 355661 285653 355779
rect 285771 355661 285787 355779
rect 285477 355619 285787 355661
rect 285477 355501 285493 355619
rect 285611 355501 285653 355619
rect 285771 355501 285787 355619
rect 283617 354819 283927 354835
rect 283617 354701 283633 354819
rect 283751 354701 283793 354819
rect 283911 354701 283927 354819
rect 283617 354659 283927 354701
rect 283617 354541 283633 354659
rect 283751 354541 283793 354659
rect 283911 354541 283927 354659
rect 281757 353859 282067 353875
rect 281757 353741 281773 353859
rect 281891 353741 281933 353859
rect 282051 353741 282067 353859
rect 281757 353699 282067 353741
rect 281757 353581 281773 353699
rect 281891 353581 281933 353699
rect 282051 353581 282067 353699
rect 276477 349189 276493 349307
rect 276611 349189 276653 349307
rect 276771 349189 276787 349307
rect 276477 349147 276787 349189
rect 276477 349029 276493 349147
rect 276611 349029 276653 349147
rect 276771 349029 276787 349147
rect 276477 331307 276787 349029
rect 276477 331189 276493 331307
rect 276611 331189 276653 331307
rect 276771 331189 276787 331307
rect 276477 331147 276787 331189
rect 276477 331029 276493 331147
rect 276611 331029 276653 331147
rect 276771 331029 276787 331147
rect 276477 313307 276787 331029
rect 276477 313189 276493 313307
rect 276611 313189 276653 313307
rect 276771 313189 276787 313307
rect 276477 313147 276787 313189
rect 276477 313029 276493 313147
rect 276611 313029 276653 313147
rect 276771 313029 276787 313147
rect 276477 295307 276787 313029
rect 276477 295189 276493 295307
rect 276611 295189 276653 295307
rect 276771 295189 276787 295307
rect 276477 295147 276787 295189
rect 276477 295029 276493 295147
rect 276611 295029 276653 295147
rect 276771 295029 276787 295147
rect 276477 277307 276787 295029
rect 276477 277189 276493 277307
rect 276611 277189 276653 277307
rect 276771 277189 276787 277307
rect 276477 277147 276787 277189
rect 276477 277029 276493 277147
rect 276611 277029 276653 277147
rect 276771 277029 276787 277147
rect 276477 259307 276787 277029
rect 276477 259189 276493 259307
rect 276611 259189 276653 259307
rect 276771 259189 276787 259307
rect 276477 259147 276787 259189
rect 276477 259029 276493 259147
rect 276611 259029 276653 259147
rect 276771 259029 276787 259147
rect 276477 241307 276787 259029
rect 276477 241189 276493 241307
rect 276611 241189 276653 241307
rect 276771 241189 276787 241307
rect 276477 241147 276787 241189
rect 276477 241029 276493 241147
rect 276611 241029 276653 241147
rect 276771 241029 276787 241147
rect 276477 223307 276787 241029
rect 276477 223189 276493 223307
rect 276611 223189 276653 223307
rect 276771 223189 276787 223307
rect 276477 223147 276787 223189
rect 276477 223029 276493 223147
rect 276611 223029 276653 223147
rect 276771 223029 276787 223147
rect 276477 205307 276787 223029
rect 276477 205189 276493 205307
rect 276611 205189 276653 205307
rect 276771 205189 276787 205307
rect 276477 205147 276787 205189
rect 276477 205029 276493 205147
rect 276611 205029 276653 205147
rect 276771 205029 276787 205147
rect 276477 187307 276787 205029
rect 276477 187189 276493 187307
rect 276611 187189 276653 187307
rect 276771 187189 276787 187307
rect 276477 187147 276787 187189
rect 276477 187029 276493 187147
rect 276611 187029 276653 187147
rect 276771 187029 276787 187147
rect 276477 169307 276787 187029
rect 276477 169189 276493 169307
rect 276611 169189 276653 169307
rect 276771 169189 276787 169307
rect 276477 169147 276787 169189
rect 276477 169029 276493 169147
rect 276611 169029 276653 169147
rect 276771 169029 276787 169147
rect 276477 151307 276787 169029
rect 276477 151189 276493 151307
rect 276611 151189 276653 151307
rect 276771 151189 276787 151307
rect 276477 151147 276787 151189
rect 276477 151029 276493 151147
rect 276611 151029 276653 151147
rect 276771 151029 276787 151147
rect 276477 133307 276787 151029
rect 276477 133189 276493 133307
rect 276611 133189 276653 133307
rect 276771 133189 276787 133307
rect 276477 133147 276787 133189
rect 276477 133029 276493 133147
rect 276611 133029 276653 133147
rect 276771 133029 276787 133147
rect 276477 115307 276787 133029
rect 276477 115189 276493 115307
rect 276611 115189 276653 115307
rect 276771 115189 276787 115307
rect 276477 115147 276787 115189
rect 276477 115029 276493 115147
rect 276611 115029 276653 115147
rect 276771 115029 276787 115147
rect 276477 97307 276787 115029
rect 276477 97189 276493 97307
rect 276611 97189 276653 97307
rect 276771 97189 276787 97307
rect 276477 97147 276787 97189
rect 276477 97029 276493 97147
rect 276611 97029 276653 97147
rect 276771 97029 276787 97147
rect 276477 79307 276787 97029
rect 276477 79189 276493 79307
rect 276611 79189 276653 79307
rect 276771 79189 276787 79307
rect 276477 79147 276787 79189
rect 276477 79029 276493 79147
rect 276611 79029 276653 79147
rect 276771 79029 276787 79147
rect 276477 61307 276787 79029
rect 276477 61189 276493 61307
rect 276611 61189 276653 61307
rect 276771 61189 276787 61307
rect 276477 61147 276787 61189
rect 276477 61029 276493 61147
rect 276611 61029 276653 61147
rect 276771 61029 276787 61147
rect 276477 43307 276787 61029
rect 276477 43189 276493 43307
rect 276611 43189 276653 43307
rect 276771 43189 276787 43307
rect 276477 43147 276787 43189
rect 276477 43029 276493 43147
rect 276611 43029 276653 43147
rect 276771 43029 276787 43147
rect 276477 25307 276787 43029
rect 276477 25189 276493 25307
rect 276611 25189 276653 25307
rect 276771 25189 276787 25307
rect 276477 25147 276787 25189
rect 276477 25029 276493 25147
rect 276611 25029 276653 25147
rect 276771 25029 276787 25147
rect 276477 7307 276787 25029
rect 276477 7189 276493 7307
rect 276611 7189 276653 7307
rect 276771 7189 276787 7307
rect 276477 7147 276787 7189
rect 276477 7029 276493 7147
rect 276611 7029 276653 7147
rect 276771 7029 276787 7147
rect 267477 -3651 267493 -3533
rect 267611 -3651 267653 -3533
rect 267771 -3651 267787 -3533
rect 267477 -3693 267787 -3651
rect 267477 -3811 267493 -3693
rect 267611 -3811 267653 -3693
rect 267771 -3811 267787 -3693
rect 267477 -3827 267787 -3811
rect 276477 -3053 276787 7029
rect 279897 352899 280207 352915
rect 279897 352781 279913 352899
rect 280031 352781 280073 352899
rect 280191 352781 280207 352899
rect 279897 352739 280207 352781
rect 279897 352621 279913 352739
rect 280031 352621 280073 352739
rect 280191 352621 280207 352739
rect 279897 334727 280207 352621
rect 279897 334609 279913 334727
rect 280031 334609 280073 334727
rect 280191 334609 280207 334727
rect 279897 334567 280207 334609
rect 279897 334449 279913 334567
rect 280031 334449 280073 334567
rect 280191 334449 280207 334567
rect 279897 316727 280207 334449
rect 279897 316609 279913 316727
rect 280031 316609 280073 316727
rect 280191 316609 280207 316727
rect 279897 316567 280207 316609
rect 279897 316449 279913 316567
rect 280031 316449 280073 316567
rect 280191 316449 280207 316567
rect 279897 298727 280207 316449
rect 279897 298609 279913 298727
rect 280031 298609 280073 298727
rect 280191 298609 280207 298727
rect 279897 298567 280207 298609
rect 279897 298449 279913 298567
rect 280031 298449 280073 298567
rect 280191 298449 280207 298567
rect 279897 280727 280207 298449
rect 279897 280609 279913 280727
rect 280031 280609 280073 280727
rect 280191 280609 280207 280727
rect 279897 280567 280207 280609
rect 279897 280449 279913 280567
rect 280031 280449 280073 280567
rect 280191 280449 280207 280567
rect 279897 262727 280207 280449
rect 279897 262609 279913 262727
rect 280031 262609 280073 262727
rect 280191 262609 280207 262727
rect 279897 262567 280207 262609
rect 279897 262449 279913 262567
rect 280031 262449 280073 262567
rect 280191 262449 280207 262567
rect 279897 244727 280207 262449
rect 279897 244609 279913 244727
rect 280031 244609 280073 244727
rect 280191 244609 280207 244727
rect 279897 244567 280207 244609
rect 279897 244449 279913 244567
rect 280031 244449 280073 244567
rect 280191 244449 280207 244567
rect 279897 226727 280207 244449
rect 279897 226609 279913 226727
rect 280031 226609 280073 226727
rect 280191 226609 280207 226727
rect 279897 226567 280207 226609
rect 279897 226449 279913 226567
rect 280031 226449 280073 226567
rect 280191 226449 280207 226567
rect 279897 208727 280207 226449
rect 279897 208609 279913 208727
rect 280031 208609 280073 208727
rect 280191 208609 280207 208727
rect 279897 208567 280207 208609
rect 279897 208449 279913 208567
rect 280031 208449 280073 208567
rect 280191 208449 280207 208567
rect 279897 190727 280207 208449
rect 279897 190609 279913 190727
rect 280031 190609 280073 190727
rect 280191 190609 280207 190727
rect 279897 190567 280207 190609
rect 279897 190449 279913 190567
rect 280031 190449 280073 190567
rect 280191 190449 280207 190567
rect 279897 172727 280207 190449
rect 279897 172609 279913 172727
rect 280031 172609 280073 172727
rect 280191 172609 280207 172727
rect 279897 172567 280207 172609
rect 279897 172449 279913 172567
rect 280031 172449 280073 172567
rect 280191 172449 280207 172567
rect 279897 154727 280207 172449
rect 279897 154609 279913 154727
rect 280031 154609 280073 154727
rect 280191 154609 280207 154727
rect 279897 154567 280207 154609
rect 279897 154449 279913 154567
rect 280031 154449 280073 154567
rect 280191 154449 280207 154567
rect 279897 136727 280207 154449
rect 279897 136609 279913 136727
rect 280031 136609 280073 136727
rect 280191 136609 280207 136727
rect 279897 136567 280207 136609
rect 279897 136449 279913 136567
rect 280031 136449 280073 136567
rect 280191 136449 280207 136567
rect 279897 118727 280207 136449
rect 279897 118609 279913 118727
rect 280031 118609 280073 118727
rect 280191 118609 280207 118727
rect 279897 118567 280207 118609
rect 279897 118449 279913 118567
rect 280031 118449 280073 118567
rect 280191 118449 280207 118567
rect 279897 100727 280207 118449
rect 279897 100609 279913 100727
rect 280031 100609 280073 100727
rect 280191 100609 280207 100727
rect 279897 100567 280207 100609
rect 279897 100449 279913 100567
rect 280031 100449 280073 100567
rect 280191 100449 280207 100567
rect 279897 82727 280207 100449
rect 279897 82609 279913 82727
rect 280031 82609 280073 82727
rect 280191 82609 280207 82727
rect 279897 82567 280207 82609
rect 279897 82449 279913 82567
rect 280031 82449 280073 82567
rect 280191 82449 280207 82567
rect 279897 64727 280207 82449
rect 279897 64609 279913 64727
rect 280031 64609 280073 64727
rect 280191 64609 280207 64727
rect 279897 64567 280207 64609
rect 279897 64449 279913 64567
rect 280031 64449 280073 64567
rect 280191 64449 280207 64567
rect 279897 46727 280207 64449
rect 279897 46609 279913 46727
rect 280031 46609 280073 46727
rect 280191 46609 280207 46727
rect 279897 46567 280207 46609
rect 279897 46449 279913 46567
rect 280031 46449 280073 46567
rect 280191 46449 280207 46567
rect 279897 28727 280207 46449
rect 279897 28609 279913 28727
rect 280031 28609 280073 28727
rect 280191 28609 280207 28727
rect 279897 28567 280207 28609
rect 279897 28449 279913 28567
rect 280031 28449 280073 28567
rect 280191 28449 280207 28567
rect 279897 10727 280207 28449
rect 279897 10609 279913 10727
rect 280031 10609 280073 10727
rect 280191 10609 280207 10727
rect 279897 10567 280207 10609
rect 279897 10449 279913 10567
rect 280031 10449 280073 10567
rect 280191 10449 280207 10567
rect 279897 -653 280207 10449
rect 279897 -771 279913 -653
rect 280031 -771 280073 -653
rect 280191 -771 280207 -653
rect 279897 -813 280207 -771
rect 279897 -931 279913 -813
rect 280031 -931 280073 -813
rect 280191 -931 280207 -813
rect 279897 -947 280207 -931
rect 281757 336587 282067 353581
rect 281757 336469 281773 336587
rect 281891 336469 281933 336587
rect 282051 336469 282067 336587
rect 281757 336427 282067 336469
rect 281757 336309 281773 336427
rect 281891 336309 281933 336427
rect 282051 336309 282067 336427
rect 281757 318587 282067 336309
rect 281757 318469 281773 318587
rect 281891 318469 281933 318587
rect 282051 318469 282067 318587
rect 281757 318427 282067 318469
rect 281757 318309 281773 318427
rect 281891 318309 281933 318427
rect 282051 318309 282067 318427
rect 281757 300587 282067 318309
rect 281757 300469 281773 300587
rect 281891 300469 281933 300587
rect 282051 300469 282067 300587
rect 281757 300427 282067 300469
rect 281757 300309 281773 300427
rect 281891 300309 281933 300427
rect 282051 300309 282067 300427
rect 281757 282587 282067 300309
rect 281757 282469 281773 282587
rect 281891 282469 281933 282587
rect 282051 282469 282067 282587
rect 281757 282427 282067 282469
rect 281757 282309 281773 282427
rect 281891 282309 281933 282427
rect 282051 282309 282067 282427
rect 281757 264587 282067 282309
rect 281757 264469 281773 264587
rect 281891 264469 281933 264587
rect 282051 264469 282067 264587
rect 281757 264427 282067 264469
rect 281757 264309 281773 264427
rect 281891 264309 281933 264427
rect 282051 264309 282067 264427
rect 281757 246587 282067 264309
rect 281757 246469 281773 246587
rect 281891 246469 281933 246587
rect 282051 246469 282067 246587
rect 281757 246427 282067 246469
rect 281757 246309 281773 246427
rect 281891 246309 281933 246427
rect 282051 246309 282067 246427
rect 281757 228587 282067 246309
rect 281757 228469 281773 228587
rect 281891 228469 281933 228587
rect 282051 228469 282067 228587
rect 281757 228427 282067 228469
rect 281757 228309 281773 228427
rect 281891 228309 281933 228427
rect 282051 228309 282067 228427
rect 281757 210587 282067 228309
rect 281757 210469 281773 210587
rect 281891 210469 281933 210587
rect 282051 210469 282067 210587
rect 281757 210427 282067 210469
rect 281757 210309 281773 210427
rect 281891 210309 281933 210427
rect 282051 210309 282067 210427
rect 281757 192587 282067 210309
rect 281757 192469 281773 192587
rect 281891 192469 281933 192587
rect 282051 192469 282067 192587
rect 281757 192427 282067 192469
rect 281757 192309 281773 192427
rect 281891 192309 281933 192427
rect 282051 192309 282067 192427
rect 281757 174587 282067 192309
rect 281757 174469 281773 174587
rect 281891 174469 281933 174587
rect 282051 174469 282067 174587
rect 281757 174427 282067 174469
rect 281757 174309 281773 174427
rect 281891 174309 281933 174427
rect 282051 174309 282067 174427
rect 281757 156587 282067 174309
rect 281757 156469 281773 156587
rect 281891 156469 281933 156587
rect 282051 156469 282067 156587
rect 281757 156427 282067 156469
rect 281757 156309 281773 156427
rect 281891 156309 281933 156427
rect 282051 156309 282067 156427
rect 281757 138587 282067 156309
rect 281757 138469 281773 138587
rect 281891 138469 281933 138587
rect 282051 138469 282067 138587
rect 281757 138427 282067 138469
rect 281757 138309 281773 138427
rect 281891 138309 281933 138427
rect 282051 138309 282067 138427
rect 281757 120587 282067 138309
rect 281757 120469 281773 120587
rect 281891 120469 281933 120587
rect 282051 120469 282067 120587
rect 281757 120427 282067 120469
rect 281757 120309 281773 120427
rect 281891 120309 281933 120427
rect 282051 120309 282067 120427
rect 281757 102587 282067 120309
rect 281757 102469 281773 102587
rect 281891 102469 281933 102587
rect 282051 102469 282067 102587
rect 281757 102427 282067 102469
rect 281757 102309 281773 102427
rect 281891 102309 281933 102427
rect 282051 102309 282067 102427
rect 281757 84587 282067 102309
rect 281757 84469 281773 84587
rect 281891 84469 281933 84587
rect 282051 84469 282067 84587
rect 281757 84427 282067 84469
rect 281757 84309 281773 84427
rect 281891 84309 281933 84427
rect 282051 84309 282067 84427
rect 281757 66587 282067 84309
rect 281757 66469 281773 66587
rect 281891 66469 281933 66587
rect 282051 66469 282067 66587
rect 281757 66427 282067 66469
rect 281757 66309 281773 66427
rect 281891 66309 281933 66427
rect 282051 66309 282067 66427
rect 281757 48587 282067 66309
rect 281757 48469 281773 48587
rect 281891 48469 281933 48587
rect 282051 48469 282067 48587
rect 281757 48427 282067 48469
rect 281757 48309 281773 48427
rect 281891 48309 281933 48427
rect 282051 48309 282067 48427
rect 281757 30587 282067 48309
rect 281757 30469 281773 30587
rect 281891 30469 281933 30587
rect 282051 30469 282067 30587
rect 281757 30427 282067 30469
rect 281757 30309 281773 30427
rect 281891 30309 281933 30427
rect 282051 30309 282067 30427
rect 281757 12587 282067 30309
rect 281757 12469 281773 12587
rect 281891 12469 281933 12587
rect 282051 12469 282067 12587
rect 281757 12427 282067 12469
rect 281757 12309 281773 12427
rect 281891 12309 281933 12427
rect 282051 12309 282067 12427
rect 281757 -1613 282067 12309
rect 281757 -1731 281773 -1613
rect 281891 -1731 281933 -1613
rect 282051 -1731 282067 -1613
rect 281757 -1773 282067 -1731
rect 281757 -1891 281773 -1773
rect 281891 -1891 281933 -1773
rect 282051 -1891 282067 -1773
rect 281757 -1907 282067 -1891
rect 283617 338447 283927 354541
rect 283617 338329 283633 338447
rect 283751 338329 283793 338447
rect 283911 338329 283927 338447
rect 283617 338287 283927 338329
rect 283617 338169 283633 338287
rect 283751 338169 283793 338287
rect 283911 338169 283927 338287
rect 283617 320447 283927 338169
rect 283617 320329 283633 320447
rect 283751 320329 283793 320447
rect 283911 320329 283927 320447
rect 283617 320287 283927 320329
rect 283617 320169 283633 320287
rect 283751 320169 283793 320287
rect 283911 320169 283927 320287
rect 283617 302447 283927 320169
rect 283617 302329 283633 302447
rect 283751 302329 283793 302447
rect 283911 302329 283927 302447
rect 283617 302287 283927 302329
rect 283617 302169 283633 302287
rect 283751 302169 283793 302287
rect 283911 302169 283927 302287
rect 283617 284447 283927 302169
rect 283617 284329 283633 284447
rect 283751 284329 283793 284447
rect 283911 284329 283927 284447
rect 283617 284287 283927 284329
rect 283617 284169 283633 284287
rect 283751 284169 283793 284287
rect 283911 284169 283927 284287
rect 283617 266447 283927 284169
rect 283617 266329 283633 266447
rect 283751 266329 283793 266447
rect 283911 266329 283927 266447
rect 283617 266287 283927 266329
rect 283617 266169 283633 266287
rect 283751 266169 283793 266287
rect 283911 266169 283927 266287
rect 283617 248447 283927 266169
rect 283617 248329 283633 248447
rect 283751 248329 283793 248447
rect 283911 248329 283927 248447
rect 283617 248287 283927 248329
rect 283617 248169 283633 248287
rect 283751 248169 283793 248287
rect 283911 248169 283927 248287
rect 283617 230447 283927 248169
rect 283617 230329 283633 230447
rect 283751 230329 283793 230447
rect 283911 230329 283927 230447
rect 283617 230287 283927 230329
rect 283617 230169 283633 230287
rect 283751 230169 283793 230287
rect 283911 230169 283927 230287
rect 283617 212447 283927 230169
rect 283617 212329 283633 212447
rect 283751 212329 283793 212447
rect 283911 212329 283927 212447
rect 283617 212287 283927 212329
rect 283617 212169 283633 212287
rect 283751 212169 283793 212287
rect 283911 212169 283927 212287
rect 283617 194447 283927 212169
rect 283617 194329 283633 194447
rect 283751 194329 283793 194447
rect 283911 194329 283927 194447
rect 283617 194287 283927 194329
rect 283617 194169 283633 194287
rect 283751 194169 283793 194287
rect 283911 194169 283927 194287
rect 283617 176447 283927 194169
rect 283617 176329 283633 176447
rect 283751 176329 283793 176447
rect 283911 176329 283927 176447
rect 283617 176287 283927 176329
rect 283617 176169 283633 176287
rect 283751 176169 283793 176287
rect 283911 176169 283927 176287
rect 283617 158447 283927 176169
rect 283617 158329 283633 158447
rect 283751 158329 283793 158447
rect 283911 158329 283927 158447
rect 283617 158287 283927 158329
rect 283617 158169 283633 158287
rect 283751 158169 283793 158287
rect 283911 158169 283927 158287
rect 283617 140447 283927 158169
rect 283617 140329 283633 140447
rect 283751 140329 283793 140447
rect 283911 140329 283927 140447
rect 283617 140287 283927 140329
rect 283617 140169 283633 140287
rect 283751 140169 283793 140287
rect 283911 140169 283927 140287
rect 283617 122447 283927 140169
rect 283617 122329 283633 122447
rect 283751 122329 283793 122447
rect 283911 122329 283927 122447
rect 283617 122287 283927 122329
rect 283617 122169 283633 122287
rect 283751 122169 283793 122287
rect 283911 122169 283927 122287
rect 283617 104447 283927 122169
rect 283617 104329 283633 104447
rect 283751 104329 283793 104447
rect 283911 104329 283927 104447
rect 283617 104287 283927 104329
rect 283617 104169 283633 104287
rect 283751 104169 283793 104287
rect 283911 104169 283927 104287
rect 283617 86447 283927 104169
rect 283617 86329 283633 86447
rect 283751 86329 283793 86447
rect 283911 86329 283927 86447
rect 283617 86287 283927 86329
rect 283617 86169 283633 86287
rect 283751 86169 283793 86287
rect 283911 86169 283927 86287
rect 283617 68447 283927 86169
rect 283617 68329 283633 68447
rect 283751 68329 283793 68447
rect 283911 68329 283927 68447
rect 283617 68287 283927 68329
rect 283617 68169 283633 68287
rect 283751 68169 283793 68287
rect 283911 68169 283927 68287
rect 283617 50447 283927 68169
rect 283617 50329 283633 50447
rect 283751 50329 283793 50447
rect 283911 50329 283927 50447
rect 283617 50287 283927 50329
rect 283617 50169 283633 50287
rect 283751 50169 283793 50287
rect 283911 50169 283927 50287
rect 283617 32447 283927 50169
rect 283617 32329 283633 32447
rect 283751 32329 283793 32447
rect 283911 32329 283927 32447
rect 283617 32287 283927 32329
rect 283617 32169 283633 32287
rect 283751 32169 283793 32287
rect 283911 32169 283927 32287
rect 283617 14447 283927 32169
rect 283617 14329 283633 14447
rect 283751 14329 283793 14447
rect 283911 14329 283927 14447
rect 283617 14287 283927 14329
rect 283617 14169 283633 14287
rect 283751 14169 283793 14287
rect 283911 14169 283927 14287
rect 283617 -2573 283927 14169
rect 283617 -2691 283633 -2573
rect 283751 -2691 283793 -2573
rect 283911 -2691 283927 -2573
rect 283617 -2733 283927 -2691
rect 283617 -2851 283633 -2733
rect 283751 -2851 283793 -2733
rect 283911 -2851 283927 -2733
rect 283617 -2867 283927 -2851
rect 285477 340307 285787 355501
rect 296015 355779 296325 355795
rect 296015 355661 296031 355779
rect 296149 355661 296191 355779
rect 296309 355661 296325 355779
rect 296015 355619 296325 355661
rect 296015 355501 296031 355619
rect 296149 355501 296191 355619
rect 296309 355501 296325 355619
rect 295535 355299 295845 355315
rect 295535 355181 295551 355299
rect 295669 355181 295711 355299
rect 295829 355181 295845 355299
rect 295535 355139 295845 355181
rect 295535 355021 295551 355139
rect 295669 355021 295711 355139
rect 295829 355021 295845 355139
rect 295055 354819 295365 354835
rect 295055 354701 295071 354819
rect 295189 354701 295231 354819
rect 295349 354701 295365 354819
rect 295055 354659 295365 354701
rect 295055 354541 295071 354659
rect 295189 354541 295231 354659
rect 295349 354541 295365 354659
rect 294575 354339 294885 354355
rect 294575 354221 294591 354339
rect 294709 354221 294751 354339
rect 294869 354221 294885 354339
rect 294575 354179 294885 354221
rect 294575 354061 294591 354179
rect 294709 354061 294751 354179
rect 294869 354061 294885 354179
rect 290757 353379 291067 353875
rect 294095 353859 294405 353875
rect 294095 353741 294111 353859
rect 294229 353741 294271 353859
rect 294389 353741 294405 353859
rect 294095 353699 294405 353741
rect 294095 353581 294111 353699
rect 294229 353581 294271 353699
rect 294389 353581 294405 353699
rect 290757 353261 290773 353379
rect 290891 353261 290933 353379
rect 291051 353261 291067 353379
rect 290757 353219 291067 353261
rect 290757 353101 290773 353219
rect 290891 353101 290933 353219
rect 291051 353101 291067 353219
rect 285477 340189 285493 340307
rect 285611 340189 285653 340307
rect 285771 340189 285787 340307
rect 285477 340147 285787 340189
rect 285477 340029 285493 340147
rect 285611 340029 285653 340147
rect 285771 340029 285787 340147
rect 285477 322307 285787 340029
rect 285477 322189 285493 322307
rect 285611 322189 285653 322307
rect 285771 322189 285787 322307
rect 285477 322147 285787 322189
rect 285477 322029 285493 322147
rect 285611 322029 285653 322147
rect 285771 322029 285787 322147
rect 285477 304307 285787 322029
rect 285477 304189 285493 304307
rect 285611 304189 285653 304307
rect 285771 304189 285787 304307
rect 285477 304147 285787 304189
rect 285477 304029 285493 304147
rect 285611 304029 285653 304147
rect 285771 304029 285787 304147
rect 285477 286307 285787 304029
rect 285477 286189 285493 286307
rect 285611 286189 285653 286307
rect 285771 286189 285787 286307
rect 285477 286147 285787 286189
rect 285477 286029 285493 286147
rect 285611 286029 285653 286147
rect 285771 286029 285787 286147
rect 285477 268307 285787 286029
rect 285477 268189 285493 268307
rect 285611 268189 285653 268307
rect 285771 268189 285787 268307
rect 285477 268147 285787 268189
rect 285477 268029 285493 268147
rect 285611 268029 285653 268147
rect 285771 268029 285787 268147
rect 285477 250307 285787 268029
rect 285477 250189 285493 250307
rect 285611 250189 285653 250307
rect 285771 250189 285787 250307
rect 285477 250147 285787 250189
rect 285477 250029 285493 250147
rect 285611 250029 285653 250147
rect 285771 250029 285787 250147
rect 285477 232307 285787 250029
rect 285477 232189 285493 232307
rect 285611 232189 285653 232307
rect 285771 232189 285787 232307
rect 285477 232147 285787 232189
rect 285477 232029 285493 232147
rect 285611 232029 285653 232147
rect 285771 232029 285787 232147
rect 285477 214307 285787 232029
rect 285477 214189 285493 214307
rect 285611 214189 285653 214307
rect 285771 214189 285787 214307
rect 285477 214147 285787 214189
rect 285477 214029 285493 214147
rect 285611 214029 285653 214147
rect 285771 214029 285787 214147
rect 285477 196307 285787 214029
rect 285477 196189 285493 196307
rect 285611 196189 285653 196307
rect 285771 196189 285787 196307
rect 285477 196147 285787 196189
rect 285477 196029 285493 196147
rect 285611 196029 285653 196147
rect 285771 196029 285787 196147
rect 285477 178307 285787 196029
rect 285477 178189 285493 178307
rect 285611 178189 285653 178307
rect 285771 178189 285787 178307
rect 285477 178147 285787 178189
rect 285477 178029 285493 178147
rect 285611 178029 285653 178147
rect 285771 178029 285787 178147
rect 285477 160307 285787 178029
rect 285477 160189 285493 160307
rect 285611 160189 285653 160307
rect 285771 160189 285787 160307
rect 285477 160147 285787 160189
rect 285477 160029 285493 160147
rect 285611 160029 285653 160147
rect 285771 160029 285787 160147
rect 285477 142307 285787 160029
rect 285477 142189 285493 142307
rect 285611 142189 285653 142307
rect 285771 142189 285787 142307
rect 285477 142147 285787 142189
rect 285477 142029 285493 142147
rect 285611 142029 285653 142147
rect 285771 142029 285787 142147
rect 285477 124307 285787 142029
rect 285477 124189 285493 124307
rect 285611 124189 285653 124307
rect 285771 124189 285787 124307
rect 285477 124147 285787 124189
rect 285477 124029 285493 124147
rect 285611 124029 285653 124147
rect 285771 124029 285787 124147
rect 285477 106307 285787 124029
rect 285477 106189 285493 106307
rect 285611 106189 285653 106307
rect 285771 106189 285787 106307
rect 285477 106147 285787 106189
rect 285477 106029 285493 106147
rect 285611 106029 285653 106147
rect 285771 106029 285787 106147
rect 285477 88307 285787 106029
rect 285477 88189 285493 88307
rect 285611 88189 285653 88307
rect 285771 88189 285787 88307
rect 285477 88147 285787 88189
rect 285477 88029 285493 88147
rect 285611 88029 285653 88147
rect 285771 88029 285787 88147
rect 285477 70307 285787 88029
rect 285477 70189 285493 70307
rect 285611 70189 285653 70307
rect 285771 70189 285787 70307
rect 285477 70147 285787 70189
rect 285477 70029 285493 70147
rect 285611 70029 285653 70147
rect 285771 70029 285787 70147
rect 285477 52307 285787 70029
rect 285477 52189 285493 52307
rect 285611 52189 285653 52307
rect 285771 52189 285787 52307
rect 285477 52147 285787 52189
rect 285477 52029 285493 52147
rect 285611 52029 285653 52147
rect 285771 52029 285787 52147
rect 285477 34307 285787 52029
rect 285477 34189 285493 34307
rect 285611 34189 285653 34307
rect 285771 34189 285787 34307
rect 285477 34147 285787 34189
rect 285477 34029 285493 34147
rect 285611 34029 285653 34147
rect 285771 34029 285787 34147
rect 285477 16307 285787 34029
rect 285477 16189 285493 16307
rect 285611 16189 285653 16307
rect 285771 16189 285787 16307
rect 285477 16147 285787 16189
rect 285477 16029 285493 16147
rect 285611 16029 285653 16147
rect 285771 16029 285787 16147
rect 276477 -3171 276493 -3053
rect 276611 -3171 276653 -3053
rect 276771 -3171 276787 -3053
rect 276477 -3213 276787 -3171
rect 276477 -3331 276493 -3213
rect 276611 -3331 276653 -3213
rect 276771 -3331 276787 -3213
rect 276477 -3827 276787 -3331
rect 285477 -3533 285787 16029
rect 288897 352419 289207 352915
rect 288897 352301 288913 352419
rect 289031 352301 289073 352419
rect 289191 352301 289207 352419
rect 288897 352259 289207 352301
rect 288897 352141 288913 352259
rect 289031 352141 289073 352259
rect 289191 352141 289207 352259
rect 288897 343727 289207 352141
rect 288897 343609 288913 343727
rect 289031 343609 289073 343727
rect 289191 343609 289207 343727
rect 288897 343567 289207 343609
rect 288897 343449 288913 343567
rect 289031 343449 289073 343567
rect 289191 343449 289207 343567
rect 288897 325727 289207 343449
rect 288897 325609 288913 325727
rect 289031 325609 289073 325727
rect 289191 325609 289207 325727
rect 288897 325567 289207 325609
rect 288897 325449 288913 325567
rect 289031 325449 289073 325567
rect 289191 325449 289207 325567
rect 288897 307727 289207 325449
rect 288897 307609 288913 307727
rect 289031 307609 289073 307727
rect 289191 307609 289207 307727
rect 288897 307567 289207 307609
rect 288897 307449 288913 307567
rect 289031 307449 289073 307567
rect 289191 307449 289207 307567
rect 288897 289727 289207 307449
rect 288897 289609 288913 289727
rect 289031 289609 289073 289727
rect 289191 289609 289207 289727
rect 288897 289567 289207 289609
rect 288897 289449 288913 289567
rect 289031 289449 289073 289567
rect 289191 289449 289207 289567
rect 288897 271727 289207 289449
rect 288897 271609 288913 271727
rect 289031 271609 289073 271727
rect 289191 271609 289207 271727
rect 288897 271567 289207 271609
rect 288897 271449 288913 271567
rect 289031 271449 289073 271567
rect 289191 271449 289207 271567
rect 288897 253727 289207 271449
rect 288897 253609 288913 253727
rect 289031 253609 289073 253727
rect 289191 253609 289207 253727
rect 288897 253567 289207 253609
rect 288897 253449 288913 253567
rect 289031 253449 289073 253567
rect 289191 253449 289207 253567
rect 288897 235727 289207 253449
rect 288897 235609 288913 235727
rect 289031 235609 289073 235727
rect 289191 235609 289207 235727
rect 288897 235567 289207 235609
rect 288897 235449 288913 235567
rect 289031 235449 289073 235567
rect 289191 235449 289207 235567
rect 288897 217727 289207 235449
rect 288897 217609 288913 217727
rect 289031 217609 289073 217727
rect 289191 217609 289207 217727
rect 288897 217567 289207 217609
rect 288897 217449 288913 217567
rect 289031 217449 289073 217567
rect 289191 217449 289207 217567
rect 288897 199727 289207 217449
rect 288897 199609 288913 199727
rect 289031 199609 289073 199727
rect 289191 199609 289207 199727
rect 288897 199567 289207 199609
rect 288897 199449 288913 199567
rect 289031 199449 289073 199567
rect 289191 199449 289207 199567
rect 288897 181727 289207 199449
rect 288897 181609 288913 181727
rect 289031 181609 289073 181727
rect 289191 181609 289207 181727
rect 288897 181567 289207 181609
rect 288897 181449 288913 181567
rect 289031 181449 289073 181567
rect 289191 181449 289207 181567
rect 288897 163727 289207 181449
rect 288897 163609 288913 163727
rect 289031 163609 289073 163727
rect 289191 163609 289207 163727
rect 288897 163567 289207 163609
rect 288897 163449 288913 163567
rect 289031 163449 289073 163567
rect 289191 163449 289207 163567
rect 288897 145727 289207 163449
rect 288897 145609 288913 145727
rect 289031 145609 289073 145727
rect 289191 145609 289207 145727
rect 288897 145567 289207 145609
rect 288897 145449 288913 145567
rect 289031 145449 289073 145567
rect 289191 145449 289207 145567
rect 288897 127727 289207 145449
rect 288897 127609 288913 127727
rect 289031 127609 289073 127727
rect 289191 127609 289207 127727
rect 288897 127567 289207 127609
rect 288897 127449 288913 127567
rect 289031 127449 289073 127567
rect 289191 127449 289207 127567
rect 288897 109727 289207 127449
rect 288897 109609 288913 109727
rect 289031 109609 289073 109727
rect 289191 109609 289207 109727
rect 288897 109567 289207 109609
rect 288897 109449 288913 109567
rect 289031 109449 289073 109567
rect 289191 109449 289207 109567
rect 288897 91727 289207 109449
rect 288897 91609 288913 91727
rect 289031 91609 289073 91727
rect 289191 91609 289207 91727
rect 288897 91567 289207 91609
rect 288897 91449 288913 91567
rect 289031 91449 289073 91567
rect 289191 91449 289207 91567
rect 288897 73727 289207 91449
rect 288897 73609 288913 73727
rect 289031 73609 289073 73727
rect 289191 73609 289207 73727
rect 288897 73567 289207 73609
rect 288897 73449 288913 73567
rect 289031 73449 289073 73567
rect 289191 73449 289207 73567
rect 288897 55727 289207 73449
rect 288897 55609 288913 55727
rect 289031 55609 289073 55727
rect 289191 55609 289207 55727
rect 288897 55567 289207 55609
rect 288897 55449 288913 55567
rect 289031 55449 289073 55567
rect 289191 55449 289207 55567
rect 288897 37727 289207 55449
rect 288897 37609 288913 37727
rect 289031 37609 289073 37727
rect 289191 37609 289207 37727
rect 288897 37567 289207 37609
rect 288897 37449 288913 37567
rect 289031 37449 289073 37567
rect 289191 37449 289207 37567
rect 288897 19727 289207 37449
rect 288897 19609 288913 19727
rect 289031 19609 289073 19727
rect 289191 19609 289207 19727
rect 288897 19567 289207 19609
rect 288897 19449 288913 19567
rect 289031 19449 289073 19567
rect 289191 19449 289207 19567
rect 288897 1727 289207 19449
rect 288897 1609 288913 1727
rect 289031 1609 289073 1727
rect 289191 1609 289207 1727
rect 288897 1567 289207 1609
rect 288897 1449 288913 1567
rect 289031 1449 289073 1567
rect 289191 1449 289207 1567
rect 288897 -173 289207 1449
rect 288897 -291 288913 -173
rect 289031 -291 289073 -173
rect 289191 -291 289207 -173
rect 288897 -333 289207 -291
rect 288897 -451 288913 -333
rect 289031 -451 289073 -333
rect 289191 -451 289207 -333
rect 288897 -947 289207 -451
rect 290757 345587 291067 353101
rect 293615 353379 293925 353395
rect 293615 353261 293631 353379
rect 293749 353261 293791 353379
rect 293909 353261 293925 353379
rect 293615 353219 293925 353261
rect 293615 353101 293631 353219
rect 293749 353101 293791 353219
rect 293909 353101 293925 353219
rect 293135 352899 293445 352915
rect 293135 352781 293151 352899
rect 293269 352781 293311 352899
rect 293429 352781 293445 352899
rect 293135 352739 293445 352781
rect 293135 352621 293151 352739
rect 293269 352621 293311 352739
rect 293429 352621 293445 352739
rect 290757 345469 290773 345587
rect 290891 345469 290933 345587
rect 291051 345469 291067 345587
rect 290757 345427 291067 345469
rect 290757 345309 290773 345427
rect 290891 345309 290933 345427
rect 291051 345309 291067 345427
rect 290757 327587 291067 345309
rect 290757 327469 290773 327587
rect 290891 327469 290933 327587
rect 291051 327469 291067 327587
rect 290757 327427 291067 327469
rect 290757 327309 290773 327427
rect 290891 327309 290933 327427
rect 291051 327309 291067 327427
rect 290757 309587 291067 327309
rect 290757 309469 290773 309587
rect 290891 309469 290933 309587
rect 291051 309469 291067 309587
rect 290757 309427 291067 309469
rect 290757 309309 290773 309427
rect 290891 309309 290933 309427
rect 291051 309309 291067 309427
rect 290757 291587 291067 309309
rect 290757 291469 290773 291587
rect 290891 291469 290933 291587
rect 291051 291469 291067 291587
rect 290757 291427 291067 291469
rect 290757 291309 290773 291427
rect 290891 291309 290933 291427
rect 291051 291309 291067 291427
rect 290757 273587 291067 291309
rect 290757 273469 290773 273587
rect 290891 273469 290933 273587
rect 291051 273469 291067 273587
rect 290757 273427 291067 273469
rect 290757 273309 290773 273427
rect 290891 273309 290933 273427
rect 291051 273309 291067 273427
rect 290757 255587 291067 273309
rect 290757 255469 290773 255587
rect 290891 255469 290933 255587
rect 291051 255469 291067 255587
rect 290757 255427 291067 255469
rect 290757 255309 290773 255427
rect 290891 255309 290933 255427
rect 291051 255309 291067 255427
rect 290757 237587 291067 255309
rect 290757 237469 290773 237587
rect 290891 237469 290933 237587
rect 291051 237469 291067 237587
rect 290757 237427 291067 237469
rect 290757 237309 290773 237427
rect 290891 237309 290933 237427
rect 291051 237309 291067 237427
rect 290757 219587 291067 237309
rect 290757 219469 290773 219587
rect 290891 219469 290933 219587
rect 291051 219469 291067 219587
rect 290757 219427 291067 219469
rect 290757 219309 290773 219427
rect 290891 219309 290933 219427
rect 291051 219309 291067 219427
rect 290757 201587 291067 219309
rect 290757 201469 290773 201587
rect 290891 201469 290933 201587
rect 291051 201469 291067 201587
rect 290757 201427 291067 201469
rect 290757 201309 290773 201427
rect 290891 201309 290933 201427
rect 291051 201309 291067 201427
rect 290757 183587 291067 201309
rect 290757 183469 290773 183587
rect 290891 183469 290933 183587
rect 291051 183469 291067 183587
rect 290757 183427 291067 183469
rect 290757 183309 290773 183427
rect 290891 183309 290933 183427
rect 291051 183309 291067 183427
rect 290757 165587 291067 183309
rect 290757 165469 290773 165587
rect 290891 165469 290933 165587
rect 291051 165469 291067 165587
rect 290757 165427 291067 165469
rect 290757 165309 290773 165427
rect 290891 165309 290933 165427
rect 291051 165309 291067 165427
rect 290757 147587 291067 165309
rect 290757 147469 290773 147587
rect 290891 147469 290933 147587
rect 291051 147469 291067 147587
rect 290757 147427 291067 147469
rect 290757 147309 290773 147427
rect 290891 147309 290933 147427
rect 291051 147309 291067 147427
rect 290757 129587 291067 147309
rect 290757 129469 290773 129587
rect 290891 129469 290933 129587
rect 291051 129469 291067 129587
rect 290757 129427 291067 129469
rect 290757 129309 290773 129427
rect 290891 129309 290933 129427
rect 291051 129309 291067 129427
rect 290757 111587 291067 129309
rect 290757 111469 290773 111587
rect 290891 111469 290933 111587
rect 291051 111469 291067 111587
rect 290757 111427 291067 111469
rect 290757 111309 290773 111427
rect 290891 111309 290933 111427
rect 291051 111309 291067 111427
rect 290757 93587 291067 111309
rect 290757 93469 290773 93587
rect 290891 93469 290933 93587
rect 291051 93469 291067 93587
rect 290757 93427 291067 93469
rect 290757 93309 290773 93427
rect 290891 93309 290933 93427
rect 291051 93309 291067 93427
rect 290757 75587 291067 93309
rect 290757 75469 290773 75587
rect 290891 75469 290933 75587
rect 291051 75469 291067 75587
rect 290757 75427 291067 75469
rect 290757 75309 290773 75427
rect 290891 75309 290933 75427
rect 291051 75309 291067 75427
rect 290757 57587 291067 75309
rect 290757 57469 290773 57587
rect 290891 57469 290933 57587
rect 291051 57469 291067 57587
rect 290757 57427 291067 57469
rect 290757 57309 290773 57427
rect 290891 57309 290933 57427
rect 291051 57309 291067 57427
rect 290757 39587 291067 57309
rect 290757 39469 290773 39587
rect 290891 39469 290933 39587
rect 291051 39469 291067 39587
rect 290757 39427 291067 39469
rect 290757 39309 290773 39427
rect 290891 39309 290933 39427
rect 291051 39309 291067 39427
rect 290757 21587 291067 39309
rect 290757 21469 290773 21587
rect 290891 21469 290933 21587
rect 291051 21469 291067 21587
rect 290757 21427 291067 21469
rect 290757 21309 290773 21427
rect 290891 21309 290933 21427
rect 291051 21309 291067 21427
rect 290757 3587 291067 21309
rect 290757 3469 290773 3587
rect 290891 3469 290933 3587
rect 291051 3469 291067 3587
rect 290757 3427 291067 3469
rect 290757 3309 290773 3427
rect 290891 3309 290933 3427
rect 291051 3309 291067 3427
rect 290757 -1133 291067 3309
rect 292655 352419 292965 352435
rect 292655 352301 292671 352419
rect 292789 352301 292831 352419
rect 292949 352301 292965 352419
rect 292655 352259 292965 352301
rect 292655 352141 292671 352259
rect 292789 352141 292831 352259
rect 292949 352141 292965 352259
rect 292655 343727 292965 352141
rect 292655 343609 292671 343727
rect 292789 343609 292831 343727
rect 292949 343609 292965 343727
rect 292655 343567 292965 343609
rect 292655 343449 292671 343567
rect 292789 343449 292831 343567
rect 292949 343449 292965 343567
rect 292655 325727 292965 343449
rect 292655 325609 292671 325727
rect 292789 325609 292831 325727
rect 292949 325609 292965 325727
rect 292655 325567 292965 325609
rect 292655 325449 292671 325567
rect 292789 325449 292831 325567
rect 292949 325449 292965 325567
rect 292655 307727 292965 325449
rect 292655 307609 292671 307727
rect 292789 307609 292831 307727
rect 292949 307609 292965 307727
rect 292655 307567 292965 307609
rect 292655 307449 292671 307567
rect 292789 307449 292831 307567
rect 292949 307449 292965 307567
rect 292655 289727 292965 307449
rect 292655 289609 292671 289727
rect 292789 289609 292831 289727
rect 292949 289609 292965 289727
rect 292655 289567 292965 289609
rect 292655 289449 292671 289567
rect 292789 289449 292831 289567
rect 292949 289449 292965 289567
rect 292655 271727 292965 289449
rect 292655 271609 292671 271727
rect 292789 271609 292831 271727
rect 292949 271609 292965 271727
rect 292655 271567 292965 271609
rect 292655 271449 292671 271567
rect 292789 271449 292831 271567
rect 292949 271449 292965 271567
rect 292655 253727 292965 271449
rect 292655 253609 292671 253727
rect 292789 253609 292831 253727
rect 292949 253609 292965 253727
rect 292655 253567 292965 253609
rect 292655 253449 292671 253567
rect 292789 253449 292831 253567
rect 292949 253449 292965 253567
rect 292655 235727 292965 253449
rect 292655 235609 292671 235727
rect 292789 235609 292831 235727
rect 292949 235609 292965 235727
rect 292655 235567 292965 235609
rect 292655 235449 292671 235567
rect 292789 235449 292831 235567
rect 292949 235449 292965 235567
rect 292655 217727 292965 235449
rect 292655 217609 292671 217727
rect 292789 217609 292831 217727
rect 292949 217609 292965 217727
rect 292655 217567 292965 217609
rect 292655 217449 292671 217567
rect 292789 217449 292831 217567
rect 292949 217449 292965 217567
rect 292655 199727 292965 217449
rect 292655 199609 292671 199727
rect 292789 199609 292831 199727
rect 292949 199609 292965 199727
rect 292655 199567 292965 199609
rect 292655 199449 292671 199567
rect 292789 199449 292831 199567
rect 292949 199449 292965 199567
rect 292655 181727 292965 199449
rect 292655 181609 292671 181727
rect 292789 181609 292831 181727
rect 292949 181609 292965 181727
rect 292655 181567 292965 181609
rect 292655 181449 292671 181567
rect 292789 181449 292831 181567
rect 292949 181449 292965 181567
rect 292655 163727 292965 181449
rect 292655 163609 292671 163727
rect 292789 163609 292831 163727
rect 292949 163609 292965 163727
rect 292655 163567 292965 163609
rect 292655 163449 292671 163567
rect 292789 163449 292831 163567
rect 292949 163449 292965 163567
rect 292655 145727 292965 163449
rect 292655 145609 292671 145727
rect 292789 145609 292831 145727
rect 292949 145609 292965 145727
rect 292655 145567 292965 145609
rect 292655 145449 292671 145567
rect 292789 145449 292831 145567
rect 292949 145449 292965 145567
rect 292655 127727 292965 145449
rect 292655 127609 292671 127727
rect 292789 127609 292831 127727
rect 292949 127609 292965 127727
rect 292655 127567 292965 127609
rect 292655 127449 292671 127567
rect 292789 127449 292831 127567
rect 292949 127449 292965 127567
rect 292655 109727 292965 127449
rect 292655 109609 292671 109727
rect 292789 109609 292831 109727
rect 292949 109609 292965 109727
rect 292655 109567 292965 109609
rect 292655 109449 292671 109567
rect 292789 109449 292831 109567
rect 292949 109449 292965 109567
rect 292655 91727 292965 109449
rect 292655 91609 292671 91727
rect 292789 91609 292831 91727
rect 292949 91609 292965 91727
rect 292655 91567 292965 91609
rect 292655 91449 292671 91567
rect 292789 91449 292831 91567
rect 292949 91449 292965 91567
rect 292655 73727 292965 91449
rect 292655 73609 292671 73727
rect 292789 73609 292831 73727
rect 292949 73609 292965 73727
rect 292655 73567 292965 73609
rect 292655 73449 292671 73567
rect 292789 73449 292831 73567
rect 292949 73449 292965 73567
rect 292655 55727 292965 73449
rect 292655 55609 292671 55727
rect 292789 55609 292831 55727
rect 292949 55609 292965 55727
rect 292655 55567 292965 55609
rect 292655 55449 292671 55567
rect 292789 55449 292831 55567
rect 292949 55449 292965 55567
rect 292655 37727 292965 55449
rect 292655 37609 292671 37727
rect 292789 37609 292831 37727
rect 292949 37609 292965 37727
rect 292655 37567 292965 37609
rect 292655 37449 292671 37567
rect 292789 37449 292831 37567
rect 292949 37449 292965 37567
rect 292655 19727 292965 37449
rect 292655 19609 292671 19727
rect 292789 19609 292831 19727
rect 292949 19609 292965 19727
rect 292655 19567 292965 19609
rect 292655 19449 292671 19567
rect 292789 19449 292831 19567
rect 292949 19449 292965 19567
rect 292655 1727 292965 19449
rect 292655 1609 292671 1727
rect 292789 1609 292831 1727
rect 292949 1609 292965 1727
rect 292655 1567 292965 1609
rect 292655 1449 292671 1567
rect 292789 1449 292831 1567
rect 292949 1449 292965 1567
rect 292655 -173 292965 1449
rect 292655 -291 292671 -173
rect 292789 -291 292831 -173
rect 292949 -291 292965 -173
rect 292655 -333 292965 -291
rect 292655 -451 292671 -333
rect 292789 -451 292831 -333
rect 292949 -451 292965 -333
rect 292655 -467 292965 -451
rect 293135 334727 293445 352621
rect 293135 334609 293151 334727
rect 293269 334609 293311 334727
rect 293429 334609 293445 334727
rect 293135 334567 293445 334609
rect 293135 334449 293151 334567
rect 293269 334449 293311 334567
rect 293429 334449 293445 334567
rect 293135 316727 293445 334449
rect 293135 316609 293151 316727
rect 293269 316609 293311 316727
rect 293429 316609 293445 316727
rect 293135 316567 293445 316609
rect 293135 316449 293151 316567
rect 293269 316449 293311 316567
rect 293429 316449 293445 316567
rect 293135 298727 293445 316449
rect 293135 298609 293151 298727
rect 293269 298609 293311 298727
rect 293429 298609 293445 298727
rect 293135 298567 293445 298609
rect 293135 298449 293151 298567
rect 293269 298449 293311 298567
rect 293429 298449 293445 298567
rect 293135 280727 293445 298449
rect 293135 280609 293151 280727
rect 293269 280609 293311 280727
rect 293429 280609 293445 280727
rect 293135 280567 293445 280609
rect 293135 280449 293151 280567
rect 293269 280449 293311 280567
rect 293429 280449 293445 280567
rect 293135 262727 293445 280449
rect 293135 262609 293151 262727
rect 293269 262609 293311 262727
rect 293429 262609 293445 262727
rect 293135 262567 293445 262609
rect 293135 262449 293151 262567
rect 293269 262449 293311 262567
rect 293429 262449 293445 262567
rect 293135 244727 293445 262449
rect 293135 244609 293151 244727
rect 293269 244609 293311 244727
rect 293429 244609 293445 244727
rect 293135 244567 293445 244609
rect 293135 244449 293151 244567
rect 293269 244449 293311 244567
rect 293429 244449 293445 244567
rect 293135 226727 293445 244449
rect 293135 226609 293151 226727
rect 293269 226609 293311 226727
rect 293429 226609 293445 226727
rect 293135 226567 293445 226609
rect 293135 226449 293151 226567
rect 293269 226449 293311 226567
rect 293429 226449 293445 226567
rect 293135 208727 293445 226449
rect 293135 208609 293151 208727
rect 293269 208609 293311 208727
rect 293429 208609 293445 208727
rect 293135 208567 293445 208609
rect 293135 208449 293151 208567
rect 293269 208449 293311 208567
rect 293429 208449 293445 208567
rect 293135 190727 293445 208449
rect 293135 190609 293151 190727
rect 293269 190609 293311 190727
rect 293429 190609 293445 190727
rect 293135 190567 293445 190609
rect 293135 190449 293151 190567
rect 293269 190449 293311 190567
rect 293429 190449 293445 190567
rect 293135 172727 293445 190449
rect 293135 172609 293151 172727
rect 293269 172609 293311 172727
rect 293429 172609 293445 172727
rect 293135 172567 293445 172609
rect 293135 172449 293151 172567
rect 293269 172449 293311 172567
rect 293429 172449 293445 172567
rect 293135 154727 293445 172449
rect 293135 154609 293151 154727
rect 293269 154609 293311 154727
rect 293429 154609 293445 154727
rect 293135 154567 293445 154609
rect 293135 154449 293151 154567
rect 293269 154449 293311 154567
rect 293429 154449 293445 154567
rect 293135 136727 293445 154449
rect 293135 136609 293151 136727
rect 293269 136609 293311 136727
rect 293429 136609 293445 136727
rect 293135 136567 293445 136609
rect 293135 136449 293151 136567
rect 293269 136449 293311 136567
rect 293429 136449 293445 136567
rect 293135 118727 293445 136449
rect 293135 118609 293151 118727
rect 293269 118609 293311 118727
rect 293429 118609 293445 118727
rect 293135 118567 293445 118609
rect 293135 118449 293151 118567
rect 293269 118449 293311 118567
rect 293429 118449 293445 118567
rect 293135 100727 293445 118449
rect 293135 100609 293151 100727
rect 293269 100609 293311 100727
rect 293429 100609 293445 100727
rect 293135 100567 293445 100609
rect 293135 100449 293151 100567
rect 293269 100449 293311 100567
rect 293429 100449 293445 100567
rect 293135 82727 293445 100449
rect 293135 82609 293151 82727
rect 293269 82609 293311 82727
rect 293429 82609 293445 82727
rect 293135 82567 293445 82609
rect 293135 82449 293151 82567
rect 293269 82449 293311 82567
rect 293429 82449 293445 82567
rect 293135 64727 293445 82449
rect 293135 64609 293151 64727
rect 293269 64609 293311 64727
rect 293429 64609 293445 64727
rect 293135 64567 293445 64609
rect 293135 64449 293151 64567
rect 293269 64449 293311 64567
rect 293429 64449 293445 64567
rect 293135 46727 293445 64449
rect 293135 46609 293151 46727
rect 293269 46609 293311 46727
rect 293429 46609 293445 46727
rect 293135 46567 293445 46609
rect 293135 46449 293151 46567
rect 293269 46449 293311 46567
rect 293429 46449 293445 46567
rect 293135 28727 293445 46449
rect 293135 28609 293151 28727
rect 293269 28609 293311 28727
rect 293429 28609 293445 28727
rect 293135 28567 293445 28609
rect 293135 28449 293151 28567
rect 293269 28449 293311 28567
rect 293429 28449 293445 28567
rect 293135 10727 293445 28449
rect 293135 10609 293151 10727
rect 293269 10609 293311 10727
rect 293429 10609 293445 10727
rect 293135 10567 293445 10609
rect 293135 10449 293151 10567
rect 293269 10449 293311 10567
rect 293429 10449 293445 10567
rect 293135 -653 293445 10449
rect 293135 -771 293151 -653
rect 293269 -771 293311 -653
rect 293429 -771 293445 -653
rect 293135 -813 293445 -771
rect 293135 -931 293151 -813
rect 293269 -931 293311 -813
rect 293429 -931 293445 -813
rect 293135 -947 293445 -931
rect 293615 345587 293925 353101
rect 293615 345469 293631 345587
rect 293749 345469 293791 345587
rect 293909 345469 293925 345587
rect 293615 345427 293925 345469
rect 293615 345309 293631 345427
rect 293749 345309 293791 345427
rect 293909 345309 293925 345427
rect 293615 327587 293925 345309
rect 293615 327469 293631 327587
rect 293749 327469 293791 327587
rect 293909 327469 293925 327587
rect 293615 327427 293925 327469
rect 293615 327309 293631 327427
rect 293749 327309 293791 327427
rect 293909 327309 293925 327427
rect 293615 309587 293925 327309
rect 293615 309469 293631 309587
rect 293749 309469 293791 309587
rect 293909 309469 293925 309587
rect 293615 309427 293925 309469
rect 293615 309309 293631 309427
rect 293749 309309 293791 309427
rect 293909 309309 293925 309427
rect 293615 291587 293925 309309
rect 293615 291469 293631 291587
rect 293749 291469 293791 291587
rect 293909 291469 293925 291587
rect 293615 291427 293925 291469
rect 293615 291309 293631 291427
rect 293749 291309 293791 291427
rect 293909 291309 293925 291427
rect 293615 273587 293925 291309
rect 293615 273469 293631 273587
rect 293749 273469 293791 273587
rect 293909 273469 293925 273587
rect 293615 273427 293925 273469
rect 293615 273309 293631 273427
rect 293749 273309 293791 273427
rect 293909 273309 293925 273427
rect 293615 255587 293925 273309
rect 293615 255469 293631 255587
rect 293749 255469 293791 255587
rect 293909 255469 293925 255587
rect 293615 255427 293925 255469
rect 293615 255309 293631 255427
rect 293749 255309 293791 255427
rect 293909 255309 293925 255427
rect 293615 237587 293925 255309
rect 293615 237469 293631 237587
rect 293749 237469 293791 237587
rect 293909 237469 293925 237587
rect 293615 237427 293925 237469
rect 293615 237309 293631 237427
rect 293749 237309 293791 237427
rect 293909 237309 293925 237427
rect 293615 219587 293925 237309
rect 293615 219469 293631 219587
rect 293749 219469 293791 219587
rect 293909 219469 293925 219587
rect 293615 219427 293925 219469
rect 293615 219309 293631 219427
rect 293749 219309 293791 219427
rect 293909 219309 293925 219427
rect 293615 201587 293925 219309
rect 293615 201469 293631 201587
rect 293749 201469 293791 201587
rect 293909 201469 293925 201587
rect 293615 201427 293925 201469
rect 293615 201309 293631 201427
rect 293749 201309 293791 201427
rect 293909 201309 293925 201427
rect 293615 183587 293925 201309
rect 293615 183469 293631 183587
rect 293749 183469 293791 183587
rect 293909 183469 293925 183587
rect 293615 183427 293925 183469
rect 293615 183309 293631 183427
rect 293749 183309 293791 183427
rect 293909 183309 293925 183427
rect 293615 165587 293925 183309
rect 293615 165469 293631 165587
rect 293749 165469 293791 165587
rect 293909 165469 293925 165587
rect 293615 165427 293925 165469
rect 293615 165309 293631 165427
rect 293749 165309 293791 165427
rect 293909 165309 293925 165427
rect 293615 147587 293925 165309
rect 293615 147469 293631 147587
rect 293749 147469 293791 147587
rect 293909 147469 293925 147587
rect 293615 147427 293925 147469
rect 293615 147309 293631 147427
rect 293749 147309 293791 147427
rect 293909 147309 293925 147427
rect 293615 129587 293925 147309
rect 293615 129469 293631 129587
rect 293749 129469 293791 129587
rect 293909 129469 293925 129587
rect 293615 129427 293925 129469
rect 293615 129309 293631 129427
rect 293749 129309 293791 129427
rect 293909 129309 293925 129427
rect 293615 111587 293925 129309
rect 293615 111469 293631 111587
rect 293749 111469 293791 111587
rect 293909 111469 293925 111587
rect 293615 111427 293925 111469
rect 293615 111309 293631 111427
rect 293749 111309 293791 111427
rect 293909 111309 293925 111427
rect 293615 93587 293925 111309
rect 293615 93469 293631 93587
rect 293749 93469 293791 93587
rect 293909 93469 293925 93587
rect 293615 93427 293925 93469
rect 293615 93309 293631 93427
rect 293749 93309 293791 93427
rect 293909 93309 293925 93427
rect 293615 75587 293925 93309
rect 293615 75469 293631 75587
rect 293749 75469 293791 75587
rect 293909 75469 293925 75587
rect 293615 75427 293925 75469
rect 293615 75309 293631 75427
rect 293749 75309 293791 75427
rect 293909 75309 293925 75427
rect 293615 57587 293925 75309
rect 293615 57469 293631 57587
rect 293749 57469 293791 57587
rect 293909 57469 293925 57587
rect 293615 57427 293925 57469
rect 293615 57309 293631 57427
rect 293749 57309 293791 57427
rect 293909 57309 293925 57427
rect 293615 39587 293925 57309
rect 293615 39469 293631 39587
rect 293749 39469 293791 39587
rect 293909 39469 293925 39587
rect 293615 39427 293925 39469
rect 293615 39309 293631 39427
rect 293749 39309 293791 39427
rect 293909 39309 293925 39427
rect 293615 21587 293925 39309
rect 293615 21469 293631 21587
rect 293749 21469 293791 21587
rect 293909 21469 293925 21587
rect 293615 21427 293925 21469
rect 293615 21309 293631 21427
rect 293749 21309 293791 21427
rect 293909 21309 293925 21427
rect 293615 3587 293925 21309
rect 293615 3469 293631 3587
rect 293749 3469 293791 3587
rect 293909 3469 293925 3587
rect 293615 3427 293925 3469
rect 293615 3309 293631 3427
rect 293749 3309 293791 3427
rect 293909 3309 293925 3427
rect 290757 -1251 290773 -1133
rect 290891 -1251 290933 -1133
rect 291051 -1251 291067 -1133
rect 290757 -1293 291067 -1251
rect 290757 -1411 290773 -1293
rect 290891 -1411 290933 -1293
rect 291051 -1411 291067 -1293
rect 290757 -1907 291067 -1411
rect 293615 -1133 293925 3309
rect 293615 -1251 293631 -1133
rect 293749 -1251 293791 -1133
rect 293909 -1251 293925 -1133
rect 293615 -1293 293925 -1251
rect 293615 -1411 293631 -1293
rect 293749 -1411 293791 -1293
rect 293909 -1411 293925 -1293
rect 293615 -1427 293925 -1411
rect 294095 336587 294405 353581
rect 294095 336469 294111 336587
rect 294229 336469 294271 336587
rect 294389 336469 294405 336587
rect 294095 336427 294405 336469
rect 294095 336309 294111 336427
rect 294229 336309 294271 336427
rect 294389 336309 294405 336427
rect 294095 318587 294405 336309
rect 294095 318469 294111 318587
rect 294229 318469 294271 318587
rect 294389 318469 294405 318587
rect 294095 318427 294405 318469
rect 294095 318309 294111 318427
rect 294229 318309 294271 318427
rect 294389 318309 294405 318427
rect 294095 300587 294405 318309
rect 294095 300469 294111 300587
rect 294229 300469 294271 300587
rect 294389 300469 294405 300587
rect 294095 300427 294405 300469
rect 294095 300309 294111 300427
rect 294229 300309 294271 300427
rect 294389 300309 294405 300427
rect 294095 282587 294405 300309
rect 294095 282469 294111 282587
rect 294229 282469 294271 282587
rect 294389 282469 294405 282587
rect 294095 282427 294405 282469
rect 294095 282309 294111 282427
rect 294229 282309 294271 282427
rect 294389 282309 294405 282427
rect 294095 264587 294405 282309
rect 294095 264469 294111 264587
rect 294229 264469 294271 264587
rect 294389 264469 294405 264587
rect 294095 264427 294405 264469
rect 294095 264309 294111 264427
rect 294229 264309 294271 264427
rect 294389 264309 294405 264427
rect 294095 246587 294405 264309
rect 294095 246469 294111 246587
rect 294229 246469 294271 246587
rect 294389 246469 294405 246587
rect 294095 246427 294405 246469
rect 294095 246309 294111 246427
rect 294229 246309 294271 246427
rect 294389 246309 294405 246427
rect 294095 228587 294405 246309
rect 294095 228469 294111 228587
rect 294229 228469 294271 228587
rect 294389 228469 294405 228587
rect 294095 228427 294405 228469
rect 294095 228309 294111 228427
rect 294229 228309 294271 228427
rect 294389 228309 294405 228427
rect 294095 210587 294405 228309
rect 294095 210469 294111 210587
rect 294229 210469 294271 210587
rect 294389 210469 294405 210587
rect 294095 210427 294405 210469
rect 294095 210309 294111 210427
rect 294229 210309 294271 210427
rect 294389 210309 294405 210427
rect 294095 192587 294405 210309
rect 294095 192469 294111 192587
rect 294229 192469 294271 192587
rect 294389 192469 294405 192587
rect 294095 192427 294405 192469
rect 294095 192309 294111 192427
rect 294229 192309 294271 192427
rect 294389 192309 294405 192427
rect 294095 174587 294405 192309
rect 294095 174469 294111 174587
rect 294229 174469 294271 174587
rect 294389 174469 294405 174587
rect 294095 174427 294405 174469
rect 294095 174309 294111 174427
rect 294229 174309 294271 174427
rect 294389 174309 294405 174427
rect 294095 156587 294405 174309
rect 294095 156469 294111 156587
rect 294229 156469 294271 156587
rect 294389 156469 294405 156587
rect 294095 156427 294405 156469
rect 294095 156309 294111 156427
rect 294229 156309 294271 156427
rect 294389 156309 294405 156427
rect 294095 138587 294405 156309
rect 294095 138469 294111 138587
rect 294229 138469 294271 138587
rect 294389 138469 294405 138587
rect 294095 138427 294405 138469
rect 294095 138309 294111 138427
rect 294229 138309 294271 138427
rect 294389 138309 294405 138427
rect 294095 120587 294405 138309
rect 294095 120469 294111 120587
rect 294229 120469 294271 120587
rect 294389 120469 294405 120587
rect 294095 120427 294405 120469
rect 294095 120309 294111 120427
rect 294229 120309 294271 120427
rect 294389 120309 294405 120427
rect 294095 102587 294405 120309
rect 294095 102469 294111 102587
rect 294229 102469 294271 102587
rect 294389 102469 294405 102587
rect 294095 102427 294405 102469
rect 294095 102309 294111 102427
rect 294229 102309 294271 102427
rect 294389 102309 294405 102427
rect 294095 84587 294405 102309
rect 294095 84469 294111 84587
rect 294229 84469 294271 84587
rect 294389 84469 294405 84587
rect 294095 84427 294405 84469
rect 294095 84309 294111 84427
rect 294229 84309 294271 84427
rect 294389 84309 294405 84427
rect 294095 66587 294405 84309
rect 294095 66469 294111 66587
rect 294229 66469 294271 66587
rect 294389 66469 294405 66587
rect 294095 66427 294405 66469
rect 294095 66309 294111 66427
rect 294229 66309 294271 66427
rect 294389 66309 294405 66427
rect 294095 48587 294405 66309
rect 294095 48469 294111 48587
rect 294229 48469 294271 48587
rect 294389 48469 294405 48587
rect 294095 48427 294405 48469
rect 294095 48309 294111 48427
rect 294229 48309 294271 48427
rect 294389 48309 294405 48427
rect 294095 30587 294405 48309
rect 294095 30469 294111 30587
rect 294229 30469 294271 30587
rect 294389 30469 294405 30587
rect 294095 30427 294405 30469
rect 294095 30309 294111 30427
rect 294229 30309 294271 30427
rect 294389 30309 294405 30427
rect 294095 12587 294405 30309
rect 294095 12469 294111 12587
rect 294229 12469 294271 12587
rect 294389 12469 294405 12587
rect 294095 12427 294405 12469
rect 294095 12309 294111 12427
rect 294229 12309 294271 12427
rect 294389 12309 294405 12427
rect 294095 -1613 294405 12309
rect 294095 -1731 294111 -1613
rect 294229 -1731 294271 -1613
rect 294389 -1731 294405 -1613
rect 294095 -1773 294405 -1731
rect 294095 -1891 294111 -1773
rect 294229 -1891 294271 -1773
rect 294389 -1891 294405 -1773
rect 294095 -1907 294405 -1891
rect 294575 347447 294885 354061
rect 294575 347329 294591 347447
rect 294709 347329 294751 347447
rect 294869 347329 294885 347447
rect 294575 347287 294885 347329
rect 294575 347169 294591 347287
rect 294709 347169 294751 347287
rect 294869 347169 294885 347287
rect 294575 329447 294885 347169
rect 294575 329329 294591 329447
rect 294709 329329 294751 329447
rect 294869 329329 294885 329447
rect 294575 329287 294885 329329
rect 294575 329169 294591 329287
rect 294709 329169 294751 329287
rect 294869 329169 294885 329287
rect 294575 311447 294885 329169
rect 294575 311329 294591 311447
rect 294709 311329 294751 311447
rect 294869 311329 294885 311447
rect 294575 311287 294885 311329
rect 294575 311169 294591 311287
rect 294709 311169 294751 311287
rect 294869 311169 294885 311287
rect 294575 293447 294885 311169
rect 294575 293329 294591 293447
rect 294709 293329 294751 293447
rect 294869 293329 294885 293447
rect 294575 293287 294885 293329
rect 294575 293169 294591 293287
rect 294709 293169 294751 293287
rect 294869 293169 294885 293287
rect 294575 275447 294885 293169
rect 294575 275329 294591 275447
rect 294709 275329 294751 275447
rect 294869 275329 294885 275447
rect 294575 275287 294885 275329
rect 294575 275169 294591 275287
rect 294709 275169 294751 275287
rect 294869 275169 294885 275287
rect 294575 257447 294885 275169
rect 294575 257329 294591 257447
rect 294709 257329 294751 257447
rect 294869 257329 294885 257447
rect 294575 257287 294885 257329
rect 294575 257169 294591 257287
rect 294709 257169 294751 257287
rect 294869 257169 294885 257287
rect 294575 239447 294885 257169
rect 294575 239329 294591 239447
rect 294709 239329 294751 239447
rect 294869 239329 294885 239447
rect 294575 239287 294885 239329
rect 294575 239169 294591 239287
rect 294709 239169 294751 239287
rect 294869 239169 294885 239287
rect 294575 221447 294885 239169
rect 294575 221329 294591 221447
rect 294709 221329 294751 221447
rect 294869 221329 294885 221447
rect 294575 221287 294885 221329
rect 294575 221169 294591 221287
rect 294709 221169 294751 221287
rect 294869 221169 294885 221287
rect 294575 203447 294885 221169
rect 294575 203329 294591 203447
rect 294709 203329 294751 203447
rect 294869 203329 294885 203447
rect 294575 203287 294885 203329
rect 294575 203169 294591 203287
rect 294709 203169 294751 203287
rect 294869 203169 294885 203287
rect 294575 185447 294885 203169
rect 294575 185329 294591 185447
rect 294709 185329 294751 185447
rect 294869 185329 294885 185447
rect 294575 185287 294885 185329
rect 294575 185169 294591 185287
rect 294709 185169 294751 185287
rect 294869 185169 294885 185287
rect 294575 167447 294885 185169
rect 294575 167329 294591 167447
rect 294709 167329 294751 167447
rect 294869 167329 294885 167447
rect 294575 167287 294885 167329
rect 294575 167169 294591 167287
rect 294709 167169 294751 167287
rect 294869 167169 294885 167287
rect 294575 149447 294885 167169
rect 294575 149329 294591 149447
rect 294709 149329 294751 149447
rect 294869 149329 294885 149447
rect 294575 149287 294885 149329
rect 294575 149169 294591 149287
rect 294709 149169 294751 149287
rect 294869 149169 294885 149287
rect 294575 131447 294885 149169
rect 294575 131329 294591 131447
rect 294709 131329 294751 131447
rect 294869 131329 294885 131447
rect 294575 131287 294885 131329
rect 294575 131169 294591 131287
rect 294709 131169 294751 131287
rect 294869 131169 294885 131287
rect 294575 113447 294885 131169
rect 294575 113329 294591 113447
rect 294709 113329 294751 113447
rect 294869 113329 294885 113447
rect 294575 113287 294885 113329
rect 294575 113169 294591 113287
rect 294709 113169 294751 113287
rect 294869 113169 294885 113287
rect 294575 95447 294885 113169
rect 294575 95329 294591 95447
rect 294709 95329 294751 95447
rect 294869 95329 294885 95447
rect 294575 95287 294885 95329
rect 294575 95169 294591 95287
rect 294709 95169 294751 95287
rect 294869 95169 294885 95287
rect 294575 77447 294885 95169
rect 294575 77329 294591 77447
rect 294709 77329 294751 77447
rect 294869 77329 294885 77447
rect 294575 77287 294885 77329
rect 294575 77169 294591 77287
rect 294709 77169 294751 77287
rect 294869 77169 294885 77287
rect 294575 59447 294885 77169
rect 294575 59329 294591 59447
rect 294709 59329 294751 59447
rect 294869 59329 294885 59447
rect 294575 59287 294885 59329
rect 294575 59169 294591 59287
rect 294709 59169 294751 59287
rect 294869 59169 294885 59287
rect 294575 41447 294885 59169
rect 294575 41329 294591 41447
rect 294709 41329 294751 41447
rect 294869 41329 294885 41447
rect 294575 41287 294885 41329
rect 294575 41169 294591 41287
rect 294709 41169 294751 41287
rect 294869 41169 294885 41287
rect 294575 23447 294885 41169
rect 294575 23329 294591 23447
rect 294709 23329 294751 23447
rect 294869 23329 294885 23447
rect 294575 23287 294885 23329
rect 294575 23169 294591 23287
rect 294709 23169 294751 23287
rect 294869 23169 294885 23287
rect 294575 5447 294885 23169
rect 294575 5329 294591 5447
rect 294709 5329 294751 5447
rect 294869 5329 294885 5447
rect 294575 5287 294885 5329
rect 294575 5169 294591 5287
rect 294709 5169 294751 5287
rect 294869 5169 294885 5287
rect 294575 -2093 294885 5169
rect 294575 -2211 294591 -2093
rect 294709 -2211 294751 -2093
rect 294869 -2211 294885 -2093
rect 294575 -2253 294885 -2211
rect 294575 -2371 294591 -2253
rect 294709 -2371 294751 -2253
rect 294869 -2371 294885 -2253
rect 294575 -2387 294885 -2371
rect 295055 338447 295365 354541
rect 295055 338329 295071 338447
rect 295189 338329 295231 338447
rect 295349 338329 295365 338447
rect 295055 338287 295365 338329
rect 295055 338169 295071 338287
rect 295189 338169 295231 338287
rect 295349 338169 295365 338287
rect 295055 320447 295365 338169
rect 295055 320329 295071 320447
rect 295189 320329 295231 320447
rect 295349 320329 295365 320447
rect 295055 320287 295365 320329
rect 295055 320169 295071 320287
rect 295189 320169 295231 320287
rect 295349 320169 295365 320287
rect 295055 302447 295365 320169
rect 295055 302329 295071 302447
rect 295189 302329 295231 302447
rect 295349 302329 295365 302447
rect 295055 302287 295365 302329
rect 295055 302169 295071 302287
rect 295189 302169 295231 302287
rect 295349 302169 295365 302287
rect 295055 284447 295365 302169
rect 295055 284329 295071 284447
rect 295189 284329 295231 284447
rect 295349 284329 295365 284447
rect 295055 284287 295365 284329
rect 295055 284169 295071 284287
rect 295189 284169 295231 284287
rect 295349 284169 295365 284287
rect 295055 266447 295365 284169
rect 295055 266329 295071 266447
rect 295189 266329 295231 266447
rect 295349 266329 295365 266447
rect 295055 266287 295365 266329
rect 295055 266169 295071 266287
rect 295189 266169 295231 266287
rect 295349 266169 295365 266287
rect 295055 248447 295365 266169
rect 295055 248329 295071 248447
rect 295189 248329 295231 248447
rect 295349 248329 295365 248447
rect 295055 248287 295365 248329
rect 295055 248169 295071 248287
rect 295189 248169 295231 248287
rect 295349 248169 295365 248287
rect 295055 230447 295365 248169
rect 295055 230329 295071 230447
rect 295189 230329 295231 230447
rect 295349 230329 295365 230447
rect 295055 230287 295365 230329
rect 295055 230169 295071 230287
rect 295189 230169 295231 230287
rect 295349 230169 295365 230287
rect 295055 212447 295365 230169
rect 295055 212329 295071 212447
rect 295189 212329 295231 212447
rect 295349 212329 295365 212447
rect 295055 212287 295365 212329
rect 295055 212169 295071 212287
rect 295189 212169 295231 212287
rect 295349 212169 295365 212287
rect 295055 194447 295365 212169
rect 295055 194329 295071 194447
rect 295189 194329 295231 194447
rect 295349 194329 295365 194447
rect 295055 194287 295365 194329
rect 295055 194169 295071 194287
rect 295189 194169 295231 194287
rect 295349 194169 295365 194287
rect 295055 176447 295365 194169
rect 295055 176329 295071 176447
rect 295189 176329 295231 176447
rect 295349 176329 295365 176447
rect 295055 176287 295365 176329
rect 295055 176169 295071 176287
rect 295189 176169 295231 176287
rect 295349 176169 295365 176287
rect 295055 158447 295365 176169
rect 295055 158329 295071 158447
rect 295189 158329 295231 158447
rect 295349 158329 295365 158447
rect 295055 158287 295365 158329
rect 295055 158169 295071 158287
rect 295189 158169 295231 158287
rect 295349 158169 295365 158287
rect 295055 140447 295365 158169
rect 295055 140329 295071 140447
rect 295189 140329 295231 140447
rect 295349 140329 295365 140447
rect 295055 140287 295365 140329
rect 295055 140169 295071 140287
rect 295189 140169 295231 140287
rect 295349 140169 295365 140287
rect 295055 122447 295365 140169
rect 295055 122329 295071 122447
rect 295189 122329 295231 122447
rect 295349 122329 295365 122447
rect 295055 122287 295365 122329
rect 295055 122169 295071 122287
rect 295189 122169 295231 122287
rect 295349 122169 295365 122287
rect 295055 104447 295365 122169
rect 295055 104329 295071 104447
rect 295189 104329 295231 104447
rect 295349 104329 295365 104447
rect 295055 104287 295365 104329
rect 295055 104169 295071 104287
rect 295189 104169 295231 104287
rect 295349 104169 295365 104287
rect 295055 86447 295365 104169
rect 295055 86329 295071 86447
rect 295189 86329 295231 86447
rect 295349 86329 295365 86447
rect 295055 86287 295365 86329
rect 295055 86169 295071 86287
rect 295189 86169 295231 86287
rect 295349 86169 295365 86287
rect 295055 68447 295365 86169
rect 295055 68329 295071 68447
rect 295189 68329 295231 68447
rect 295349 68329 295365 68447
rect 295055 68287 295365 68329
rect 295055 68169 295071 68287
rect 295189 68169 295231 68287
rect 295349 68169 295365 68287
rect 295055 50447 295365 68169
rect 295055 50329 295071 50447
rect 295189 50329 295231 50447
rect 295349 50329 295365 50447
rect 295055 50287 295365 50329
rect 295055 50169 295071 50287
rect 295189 50169 295231 50287
rect 295349 50169 295365 50287
rect 295055 32447 295365 50169
rect 295055 32329 295071 32447
rect 295189 32329 295231 32447
rect 295349 32329 295365 32447
rect 295055 32287 295365 32329
rect 295055 32169 295071 32287
rect 295189 32169 295231 32287
rect 295349 32169 295365 32287
rect 295055 14447 295365 32169
rect 295055 14329 295071 14447
rect 295189 14329 295231 14447
rect 295349 14329 295365 14447
rect 295055 14287 295365 14329
rect 295055 14169 295071 14287
rect 295189 14169 295231 14287
rect 295349 14169 295365 14287
rect 295055 -2573 295365 14169
rect 295055 -2691 295071 -2573
rect 295189 -2691 295231 -2573
rect 295349 -2691 295365 -2573
rect 295055 -2733 295365 -2691
rect 295055 -2851 295071 -2733
rect 295189 -2851 295231 -2733
rect 295349 -2851 295365 -2733
rect 295055 -2867 295365 -2851
rect 295535 349307 295845 355021
rect 295535 349189 295551 349307
rect 295669 349189 295711 349307
rect 295829 349189 295845 349307
rect 295535 349147 295845 349189
rect 295535 349029 295551 349147
rect 295669 349029 295711 349147
rect 295829 349029 295845 349147
rect 295535 331307 295845 349029
rect 295535 331189 295551 331307
rect 295669 331189 295711 331307
rect 295829 331189 295845 331307
rect 295535 331147 295845 331189
rect 295535 331029 295551 331147
rect 295669 331029 295711 331147
rect 295829 331029 295845 331147
rect 295535 313307 295845 331029
rect 295535 313189 295551 313307
rect 295669 313189 295711 313307
rect 295829 313189 295845 313307
rect 295535 313147 295845 313189
rect 295535 313029 295551 313147
rect 295669 313029 295711 313147
rect 295829 313029 295845 313147
rect 295535 295307 295845 313029
rect 295535 295189 295551 295307
rect 295669 295189 295711 295307
rect 295829 295189 295845 295307
rect 295535 295147 295845 295189
rect 295535 295029 295551 295147
rect 295669 295029 295711 295147
rect 295829 295029 295845 295147
rect 295535 277307 295845 295029
rect 295535 277189 295551 277307
rect 295669 277189 295711 277307
rect 295829 277189 295845 277307
rect 295535 277147 295845 277189
rect 295535 277029 295551 277147
rect 295669 277029 295711 277147
rect 295829 277029 295845 277147
rect 295535 259307 295845 277029
rect 295535 259189 295551 259307
rect 295669 259189 295711 259307
rect 295829 259189 295845 259307
rect 295535 259147 295845 259189
rect 295535 259029 295551 259147
rect 295669 259029 295711 259147
rect 295829 259029 295845 259147
rect 295535 241307 295845 259029
rect 295535 241189 295551 241307
rect 295669 241189 295711 241307
rect 295829 241189 295845 241307
rect 295535 241147 295845 241189
rect 295535 241029 295551 241147
rect 295669 241029 295711 241147
rect 295829 241029 295845 241147
rect 295535 223307 295845 241029
rect 295535 223189 295551 223307
rect 295669 223189 295711 223307
rect 295829 223189 295845 223307
rect 295535 223147 295845 223189
rect 295535 223029 295551 223147
rect 295669 223029 295711 223147
rect 295829 223029 295845 223147
rect 295535 205307 295845 223029
rect 295535 205189 295551 205307
rect 295669 205189 295711 205307
rect 295829 205189 295845 205307
rect 295535 205147 295845 205189
rect 295535 205029 295551 205147
rect 295669 205029 295711 205147
rect 295829 205029 295845 205147
rect 295535 187307 295845 205029
rect 295535 187189 295551 187307
rect 295669 187189 295711 187307
rect 295829 187189 295845 187307
rect 295535 187147 295845 187189
rect 295535 187029 295551 187147
rect 295669 187029 295711 187147
rect 295829 187029 295845 187147
rect 295535 169307 295845 187029
rect 295535 169189 295551 169307
rect 295669 169189 295711 169307
rect 295829 169189 295845 169307
rect 295535 169147 295845 169189
rect 295535 169029 295551 169147
rect 295669 169029 295711 169147
rect 295829 169029 295845 169147
rect 295535 151307 295845 169029
rect 295535 151189 295551 151307
rect 295669 151189 295711 151307
rect 295829 151189 295845 151307
rect 295535 151147 295845 151189
rect 295535 151029 295551 151147
rect 295669 151029 295711 151147
rect 295829 151029 295845 151147
rect 295535 133307 295845 151029
rect 295535 133189 295551 133307
rect 295669 133189 295711 133307
rect 295829 133189 295845 133307
rect 295535 133147 295845 133189
rect 295535 133029 295551 133147
rect 295669 133029 295711 133147
rect 295829 133029 295845 133147
rect 295535 115307 295845 133029
rect 295535 115189 295551 115307
rect 295669 115189 295711 115307
rect 295829 115189 295845 115307
rect 295535 115147 295845 115189
rect 295535 115029 295551 115147
rect 295669 115029 295711 115147
rect 295829 115029 295845 115147
rect 295535 97307 295845 115029
rect 295535 97189 295551 97307
rect 295669 97189 295711 97307
rect 295829 97189 295845 97307
rect 295535 97147 295845 97189
rect 295535 97029 295551 97147
rect 295669 97029 295711 97147
rect 295829 97029 295845 97147
rect 295535 79307 295845 97029
rect 295535 79189 295551 79307
rect 295669 79189 295711 79307
rect 295829 79189 295845 79307
rect 295535 79147 295845 79189
rect 295535 79029 295551 79147
rect 295669 79029 295711 79147
rect 295829 79029 295845 79147
rect 295535 61307 295845 79029
rect 295535 61189 295551 61307
rect 295669 61189 295711 61307
rect 295829 61189 295845 61307
rect 295535 61147 295845 61189
rect 295535 61029 295551 61147
rect 295669 61029 295711 61147
rect 295829 61029 295845 61147
rect 295535 43307 295845 61029
rect 295535 43189 295551 43307
rect 295669 43189 295711 43307
rect 295829 43189 295845 43307
rect 295535 43147 295845 43189
rect 295535 43029 295551 43147
rect 295669 43029 295711 43147
rect 295829 43029 295845 43147
rect 295535 25307 295845 43029
rect 295535 25189 295551 25307
rect 295669 25189 295711 25307
rect 295829 25189 295845 25307
rect 295535 25147 295845 25189
rect 295535 25029 295551 25147
rect 295669 25029 295711 25147
rect 295829 25029 295845 25147
rect 295535 7307 295845 25029
rect 295535 7189 295551 7307
rect 295669 7189 295711 7307
rect 295829 7189 295845 7307
rect 295535 7147 295845 7189
rect 295535 7029 295551 7147
rect 295669 7029 295711 7147
rect 295829 7029 295845 7147
rect 295535 -3053 295845 7029
rect 295535 -3171 295551 -3053
rect 295669 -3171 295711 -3053
rect 295829 -3171 295845 -3053
rect 295535 -3213 295845 -3171
rect 295535 -3331 295551 -3213
rect 295669 -3331 295711 -3213
rect 295829 -3331 295845 -3213
rect 295535 -3347 295845 -3331
rect 296015 340307 296325 355501
rect 296015 340189 296031 340307
rect 296149 340189 296191 340307
rect 296309 340189 296325 340307
rect 296015 340147 296325 340189
rect 296015 340029 296031 340147
rect 296149 340029 296191 340147
rect 296309 340029 296325 340147
rect 296015 322307 296325 340029
rect 296015 322189 296031 322307
rect 296149 322189 296191 322307
rect 296309 322189 296325 322307
rect 296015 322147 296325 322189
rect 296015 322029 296031 322147
rect 296149 322029 296191 322147
rect 296309 322029 296325 322147
rect 296015 304307 296325 322029
rect 296015 304189 296031 304307
rect 296149 304189 296191 304307
rect 296309 304189 296325 304307
rect 296015 304147 296325 304189
rect 296015 304029 296031 304147
rect 296149 304029 296191 304147
rect 296309 304029 296325 304147
rect 296015 286307 296325 304029
rect 296015 286189 296031 286307
rect 296149 286189 296191 286307
rect 296309 286189 296325 286307
rect 296015 286147 296325 286189
rect 296015 286029 296031 286147
rect 296149 286029 296191 286147
rect 296309 286029 296325 286147
rect 296015 268307 296325 286029
rect 296015 268189 296031 268307
rect 296149 268189 296191 268307
rect 296309 268189 296325 268307
rect 296015 268147 296325 268189
rect 296015 268029 296031 268147
rect 296149 268029 296191 268147
rect 296309 268029 296325 268147
rect 296015 250307 296325 268029
rect 296015 250189 296031 250307
rect 296149 250189 296191 250307
rect 296309 250189 296325 250307
rect 296015 250147 296325 250189
rect 296015 250029 296031 250147
rect 296149 250029 296191 250147
rect 296309 250029 296325 250147
rect 296015 232307 296325 250029
rect 296015 232189 296031 232307
rect 296149 232189 296191 232307
rect 296309 232189 296325 232307
rect 296015 232147 296325 232189
rect 296015 232029 296031 232147
rect 296149 232029 296191 232147
rect 296309 232029 296325 232147
rect 296015 214307 296325 232029
rect 296015 214189 296031 214307
rect 296149 214189 296191 214307
rect 296309 214189 296325 214307
rect 296015 214147 296325 214189
rect 296015 214029 296031 214147
rect 296149 214029 296191 214147
rect 296309 214029 296325 214147
rect 296015 196307 296325 214029
rect 296015 196189 296031 196307
rect 296149 196189 296191 196307
rect 296309 196189 296325 196307
rect 296015 196147 296325 196189
rect 296015 196029 296031 196147
rect 296149 196029 296191 196147
rect 296309 196029 296325 196147
rect 296015 178307 296325 196029
rect 296015 178189 296031 178307
rect 296149 178189 296191 178307
rect 296309 178189 296325 178307
rect 296015 178147 296325 178189
rect 296015 178029 296031 178147
rect 296149 178029 296191 178147
rect 296309 178029 296325 178147
rect 296015 160307 296325 178029
rect 296015 160189 296031 160307
rect 296149 160189 296191 160307
rect 296309 160189 296325 160307
rect 296015 160147 296325 160189
rect 296015 160029 296031 160147
rect 296149 160029 296191 160147
rect 296309 160029 296325 160147
rect 296015 142307 296325 160029
rect 296015 142189 296031 142307
rect 296149 142189 296191 142307
rect 296309 142189 296325 142307
rect 296015 142147 296325 142189
rect 296015 142029 296031 142147
rect 296149 142029 296191 142147
rect 296309 142029 296325 142147
rect 296015 124307 296325 142029
rect 296015 124189 296031 124307
rect 296149 124189 296191 124307
rect 296309 124189 296325 124307
rect 296015 124147 296325 124189
rect 296015 124029 296031 124147
rect 296149 124029 296191 124147
rect 296309 124029 296325 124147
rect 296015 106307 296325 124029
rect 296015 106189 296031 106307
rect 296149 106189 296191 106307
rect 296309 106189 296325 106307
rect 296015 106147 296325 106189
rect 296015 106029 296031 106147
rect 296149 106029 296191 106147
rect 296309 106029 296325 106147
rect 296015 88307 296325 106029
rect 296015 88189 296031 88307
rect 296149 88189 296191 88307
rect 296309 88189 296325 88307
rect 296015 88147 296325 88189
rect 296015 88029 296031 88147
rect 296149 88029 296191 88147
rect 296309 88029 296325 88147
rect 296015 70307 296325 88029
rect 296015 70189 296031 70307
rect 296149 70189 296191 70307
rect 296309 70189 296325 70307
rect 296015 70147 296325 70189
rect 296015 70029 296031 70147
rect 296149 70029 296191 70147
rect 296309 70029 296325 70147
rect 296015 52307 296325 70029
rect 296015 52189 296031 52307
rect 296149 52189 296191 52307
rect 296309 52189 296325 52307
rect 296015 52147 296325 52189
rect 296015 52029 296031 52147
rect 296149 52029 296191 52147
rect 296309 52029 296325 52147
rect 296015 34307 296325 52029
rect 296015 34189 296031 34307
rect 296149 34189 296191 34307
rect 296309 34189 296325 34307
rect 296015 34147 296325 34189
rect 296015 34029 296031 34147
rect 296149 34029 296191 34147
rect 296309 34029 296325 34147
rect 296015 16307 296325 34029
rect 296015 16189 296031 16307
rect 296149 16189 296191 16307
rect 296309 16189 296325 16307
rect 296015 16147 296325 16189
rect 296015 16029 296031 16147
rect 296149 16029 296191 16147
rect 296309 16029 296325 16147
rect 285477 -3651 285493 -3533
rect 285611 -3651 285653 -3533
rect 285771 -3651 285787 -3533
rect 285477 -3693 285787 -3651
rect 285477 -3811 285493 -3693
rect 285611 -3811 285653 -3693
rect 285771 -3811 285787 -3693
rect 285477 -3827 285787 -3811
rect 296015 -3533 296325 16029
rect 296015 -3651 296031 -3533
rect 296149 -3651 296191 -3533
rect 296309 -3651 296325 -3533
rect 296015 -3693 296325 -3651
rect 296015 -3811 296031 -3693
rect 296149 -3811 296191 -3693
rect 296309 -3811 296325 -3693
rect 296015 -3827 296325 -3811
<< via4 >>
rect -4347 355661 -4229 355779
rect -4187 355661 -4069 355779
rect -4347 355501 -4229 355619
rect -4187 355501 -4069 355619
rect -4347 340189 -4229 340307
rect -4187 340189 -4069 340307
rect -4347 340029 -4229 340147
rect -4187 340029 -4069 340147
rect -4347 322189 -4229 322307
rect -4187 322189 -4069 322307
rect -4347 322029 -4229 322147
rect -4187 322029 -4069 322147
rect -4347 304189 -4229 304307
rect -4187 304189 -4069 304307
rect -4347 304029 -4229 304147
rect -4187 304029 -4069 304147
rect -4347 286189 -4229 286307
rect -4187 286189 -4069 286307
rect -4347 286029 -4229 286147
rect -4187 286029 -4069 286147
rect -4347 268189 -4229 268307
rect -4187 268189 -4069 268307
rect -4347 268029 -4229 268147
rect -4187 268029 -4069 268147
rect -4347 250189 -4229 250307
rect -4187 250189 -4069 250307
rect -4347 250029 -4229 250147
rect -4187 250029 -4069 250147
rect -4347 232189 -4229 232307
rect -4187 232189 -4069 232307
rect -4347 232029 -4229 232147
rect -4187 232029 -4069 232147
rect -4347 214189 -4229 214307
rect -4187 214189 -4069 214307
rect -4347 214029 -4229 214147
rect -4187 214029 -4069 214147
rect -4347 196189 -4229 196307
rect -4187 196189 -4069 196307
rect -4347 196029 -4229 196147
rect -4187 196029 -4069 196147
rect -4347 178189 -4229 178307
rect -4187 178189 -4069 178307
rect -4347 178029 -4229 178147
rect -4187 178029 -4069 178147
rect -4347 160189 -4229 160307
rect -4187 160189 -4069 160307
rect -4347 160029 -4229 160147
rect -4187 160029 -4069 160147
rect -4347 142189 -4229 142307
rect -4187 142189 -4069 142307
rect -4347 142029 -4229 142147
rect -4187 142029 -4069 142147
rect -4347 124189 -4229 124307
rect -4187 124189 -4069 124307
rect -4347 124029 -4229 124147
rect -4187 124029 -4069 124147
rect -4347 106189 -4229 106307
rect -4187 106189 -4069 106307
rect -4347 106029 -4229 106147
rect -4187 106029 -4069 106147
rect -4347 88189 -4229 88307
rect -4187 88189 -4069 88307
rect -4347 88029 -4229 88147
rect -4187 88029 -4069 88147
rect -4347 70189 -4229 70307
rect -4187 70189 -4069 70307
rect -4347 70029 -4229 70147
rect -4187 70029 -4069 70147
rect -4347 52189 -4229 52307
rect -4187 52189 -4069 52307
rect -4347 52029 -4229 52147
rect -4187 52029 -4069 52147
rect -4347 34189 -4229 34307
rect -4187 34189 -4069 34307
rect -4347 34029 -4229 34147
rect -4187 34029 -4069 34147
rect -4347 16189 -4229 16307
rect -4187 16189 -4069 16307
rect -4347 16029 -4229 16147
rect -4187 16029 -4069 16147
rect -3867 355181 -3749 355299
rect -3707 355181 -3589 355299
rect -3867 355021 -3749 355139
rect -3707 355021 -3589 355139
rect 6493 355181 6611 355299
rect 6653 355181 6771 355299
rect 6493 355021 6611 355139
rect 6653 355021 6771 355139
rect -3867 349189 -3749 349307
rect -3707 349189 -3589 349307
rect -3867 349029 -3749 349147
rect -3707 349029 -3589 349147
rect -3867 331189 -3749 331307
rect -3707 331189 -3589 331307
rect -3867 331029 -3749 331147
rect -3707 331029 -3589 331147
rect -3867 313189 -3749 313307
rect -3707 313189 -3589 313307
rect -3867 313029 -3749 313147
rect -3707 313029 -3589 313147
rect -3867 295189 -3749 295307
rect -3707 295189 -3589 295307
rect -3867 295029 -3749 295147
rect -3707 295029 -3589 295147
rect -3867 277189 -3749 277307
rect -3707 277189 -3589 277307
rect -3867 277029 -3749 277147
rect -3707 277029 -3589 277147
rect -3867 259189 -3749 259307
rect -3707 259189 -3589 259307
rect -3867 259029 -3749 259147
rect -3707 259029 -3589 259147
rect -3867 241189 -3749 241307
rect -3707 241189 -3589 241307
rect -3867 241029 -3749 241147
rect -3707 241029 -3589 241147
rect -3867 223189 -3749 223307
rect -3707 223189 -3589 223307
rect -3867 223029 -3749 223147
rect -3707 223029 -3589 223147
rect -3867 205189 -3749 205307
rect -3707 205189 -3589 205307
rect -3867 205029 -3749 205147
rect -3707 205029 -3589 205147
rect -3867 187189 -3749 187307
rect -3707 187189 -3589 187307
rect -3867 187029 -3749 187147
rect -3707 187029 -3589 187147
rect -3867 169189 -3749 169307
rect -3707 169189 -3589 169307
rect -3867 169029 -3749 169147
rect -3707 169029 -3589 169147
rect -3867 151189 -3749 151307
rect -3707 151189 -3589 151307
rect -3867 151029 -3749 151147
rect -3707 151029 -3589 151147
rect -3867 133189 -3749 133307
rect -3707 133189 -3589 133307
rect -3867 133029 -3749 133147
rect -3707 133029 -3589 133147
rect -3867 115189 -3749 115307
rect -3707 115189 -3589 115307
rect -3867 115029 -3749 115147
rect -3707 115029 -3589 115147
rect -3867 97189 -3749 97307
rect -3707 97189 -3589 97307
rect -3867 97029 -3749 97147
rect -3707 97029 -3589 97147
rect -3867 79189 -3749 79307
rect -3707 79189 -3589 79307
rect -3867 79029 -3749 79147
rect -3707 79029 -3589 79147
rect -3867 61189 -3749 61307
rect -3707 61189 -3589 61307
rect -3867 61029 -3749 61147
rect -3707 61029 -3589 61147
rect -3867 43189 -3749 43307
rect -3707 43189 -3589 43307
rect -3867 43029 -3749 43147
rect -3707 43029 -3589 43147
rect -3867 25189 -3749 25307
rect -3707 25189 -3589 25307
rect -3867 25029 -3749 25147
rect -3707 25029 -3589 25147
rect -3867 7189 -3749 7307
rect -3707 7189 -3589 7307
rect -3867 7029 -3749 7147
rect -3707 7029 -3589 7147
rect -3387 354701 -3269 354819
rect -3227 354701 -3109 354819
rect -3387 354541 -3269 354659
rect -3227 354541 -3109 354659
rect -3387 338329 -3269 338447
rect -3227 338329 -3109 338447
rect -3387 338169 -3269 338287
rect -3227 338169 -3109 338287
rect -3387 320329 -3269 320447
rect -3227 320329 -3109 320447
rect -3387 320169 -3269 320287
rect -3227 320169 -3109 320287
rect -3387 302329 -3269 302447
rect -3227 302329 -3109 302447
rect -3387 302169 -3269 302287
rect -3227 302169 -3109 302287
rect -3387 284329 -3269 284447
rect -3227 284329 -3109 284447
rect -3387 284169 -3269 284287
rect -3227 284169 -3109 284287
rect -3387 266329 -3269 266447
rect -3227 266329 -3109 266447
rect -3387 266169 -3269 266287
rect -3227 266169 -3109 266287
rect -3387 248329 -3269 248447
rect -3227 248329 -3109 248447
rect -3387 248169 -3269 248287
rect -3227 248169 -3109 248287
rect -3387 230329 -3269 230447
rect -3227 230329 -3109 230447
rect -3387 230169 -3269 230287
rect -3227 230169 -3109 230287
rect -3387 212329 -3269 212447
rect -3227 212329 -3109 212447
rect -3387 212169 -3269 212287
rect -3227 212169 -3109 212287
rect -3387 194329 -3269 194447
rect -3227 194329 -3109 194447
rect -3387 194169 -3269 194287
rect -3227 194169 -3109 194287
rect -3387 176329 -3269 176447
rect -3227 176329 -3109 176447
rect -3387 176169 -3269 176287
rect -3227 176169 -3109 176287
rect -3387 158329 -3269 158447
rect -3227 158329 -3109 158447
rect -3387 158169 -3269 158287
rect -3227 158169 -3109 158287
rect -3387 140329 -3269 140447
rect -3227 140329 -3109 140447
rect -3387 140169 -3269 140287
rect -3227 140169 -3109 140287
rect -3387 122329 -3269 122447
rect -3227 122329 -3109 122447
rect -3387 122169 -3269 122287
rect -3227 122169 -3109 122287
rect -3387 104329 -3269 104447
rect -3227 104329 -3109 104447
rect -3387 104169 -3269 104287
rect -3227 104169 -3109 104287
rect -3387 86329 -3269 86447
rect -3227 86329 -3109 86447
rect -3387 86169 -3269 86287
rect -3227 86169 -3109 86287
rect -3387 68329 -3269 68447
rect -3227 68329 -3109 68447
rect -3387 68169 -3269 68287
rect -3227 68169 -3109 68287
rect -3387 50329 -3269 50447
rect -3227 50329 -3109 50447
rect -3387 50169 -3269 50287
rect -3227 50169 -3109 50287
rect -3387 32329 -3269 32447
rect -3227 32329 -3109 32447
rect -3387 32169 -3269 32287
rect -3227 32169 -3109 32287
rect -3387 14329 -3269 14447
rect -3227 14329 -3109 14447
rect -3387 14169 -3269 14287
rect -3227 14169 -3109 14287
rect -2907 354221 -2789 354339
rect -2747 354221 -2629 354339
rect -2907 354061 -2789 354179
rect -2747 354061 -2629 354179
rect 4633 354221 4751 354339
rect 4793 354221 4911 354339
rect 4633 354061 4751 354179
rect 4793 354061 4911 354179
rect -2907 347329 -2789 347447
rect -2747 347329 -2629 347447
rect -2907 347169 -2789 347287
rect -2747 347169 -2629 347287
rect -2907 329329 -2789 329447
rect -2747 329329 -2629 329447
rect -2907 329169 -2789 329287
rect -2747 329169 -2629 329287
rect -2907 311329 -2789 311447
rect -2747 311329 -2629 311447
rect -2907 311169 -2789 311287
rect -2747 311169 -2629 311287
rect -2907 293329 -2789 293447
rect -2747 293329 -2629 293447
rect -2907 293169 -2789 293287
rect -2747 293169 -2629 293287
rect -2907 275329 -2789 275447
rect -2747 275329 -2629 275447
rect -2907 275169 -2789 275287
rect -2747 275169 -2629 275287
rect -2907 257329 -2789 257447
rect -2747 257329 -2629 257447
rect -2907 257169 -2789 257287
rect -2747 257169 -2629 257287
rect -2907 239329 -2789 239447
rect -2747 239329 -2629 239447
rect -2907 239169 -2789 239287
rect -2747 239169 -2629 239287
rect -2907 221329 -2789 221447
rect -2747 221329 -2629 221447
rect -2907 221169 -2789 221287
rect -2747 221169 -2629 221287
rect -2907 203329 -2789 203447
rect -2747 203329 -2629 203447
rect -2907 203169 -2789 203287
rect -2747 203169 -2629 203287
rect -2907 185329 -2789 185447
rect -2747 185329 -2629 185447
rect -2907 185169 -2789 185287
rect -2747 185169 -2629 185287
rect -2907 167329 -2789 167447
rect -2747 167329 -2629 167447
rect -2907 167169 -2789 167287
rect -2747 167169 -2629 167287
rect -2907 149329 -2789 149447
rect -2747 149329 -2629 149447
rect -2907 149169 -2789 149287
rect -2747 149169 -2629 149287
rect -2907 131329 -2789 131447
rect -2747 131329 -2629 131447
rect -2907 131169 -2789 131287
rect -2747 131169 -2629 131287
rect -2907 113329 -2789 113447
rect -2747 113329 -2629 113447
rect -2907 113169 -2789 113287
rect -2747 113169 -2629 113287
rect -2907 95329 -2789 95447
rect -2747 95329 -2629 95447
rect -2907 95169 -2789 95287
rect -2747 95169 -2629 95287
rect -2907 77329 -2789 77447
rect -2747 77329 -2629 77447
rect -2907 77169 -2789 77287
rect -2747 77169 -2629 77287
rect -2907 59329 -2789 59447
rect -2747 59329 -2629 59447
rect -2907 59169 -2789 59287
rect -2747 59169 -2629 59287
rect -2907 41329 -2789 41447
rect -2747 41329 -2629 41447
rect -2907 41169 -2789 41287
rect -2747 41169 -2629 41287
rect -2907 23329 -2789 23447
rect -2747 23329 -2629 23447
rect -2907 23169 -2789 23287
rect -2747 23169 -2629 23287
rect -2907 5329 -2789 5447
rect -2747 5329 -2629 5447
rect -2907 5169 -2789 5287
rect -2747 5169 -2629 5287
rect -2427 353741 -2309 353859
rect -2267 353741 -2149 353859
rect -2427 353581 -2309 353699
rect -2267 353581 -2149 353699
rect -2427 336469 -2309 336587
rect -2267 336469 -2149 336587
rect -2427 336309 -2309 336427
rect -2267 336309 -2149 336427
rect -2427 318469 -2309 318587
rect -2267 318469 -2149 318587
rect -2427 318309 -2309 318427
rect -2267 318309 -2149 318427
rect -2427 300469 -2309 300587
rect -2267 300469 -2149 300587
rect -2427 300309 -2309 300427
rect -2267 300309 -2149 300427
rect -2427 282469 -2309 282587
rect -2267 282469 -2149 282587
rect -2427 282309 -2309 282427
rect -2267 282309 -2149 282427
rect -2427 264469 -2309 264587
rect -2267 264469 -2149 264587
rect -2427 264309 -2309 264427
rect -2267 264309 -2149 264427
rect -2427 246469 -2309 246587
rect -2267 246469 -2149 246587
rect -2427 246309 -2309 246427
rect -2267 246309 -2149 246427
rect -2427 228469 -2309 228587
rect -2267 228469 -2149 228587
rect -2427 228309 -2309 228427
rect -2267 228309 -2149 228427
rect -2427 210469 -2309 210587
rect -2267 210469 -2149 210587
rect -2427 210309 -2309 210427
rect -2267 210309 -2149 210427
rect -2427 192469 -2309 192587
rect -2267 192469 -2149 192587
rect -2427 192309 -2309 192427
rect -2267 192309 -2149 192427
rect -2427 174469 -2309 174587
rect -2267 174469 -2149 174587
rect -2427 174309 -2309 174427
rect -2267 174309 -2149 174427
rect -2427 156469 -2309 156587
rect -2267 156469 -2149 156587
rect -2427 156309 -2309 156427
rect -2267 156309 -2149 156427
rect -2427 138469 -2309 138587
rect -2267 138469 -2149 138587
rect -2427 138309 -2309 138427
rect -2267 138309 -2149 138427
rect -2427 120469 -2309 120587
rect -2267 120469 -2149 120587
rect -2427 120309 -2309 120427
rect -2267 120309 -2149 120427
rect -2427 102469 -2309 102587
rect -2267 102469 -2149 102587
rect -2427 102309 -2309 102427
rect -2267 102309 -2149 102427
rect -2427 84469 -2309 84587
rect -2267 84469 -2149 84587
rect -2427 84309 -2309 84427
rect -2267 84309 -2149 84427
rect -2427 66469 -2309 66587
rect -2267 66469 -2149 66587
rect -2427 66309 -2309 66427
rect -2267 66309 -2149 66427
rect -2427 48469 -2309 48587
rect -2267 48469 -2149 48587
rect -2427 48309 -2309 48427
rect -2267 48309 -2149 48427
rect -2427 30469 -2309 30587
rect -2267 30469 -2149 30587
rect -2427 30309 -2309 30427
rect -2267 30309 -2149 30427
rect -2427 12469 -2309 12587
rect -2267 12469 -2149 12587
rect -2427 12309 -2309 12427
rect -2267 12309 -2149 12427
rect -1947 353261 -1829 353379
rect -1787 353261 -1669 353379
rect -1947 353101 -1829 353219
rect -1787 353101 -1669 353219
rect 2773 353261 2891 353379
rect 2933 353261 3051 353379
rect 2773 353101 2891 353219
rect 2933 353101 3051 353219
rect -1947 345469 -1829 345587
rect -1787 345469 -1669 345587
rect -1947 345309 -1829 345427
rect -1787 345309 -1669 345427
rect -1947 327469 -1829 327587
rect -1787 327469 -1669 327587
rect -1947 327309 -1829 327427
rect -1787 327309 -1669 327427
rect -1947 309469 -1829 309587
rect -1787 309469 -1669 309587
rect -1947 309309 -1829 309427
rect -1787 309309 -1669 309427
rect -1947 291469 -1829 291587
rect -1787 291469 -1669 291587
rect -1947 291309 -1829 291427
rect -1787 291309 -1669 291427
rect -1947 273469 -1829 273587
rect -1787 273469 -1669 273587
rect -1947 273309 -1829 273427
rect -1787 273309 -1669 273427
rect -1947 255469 -1829 255587
rect -1787 255469 -1669 255587
rect -1947 255309 -1829 255427
rect -1787 255309 -1669 255427
rect -1947 237469 -1829 237587
rect -1787 237469 -1669 237587
rect -1947 237309 -1829 237427
rect -1787 237309 -1669 237427
rect -1947 219469 -1829 219587
rect -1787 219469 -1669 219587
rect -1947 219309 -1829 219427
rect -1787 219309 -1669 219427
rect -1947 201469 -1829 201587
rect -1787 201469 -1669 201587
rect -1947 201309 -1829 201427
rect -1787 201309 -1669 201427
rect -1947 183469 -1829 183587
rect -1787 183469 -1669 183587
rect -1947 183309 -1829 183427
rect -1787 183309 -1669 183427
rect -1947 165469 -1829 165587
rect -1787 165469 -1669 165587
rect -1947 165309 -1829 165427
rect -1787 165309 -1669 165427
rect -1947 147469 -1829 147587
rect -1787 147469 -1669 147587
rect -1947 147309 -1829 147427
rect -1787 147309 -1669 147427
rect -1947 129469 -1829 129587
rect -1787 129469 -1669 129587
rect -1947 129309 -1829 129427
rect -1787 129309 -1669 129427
rect -1947 111469 -1829 111587
rect -1787 111469 -1669 111587
rect -1947 111309 -1829 111427
rect -1787 111309 -1669 111427
rect -1947 93469 -1829 93587
rect -1787 93469 -1669 93587
rect -1947 93309 -1829 93427
rect -1787 93309 -1669 93427
rect -1947 75469 -1829 75587
rect -1787 75469 -1669 75587
rect -1947 75309 -1829 75427
rect -1787 75309 -1669 75427
rect -1947 57469 -1829 57587
rect -1787 57469 -1669 57587
rect -1947 57309 -1829 57427
rect -1787 57309 -1669 57427
rect -1947 39469 -1829 39587
rect -1787 39469 -1669 39587
rect -1947 39309 -1829 39427
rect -1787 39309 -1669 39427
rect -1947 21469 -1829 21587
rect -1787 21469 -1669 21587
rect -1947 21309 -1829 21427
rect -1787 21309 -1669 21427
rect -1947 3469 -1829 3587
rect -1787 3469 -1669 3587
rect -1947 3309 -1829 3427
rect -1787 3309 -1669 3427
rect -1467 352781 -1349 352899
rect -1307 352781 -1189 352899
rect -1467 352621 -1349 352739
rect -1307 352621 -1189 352739
rect -1467 334609 -1349 334727
rect -1307 334609 -1189 334727
rect -1467 334449 -1349 334567
rect -1307 334449 -1189 334567
rect -1467 316609 -1349 316727
rect -1307 316609 -1189 316727
rect -1467 316449 -1349 316567
rect -1307 316449 -1189 316567
rect -1467 298609 -1349 298727
rect -1307 298609 -1189 298727
rect -1467 298449 -1349 298567
rect -1307 298449 -1189 298567
rect -1467 280609 -1349 280727
rect -1307 280609 -1189 280727
rect -1467 280449 -1349 280567
rect -1307 280449 -1189 280567
rect -1467 262609 -1349 262727
rect -1307 262609 -1189 262727
rect -1467 262449 -1349 262567
rect -1307 262449 -1189 262567
rect -1467 244609 -1349 244727
rect -1307 244609 -1189 244727
rect -1467 244449 -1349 244567
rect -1307 244449 -1189 244567
rect -1467 226609 -1349 226727
rect -1307 226609 -1189 226727
rect -1467 226449 -1349 226567
rect -1307 226449 -1189 226567
rect -1467 208609 -1349 208727
rect -1307 208609 -1189 208727
rect -1467 208449 -1349 208567
rect -1307 208449 -1189 208567
rect -1467 190609 -1349 190727
rect -1307 190609 -1189 190727
rect -1467 190449 -1349 190567
rect -1307 190449 -1189 190567
rect -1467 172609 -1349 172727
rect -1307 172609 -1189 172727
rect -1467 172449 -1349 172567
rect -1307 172449 -1189 172567
rect -1467 154609 -1349 154727
rect -1307 154609 -1189 154727
rect -1467 154449 -1349 154567
rect -1307 154449 -1189 154567
rect -1467 136609 -1349 136727
rect -1307 136609 -1189 136727
rect -1467 136449 -1349 136567
rect -1307 136449 -1189 136567
rect -1467 118609 -1349 118727
rect -1307 118609 -1189 118727
rect -1467 118449 -1349 118567
rect -1307 118449 -1189 118567
rect -1467 100609 -1349 100727
rect -1307 100609 -1189 100727
rect -1467 100449 -1349 100567
rect -1307 100449 -1189 100567
rect -1467 82609 -1349 82727
rect -1307 82609 -1189 82727
rect -1467 82449 -1349 82567
rect -1307 82449 -1189 82567
rect -1467 64609 -1349 64727
rect -1307 64609 -1189 64727
rect -1467 64449 -1349 64567
rect -1307 64449 -1189 64567
rect -1467 46609 -1349 46727
rect -1307 46609 -1189 46727
rect -1467 46449 -1349 46567
rect -1307 46449 -1189 46567
rect -1467 28609 -1349 28727
rect -1307 28609 -1189 28727
rect -1467 28449 -1349 28567
rect -1307 28449 -1189 28567
rect -1467 10609 -1349 10727
rect -1307 10609 -1189 10727
rect -1467 10449 -1349 10567
rect -1307 10449 -1189 10567
rect -987 352301 -869 352419
rect -827 352301 -709 352419
rect -987 352141 -869 352259
rect -827 352141 -709 352259
rect -987 343609 -869 343727
rect -827 343609 -709 343727
rect -987 343449 -869 343567
rect -827 343449 -709 343567
rect -987 325609 -869 325727
rect -827 325609 -709 325727
rect -987 325449 -869 325567
rect -827 325449 -709 325567
rect -987 307609 -869 307727
rect -827 307609 -709 307727
rect -987 307449 -869 307567
rect -827 307449 -709 307567
rect -987 289609 -869 289727
rect -827 289609 -709 289727
rect -987 289449 -869 289567
rect -827 289449 -709 289567
rect -987 271609 -869 271727
rect -827 271609 -709 271727
rect -987 271449 -869 271567
rect -827 271449 -709 271567
rect -987 253609 -869 253727
rect -827 253609 -709 253727
rect -987 253449 -869 253567
rect -827 253449 -709 253567
rect -987 235609 -869 235727
rect -827 235609 -709 235727
rect -987 235449 -869 235567
rect -827 235449 -709 235567
rect -987 217609 -869 217727
rect -827 217609 -709 217727
rect -987 217449 -869 217567
rect -827 217449 -709 217567
rect -987 199609 -869 199727
rect -827 199609 -709 199727
rect -987 199449 -869 199567
rect -827 199449 -709 199567
rect -987 181609 -869 181727
rect -827 181609 -709 181727
rect -987 181449 -869 181567
rect -827 181449 -709 181567
rect -987 163609 -869 163727
rect -827 163609 -709 163727
rect -987 163449 -869 163567
rect -827 163449 -709 163567
rect -987 145609 -869 145727
rect -827 145609 -709 145727
rect -987 145449 -869 145567
rect -827 145449 -709 145567
rect -987 127609 -869 127727
rect -827 127609 -709 127727
rect -987 127449 -869 127567
rect -827 127449 -709 127567
rect -987 109609 -869 109727
rect -827 109609 -709 109727
rect -987 109449 -869 109567
rect -827 109449 -709 109567
rect -987 91609 -869 91727
rect -827 91609 -709 91727
rect -987 91449 -869 91567
rect -827 91449 -709 91567
rect -987 73609 -869 73727
rect -827 73609 -709 73727
rect -987 73449 -869 73567
rect -827 73449 -709 73567
rect -987 55609 -869 55727
rect -827 55609 -709 55727
rect -987 55449 -869 55567
rect -827 55449 -709 55567
rect -987 37609 -869 37727
rect -827 37609 -709 37727
rect -987 37449 -869 37567
rect -827 37449 -709 37567
rect -987 19609 -869 19727
rect -827 19609 -709 19727
rect -987 19449 -869 19567
rect -827 19449 -709 19567
rect -987 1609 -869 1727
rect -827 1609 -709 1727
rect -987 1449 -869 1567
rect -827 1449 -709 1567
rect -987 -291 -869 -173
rect -827 -291 -709 -173
rect -987 -451 -869 -333
rect -827 -451 -709 -333
rect 913 352301 1031 352419
rect 1073 352301 1191 352419
rect 913 352141 1031 352259
rect 1073 352141 1191 352259
rect 913 343609 1031 343727
rect 1073 343609 1191 343727
rect 913 343449 1031 343567
rect 1073 343449 1191 343567
rect 913 325609 1031 325727
rect 1073 325609 1191 325727
rect 913 325449 1031 325567
rect 1073 325449 1191 325567
rect 913 307609 1031 307727
rect 1073 307609 1191 307727
rect 913 307449 1031 307567
rect 1073 307449 1191 307567
rect 913 289609 1031 289727
rect 1073 289609 1191 289727
rect 913 289449 1031 289567
rect 1073 289449 1191 289567
rect 913 271609 1031 271727
rect 1073 271609 1191 271727
rect 913 271449 1031 271567
rect 1073 271449 1191 271567
rect 913 253609 1031 253727
rect 1073 253609 1191 253727
rect 913 253449 1031 253567
rect 1073 253449 1191 253567
rect 913 235609 1031 235727
rect 1073 235609 1191 235727
rect 913 235449 1031 235567
rect 1073 235449 1191 235567
rect 913 217609 1031 217727
rect 1073 217609 1191 217727
rect 913 217449 1031 217567
rect 1073 217449 1191 217567
rect 913 199609 1031 199727
rect 1073 199609 1191 199727
rect 913 199449 1031 199567
rect 1073 199449 1191 199567
rect 913 181609 1031 181727
rect 1073 181609 1191 181727
rect 913 181449 1031 181567
rect 1073 181449 1191 181567
rect 913 163609 1031 163727
rect 1073 163609 1191 163727
rect 913 163449 1031 163567
rect 1073 163449 1191 163567
rect 913 145609 1031 145727
rect 1073 145609 1191 145727
rect 913 145449 1031 145567
rect 1073 145449 1191 145567
rect 913 127609 1031 127727
rect 1073 127609 1191 127727
rect 913 127449 1031 127567
rect 1073 127449 1191 127567
rect 913 109609 1031 109727
rect 1073 109609 1191 109727
rect 913 109449 1031 109567
rect 1073 109449 1191 109567
rect 913 91609 1031 91727
rect 1073 91609 1191 91727
rect 913 91449 1031 91567
rect 1073 91449 1191 91567
rect 913 73609 1031 73727
rect 1073 73609 1191 73727
rect 913 73449 1031 73567
rect 1073 73449 1191 73567
rect 913 55609 1031 55727
rect 1073 55609 1191 55727
rect 913 55449 1031 55567
rect 1073 55449 1191 55567
rect 913 37609 1031 37727
rect 1073 37609 1191 37727
rect 913 37449 1031 37567
rect 1073 37449 1191 37567
rect 913 19609 1031 19727
rect 1073 19609 1191 19727
rect 913 19449 1031 19567
rect 1073 19449 1191 19567
rect 913 1609 1031 1727
rect 1073 1609 1191 1727
rect 913 1449 1031 1567
rect 1073 1449 1191 1567
rect 913 -291 1031 -173
rect 1073 -291 1191 -173
rect 913 -451 1031 -333
rect 1073 -451 1191 -333
rect -1467 -771 -1349 -653
rect -1307 -771 -1189 -653
rect -1467 -931 -1349 -813
rect -1307 -931 -1189 -813
rect 2773 345469 2891 345587
rect 2933 345469 3051 345587
rect 2773 345309 2891 345427
rect 2933 345309 3051 345427
rect 2773 327469 2891 327587
rect 2933 327469 3051 327587
rect 2773 327309 2891 327427
rect 2933 327309 3051 327427
rect 2773 309469 2891 309587
rect 2933 309469 3051 309587
rect 2773 309309 2891 309427
rect 2933 309309 3051 309427
rect 2773 291469 2891 291587
rect 2933 291469 3051 291587
rect 2773 291309 2891 291427
rect 2933 291309 3051 291427
rect 2773 273469 2891 273587
rect 2933 273469 3051 273587
rect 2773 273309 2891 273427
rect 2933 273309 3051 273427
rect 2773 255469 2891 255587
rect 2933 255469 3051 255587
rect 2773 255309 2891 255427
rect 2933 255309 3051 255427
rect 2773 237469 2891 237587
rect 2933 237469 3051 237587
rect 2773 237309 2891 237427
rect 2933 237309 3051 237427
rect 2773 219469 2891 219587
rect 2933 219469 3051 219587
rect 2773 219309 2891 219427
rect 2933 219309 3051 219427
rect 2773 201469 2891 201587
rect 2933 201469 3051 201587
rect 2773 201309 2891 201427
rect 2933 201309 3051 201427
rect 2773 183469 2891 183587
rect 2933 183469 3051 183587
rect 2773 183309 2891 183427
rect 2933 183309 3051 183427
rect 2773 165469 2891 165587
rect 2933 165469 3051 165587
rect 2773 165309 2891 165427
rect 2933 165309 3051 165427
rect 2773 147469 2891 147587
rect 2933 147469 3051 147587
rect 2773 147309 2891 147427
rect 2933 147309 3051 147427
rect 2773 129469 2891 129587
rect 2933 129469 3051 129587
rect 2773 129309 2891 129427
rect 2933 129309 3051 129427
rect 2773 111469 2891 111587
rect 2933 111469 3051 111587
rect 2773 111309 2891 111427
rect 2933 111309 3051 111427
rect 2773 93469 2891 93587
rect 2933 93469 3051 93587
rect 2773 93309 2891 93427
rect 2933 93309 3051 93427
rect 2773 75469 2891 75587
rect 2933 75469 3051 75587
rect 2773 75309 2891 75427
rect 2933 75309 3051 75427
rect 2773 57469 2891 57587
rect 2933 57469 3051 57587
rect 2773 57309 2891 57427
rect 2933 57309 3051 57427
rect 2773 39469 2891 39587
rect 2933 39469 3051 39587
rect 2773 39309 2891 39427
rect 2933 39309 3051 39427
rect 2773 21469 2891 21587
rect 2933 21469 3051 21587
rect 2773 21309 2891 21427
rect 2933 21309 3051 21427
rect 2773 3469 2891 3587
rect 2933 3469 3051 3587
rect 2773 3309 2891 3427
rect 2933 3309 3051 3427
rect -1947 -1251 -1829 -1133
rect -1787 -1251 -1669 -1133
rect -1947 -1411 -1829 -1293
rect -1787 -1411 -1669 -1293
rect 2773 -1251 2891 -1133
rect 2933 -1251 3051 -1133
rect 2773 -1411 2891 -1293
rect 2933 -1411 3051 -1293
rect -2427 -1731 -2309 -1613
rect -2267 -1731 -2149 -1613
rect -2427 -1891 -2309 -1773
rect -2267 -1891 -2149 -1773
rect 4633 347329 4751 347447
rect 4793 347329 4911 347447
rect 4633 347169 4751 347287
rect 4793 347169 4911 347287
rect 4633 329329 4751 329447
rect 4793 329329 4911 329447
rect 4633 329169 4751 329287
rect 4793 329169 4911 329287
rect 4633 311329 4751 311447
rect 4793 311329 4911 311447
rect 4633 311169 4751 311287
rect 4793 311169 4911 311287
rect 4633 293329 4751 293447
rect 4793 293329 4911 293447
rect 4633 293169 4751 293287
rect 4793 293169 4911 293287
rect 4633 275329 4751 275447
rect 4793 275329 4911 275447
rect 4633 275169 4751 275287
rect 4793 275169 4911 275287
rect 4633 257329 4751 257447
rect 4793 257329 4911 257447
rect 4633 257169 4751 257287
rect 4793 257169 4911 257287
rect 4633 239329 4751 239447
rect 4793 239329 4911 239447
rect 4633 239169 4751 239287
rect 4793 239169 4911 239287
rect 4633 221329 4751 221447
rect 4793 221329 4911 221447
rect 4633 221169 4751 221287
rect 4793 221169 4911 221287
rect 4633 203329 4751 203447
rect 4793 203329 4911 203447
rect 4633 203169 4751 203287
rect 4793 203169 4911 203287
rect 4633 185329 4751 185447
rect 4793 185329 4911 185447
rect 4633 185169 4751 185287
rect 4793 185169 4911 185287
rect 4633 167329 4751 167447
rect 4793 167329 4911 167447
rect 4633 167169 4751 167287
rect 4793 167169 4911 167287
rect 4633 149329 4751 149447
rect 4793 149329 4911 149447
rect 4633 149169 4751 149287
rect 4793 149169 4911 149287
rect 4633 131329 4751 131447
rect 4793 131329 4911 131447
rect 4633 131169 4751 131287
rect 4793 131169 4911 131287
rect 4633 113329 4751 113447
rect 4793 113329 4911 113447
rect 4633 113169 4751 113287
rect 4793 113169 4911 113287
rect 4633 95329 4751 95447
rect 4793 95329 4911 95447
rect 4633 95169 4751 95287
rect 4793 95169 4911 95287
rect 4633 77329 4751 77447
rect 4793 77329 4911 77447
rect 4633 77169 4751 77287
rect 4793 77169 4911 77287
rect 4633 59329 4751 59447
rect 4793 59329 4911 59447
rect 4633 59169 4751 59287
rect 4793 59169 4911 59287
rect 4633 41329 4751 41447
rect 4793 41329 4911 41447
rect 4633 41169 4751 41287
rect 4793 41169 4911 41287
rect 4633 23329 4751 23447
rect 4793 23329 4911 23447
rect 4633 23169 4751 23287
rect 4793 23169 4911 23287
rect 4633 5329 4751 5447
rect 4793 5329 4911 5447
rect 4633 5169 4751 5287
rect 4793 5169 4911 5287
rect -2907 -2211 -2789 -2093
rect -2747 -2211 -2629 -2093
rect -2907 -2371 -2789 -2253
rect -2747 -2371 -2629 -2253
rect 4633 -2211 4751 -2093
rect 4793 -2211 4911 -2093
rect 4633 -2371 4751 -2253
rect 4793 -2371 4911 -2253
rect -3387 -2691 -3269 -2573
rect -3227 -2691 -3109 -2573
rect -3387 -2851 -3269 -2733
rect -3227 -2851 -3109 -2733
rect 15493 355661 15611 355779
rect 15653 355661 15771 355779
rect 15493 355501 15611 355619
rect 15653 355501 15771 355619
rect 13633 354701 13751 354819
rect 13793 354701 13911 354819
rect 13633 354541 13751 354659
rect 13793 354541 13911 354659
rect 11773 353741 11891 353859
rect 11933 353741 12051 353859
rect 11773 353581 11891 353699
rect 11933 353581 12051 353699
rect 6493 349189 6611 349307
rect 6653 349189 6771 349307
rect 6493 349029 6611 349147
rect 6653 349029 6771 349147
rect 6493 331189 6611 331307
rect 6653 331189 6771 331307
rect 6493 331029 6611 331147
rect 6653 331029 6771 331147
rect 6493 313189 6611 313307
rect 6653 313189 6771 313307
rect 6493 313029 6611 313147
rect 6653 313029 6771 313147
rect 6493 295189 6611 295307
rect 6653 295189 6771 295307
rect 6493 295029 6611 295147
rect 6653 295029 6771 295147
rect 6493 277189 6611 277307
rect 6653 277189 6771 277307
rect 6493 277029 6611 277147
rect 6653 277029 6771 277147
rect 6493 259189 6611 259307
rect 6653 259189 6771 259307
rect 6493 259029 6611 259147
rect 6653 259029 6771 259147
rect 6493 241189 6611 241307
rect 6653 241189 6771 241307
rect 6493 241029 6611 241147
rect 6653 241029 6771 241147
rect 6493 223189 6611 223307
rect 6653 223189 6771 223307
rect 6493 223029 6611 223147
rect 6653 223029 6771 223147
rect 6493 205189 6611 205307
rect 6653 205189 6771 205307
rect 6493 205029 6611 205147
rect 6653 205029 6771 205147
rect 6493 187189 6611 187307
rect 6653 187189 6771 187307
rect 6493 187029 6611 187147
rect 6653 187029 6771 187147
rect 6493 169189 6611 169307
rect 6653 169189 6771 169307
rect 6493 169029 6611 169147
rect 6653 169029 6771 169147
rect 6493 151189 6611 151307
rect 6653 151189 6771 151307
rect 6493 151029 6611 151147
rect 6653 151029 6771 151147
rect 6493 133189 6611 133307
rect 6653 133189 6771 133307
rect 6493 133029 6611 133147
rect 6653 133029 6771 133147
rect 6493 115189 6611 115307
rect 6653 115189 6771 115307
rect 6493 115029 6611 115147
rect 6653 115029 6771 115147
rect 6493 97189 6611 97307
rect 6653 97189 6771 97307
rect 6493 97029 6611 97147
rect 6653 97029 6771 97147
rect 6493 79189 6611 79307
rect 6653 79189 6771 79307
rect 6493 79029 6611 79147
rect 6653 79029 6771 79147
rect 6493 61189 6611 61307
rect 6653 61189 6771 61307
rect 6493 61029 6611 61147
rect 6653 61029 6771 61147
rect 6493 43189 6611 43307
rect 6653 43189 6771 43307
rect 6493 43029 6611 43147
rect 6653 43029 6771 43147
rect 6493 25189 6611 25307
rect 6653 25189 6771 25307
rect 6493 25029 6611 25147
rect 6653 25029 6771 25147
rect 6493 7189 6611 7307
rect 6653 7189 6771 7307
rect 6493 7029 6611 7147
rect 6653 7029 6771 7147
rect -3867 -3171 -3749 -3053
rect -3707 -3171 -3589 -3053
rect -3867 -3331 -3749 -3213
rect -3707 -3331 -3589 -3213
rect 9913 352781 10031 352899
rect 10073 352781 10191 352899
rect 9913 352621 10031 352739
rect 10073 352621 10191 352739
rect 9913 334609 10031 334727
rect 10073 334609 10191 334727
rect 9913 334449 10031 334567
rect 10073 334449 10191 334567
rect 9913 316609 10031 316727
rect 10073 316609 10191 316727
rect 9913 316449 10031 316567
rect 10073 316449 10191 316567
rect 9913 298609 10031 298727
rect 10073 298609 10191 298727
rect 9913 298449 10031 298567
rect 10073 298449 10191 298567
rect 9913 280609 10031 280727
rect 10073 280609 10191 280727
rect 9913 280449 10031 280567
rect 10073 280449 10191 280567
rect 9913 262609 10031 262727
rect 10073 262609 10191 262727
rect 9913 262449 10031 262567
rect 10073 262449 10191 262567
rect 9913 244609 10031 244727
rect 10073 244609 10191 244727
rect 9913 244449 10031 244567
rect 10073 244449 10191 244567
rect 9913 226609 10031 226727
rect 10073 226609 10191 226727
rect 9913 226449 10031 226567
rect 10073 226449 10191 226567
rect 9913 208609 10031 208727
rect 10073 208609 10191 208727
rect 9913 208449 10031 208567
rect 10073 208449 10191 208567
rect 9913 190609 10031 190727
rect 10073 190609 10191 190727
rect 9913 190449 10031 190567
rect 10073 190449 10191 190567
rect 9913 172609 10031 172727
rect 10073 172609 10191 172727
rect 9913 172449 10031 172567
rect 10073 172449 10191 172567
rect 9913 154609 10031 154727
rect 10073 154609 10191 154727
rect 9913 154449 10031 154567
rect 10073 154449 10191 154567
rect 9913 136609 10031 136727
rect 10073 136609 10191 136727
rect 9913 136449 10031 136567
rect 10073 136449 10191 136567
rect 9913 118609 10031 118727
rect 10073 118609 10191 118727
rect 9913 118449 10031 118567
rect 10073 118449 10191 118567
rect 9913 100609 10031 100727
rect 10073 100609 10191 100727
rect 9913 100449 10031 100567
rect 10073 100449 10191 100567
rect 9913 82609 10031 82727
rect 10073 82609 10191 82727
rect 9913 82449 10031 82567
rect 10073 82449 10191 82567
rect 9913 64609 10031 64727
rect 10073 64609 10191 64727
rect 9913 64449 10031 64567
rect 10073 64449 10191 64567
rect 9913 46609 10031 46727
rect 10073 46609 10191 46727
rect 9913 46449 10031 46567
rect 10073 46449 10191 46567
rect 9913 28609 10031 28727
rect 10073 28609 10191 28727
rect 9913 28449 10031 28567
rect 10073 28449 10191 28567
rect 9913 10609 10031 10727
rect 10073 10609 10191 10727
rect 9913 10449 10031 10567
rect 10073 10449 10191 10567
rect 9913 -771 10031 -653
rect 10073 -771 10191 -653
rect 9913 -931 10031 -813
rect 10073 -931 10191 -813
rect 11773 336469 11891 336587
rect 11933 336469 12051 336587
rect 11773 336309 11891 336427
rect 11933 336309 12051 336427
rect 11773 318469 11891 318587
rect 11933 318469 12051 318587
rect 11773 318309 11891 318427
rect 11933 318309 12051 318427
rect 11773 300469 11891 300587
rect 11933 300469 12051 300587
rect 11773 300309 11891 300427
rect 11933 300309 12051 300427
rect 11773 282469 11891 282587
rect 11933 282469 12051 282587
rect 11773 282309 11891 282427
rect 11933 282309 12051 282427
rect 11773 264469 11891 264587
rect 11933 264469 12051 264587
rect 11773 264309 11891 264427
rect 11933 264309 12051 264427
rect 11773 246469 11891 246587
rect 11933 246469 12051 246587
rect 11773 246309 11891 246427
rect 11933 246309 12051 246427
rect 11773 228469 11891 228587
rect 11933 228469 12051 228587
rect 11773 228309 11891 228427
rect 11933 228309 12051 228427
rect 11773 210469 11891 210587
rect 11933 210469 12051 210587
rect 11773 210309 11891 210427
rect 11933 210309 12051 210427
rect 11773 192469 11891 192587
rect 11933 192469 12051 192587
rect 11773 192309 11891 192427
rect 11933 192309 12051 192427
rect 11773 174469 11891 174587
rect 11933 174469 12051 174587
rect 11773 174309 11891 174427
rect 11933 174309 12051 174427
rect 11773 156469 11891 156587
rect 11933 156469 12051 156587
rect 11773 156309 11891 156427
rect 11933 156309 12051 156427
rect 11773 138469 11891 138587
rect 11933 138469 12051 138587
rect 11773 138309 11891 138427
rect 11933 138309 12051 138427
rect 11773 120469 11891 120587
rect 11933 120469 12051 120587
rect 11773 120309 11891 120427
rect 11933 120309 12051 120427
rect 11773 102469 11891 102587
rect 11933 102469 12051 102587
rect 11773 102309 11891 102427
rect 11933 102309 12051 102427
rect 11773 84469 11891 84587
rect 11933 84469 12051 84587
rect 11773 84309 11891 84427
rect 11933 84309 12051 84427
rect 11773 66469 11891 66587
rect 11933 66469 12051 66587
rect 11773 66309 11891 66427
rect 11933 66309 12051 66427
rect 11773 48469 11891 48587
rect 11933 48469 12051 48587
rect 11773 48309 11891 48427
rect 11933 48309 12051 48427
rect 11773 30469 11891 30587
rect 11933 30469 12051 30587
rect 11773 30309 11891 30427
rect 11933 30309 12051 30427
rect 11773 12469 11891 12587
rect 11933 12469 12051 12587
rect 11773 12309 11891 12427
rect 11933 12309 12051 12427
rect 11773 -1731 11891 -1613
rect 11933 -1731 12051 -1613
rect 11773 -1891 11891 -1773
rect 11933 -1891 12051 -1773
rect 13633 338329 13751 338447
rect 13793 338329 13911 338447
rect 13633 338169 13751 338287
rect 13793 338169 13911 338287
rect 13633 320329 13751 320447
rect 13793 320329 13911 320447
rect 13633 320169 13751 320287
rect 13793 320169 13911 320287
rect 13633 302329 13751 302447
rect 13793 302329 13911 302447
rect 13633 302169 13751 302287
rect 13793 302169 13911 302287
rect 13633 284329 13751 284447
rect 13793 284329 13911 284447
rect 13633 284169 13751 284287
rect 13793 284169 13911 284287
rect 13633 266329 13751 266447
rect 13793 266329 13911 266447
rect 13633 266169 13751 266287
rect 13793 266169 13911 266287
rect 13633 248329 13751 248447
rect 13793 248329 13911 248447
rect 13633 248169 13751 248287
rect 13793 248169 13911 248287
rect 13633 230329 13751 230447
rect 13793 230329 13911 230447
rect 13633 230169 13751 230287
rect 13793 230169 13911 230287
rect 13633 212329 13751 212447
rect 13793 212329 13911 212447
rect 13633 212169 13751 212287
rect 13793 212169 13911 212287
rect 13633 194329 13751 194447
rect 13793 194329 13911 194447
rect 13633 194169 13751 194287
rect 13793 194169 13911 194287
rect 13633 176329 13751 176447
rect 13793 176329 13911 176447
rect 13633 176169 13751 176287
rect 13793 176169 13911 176287
rect 13633 158329 13751 158447
rect 13793 158329 13911 158447
rect 13633 158169 13751 158287
rect 13793 158169 13911 158287
rect 13633 140329 13751 140447
rect 13793 140329 13911 140447
rect 13633 140169 13751 140287
rect 13793 140169 13911 140287
rect 13633 122329 13751 122447
rect 13793 122329 13911 122447
rect 13633 122169 13751 122287
rect 13793 122169 13911 122287
rect 13633 104329 13751 104447
rect 13793 104329 13911 104447
rect 13633 104169 13751 104287
rect 13793 104169 13911 104287
rect 13633 86329 13751 86447
rect 13793 86329 13911 86447
rect 13633 86169 13751 86287
rect 13793 86169 13911 86287
rect 13633 68329 13751 68447
rect 13793 68329 13911 68447
rect 13633 68169 13751 68287
rect 13793 68169 13911 68287
rect 13633 50329 13751 50447
rect 13793 50329 13911 50447
rect 13633 50169 13751 50287
rect 13793 50169 13911 50287
rect 13633 32329 13751 32447
rect 13793 32329 13911 32447
rect 13633 32169 13751 32287
rect 13793 32169 13911 32287
rect 13633 14329 13751 14447
rect 13793 14329 13911 14447
rect 13633 14169 13751 14287
rect 13793 14169 13911 14287
rect 13633 -2691 13751 -2573
rect 13793 -2691 13911 -2573
rect 13633 -2851 13751 -2733
rect 13793 -2851 13911 -2733
rect 24493 355181 24611 355299
rect 24653 355181 24771 355299
rect 24493 355021 24611 355139
rect 24653 355021 24771 355139
rect 22633 354221 22751 354339
rect 22793 354221 22911 354339
rect 22633 354061 22751 354179
rect 22793 354061 22911 354179
rect 20773 353261 20891 353379
rect 20933 353261 21051 353379
rect 20773 353101 20891 353219
rect 20933 353101 21051 353219
rect 15493 340189 15611 340307
rect 15653 340189 15771 340307
rect 15493 340029 15611 340147
rect 15653 340029 15771 340147
rect 15493 322189 15611 322307
rect 15653 322189 15771 322307
rect 15493 322029 15611 322147
rect 15653 322029 15771 322147
rect 15493 304189 15611 304307
rect 15653 304189 15771 304307
rect 15493 304029 15611 304147
rect 15653 304029 15771 304147
rect 15493 286189 15611 286307
rect 15653 286189 15771 286307
rect 15493 286029 15611 286147
rect 15653 286029 15771 286147
rect 15493 268189 15611 268307
rect 15653 268189 15771 268307
rect 15493 268029 15611 268147
rect 15653 268029 15771 268147
rect 15493 250189 15611 250307
rect 15653 250189 15771 250307
rect 15493 250029 15611 250147
rect 15653 250029 15771 250147
rect 15493 232189 15611 232307
rect 15653 232189 15771 232307
rect 15493 232029 15611 232147
rect 15653 232029 15771 232147
rect 15493 214189 15611 214307
rect 15653 214189 15771 214307
rect 15493 214029 15611 214147
rect 15653 214029 15771 214147
rect 15493 196189 15611 196307
rect 15653 196189 15771 196307
rect 15493 196029 15611 196147
rect 15653 196029 15771 196147
rect 15493 178189 15611 178307
rect 15653 178189 15771 178307
rect 15493 178029 15611 178147
rect 15653 178029 15771 178147
rect 15493 160189 15611 160307
rect 15653 160189 15771 160307
rect 15493 160029 15611 160147
rect 15653 160029 15771 160147
rect 15493 142189 15611 142307
rect 15653 142189 15771 142307
rect 15493 142029 15611 142147
rect 15653 142029 15771 142147
rect 15493 124189 15611 124307
rect 15653 124189 15771 124307
rect 15493 124029 15611 124147
rect 15653 124029 15771 124147
rect 15493 106189 15611 106307
rect 15653 106189 15771 106307
rect 15493 106029 15611 106147
rect 15653 106029 15771 106147
rect 15493 88189 15611 88307
rect 15653 88189 15771 88307
rect 15493 88029 15611 88147
rect 15653 88029 15771 88147
rect 15493 70189 15611 70307
rect 15653 70189 15771 70307
rect 15493 70029 15611 70147
rect 15653 70029 15771 70147
rect 15493 52189 15611 52307
rect 15653 52189 15771 52307
rect 15493 52029 15611 52147
rect 15653 52029 15771 52147
rect 15493 34189 15611 34307
rect 15653 34189 15771 34307
rect 15493 34029 15611 34147
rect 15653 34029 15771 34147
rect 15493 16189 15611 16307
rect 15653 16189 15771 16307
rect 15493 16029 15611 16147
rect 15653 16029 15771 16147
rect 6493 -3171 6611 -3053
rect 6653 -3171 6771 -3053
rect 6493 -3331 6611 -3213
rect 6653 -3331 6771 -3213
rect -4347 -3651 -4229 -3533
rect -4187 -3651 -4069 -3533
rect -4347 -3811 -4229 -3693
rect -4187 -3811 -4069 -3693
rect 18913 352301 19031 352419
rect 19073 352301 19191 352419
rect 18913 352141 19031 352259
rect 19073 352141 19191 352259
rect 18913 343609 19031 343727
rect 19073 343609 19191 343727
rect 18913 343449 19031 343567
rect 19073 343449 19191 343567
rect 18913 325609 19031 325727
rect 19073 325609 19191 325727
rect 18913 325449 19031 325567
rect 19073 325449 19191 325567
rect 18913 307609 19031 307727
rect 19073 307609 19191 307727
rect 18913 307449 19031 307567
rect 19073 307449 19191 307567
rect 18913 289609 19031 289727
rect 19073 289609 19191 289727
rect 18913 289449 19031 289567
rect 19073 289449 19191 289567
rect 18913 271609 19031 271727
rect 19073 271609 19191 271727
rect 18913 271449 19031 271567
rect 19073 271449 19191 271567
rect 18913 253609 19031 253727
rect 19073 253609 19191 253727
rect 18913 253449 19031 253567
rect 19073 253449 19191 253567
rect 18913 235609 19031 235727
rect 19073 235609 19191 235727
rect 18913 235449 19031 235567
rect 19073 235449 19191 235567
rect 18913 217609 19031 217727
rect 19073 217609 19191 217727
rect 18913 217449 19031 217567
rect 19073 217449 19191 217567
rect 18913 199609 19031 199727
rect 19073 199609 19191 199727
rect 18913 199449 19031 199567
rect 19073 199449 19191 199567
rect 18913 181609 19031 181727
rect 19073 181609 19191 181727
rect 18913 181449 19031 181567
rect 19073 181449 19191 181567
rect 18913 163609 19031 163727
rect 19073 163609 19191 163727
rect 18913 163449 19031 163567
rect 19073 163449 19191 163567
rect 18913 145609 19031 145727
rect 19073 145609 19191 145727
rect 18913 145449 19031 145567
rect 19073 145449 19191 145567
rect 18913 127609 19031 127727
rect 19073 127609 19191 127727
rect 18913 127449 19031 127567
rect 19073 127449 19191 127567
rect 18913 109609 19031 109727
rect 19073 109609 19191 109727
rect 18913 109449 19031 109567
rect 19073 109449 19191 109567
rect 18913 91609 19031 91727
rect 19073 91609 19191 91727
rect 18913 91449 19031 91567
rect 19073 91449 19191 91567
rect 18913 73609 19031 73727
rect 19073 73609 19191 73727
rect 18913 73449 19031 73567
rect 19073 73449 19191 73567
rect 18913 55609 19031 55727
rect 19073 55609 19191 55727
rect 18913 55449 19031 55567
rect 19073 55449 19191 55567
rect 18913 37609 19031 37727
rect 19073 37609 19191 37727
rect 18913 37449 19031 37567
rect 19073 37449 19191 37567
rect 18913 19609 19031 19727
rect 19073 19609 19191 19727
rect 18913 19449 19031 19567
rect 19073 19449 19191 19567
rect 18913 1609 19031 1727
rect 19073 1609 19191 1727
rect 18913 1449 19031 1567
rect 19073 1449 19191 1567
rect 18913 -291 19031 -173
rect 19073 -291 19191 -173
rect 18913 -451 19031 -333
rect 19073 -451 19191 -333
rect 20773 345469 20891 345587
rect 20933 345469 21051 345587
rect 20773 345309 20891 345427
rect 20933 345309 21051 345427
rect 20773 327469 20891 327587
rect 20933 327469 21051 327587
rect 20773 327309 20891 327427
rect 20933 327309 21051 327427
rect 20773 309469 20891 309587
rect 20933 309469 21051 309587
rect 20773 309309 20891 309427
rect 20933 309309 21051 309427
rect 20773 291469 20891 291587
rect 20933 291469 21051 291587
rect 20773 291309 20891 291427
rect 20933 291309 21051 291427
rect 20773 273469 20891 273587
rect 20933 273469 21051 273587
rect 20773 273309 20891 273427
rect 20933 273309 21051 273427
rect 20773 255469 20891 255587
rect 20933 255469 21051 255587
rect 20773 255309 20891 255427
rect 20933 255309 21051 255427
rect 20773 237469 20891 237587
rect 20933 237469 21051 237587
rect 20773 237309 20891 237427
rect 20933 237309 21051 237427
rect 20773 219469 20891 219587
rect 20933 219469 21051 219587
rect 20773 219309 20891 219427
rect 20933 219309 21051 219427
rect 20773 201469 20891 201587
rect 20933 201469 21051 201587
rect 20773 201309 20891 201427
rect 20933 201309 21051 201427
rect 20773 183469 20891 183587
rect 20933 183469 21051 183587
rect 20773 183309 20891 183427
rect 20933 183309 21051 183427
rect 20773 165469 20891 165587
rect 20933 165469 21051 165587
rect 20773 165309 20891 165427
rect 20933 165309 21051 165427
rect 20773 147469 20891 147587
rect 20933 147469 21051 147587
rect 20773 147309 20891 147427
rect 20933 147309 21051 147427
rect 20773 129469 20891 129587
rect 20933 129469 21051 129587
rect 20773 129309 20891 129427
rect 20933 129309 21051 129427
rect 20773 111469 20891 111587
rect 20933 111469 21051 111587
rect 20773 111309 20891 111427
rect 20933 111309 21051 111427
rect 20773 93469 20891 93587
rect 20933 93469 21051 93587
rect 20773 93309 20891 93427
rect 20933 93309 21051 93427
rect 20773 75469 20891 75587
rect 20933 75469 21051 75587
rect 20773 75309 20891 75427
rect 20933 75309 21051 75427
rect 20773 57469 20891 57587
rect 20933 57469 21051 57587
rect 20773 57309 20891 57427
rect 20933 57309 21051 57427
rect 20773 39469 20891 39587
rect 20933 39469 21051 39587
rect 20773 39309 20891 39427
rect 20933 39309 21051 39427
rect 20773 21469 20891 21587
rect 20933 21469 21051 21587
rect 20773 21309 20891 21427
rect 20933 21309 21051 21427
rect 20773 3469 20891 3587
rect 20933 3469 21051 3587
rect 20773 3309 20891 3427
rect 20933 3309 21051 3427
rect 20773 -1251 20891 -1133
rect 20933 -1251 21051 -1133
rect 20773 -1411 20891 -1293
rect 20933 -1411 21051 -1293
rect 22633 347329 22751 347447
rect 22793 347329 22911 347447
rect 22633 347169 22751 347287
rect 22793 347169 22911 347287
rect 22633 329329 22751 329447
rect 22793 329329 22911 329447
rect 22633 329169 22751 329287
rect 22793 329169 22911 329287
rect 22633 311329 22751 311447
rect 22793 311329 22911 311447
rect 22633 311169 22751 311287
rect 22793 311169 22911 311287
rect 22633 293329 22751 293447
rect 22793 293329 22911 293447
rect 22633 293169 22751 293287
rect 22793 293169 22911 293287
rect 22633 275329 22751 275447
rect 22793 275329 22911 275447
rect 22633 275169 22751 275287
rect 22793 275169 22911 275287
rect 22633 257329 22751 257447
rect 22793 257329 22911 257447
rect 22633 257169 22751 257287
rect 22793 257169 22911 257287
rect 22633 239329 22751 239447
rect 22793 239329 22911 239447
rect 22633 239169 22751 239287
rect 22793 239169 22911 239287
rect 22633 221329 22751 221447
rect 22793 221329 22911 221447
rect 22633 221169 22751 221287
rect 22793 221169 22911 221287
rect 22633 203329 22751 203447
rect 22793 203329 22911 203447
rect 22633 203169 22751 203287
rect 22793 203169 22911 203287
rect 22633 185329 22751 185447
rect 22793 185329 22911 185447
rect 22633 185169 22751 185287
rect 22793 185169 22911 185287
rect 22633 167329 22751 167447
rect 22793 167329 22911 167447
rect 22633 167169 22751 167287
rect 22793 167169 22911 167287
rect 22633 149329 22751 149447
rect 22793 149329 22911 149447
rect 22633 149169 22751 149287
rect 22793 149169 22911 149287
rect 22633 131329 22751 131447
rect 22793 131329 22911 131447
rect 22633 131169 22751 131287
rect 22793 131169 22911 131287
rect 22633 113329 22751 113447
rect 22793 113329 22911 113447
rect 22633 113169 22751 113287
rect 22793 113169 22911 113287
rect 22633 95329 22751 95447
rect 22793 95329 22911 95447
rect 22633 95169 22751 95287
rect 22793 95169 22911 95287
rect 22633 77329 22751 77447
rect 22793 77329 22911 77447
rect 22633 77169 22751 77287
rect 22793 77169 22911 77287
rect 22633 59329 22751 59447
rect 22793 59329 22911 59447
rect 22633 59169 22751 59287
rect 22793 59169 22911 59287
rect 22633 41329 22751 41447
rect 22793 41329 22911 41447
rect 22633 41169 22751 41287
rect 22793 41169 22911 41287
rect 22633 23329 22751 23447
rect 22793 23329 22911 23447
rect 22633 23169 22751 23287
rect 22793 23169 22911 23287
rect 22633 5329 22751 5447
rect 22793 5329 22911 5447
rect 22633 5169 22751 5287
rect 22793 5169 22911 5287
rect 22633 -2211 22751 -2093
rect 22793 -2211 22911 -2093
rect 22633 -2371 22751 -2253
rect 22793 -2371 22911 -2253
rect 33493 355661 33611 355779
rect 33653 355661 33771 355779
rect 33493 355501 33611 355619
rect 33653 355501 33771 355619
rect 31633 354701 31751 354819
rect 31793 354701 31911 354819
rect 31633 354541 31751 354659
rect 31793 354541 31911 354659
rect 29773 353741 29891 353859
rect 29933 353741 30051 353859
rect 29773 353581 29891 353699
rect 29933 353581 30051 353699
rect 24493 349189 24611 349307
rect 24653 349189 24771 349307
rect 24493 349029 24611 349147
rect 24653 349029 24771 349147
rect 24493 331189 24611 331307
rect 24653 331189 24771 331307
rect 24493 331029 24611 331147
rect 24653 331029 24771 331147
rect 24493 313189 24611 313307
rect 24653 313189 24771 313307
rect 24493 313029 24611 313147
rect 24653 313029 24771 313147
rect 24493 295189 24611 295307
rect 24653 295189 24771 295307
rect 24493 295029 24611 295147
rect 24653 295029 24771 295147
rect 24493 277189 24611 277307
rect 24653 277189 24771 277307
rect 24493 277029 24611 277147
rect 24653 277029 24771 277147
rect 24493 259189 24611 259307
rect 24653 259189 24771 259307
rect 24493 259029 24611 259147
rect 24653 259029 24771 259147
rect 24493 241189 24611 241307
rect 24653 241189 24771 241307
rect 24493 241029 24611 241147
rect 24653 241029 24771 241147
rect 24493 223189 24611 223307
rect 24653 223189 24771 223307
rect 24493 223029 24611 223147
rect 24653 223029 24771 223147
rect 24493 205189 24611 205307
rect 24653 205189 24771 205307
rect 24493 205029 24611 205147
rect 24653 205029 24771 205147
rect 24493 187189 24611 187307
rect 24653 187189 24771 187307
rect 24493 187029 24611 187147
rect 24653 187029 24771 187147
rect 24493 169189 24611 169307
rect 24653 169189 24771 169307
rect 24493 169029 24611 169147
rect 24653 169029 24771 169147
rect 24493 151189 24611 151307
rect 24653 151189 24771 151307
rect 24493 151029 24611 151147
rect 24653 151029 24771 151147
rect 24493 133189 24611 133307
rect 24653 133189 24771 133307
rect 24493 133029 24611 133147
rect 24653 133029 24771 133147
rect 24493 115189 24611 115307
rect 24653 115189 24771 115307
rect 24493 115029 24611 115147
rect 24653 115029 24771 115147
rect 24493 97189 24611 97307
rect 24653 97189 24771 97307
rect 24493 97029 24611 97147
rect 24653 97029 24771 97147
rect 24493 79189 24611 79307
rect 24653 79189 24771 79307
rect 24493 79029 24611 79147
rect 24653 79029 24771 79147
rect 24493 61189 24611 61307
rect 24653 61189 24771 61307
rect 24493 61029 24611 61147
rect 24653 61029 24771 61147
rect 24493 43189 24611 43307
rect 24653 43189 24771 43307
rect 24493 43029 24611 43147
rect 24653 43029 24771 43147
rect 24493 25189 24611 25307
rect 24653 25189 24771 25307
rect 24493 25029 24611 25147
rect 24653 25029 24771 25147
rect 24493 7189 24611 7307
rect 24653 7189 24771 7307
rect 24493 7029 24611 7147
rect 24653 7029 24771 7147
rect 15493 -3651 15611 -3533
rect 15653 -3651 15771 -3533
rect 15493 -3811 15611 -3693
rect 15653 -3811 15771 -3693
rect 27913 352781 28031 352899
rect 28073 352781 28191 352899
rect 27913 352621 28031 352739
rect 28073 352621 28191 352739
rect 27913 334609 28031 334727
rect 28073 334609 28191 334727
rect 27913 334449 28031 334567
rect 28073 334449 28191 334567
rect 27913 316609 28031 316727
rect 28073 316609 28191 316727
rect 27913 316449 28031 316567
rect 28073 316449 28191 316567
rect 27913 298609 28031 298727
rect 28073 298609 28191 298727
rect 27913 298449 28031 298567
rect 28073 298449 28191 298567
rect 27913 280609 28031 280727
rect 28073 280609 28191 280727
rect 27913 280449 28031 280567
rect 28073 280449 28191 280567
rect 27913 262609 28031 262727
rect 28073 262609 28191 262727
rect 27913 262449 28031 262567
rect 28073 262449 28191 262567
rect 27913 244609 28031 244727
rect 28073 244609 28191 244727
rect 27913 244449 28031 244567
rect 28073 244449 28191 244567
rect 27913 226609 28031 226727
rect 28073 226609 28191 226727
rect 27913 226449 28031 226567
rect 28073 226449 28191 226567
rect 27913 208609 28031 208727
rect 28073 208609 28191 208727
rect 27913 208449 28031 208567
rect 28073 208449 28191 208567
rect 27913 190609 28031 190727
rect 28073 190609 28191 190727
rect 27913 190449 28031 190567
rect 28073 190449 28191 190567
rect 27913 172609 28031 172727
rect 28073 172609 28191 172727
rect 27913 172449 28031 172567
rect 28073 172449 28191 172567
rect 27913 154609 28031 154727
rect 28073 154609 28191 154727
rect 27913 154449 28031 154567
rect 28073 154449 28191 154567
rect 27913 136609 28031 136727
rect 28073 136609 28191 136727
rect 27913 136449 28031 136567
rect 28073 136449 28191 136567
rect 27913 118609 28031 118727
rect 28073 118609 28191 118727
rect 27913 118449 28031 118567
rect 28073 118449 28191 118567
rect 27913 100609 28031 100727
rect 28073 100609 28191 100727
rect 27913 100449 28031 100567
rect 28073 100449 28191 100567
rect 27913 82609 28031 82727
rect 28073 82609 28191 82727
rect 27913 82449 28031 82567
rect 28073 82449 28191 82567
rect 27913 64609 28031 64727
rect 28073 64609 28191 64727
rect 27913 64449 28031 64567
rect 28073 64449 28191 64567
rect 27913 46609 28031 46727
rect 28073 46609 28191 46727
rect 27913 46449 28031 46567
rect 28073 46449 28191 46567
rect 27913 28609 28031 28727
rect 28073 28609 28191 28727
rect 27913 28449 28031 28567
rect 28073 28449 28191 28567
rect 27913 10609 28031 10727
rect 28073 10609 28191 10727
rect 27913 10449 28031 10567
rect 28073 10449 28191 10567
rect 27913 -771 28031 -653
rect 28073 -771 28191 -653
rect 27913 -931 28031 -813
rect 28073 -931 28191 -813
rect 29773 336469 29891 336587
rect 29933 336469 30051 336587
rect 29773 336309 29891 336427
rect 29933 336309 30051 336427
rect 29773 318469 29891 318587
rect 29933 318469 30051 318587
rect 29773 318309 29891 318427
rect 29933 318309 30051 318427
rect 29773 300469 29891 300587
rect 29933 300469 30051 300587
rect 29773 300309 29891 300427
rect 29933 300309 30051 300427
rect 29773 282469 29891 282587
rect 29933 282469 30051 282587
rect 29773 282309 29891 282427
rect 29933 282309 30051 282427
rect 29773 264469 29891 264587
rect 29933 264469 30051 264587
rect 29773 264309 29891 264427
rect 29933 264309 30051 264427
rect 29773 246469 29891 246587
rect 29933 246469 30051 246587
rect 29773 246309 29891 246427
rect 29933 246309 30051 246427
rect 29773 228469 29891 228587
rect 29933 228469 30051 228587
rect 29773 228309 29891 228427
rect 29933 228309 30051 228427
rect 29773 210469 29891 210587
rect 29933 210469 30051 210587
rect 29773 210309 29891 210427
rect 29933 210309 30051 210427
rect 29773 192469 29891 192587
rect 29933 192469 30051 192587
rect 29773 192309 29891 192427
rect 29933 192309 30051 192427
rect 29773 174469 29891 174587
rect 29933 174469 30051 174587
rect 29773 174309 29891 174427
rect 29933 174309 30051 174427
rect 29773 156469 29891 156587
rect 29933 156469 30051 156587
rect 29773 156309 29891 156427
rect 29933 156309 30051 156427
rect 29773 138469 29891 138587
rect 29933 138469 30051 138587
rect 29773 138309 29891 138427
rect 29933 138309 30051 138427
rect 29773 120469 29891 120587
rect 29933 120469 30051 120587
rect 29773 120309 29891 120427
rect 29933 120309 30051 120427
rect 29773 102469 29891 102587
rect 29933 102469 30051 102587
rect 29773 102309 29891 102427
rect 29933 102309 30051 102427
rect 29773 84469 29891 84587
rect 29933 84469 30051 84587
rect 29773 84309 29891 84427
rect 29933 84309 30051 84427
rect 29773 66469 29891 66587
rect 29933 66469 30051 66587
rect 29773 66309 29891 66427
rect 29933 66309 30051 66427
rect 29773 48469 29891 48587
rect 29933 48469 30051 48587
rect 29773 48309 29891 48427
rect 29933 48309 30051 48427
rect 29773 30469 29891 30587
rect 29933 30469 30051 30587
rect 29773 30309 29891 30427
rect 29933 30309 30051 30427
rect 29773 12469 29891 12587
rect 29933 12469 30051 12587
rect 29773 12309 29891 12427
rect 29933 12309 30051 12427
rect 29773 -1731 29891 -1613
rect 29933 -1731 30051 -1613
rect 29773 -1891 29891 -1773
rect 29933 -1891 30051 -1773
rect 31633 338329 31751 338447
rect 31793 338329 31911 338447
rect 31633 338169 31751 338287
rect 31793 338169 31911 338287
rect 31633 320329 31751 320447
rect 31793 320329 31911 320447
rect 31633 320169 31751 320287
rect 31793 320169 31911 320287
rect 31633 302329 31751 302447
rect 31793 302329 31911 302447
rect 31633 302169 31751 302287
rect 31793 302169 31911 302287
rect 31633 284329 31751 284447
rect 31793 284329 31911 284447
rect 31633 284169 31751 284287
rect 31793 284169 31911 284287
rect 31633 266329 31751 266447
rect 31793 266329 31911 266447
rect 31633 266169 31751 266287
rect 31793 266169 31911 266287
rect 31633 248329 31751 248447
rect 31793 248329 31911 248447
rect 31633 248169 31751 248287
rect 31793 248169 31911 248287
rect 31633 230329 31751 230447
rect 31793 230329 31911 230447
rect 31633 230169 31751 230287
rect 31793 230169 31911 230287
rect 31633 212329 31751 212447
rect 31793 212329 31911 212447
rect 31633 212169 31751 212287
rect 31793 212169 31911 212287
rect 31633 194329 31751 194447
rect 31793 194329 31911 194447
rect 31633 194169 31751 194287
rect 31793 194169 31911 194287
rect 31633 176329 31751 176447
rect 31793 176329 31911 176447
rect 31633 176169 31751 176287
rect 31793 176169 31911 176287
rect 31633 158329 31751 158447
rect 31793 158329 31911 158447
rect 31633 158169 31751 158287
rect 31793 158169 31911 158287
rect 31633 140329 31751 140447
rect 31793 140329 31911 140447
rect 31633 140169 31751 140287
rect 31793 140169 31911 140287
rect 31633 122329 31751 122447
rect 31793 122329 31911 122447
rect 31633 122169 31751 122287
rect 31793 122169 31911 122287
rect 31633 104329 31751 104447
rect 31793 104329 31911 104447
rect 31633 104169 31751 104287
rect 31793 104169 31911 104287
rect 31633 86329 31751 86447
rect 31793 86329 31911 86447
rect 31633 86169 31751 86287
rect 31793 86169 31911 86287
rect 31633 68329 31751 68447
rect 31793 68329 31911 68447
rect 31633 68169 31751 68287
rect 31793 68169 31911 68287
rect 31633 50329 31751 50447
rect 31793 50329 31911 50447
rect 31633 50169 31751 50287
rect 31793 50169 31911 50287
rect 31633 32329 31751 32447
rect 31793 32329 31911 32447
rect 31633 32169 31751 32287
rect 31793 32169 31911 32287
rect 31633 14329 31751 14447
rect 31793 14329 31911 14447
rect 31633 14169 31751 14287
rect 31793 14169 31911 14287
rect 31633 -2691 31751 -2573
rect 31793 -2691 31911 -2573
rect 31633 -2851 31751 -2733
rect 31793 -2851 31911 -2733
rect 42493 355181 42611 355299
rect 42653 355181 42771 355299
rect 42493 355021 42611 355139
rect 42653 355021 42771 355139
rect 40633 354221 40751 354339
rect 40793 354221 40911 354339
rect 40633 354061 40751 354179
rect 40793 354061 40911 354179
rect 38773 353261 38891 353379
rect 38933 353261 39051 353379
rect 38773 353101 38891 353219
rect 38933 353101 39051 353219
rect 33493 340189 33611 340307
rect 33653 340189 33771 340307
rect 33493 340029 33611 340147
rect 33653 340029 33771 340147
rect 33493 322189 33611 322307
rect 33653 322189 33771 322307
rect 33493 322029 33611 322147
rect 33653 322029 33771 322147
rect 33493 304189 33611 304307
rect 33653 304189 33771 304307
rect 33493 304029 33611 304147
rect 33653 304029 33771 304147
rect 33493 286189 33611 286307
rect 33653 286189 33771 286307
rect 33493 286029 33611 286147
rect 33653 286029 33771 286147
rect 33493 268189 33611 268307
rect 33653 268189 33771 268307
rect 33493 268029 33611 268147
rect 33653 268029 33771 268147
rect 33493 250189 33611 250307
rect 33653 250189 33771 250307
rect 33493 250029 33611 250147
rect 33653 250029 33771 250147
rect 33493 232189 33611 232307
rect 33653 232189 33771 232307
rect 33493 232029 33611 232147
rect 33653 232029 33771 232147
rect 33493 214189 33611 214307
rect 33653 214189 33771 214307
rect 33493 214029 33611 214147
rect 33653 214029 33771 214147
rect 33493 196189 33611 196307
rect 33653 196189 33771 196307
rect 33493 196029 33611 196147
rect 33653 196029 33771 196147
rect 33493 178189 33611 178307
rect 33653 178189 33771 178307
rect 33493 178029 33611 178147
rect 33653 178029 33771 178147
rect 33493 160189 33611 160307
rect 33653 160189 33771 160307
rect 33493 160029 33611 160147
rect 33653 160029 33771 160147
rect 33493 142189 33611 142307
rect 33653 142189 33771 142307
rect 33493 142029 33611 142147
rect 33653 142029 33771 142147
rect 33493 124189 33611 124307
rect 33653 124189 33771 124307
rect 33493 124029 33611 124147
rect 33653 124029 33771 124147
rect 33493 106189 33611 106307
rect 33653 106189 33771 106307
rect 33493 106029 33611 106147
rect 33653 106029 33771 106147
rect 33493 88189 33611 88307
rect 33653 88189 33771 88307
rect 33493 88029 33611 88147
rect 33653 88029 33771 88147
rect 33493 70189 33611 70307
rect 33653 70189 33771 70307
rect 33493 70029 33611 70147
rect 33653 70029 33771 70147
rect 33493 52189 33611 52307
rect 33653 52189 33771 52307
rect 33493 52029 33611 52147
rect 33653 52029 33771 52147
rect 33493 34189 33611 34307
rect 33653 34189 33771 34307
rect 33493 34029 33611 34147
rect 33653 34029 33771 34147
rect 33493 16189 33611 16307
rect 33653 16189 33771 16307
rect 33493 16029 33611 16147
rect 33653 16029 33771 16147
rect 24493 -3171 24611 -3053
rect 24653 -3171 24771 -3053
rect 24493 -3331 24611 -3213
rect 24653 -3331 24771 -3213
rect 36913 352301 37031 352419
rect 37073 352301 37191 352419
rect 36913 352141 37031 352259
rect 37073 352141 37191 352259
rect 36913 343609 37031 343727
rect 37073 343609 37191 343727
rect 36913 343449 37031 343567
rect 37073 343449 37191 343567
rect 36913 325609 37031 325727
rect 37073 325609 37191 325727
rect 36913 325449 37031 325567
rect 37073 325449 37191 325567
rect 36913 307609 37031 307727
rect 37073 307609 37191 307727
rect 36913 307449 37031 307567
rect 37073 307449 37191 307567
rect 36913 289609 37031 289727
rect 37073 289609 37191 289727
rect 36913 289449 37031 289567
rect 37073 289449 37191 289567
rect 36913 271609 37031 271727
rect 37073 271609 37191 271727
rect 36913 271449 37031 271567
rect 37073 271449 37191 271567
rect 36913 253609 37031 253727
rect 37073 253609 37191 253727
rect 36913 253449 37031 253567
rect 37073 253449 37191 253567
rect 36913 235609 37031 235727
rect 37073 235609 37191 235727
rect 36913 235449 37031 235567
rect 37073 235449 37191 235567
rect 36913 217609 37031 217727
rect 37073 217609 37191 217727
rect 36913 217449 37031 217567
rect 37073 217449 37191 217567
rect 36913 199609 37031 199727
rect 37073 199609 37191 199727
rect 36913 199449 37031 199567
rect 37073 199449 37191 199567
rect 36913 181609 37031 181727
rect 37073 181609 37191 181727
rect 36913 181449 37031 181567
rect 37073 181449 37191 181567
rect 36913 163609 37031 163727
rect 37073 163609 37191 163727
rect 36913 163449 37031 163567
rect 37073 163449 37191 163567
rect 36913 145609 37031 145727
rect 37073 145609 37191 145727
rect 36913 145449 37031 145567
rect 37073 145449 37191 145567
rect 36913 127609 37031 127727
rect 37073 127609 37191 127727
rect 36913 127449 37031 127567
rect 37073 127449 37191 127567
rect 36913 109609 37031 109727
rect 37073 109609 37191 109727
rect 36913 109449 37031 109567
rect 37073 109449 37191 109567
rect 36913 91609 37031 91727
rect 37073 91609 37191 91727
rect 36913 91449 37031 91567
rect 37073 91449 37191 91567
rect 36913 73609 37031 73727
rect 37073 73609 37191 73727
rect 36913 73449 37031 73567
rect 37073 73449 37191 73567
rect 36913 55609 37031 55727
rect 37073 55609 37191 55727
rect 36913 55449 37031 55567
rect 37073 55449 37191 55567
rect 36913 37609 37031 37727
rect 37073 37609 37191 37727
rect 36913 37449 37031 37567
rect 37073 37449 37191 37567
rect 36913 19609 37031 19727
rect 37073 19609 37191 19727
rect 36913 19449 37031 19567
rect 37073 19449 37191 19567
rect 36913 1609 37031 1727
rect 37073 1609 37191 1727
rect 36913 1449 37031 1567
rect 37073 1449 37191 1567
rect 36913 -291 37031 -173
rect 37073 -291 37191 -173
rect 36913 -451 37031 -333
rect 37073 -451 37191 -333
rect 38773 345469 38891 345587
rect 38933 345469 39051 345587
rect 38773 345309 38891 345427
rect 38933 345309 39051 345427
rect 38773 327469 38891 327587
rect 38933 327469 39051 327587
rect 38773 327309 38891 327427
rect 38933 327309 39051 327427
rect 38773 309469 38891 309587
rect 38933 309469 39051 309587
rect 38773 309309 38891 309427
rect 38933 309309 39051 309427
rect 38773 291469 38891 291587
rect 38933 291469 39051 291587
rect 38773 291309 38891 291427
rect 38933 291309 39051 291427
rect 38773 273469 38891 273587
rect 38933 273469 39051 273587
rect 38773 273309 38891 273427
rect 38933 273309 39051 273427
rect 38773 255469 38891 255587
rect 38933 255469 39051 255587
rect 38773 255309 38891 255427
rect 38933 255309 39051 255427
rect 38773 237469 38891 237587
rect 38933 237469 39051 237587
rect 38773 237309 38891 237427
rect 38933 237309 39051 237427
rect 38773 219469 38891 219587
rect 38933 219469 39051 219587
rect 38773 219309 38891 219427
rect 38933 219309 39051 219427
rect 38773 201469 38891 201587
rect 38933 201469 39051 201587
rect 38773 201309 38891 201427
rect 38933 201309 39051 201427
rect 38773 183469 38891 183587
rect 38933 183469 39051 183587
rect 38773 183309 38891 183427
rect 38933 183309 39051 183427
rect 38773 165469 38891 165587
rect 38933 165469 39051 165587
rect 38773 165309 38891 165427
rect 38933 165309 39051 165427
rect 38773 147469 38891 147587
rect 38933 147469 39051 147587
rect 38773 147309 38891 147427
rect 38933 147309 39051 147427
rect 38773 129469 38891 129587
rect 38933 129469 39051 129587
rect 38773 129309 38891 129427
rect 38933 129309 39051 129427
rect 38773 111469 38891 111587
rect 38933 111469 39051 111587
rect 38773 111309 38891 111427
rect 38933 111309 39051 111427
rect 38773 93469 38891 93587
rect 38933 93469 39051 93587
rect 38773 93309 38891 93427
rect 38933 93309 39051 93427
rect 38773 75469 38891 75587
rect 38933 75469 39051 75587
rect 38773 75309 38891 75427
rect 38933 75309 39051 75427
rect 38773 57469 38891 57587
rect 38933 57469 39051 57587
rect 38773 57309 38891 57427
rect 38933 57309 39051 57427
rect 38773 39469 38891 39587
rect 38933 39469 39051 39587
rect 38773 39309 38891 39427
rect 38933 39309 39051 39427
rect 38773 21469 38891 21587
rect 38933 21469 39051 21587
rect 38773 21309 38891 21427
rect 38933 21309 39051 21427
rect 38773 3469 38891 3587
rect 38933 3469 39051 3587
rect 38773 3309 38891 3427
rect 38933 3309 39051 3427
rect 38773 -1251 38891 -1133
rect 38933 -1251 39051 -1133
rect 38773 -1411 38891 -1293
rect 38933 -1411 39051 -1293
rect 40633 347329 40751 347447
rect 40793 347329 40911 347447
rect 40633 347169 40751 347287
rect 40793 347169 40911 347287
rect 40633 329329 40751 329447
rect 40793 329329 40911 329447
rect 40633 329169 40751 329287
rect 40793 329169 40911 329287
rect 40633 311329 40751 311447
rect 40793 311329 40911 311447
rect 40633 311169 40751 311287
rect 40793 311169 40911 311287
rect 40633 293329 40751 293447
rect 40793 293329 40911 293447
rect 40633 293169 40751 293287
rect 40793 293169 40911 293287
rect 40633 275329 40751 275447
rect 40793 275329 40911 275447
rect 40633 275169 40751 275287
rect 40793 275169 40911 275287
rect 40633 257329 40751 257447
rect 40793 257329 40911 257447
rect 40633 257169 40751 257287
rect 40793 257169 40911 257287
rect 40633 239329 40751 239447
rect 40793 239329 40911 239447
rect 40633 239169 40751 239287
rect 40793 239169 40911 239287
rect 40633 221329 40751 221447
rect 40793 221329 40911 221447
rect 40633 221169 40751 221287
rect 40793 221169 40911 221287
rect 40633 203329 40751 203447
rect 40793 203329 40911 203447
rect 40633 203169 40751 203287
rect 40793 203169 40911 203287
rect 40633 185329 40751 185447
rect 40793 185329 40911 185447
rect 40633 185169 40751 185287
rect 40793 185169 40911 185287
rect 40633 167329 40751 167447
rect 40793 167329 40911 167447
rect 40633 167169 40751 167287
rect 40793 167169 40911 167287
rect 40633 149329 40751 149447
rect 40793 149329 40911 149447
rect 40633 149169 40751 149287
rect 40793 149169 40911 149287
rect 40633 131329 40751 131447
rect 40793 131329 40911 131447
rect 40633 131169 40751 131287
rect 40793 131169 40911 131287
rect 40633 113329 40751 113447
rect 40793 113329 40911 113447
rect 40633 113169 40751 113287
rect 40793 113169 40911 113287
rect 40633 95329 40751 95447
rect 40793 95329 40911 95447
rect 40633 95169 40751 95287
rect 40793 95169 40911 95287
rect 40633 77329 40751 77447
rect 40793 77329 40911 77447
rect 40633 77169 40751 77287
rect 40793 77169 40911 77287
rect 40633 59329 40751 59447
rect 40793 59329 40911 59447
rect 40633 59169 40751 59287
rect 40793 59169 40911 59287
rect 40633 41329 40751 41447
rect 40793 41329 40911 41447
rect 40633 41169 40751 41287
rect 40793 41169 40911 41287
rect 40633 23329 40751 23447
rect 40793 23329 40911 23447
rect 40633 23169 40751 23287
rect 40793 23169 40911 23287
rect 40633 5329 40751 5447
rect 40793 5329 40911 5447
rect 40633 5169 40751 5287
rect 40793 5169 40911 5287
rect 40633 -2211 40751 -2093
rect 40793 -2211 40911 -2093
rect 40633 -2371 40751 -2253
rect 40793 -2371 40911 -2253
rect 51493 355661 51611 355779
rect 51653 355661 51771 355779
rect 51493 355501 51611 355619
rect 51653 355501 51771 355619
rect 49633 354701 49751 354819
rect 49793 354701 49911 354819
rect 49633 354541 49751 354659
rect 49793 354541 49911 354659
rect 47773 353741 47891 353859
rect 47933 353741 48051 353859
rect 47773 353581 47891 353699
rect 47933 353581 48051 353699
rect 42493 349189 42611 349307
rect 42653 349189 42771 349307
rect 42493 349029 42611 349147
rect 42653 349029 42771 349147
rect 42493 331189 42611 331307
rect 42653 331189 42771 331307
rect 42493 331029 42611 331147
rect 42653 331029 42771 331147
rect 42493 313189 42611 313307
rect 42653 313189 42771 313307
rect 42493 313029 42611 313147
rect 42653 313029 42771 313147
rect 42493 295189 42611 295307
rect 42653 295189 42771 295307
rect 42493 295029 42611 295147
rect 42653 295029 42771 295147
rect 42493 277189 42611 277307
rect 42653 277189 42771 277307
rect 42493 277029 42611 277147
rect 42653 277029 42771 277147
rect 42493 259189 42611 259307
rect 42653 259189 42771 259307
rect 42493 259029 42611 259147
rect 42653 259029 42771 259147
rect 42493 241189 42611 241307
rect 42653 241189 42771 241307
rect 42493 241029 42611 241147
rect 42653 241029 42771 241147
rect 42493 223189 42611 223307
rect 42653 223189 42771 223307
rect 42493 223029 42611 223147
rect 42653 223029 42771 223147
rect 42493 205189 42611 205307
rect 42653 205189 42771 205307
rect 42493 205029 42611 205147
rect 42653 205029 42771 205147
rect 42493 187189 42611 187307
rect 42653 187189 42771 187307
rect 42493 187029 42611 187147
rect 42653 187029 42771 187147
rect 42493 169189 42611 169307
rect 42653 169189 42771 169307
rect 42493 169029 42611 169147
rect 42653 169029 42771 169147
rect 42493 151189 42611 151307
rect 42653 151189 42771 151307
rect 42493 151029 42611 151147
rect 42653 151029 42771 151147
rect 42493 133189 42611 133307
rect 42653 133189 42771 133307
rect 42493 133029 42611 133147
rect 42653 133029 42771 133147
rect 42493 115189 42611 115307
rect 42653 115189 42771 115307
rect 42493 115029 42611 115147
rect 42653 115029 42771 115147
rect 42493 97189 42611 97307
rect 42653 97189 42771 97307
rect 42493 97029 42611 97147
rect 42653 97029 42771 97147
rect 42493 79189 42611 79307
rect 42653 79189 42771 79307
rect 42493 79029 42611 79147
rect 42653 79029 42771 79147
rect 42493 61189 42611 61307
rect 42653 61189 42771 61307
rect 42493 61029 42611 61147
rect 42653 61029 42771 61147
rect 42493 43189 42611 43307
rect 42653 43189 42771 43307
rect 42493 43029 42611 43147
rect 42653 43029 42771 43147
rect 42493 25189 42611 25307
rect 42653 25189 42771 25307
rect 42493 25029 42611 25147
rect 42653 25029 42771 25147
rect 42493 7189 42611 7307
rect 42653 7189 42771 7307
rect 42493 7029 42611 7147
rect 42653 7029 42771 7147
rect 33493 -3651 33611 -3533
rect 33653 -3651 33771 -3533
rect 33493 -3811 33611 -3693
rect 33653 -3811 33771 -3693
rect 45913 352781 46031 352899
rect 46073 352781 46191 352899
rect 45913 352621 46031 352739
rect 46073 352621 46191 352739
rect 45913 334609 46031 334727
rect 46073 334609 46191 334727
rect 45913 334449 46031 334567
rect 46073 334449 46191 334567
rect 45913 316609 46031 316727
rect 46073 316609 46191 316727
rect 45913 316449 46031 316567
rect 46073 316449 46191 316567
rect 45913 298609 46031 298727
rect 46073 298609 46191 298727
rect 45913 298449 46031 298567
rect 46073 298449 46191 298567
rect 45913 280609 46031 280727
rect 46073 280609 46191 280727
rect 45913 280449 46031 280567
rect 46073 280449 46191 280567
rect 45913 262609 46031 262727
rect 46073 262609 46191 262727
rect 45913 262449 46031 262567
rect 46073 262449 46191 262567
rect 45913 244609 46031 244727
rect 46073 244609 46191 244727
rect 45913 244449 46031 244567
rect 46073 244449 46191 244567
rect 45913 226609 46031 226727
rect 46073 226609 46191 226727
rect 45913 226449 46031 226567
rect 46073 226449 46191 226567
rect 45913 208609 46031 208727
rect 46073 208609 46191 208727
rect 45913 208449 46031 208567
rect 46073 208449 46191 208567
rect 45913 190609 46031 190727
rect 46073 190609 46191 190727
rect 45913 190449 46031 190567
rect 46073 190449 46191 190567
rect 45913 172609 46031 172727
rect 46073 172609 46191 172727
rect 45913 172449 46031 172567
rect 46073 172449 46191 172567
rect 45913 154609 46031 154727
rect 46073 154609 46191 154727
rect 45913 154449 46031 154567
rect 46073 154449 46191 154567
rect 45913 136609 46031 136727
rect 46073 136609 46191 136727
rect 45913 136449 46031 136567
rect 46073 136449 46191 136567
rect 45913 118609 46031 118727
rect 46073 118609 46191 118727
rect 45913 118449 46031 118567
rect 46073 118449 46191 118567
rect 45913 100609 46031 100727
rect 46073 100609 46191 100727
rect 45913 100449 46031 100567
rect 46073 100449 46191 100567
rect 45913 82609 46031 82727
rect 46073 82609 46191 82727
rect 45913 82449 46031 82567
rect 46073 82449 46191 82567
rect 45913 64609 46031 64727
rect 46073 64609 46191 64727
rect 45913 64449 46031 64567
rect 46073 64449 46191 64567
rect 45913 46609 46031 46727
rect 46073 46609 46191 46727
rect 45913 46449 46031 46567
rect 46073 46449 46191 46567
rect 45913 28609 46031 28727
rect 46073 28609 46191 28727
rect 45913 28449 46031 28567
rect 46073 28449 46191 28567
rect 45913 10609 46031 10727
rect 46073 10609 46191 10727
rect 45913 10449 46031 10567
rect 46073 10449 46191 10567
rect 45913 -771 46031 -653
rect 46073 -771 46191 -653
rect 45913 -931 46031 -813
rect 46073 -931 46191 -813
rect 47773 336469 47891 336587
rect 47933 336469 48051 336587
rect 47773 336309 47891 336427
rect 47933 336309 48051 336427
rect 47773 318469 47891 318587
rect 47933 318469 48051 318587
rect 47773 318309 47891 318427
rect 47933 318309 48051 318427
rect 47773 300469 47891 300587
rect 47933 300469 48051 300587
rect 47773 300309 47891 300427
rect 47933 300309 48051 300427
rect 47773 282469 47891 282587
rect 47933 282469 48051 282587
rect 47773 282309 47891 282427
rect 47933 282309 48051 282427
rect 47773 264469 47891 264587
rect 47933 264469 48051 264587
rect 47773 264309 47891 264427
rect 47933 264309 48051 264427
rect 47773 246469 47891 246587
rect 47933 246469 48051 246587
rect 47773 246309 47891 246427
rect 47933 246309 48051 246427
rect 47773 228469 47891 228587
rect 47933 228469 48051 228587
rect 47773 228309 47891 228427
rect 47933 228309 48051 228427
rect 47773 210469 47891 210587
rect 47933 210469 48051 210587
rect 47773 210309 47891 210427
rect 47933 210309 48051 210427
rect 47773 192469 47891 192587
rect 47933 192469 48051 192587
rect 47773 192309 47891 192427
rect 47933 192309 48051 192427
rect 47773 174469 47891 174587
rect 47933 174469 48051 174587
rect 47773 174309 47891 174427
rect 47933 174309 48051 174427
rect 47773 156469 47891 156587
rect 47933 156469 48051 156587
rect 47773 156309 47891 156427
rect 47933 156309 48051 156427
rect 47773 138469 47891 138587
rect 47933 138469 48051 138587
rect 47773 138309 47891 138427
rect 47933 138309 48051 138427
rect 47773 120469 47891 120587
rect 47933 120469 48051 120587
rect 47773 120309 47891 120427
rect 47933 120309 48051 120427
rect 47773 102469 47891 102587
rect 47933 102469 48051 102587
rect 47773 102309 47891 102427
rect 47933 102309 48051 102427
rect 47773 84469 47891 84587
rect 47933 84469 48051 84587
rect 47773 84309 47891 84427
rect 47933 84309 48051 84427
rect 47773 66469 47891 66587
rect 47933 66469 48051 66587
rect 47773 66309 47891 66427
rect 47933 66309 48051 66427
rect 47773 48469 47891 48587
rect 47933 48469 48051 48587
rect 47773 48309 47891 48427
rect 47933 48309 48051 48427
rect 47773 30469 47891 30587
rect 47933 30469 48051 30587
rect 47773 30309 47891 30427
rect 47933 30309 48051 30427
rect 47773 12469 47891 12587
rect 47933 12469 48051 12587
rect 47773 12309 47891 12427
rect 47933 12309 48051 12427
rect 47773 -1731 47891 -1613
rect 47933 -1731 48051 -1613
rect 47773 -1891 47891 -1773
rect 47933 -1891 48051 -1773
rect 49633 338329 49751 338447
rect 49793 338329 49911 338447
rect 49633 338169 49751 338287
rect 49793 338169 49911 338287
rect 49633 320329 49751 320447
rect 49793 320329 49911 320447
rect 49633 320169 49751 320287
rect 49793 320169 49911 320287
rect 49633 302329 49751 302447
rect 49793 302329 49911 302447
rect 49633 302169 49751 302287
rect 49793 302169 49911 302287
rect 49633 284329 49751 284447
rect 49793 284329 49911 284447
rect 49633 284169 49751 284287
rect 49793 284169 49911 284287
rect 49633 266329 49751 266447
rect 49793 266329 49911 266447
rect 49633 266169 49751 266287
rect 49793 266169 49911 266287
rect 49633 248329 49751 248447
rect 49793 248329 49911 248447
rect 49633 248169 49751 248287
rect 49793 248169 49911 248287
rect 49633 230329 49751 230447
rect 49793 230329 49911 230447
rect 49633 230169 49751 230287
rect 49793 230169 49911 230287
rect 49633 212329 49751 212447
rect 49793 212329 49911 212447
rect 49633 212169 49751 212287
rect 49793 212169 49911 212287
rect 49633 194329 49751 194447
rect 49793 194329 49911 194447
rect 49633 194169 49751 194287
rect 49793 194169 49911 194287
rect 49633 176329 49751 176447
rect 49793 176329 49911 176447
rect 49633 176169 49751 176287
rect 49793 176169 49911 176287
rect 49633 158329 49751 158447
rect 49793 158329 49911 158447
rect 49633 158169 49751 158287
rect 49793 158169 49911 158287
rect 49633 140329 49751 140447
rect 49793 140329 49911 140447
rect 49633 140169 49751 140287
rect 49793 140169 49911 140287
rect 49633 122329 49751 122447
rect 49793 122329 49911 122447
rect 49633 122169 49751 122287
rect 49793 122169 49911 122287
rect 49633 104329 49751 104447
rect 49793 104329 49911 104447
rect 49633 104169 49751 104287
rect 49793 104169 49911 104287
rect 49633 86329 49751 86447
rect 49793 86329 49911 86447
rect 49633 86169 49751 86287
rect 49793 86169 49911 86287
rect 49633 68329 49751 68447
rect 49793 68329 49911 68447
rect 49633 68169 49751 68287
rect 49793 68169 49911 68287
rect 49633 50329 49751 50447
rect 49793 50329 49911 50447
rect 49633 50169 49751 50287
rect 49793 50169 49911 50287
rect 49633 32329 49751 32447
rect 49793 32329 49911 32447
rect 49633 32169 49751 32287
rect 49793 32169 49911 32287
rect 49633 14329 49751 14447
rect 49793 14329 49911 14447
rect 49633 14169 49751 14287
rect 49793 14169 49911 14287
rect 49633 -2691 49751 -2573
rect 49793 -2691 49911 -2573
rect 49633 -2851 49751 -2733
rect 49793 -2851 49911 -2733
rect 60493 355181 60611 355299
rect 60653 355181 60771 355299
rect 60493 355021 60611 355139
rect 60653 355021 60771 355139
rect 58633 354221 58751 354339
rect 58793 354221 58911 354339
rect 58633 354061 58751 354179
rect 58793 354061 58911 354179
rect 56773 353261 56891 353379
rect 56933 353261 57051 353379
rect 56773 353101 56891 353219
rect 56933 353101 57051 353219
rect 51493 340189 51611 340307
rect 51653 340189 51771 340307
rect 51493 340029 51611 340147
rect 51653 340029 51771 340147
rect 51493 322189 51611 322307
rect 51653 322189 51771 322307
rect 51493 322029 51611 322147
rect 51653 322029 51771 322147
rect 51493 304189 51611 304307
rect 51653 304189 51771 304307
rect 51493 304029 51611 304147
rect 51653 304029 51771 304147
rect 51493 286189 51611 286307
rect 51653 286189 51771 286307
rect 51493 286029 51611 286147
rect 51653 286029 51771 286147
rect 51493 268189 51611 268307
rect 51653 268189 51771 268307
rect 51493 268029 51611 268147
rect 51653 268029 51771 268147
rect 51493 250189 51611 250307
rect 51653 250189 51771 250307
rect 51493 250029 51611 250147
rect 51653 250029 51771 250147
rect 51493 232189 51611 232307
rect 51653 232189 51771 232307
rect 51493 232029 51611 232147
rect 51653 232029 51771 232147
rect 51493 214189 51611 214307
rect 51653 214189 51771 214307
rect 51493 214029 51611 214147
rect 51653 214029 51771 214147
rect 51493 196189 51611 196307
rect 51653 196189 51771 196307
rect 51493 196029 51611 196147
rect 51653 196029 51771 196147
rect 51493 178189 51611 178307
rect 51653 178189 51771 178307
rect 51493 178029 51611 178147
rect 51653 178029 51771 178147
rect 51493 160189 51611 160307
rect 51653 160189 51771 160307
rect 51493 160029 51611 160147
rect 51653 160029 51771 160147
rect 51493 142189 51611 142307
rect 51653 142189 51771 142307
rect 51493 142029 51611 142147
rect 51653 142029 51771 142147
rect 51493 124189 51611 124307
rect 51653 124189 51771 124307
rect 51493 124029 51611 124147
rect 51653 124029 51771 124147
rect 51493 106189 51611 106307
rect 51653 106189 51771 106307
rect 51493 106029 51611 106147
rect 51653 106029 51771 106147
rect 51493 88189 51611 88307
rect 51653 88189 51771 88307
rect 51493 88029 51611 88147
rect 51653 88029 51771 88147
rect 51493 70189 51611 70307
rect 51653 70189 51771 70307
rect 51493 70029 51611 70147
rect 51653 70029 51771 70147
rect 51493 52189 51611 52307
rect 51653 52189 51771 52307
rect 51493 52029 51611 52147
rect 51653 52029 51771 52147
rect 51493 34189 51611 34307
rect 51653 34189 51771 34307
rect 51493 34029 51611 34147
rect 51653 34029 51771 34147
rect 51493 16189 51611 16307
rect 51653 16189 51771 16307
rect 51493 16029 51611 16147
rect 51653 16029 51771 16147
rect 42493 -3171 42611 -3053
rect 42653 -3171 42771 -3053
rect 42493 -3331 42611 -3213
rect 42653 -3331 42771 -3213
rect 54913 352301 55031 352419
rect 55073 352301 55191 352419
rect 54913 352141 55031 352259
rect 55073 352141 55191 352259
rect 54913 343609 55031 343727
rect 55073 343609 55191 343727
rect 54913 343449 55031 343567
rect 55073 343449 55191 343567
rect 54913 325609 55031 325727
rect 55073 325609 55191 325727
rect 54913 325449 55031 325567
rect 55073 325449 55191 325567
rect 54913 307609 55031 307727
rect 55073 307609 55191 307727
rect 54913 307449 55031 307567
rect 55073 307449 55191 307567
rect 54913 289609 55031 289727
rect 55073 289609 55191 289727
rect 54913 289449 55031 289567
rect 55073 289449 55191 289567
rect 54913 271609 55031 271727
rect 55073 271609 55191 271727
rect 54913 271449 55031 271567
rect 55073 271449 55191 271567
rect 54913 253609 55031 253727
rect 55073 253609 55191 253727
rect 54913 253449 55031 253567
rect 55073 253449 55191 253567
rect 54913 235609 55031 235727
rect 55073 235609 55191 235727
rect 54913 235449 55031 235567
rect 55073 235449 55191 235567
rect 54913 217609 55031 217727
rect 55073 217609 55191 217727
rect 54913 217449 55031 217567
rect 55073 217449 55191 217567
rect 54913 199609 55031 199727
rect 55073 199609 55191 199727
rect 54913 199449 55031 199567
rect 55073 199449 55191 199567
rect 54913 181609 55031 181727
rect 55073 181609 55191 181727
rect 54913 181449 55031 181567
rect 55073 181449 55191 181567
rect 54913 163609 55031 163727
rect 55073 163609 55191 163727
rect 54913 163449 55031 163567
rect 55073 163449 55191 163567
rect 54913 145609 55031 145727
rect 55073 145609 55191 145727
rect 54913 145449 55031 145567
rect 55073 145449 55191 145567
rect 54913 127609 55031 127727
rect 55073 127609 55191 127727
rect 54913 127449 55031 127567
rect 55073 127449 55191 127567
rect 54913 109609 55031 109727
rect 55073 109609 55191 109727
rect 54913 109449 55031 109567
rect 55073 109449 55191 109567
rect 54913 91609 55031 91727
rect 55073 91609 55191 91727
rect 54913 91449 55031 91567
rect 55073 91449 55191 91567
rect 54913 73609 55031 73727
rect 55073 73609 55191 73727
rect 54913 73449 55031 73567
rect 55073 73449 55191 73567
rect 54913 55609 55031 55727
rect 55073 55609 55191 55727
rect 54913 55449 55031 55567
rect 55073 55449 55191 55567
rect 54913 37609 55031 37727
rect 55073 37609 55191 37727
rect 54913 37449 55031 37567
rect 55073 37449 55191 37567
rect 54913 19609 55031 19727
rect 55073 19609 55191 19727
rect 54913 19449 55031 19567
rect 55073 19449 55191 19567
rect 54913 1609 55031 1727
rect 55073 1609 55191 1727
rect 54913 1449 55031 1567
rect 55073 1449 55191 1567
rect 54913 -291 55031 -173
rect 55073 -291 55191 -173
rect 54913 -451 55031 -333
rect 55073 -451 55191 -333
rect 56773 345469 56891 345587
rect 56933 345469 57051 345587
rect 56773 345309 56891 345427
rect 56933 345309 57051 345427
rect 56773 327469 56891 327587
rect 56933 327469 57051 327587
rect 56773 327309 56891 327427
rect 56933 327309 57051 327427
rect 56773 309469 56891 309587
rect 56933 309469 57051 309587
rect 56773 309309 56891 309427
rect 56933 309309 57051 309427
rect 56773 291469 56891 291587
rect 56933 291469 57051 291587
rect 56773 291309 56891 291427
rect 56933 291309 57051 291427
rect 56773 273469 56891 273587
rect 56933 273469 57051 273587
rect 56773 273309 56891 273427
rect 56933 273309 57051 273427
rect 56773 255469 56891 255587
rect 56933 255469 57051 255587
rect 56773 255309 56891 255427
rect 56933 255309 57051 255427
rect 56773 237469 56891 237587
rect 56933 237469 57051 237587
rect 56773 237309 56891 237427
rect 56933 237309 57051 237427
rect 56773 219469 56891 219587
rect 56933 219469 57051 219587
rect 56773 219309 56891 219427
rect 56933 219309 57051 219427
rect 56773 201469 56891 201587
rect 56933 201469 57051 201587
rect 56773 201309 56891 201427
rect 56933 201309 57051 201427
rect 56773 183469 56891 183587
rect 56933 183469 57051 183587
rect 56773 183309 56891 183427
rect 56933 183309 57051 183427
rect 56773 165469 56891 165587
rect 56933 165469 57051 165587
rect 56773 165309 56891 165427
rect 56933 165309 57051 165427
rect 56773 147469 56891 147587
rect 56933 147469 57051 147587
rect 56773 147309 56891 147427
rect 56933 147309 57051 147427
rect 56773 129469 56891 129587
rect 56933 129469 57051 129587
rect 56773 129309 56891 129427
rect 56933 129309 57051 129427
rect 56773 111469 56891 111587
rect 56933 111469 57051 111587
rect 56773 111309 56891 111427
rect 56933 111309 57051 111427
rect 56773 93469 56891 93587
rect 56933 93469 57051 93587
rect 56773 93309 56891 93427
rect 56933 93309 57051 93427
rect 56773 75469 56891 75587
rect 56933 75469 57051 75587
rect 56773 75309 56891 75427
rect 56933 75309 57051 75427
rect 56773 57469 56891 57587
rect 56933 57469 57051 57587
rect 56773 57309 56891 57427
rect 56933 57309 57051 57427
rect 56773 39469 56891 39587
rect 56933 39469 57051 39587
rect 56773 39309 56891 39427
rect 56933 39309 57051 39427
rect 56773 21469 56891 21587
rect 56933 21469 57051 21587
rect 56773 21309 56891 21427
rect 56933 21309 57051 21427
rect 56773 3469 56891 3587
rect 56933 3469 57051 3587
rect 56773 3309 56891 3427
rect 56933 3309 57051 3427
rect 56773 -1251 56891 -1133
rect 56933 -1251 57051 -1133
rect 56773 -1411 56891 -1293
rect 56933 -1411 57051 -1293
rect 58633 347329 58751 347447
rect 58793 347329 58911 347447
rect 58633 347169 58751 347287
rect 58793 347169 58911 347287
rect 58633 329329 58751 329447
rect 58793 329329 58911 329447
rect 58633 329169 58751 329287
rect 58793 329169 58911 329287
rect 58633 311329 58751 311447
rect 58793 311329 58911 311447
rect 58633 311169 58751 311287
rect 58793 311169 58911 311287
rect 58633 293329 58751 293447
rect 58793 293329 58911 293447
rect 58633 293169 58751 293287
rect 58793 293169 58911 293287
rect 58633 275329 58751 275447
rect 58793 275329 58911 275447
rect 58633 275169 58751 275287
rect 58793 275169 58911 275287
rect 58633 257329 58751 257447
rect 58793 257329 58911 257447
rect 58633 257169 58751 257287
rect 58793 257169 58911 257287
rect 58633 239329 58751 239447
rect 58793 239329 58911 239447
rect 58633 239169 58751 239287
rect 58793 239169 58911 239287
rect 58633 221329 58751 221447
rect 58793 221329 58911 221447
rect 58633 221169 58751 221287
rect 58793 221169 58911 221287
rect 58633 203329 58751 203447
rect 58793 203329 58911 203447
rect 58633 203169 58751 203287
rect 58793 203169 58911 203287
rect 58633 185329 58751 185447
rect 58793 185329 58911 185447
rect 58633 185169 58751 185287
rect 58793 185169 58911 185287
rect 58633 167329 58751 167447
rect 58793 167329 58911 167447
rect 58633 167169 58751 167287
rect 58793 167169 58911 167287
rect 58633 149329 58751 149447
rect 58793 149329 58911 149447
rect 58633 149169 58751 149287
rect 58793 149169 58911 149287
rect 58633 131329 58751 131447
rect 58793 131329 58911 131447
rect 58633 131169 58751 131287
rect 58793 131169 58911 131287
rect 58633 113329 58751 113447
rect 58793 113329 58911 113447
rect 58633 113169 58751 113287
rect 58793 113169 58911 113287
rect 58633 95329 58751 95447
rect 58793 95329 58911 95447
rect 58633 95169 58751 95287
rect 58793 95169 58911 95287
rect 58633 77329 58751 77447
rect 58793 77329 58911 77447
rect 58633 77169 58751 77287
rect 58793 77169 58911 77287
rect 58633 59329 58751 59447
rect 58793 59329 58911 59447
rect 58633 59169 58751 59287
rect 58793 59169 58911 59287
rect 58633 41329 58751 41447
rect 58793 41329 58911 41447
rect 58633 41169 58751 41287
rect 58793 41169 58911 41287
rect 58633 23329 58751 23447
rect 58793 23329 58911 23447
rect 58633 23169 58751 23287
rect 58793 23169 58911 23287
rect 58633 5329 58751 5447
rect 58793 5329 58911 5447
rect 58633 5169 58751 5287
rect 58793 5169 58911 5287
rect 58633 -2211 58751 -2093
rect 58793 -2211 58911 -2093
rect 58633 -2371 58751 -2253
rect 58793 -2371 58911 -2253
rect 69493 355661 69611 355779
rect 69653 355661 69771 355779
rect 69493 355501 69611 355619
rect 69653 355501 69771 355619
rect 67633 354701 67751 354819
rect 67793 354701 67911 354819
rect 67633 354541 67751 354659
rect 67793 354541 67911 354659
rect 65773 353741 65891 353859
rect 65933 353741 66051 353859
rect 65773 353581 65891 353699
rect 65933 353581 66051 353699
rect 60493 349189 60611 349307
rect 60653 349189 60771 349307
rect 60493 349029 60611 349147
rect 60653 349029 60771 349147
rect 60493 331189 60611 331307
rect 60653 331189 60771 331307
rect 60493 331029 60611 331147
rect 60653 331029 60771 331147
rect 60493 313189 60611 313307
rect 60653 313189 60771 313307
rect 60493 313029 60611 313147
rect 60653 313029 60771 313147
rect 60493 295189 60611 295307
rect 60653 295189 60771 295307
rect 60493 295029 60611 295147
rect 60653 295029 60771 295147
rect 60493 277189 60611 277307
rect 60653 277189 60771 277307
rect 60493 277029 60611 277147
rect 60653 277029 60771 277147
rect 60493 259189 60611 259307
rect 60653 259189 60771 259307
rect 60493 259029 60611 259147
rect 60653 259029 60771 259147
rect 60493 241189 60611 241307
rect 60653 241189 60771 241307
rect 60493 241029 60611 241147
rect 60653 241029 60771 241147
rect 60493 223189 60611 223307
rect 60653 223189 60771 223307
rect 60493 223029 60611 223147
rect 60653 223029 60771 223147
rect 60493 205189 60611 205307
rect 60653 205189 60771 205307
rect 60493 205029 60611 205147
rect 60653 205029 60771 205147
rect 60493 187189 60611 187307
rect 60653 187189 60771 187307
rect 60493 187029 60611 187147
rect 60653 187029 60771 187147
rect 60493 169189 60611 169307
rect 60653 169189 60771 169307
rect 60493 169029 60611 169147
rect 60653 169029 60771 169147
rect 60493 151189 60611 151307
rect 60653 151189 60771 151307
rect 60493 151029 60611 151147
rect 60653 151029 60771 151147
rect 60493 133189 60611 133307
rect 60653 133189 60771 133307
rect 60493 133029 60611 133147
rect 60653 133029 60771 133147
rect 60493 115189 60611 115307
rect 60653 115189 60771 115307
rect 60493 115029 60611 115147
rect 60653 115029 60771 115147
rect 60493 97189 60611 97307
rect 60653 97189 60771 97307
rect 60493 97029 60611 97147
rect 60653 97029 60771 97147
rect 60493 79189 60611 79307
rect 60653 79189 60771 79307
rect 60493 79029 60611 79147
rect 60653 79029 60771 79147
rect 60493 61189 60611 61307
rect 60653 61189 60771 61307
rect 60493 61029 60611 61147
rect 60653 61029 60771 61147
rect 60493 43189 60611 43307
rect 60653 43189 60771 43307
rect 60493 43029 60611 43147
rect 60653 43029 60771 43147
rect 60493 25189 60611 25307
rect 60653 25189 60771 25307
rect 60493 25029 60611 25147
rect 60653 25029 60771 25147
rect 60493 7189 60611 7307
rect 60653 7189 60771 7307
rect 60493 7029 60611 7147
rect 60653 7029 60771 7147
rect 51493 -3651 51611 -3533
rect 51653 -3651 51771 -3533
rect 51493 -3811 51611 -3693
rect 51653 -3811 51771 -3693
rect 63913 352781 64031 352899
rect 64073 352781 64191 352899
rect 63913 352621 64031 352739
rect 64073 352621 64191 352739
rect 63913 334609 64031 334727
rect 64073 334609 64191 334727
rect 63913 334449 64031 334567
rect 64073 334449 64191 334567
rect 63913 316609 64031 316727
rect 64073 316609 64191 316727
rect 63913 316449 64031 316567
rect 64073 316449 64191 316567
rect 63913 298609 64031 298727
rect 64073 298609 64191 298727
rect 63913 298449 64031 298567
rect 64073 298449 64191 298567
rect 63913 280609 64031 280727
rect 64073 280609 64191 280727
rect 63913 280449 64031 280567
rect 64073 280449 64191 280567
rect 63913 262609 64031 262727
rect 64073 262609 64191 262727
rect 63913 262449 64031 262567
rect 64073 262449 64191 262567
rect 63913 244609 64031 244727
rect 64073 244609 64191 244727
rect 63913 244449 64031 244567
rect 64073 244449 64191 244567
rect 63913 226609 64031 226727
rect 64073 226609 64191 226727
rect 63913 226449 64031 226567
rect 64073 226449 64191 226567
rect 63913 208609 64031 208727
rect 64073 208609 64191 208727
rect 63913 208449 64031 208567
rect 64073 208449 64191 208567
rect 63913 190609 64031 190727
rect 64073 190609 64191 190727
rect 63913 190449 64031 190567
rect 64073 190449 64191 190567
rect 63913 172609 64031 172727
rect 64073 172609 64191 172727
rect 63913 172449 64031 172567
rect 64073 172449 64191 172567
rect 63913 154609 64031 154727
rect 64073 154609 64191 154727
rect 63913 154449 64031 154567
rect 64073 154449 64191 154567
rect 63913 136609 64031 136727
rect 64073 136609 64191 136727
rect 63913 136449 64031 136567
rect 64073 136449 64191 136567
rect 63913 118609 64031 118727
rect 64073 118609 64191 118727
rect 63913 118449 64031 118567
rect 64073 118449 64191 118567
rect 63913 100609 64031 100727
rect 64073 100609 64191 100727
rect 63913 100449 64031 100567
rect 64073 100449 64191 100567
rect 63913 82609 64031 82727
rect 64073 82609 64191 82727
rect 63913 82449 64031 82567
rect 64073 82449 64191 82567
rect 63913 64609 64031 64727
rect 64073 64609 64191 64727
rect 63913 64449 64031 64567
rect 64073 64449 64191 64567
rect 63913 46609 64031 46727
rect 64073 46609 64191 46727
rect 63913 46449 64031 46567
rect 64073 46449 64191 46567
rect 63913 28609 64031 28727
rect 64073 28609 64191 28727
rect 63913 28449 64031 28567
rect 64073 28449 64191 28567
rect 63913 10609 64031 10727
rect 64073 10609 64191 10727
rect 63913 10449 64031 10567
rect 64073 10449 64191 10567
rect 63913 -771 64031 -653
rect 64073 -771 64191 -653
rect 63913 -931 64031 -813
rect 64073 -931 64191 -813
rect 65773 336469 65891 336587
rect 65933 336469 66051 336587
rect 65773 336309 65891 336427
rect 65933 336309 66051 336427
rect 65773 318469 65891 318587
rect 65933 318469 66051 318587
rect 65773 318309 65891 318427
rect 65933 318309 66051 318427
rect 65773 300469 65891 300587
rect 65933 300469 66051 300587
rect 65773 300309 65891 300427
rect 65933 300309 66051 300427
rect 65773 282469 65891 282587
rect 65933 282469 66051 282587
rect 65773 282309 65891 282427
rect 65933 282309 66051 282427
rect 65773 264469 65891 264587
rect 65933 264469 66051 264587
rect 65773 264309 65891 264427
rect 65933 264309 66051 264427
rect 65773 246469 65891 246587
rect 65933 246469 66051 246587
rect 65773 246309 65891 246427
rect 65933 246309 66051 246427
rect 65773 228469 65891 228587
rect 65933 228469 66051 228587
rect 65773 228309 65891 228427
rect 65933 228309 66051 228427
rect 65773 210469 65891 210587
rect 65933 210469 66051 210587
rect 65773 210309 65891 210427
rect 65933 210309 66051 210427
rect 65773 192469 65891 192587
rect 65933 192469 66051 192587
rect 65773 192309 65891 192427
rect 65933 192309 66051 192427
rect 65773 174469 65891 174587
rect 65933 174469 66051 174587
rect 65773 174309 65891 174427
rect 65933 174309 66051 174427
rect 65773 156469 65891 156587
rect 65933 156469 66051 156587
rect 65773 156309 65891 156427
rect 65933 156309 66051 156427
rect 65773 138469 65891 138587
rect 65933 138469 66051 138587
rect 65773 138309 65891 138427
rect 65933 138309 66051 138427
rect 65773 120469 65891 120587
rect 65933 120469 66051 120587
rect 65773 120309 65891 120427
rect 65933 120309 66051 120427
rect 65773 102469 65891 102587
rect 65933 102469 66051 102587
rect 65773 102309 65891 102427
rect 65933 102309 66051 102427
rect 65773 84469 65891 84587
rect 65933 84469 66051 84587
rect 65773 84309 65891 84427
rect 65933 84309 66051 84427
rect 65773 66469 65891 66587
rect 65933 66469 66051 66587
rect 65773 66309 65891 66427
rect 65933 66309 66051 66427
rect 65773 48469 65891 48587
rect 65933 48469 66051 48587
rect 65773 48309 65891 48427
rect 65933 48309 66051 48427
rect 65773 30469 65891 30587
rect 65933 30469 66051 30587
rect 65773 30309 65891 30427
rect 65933 30309 66051 30427
rect 65773 12469 65891 12587
rect 65933 12469 66051 12587
rect 65773 12309 65891 12427
rect 65933 12309 66051 12427
rect 65773 -1731 65891 -1613
rect 65933 -1731 66051 -1613
rect 65773 -1891 65891 -1773
rect 65933 -1891 66051 -1773
rect 67633 338329 67751 338447
rect 67793 338329 67911 338447
rect 67633 338169 67751 338287
rect 67793 338169 67911 338287
rect 67633 320329 67751 320447
rect 67793 320329 67911 320447
rect 67633 320169 67751 320287
rect 67793 320169 67911 320287
rect 67633 302329 67751 302447
rect 67793 302329 67911 302447
rect 67633 302169 67751 302287
rect 67793 302169 67911 302287
rect 67633 284329 67751 284447
rect 67793 284329 67911 284447
rect 67633 284169 67751 284287
rect 67793 284169 67911 284287
rect 67633 266329 67751 266447
rect 67793 266329 67911 266447
rect 67633 266169 67751 266287
rect 67793 266169 67911 266287
rect 67633 248329 67751 248447
rect 67793 248329 67911 248447
rect 67633 248169 67751 248287
rect 67793 248169 67911 248287
rect 67633 230329 67751 230447
rect 67793 230329 67911 230447
rect 67633 230169 67751 230287
rect 67793 230169 67911 230287
rect 67633 212329 67751 212447
rect 67793 212329 67911 212447
rect 67633 212169 67751 212287
rect 67793 212169 67911 212287
rect 67633 194329 67751 194447
rect 67793 194329 67911 194447
rect 67633 194169 67751 194287
rect 67793 194169 67911 194287
rect 67633 176329 67751 176447
rect 67793 176329 67911 176447
rect 67633 176169 67751 176287
rect 67793 176169 67911 176287
rect 67633 158329 67751 158447
rect 67793 158329 67911 158447
rect 67633 158169 67751 158287
rect 67793 158169 67911 158287
rect 67633 140329 67751 140447
rect 67793 140329 67911 140447
rect 67633 140169 67751 140287
rect 67793 140169 67911 140287
rect 67633 122329 67751 122447
rect 67793 122329 67911 122447
rect 67633 122169 67751 122287
rect 67793 122169 67911 122287
rect 67633 104329 67751 104447
rect 67793 104329 67911 104447
rect 67633 104169 67751 104287
rect 67793 104169 67911 104287
rect 67633 86329 67751 86447
rect 67793 86329 67911 86447
rect 67633 86169 67751 86287
rect 67793 86169 67911 86287
rect 67633 68329 67751 68447
rect 67793 68329 67911 68447
rect 67633 68169 67751 68287
rect 67793 68169 67911 68287
rect 67633 50329 67751 50447
rect 67793 50329 67911 50447
rect 67633 50169 67751 50287
rect 67793 50169 67911 50287
rect 67633 32329 67751 32447
rect 67793 32329 67911 32447
rect 67633 32169 67751 32287
rect 67793 32169 67911 32287
rect 67633 14329 67751 14447
rect 67793 14329 67911 14447
rect 67633 14169 67751 14287
rect 67793 14169 67911 14287
rect 67633 -2691 67751 -2573
rect 67793 -2691 67911 -2573
rect 67633 -2851 67751 -2733
rect 67793 -2851 67911 -2733
rect 78493 355181 78611 355299
rect 78653 355181 78771 355299
rect 78493 355021 78611 355139
rect 78653 355021 78771 355139
rect 76633 354221 76751 354339
rect 76793 354221 76911 354339
rect 76633 354061 76751 354179
rect 76793 354061 76911 354179
rect 74773 353261 74891 353379
rect 74933 353261 75051 353379
rect 74773 353101 74891 353219
rect 74933 353101 75051 353219
rect 69493 340189 69611 340307
rect 69653 340189 69771 340307
rect 69493 340029 69611 340147
rect 69653 340029 69771 340147
rect 69493 322189 69611 322307
rect 69653 322189 69771 322307
rect 69493 322029 69611 322147
rect 69653 322029 69771 322147
rect 69493 304189 69611 304307
rect 69653 304189 69771 304307
rect 69493 304029 69611 304147
rect 69653 304029 69771 304147
rect 69493 286189 69611 286307
rect 69653 286189 69771 286307
rect 69493 286029 69611 286147
rect 69653 286029 69771 286147
rect 69493 268189 69611 268307
rect 69653 268189 69771 268307
rect 69493 268029 69611 268147
rect 69653 268029 69771 268147
rect 69493 250189 69611 250307
rect 69653 250189 69771 250307
rect 69493 250029 69611 250147
rect 69653 250029 69771 250147
rect 69493 232189 69611 232307
rect 69653 232189 69771 232307
rect 69493 232029 69611 232147
rect 69653 232029 69771 232147
rect 69493 214189 69611 214307
rect 69653 214189 69771 214307
rect 69493 214029 69611 214147
rect 69653 214029 69771 214147
rect 69493 196189 69611 196307
rect 69653 196189 69771 196307
rect 69493 196029 69611 196147
rect 69653 196029 69771 196147
rect 69493 178189 69611 178307
rect 69653 178189 69771 178307
rect 69493 178029 69611 178147
rect 69653 178029 69771 178147
rect 69493 160189 69611 160307
rect 69653 160189 69771 160307
rect 69493 160029 69611 160147
rect 69653 160029 69771 160147
rect 69493 142189 69611 142307
rect 69653 142189 69771 142307
rect 69493 142029 69611 142147
rect 69653 142029 69771 142147
rect 69493 124189 69611 124307
rect 69653 124189 69771 124307
rect 69493 124029 69611 124147
rect 69653 124029 69771 124147
rect 69493 106189 69611 106307
rect 69653 106189 69771 106307
rect 69493 106029 69611 106147
rect 69653 106029 69771 106147
rect 69493 88189 69611 88307
rect 69653 88189 69771 88307
rect 69493 88029 69611 88147
rect 69653 88029 69771 88147
rect 69493 70189 69611 70307
rect 69653 70189 69771 70307
rect 69493 70029 69611 70147
rect 69653 70029 69771 70147
rect 69493 52189 69611 52307
rect 69653 52189 69771 52307
rect 69493 52029 69611 52147
rect 69653 52029 69771 52147
rect 69493 34189 69611 34307
rect 69653 34189 69771 34307
rect 69493 34029 69611 34147
rect 69653 34029 69771 34147
rect 69493 16189 69611 16307
rect 69653 16189 69771 16307
rect 69493 16029 69611 16147
rect 69653 16029 69771 16147
rect 60493 -3171 60611 -3053
rect 60653 -3171 60771 -3053
rect 60493 -3331 60611 -3213
rect 60653 -3331 60771 -3213
rect 72913 352301 73031 352419
rect 73073 352301 73191 352419
rect 72913 352141 73031 352259
rect 73073 352141 73191 352259
rect 72913 343609 73031 343727
rect 73073 343609 73191 343727
rect 72913 343449 73031 343567
rect 73073 343449 73191 343567
rect 72913 325609 73031 325727
rect 73073 325609 73191 325727
rect 72913 325449 73031 325567
rect 73073 325449 73191 325567
rect 72913 307609 73031 307727
rect 73073 307609 73191 307727
rect 72913 307449 73031 307567
rect 73073 307449 73191 307567
rect 72913 289609 73031 289727
rect 73073 289609 73191 289727
rect 72913 289449 73031 289567
rect 73073 289449 73191 289567
rect 72913 271609 73031 271727
rect 73073 271609 73191 271727
rect 72913 271449 73031 271567
rect 73073 271449 73191 271567
rect 72913 253609 73031 253727
rect 73073 253609 73191 253727
rect 72913 253449 73031 253567
rect 73073 253449 73191 253567
rect 72913 235609 73031 235727
rect 73073 235609 73191 235727
rect 72913 235449 73031 235567
rect 73073 235449 73191 235567
rect 72913 217609 73031 217727
rect 73073 217609 73191 217727
rect 72913 217449 73031 217567
rect 73073 217449 73191 217567
rect 72913 199609 73031 199727
rect 73073 199609 73191 199727
rect 72913 199449 73031 199567
rect 73073 199449 73191 199567
rect 72913 181609 73031 181727
rect 73073 181609 73191 181727
rect 72913 181449 73031 181567
rect 73073 181449 73191 181567
rect 72913 163609 73031 163727
rect 73073 163609 73191 163727
rect 72913 163449 73031 163567
rect 73073 163449 73191 163567
rect 72913 145609 73031 145727
rect 73073 145609 73191 145727
rect 72913 145449 73031 145567
rect 73073 145449 73191 145567
rect 72913 127609 73031 127727
rect 73073 127609 73191 127727
rect 72913 127449 73031 127567
rect 73073 127449 73191 127567
rect 72913 109609 73031 109727
rect 73073 109609 73191 109727
rect 72913 109449 73031 109567
rect 73073 109449 73191 109567
rect 72913 91609 73031 91727
rect 73073 91609 73191 91727
rect 72913 91449 73031 91567
rect 73073 91449 73191 91567
rect 72913 73609 73031 73727
rect 73073 73609 73191 73727
rect 72913 73449 73031 73567
rect 73073 73449 73191 73567
rect 72913 55609 73031 55727
rect 73073 55609 73191 55727
rect 72913 55449 73031 55567
rect 73073 55449 73191 55567
rect 72913 37609 73031 37727
rect 73073 37609 73191 37727
rect 72913 37449 73031 37567
rect 73073 37449 73191 37567
rect 72913 19609 73031 19727
rect 73073 19609 73191 19727
rect 72913 19449 73031 19567
rect 73073 19449 73191 19567
rect 72913 1609 73031 1727
rect 73073 1609 73191 1727
rect 72913 1449 73031 1567
rect 73073 1449 73191 1567
rect 72913 -291 73031 -173
rect 73073 -291 73191 -173
rect 72913 -451 73031 -333
rect 73073 -451 73191 -333
rect 74773 345469 74891 345587
rect 74933 345469 75051 345587
rect 74773 345309 74891 345427
rect 74933 345309 75051 345427
rect 74773 327469 74891 327587
rect 74933 327469 75051 327587
rect 74773 327309 74891 327427
rect 74933 327309 75051 327427
rect 74773 309469 74891 309587
rect 74933 309469 75051 309587
rect 74773 309309 74891 309427
rect 74933 309309 75051 309427
rect 74773 291469 74891 291587
rect 74933 291469 75051 291587
rect 74773 291309 74891 291427
rect 74933 291309 75051 291427
rect 74773 273469 74891 273587
rect 74933 273469 75051 273587
rect 74773 273309 74891 273427
rect 74933 273309 75051 273427
rect 74773 255469 74891 255587
rect 74933 255469 75051 255587
rect 74773 255309 74891 255427
rect 74933 255309 75051 255427
rect 74773 237469 74891 237587
rect 74933 237469 75051 237587
rect 74773 237309 74891 237427
rect 74933 237309 75051 237427
rect 74773 219469 74891 219587
rect 74933 219469 75051 219587
rect 74773 219309 74891 219427
rect 74933 219309 75051 219427
rect 74773 201469 74891 201587
rect 74933 201469 75051 201587
rect 74773 201309 74891 201427
rect 74933 201309 75051 201427
rect 74773 183469 74891 183587
rect 74933 183469 75051 183587
rect 74773 183309 74891 183427
rect 74933 183309 75051 183427
rect 74773 165469 74891 165587
rect 74933 165469 75051 165587
rect 74773 165309 74891 165427
rect 74933 165309 75051 165427
rect 74773 147469 74891 147587
rect 74933 147469 75051 147587
rect 74773 147309 74891 147427
rect 74933 147309 75051 147427
rect 74773 129469 74891 129587
rect 74933 129469 75051 129587
rect 74773 129309 74891 129427
rect 74933 129309 75051 129427
rect 74773 111469 74891 111587
rect 74933 111469 75051 111587
rect 74773 111309 74891 111427
rect 74933 111309 75051 111427
rect 74773 93469 74891 93587
rect 74933 93469 75051 93587
rect 74773 93309 74891 93427
rect 74933 93309 75051 93427
rect 74773 75469 74891 75587
rect 74933 75469 75051 75587
rect 74773 75309 74891 75427
rect 74933 75309 75051 75427
rect 74773 57469 74891 57587
rect 74933 57469 75051 57587
rect 74773 57309 74891 57427
rect 74933 57309 75051 57427
rect 74773 39469 74891 39587
rect 74933 39469 75051 39587
rect 74773 39309 74891 39427
rect 74933 39309 75051 39427
rect 74773 21469 74891 21587
rect 74933 21469 75051 21587
rect 74773 21309 74891 21427
rect 74933 21309 75051 21427
rect 74773 3469 74891 3587
rect 74933 3469 75051 3587
rect 74773 3309 74891 3427
rect 74933 3309 75051 3427
rect 74773 -1251 74891 -1133
rect 74933 -1251 75051 -1133
rect 74773 -1411 74891 -1293
rect 74933 -1411 75051 -1293
rect 76633 347329 76751 347447
rect 76793 347329 76911 347447
rect 76633 347169 76751 347287
rect 76793 347169 76911 347287
rect 76633 329329 76751 329447
rect 76793 329329 76911 329447
rect 76633 329169 76751 329287
rect 76793 329169 76911 329287
rect 76633 311329 76751 311447
rect 76793 311329 76911 311447
rect 76633 311169 76751 311287
rect 76793 311169 76911 311287
rect 76633 293329 76751 293447
rect 76793 293329 76911 293447
rect 76633 293169 76751 293287
rect 76793 293169 76911 293287
rect 76633 275329 76751 275447
rect 76793 275329 76911 275447
rect 76633 275169 76751 275287
rect 76793 275169 76911 275287
rect 76633 257329 76751 257447
rect 76793 257329 76911 257447
rect 76633 257169 76751 257287
rect 76793 257169 76911 257287
rect 76633 239329 76751 239447
rect 76793 239329 76911 239447
rect 76633 239169 76751 239287
rect 76793 239169 76911 239287
rect 76633 221329 76751 221447
rect 76793 221329 76911 221447
rect 76633 221169 76751 221287
rect 76793 221169 76911 221287
rect 76633 203329 76751 203447
rect 76793 203329 76911 203447
rect 76633 203169 76751 203287
rect 76793 203169 76911 203287
rect 76633 185329 76751 185447
rect 76793 185329 76911 185447
rect 76633 185169 76751 185287
rect 76793 185169 76911 185287
rect 76633 167329 76751 167447
rect 76793 167329 76911 167447
rect 76633 167169 76751 167287
rect 76793 167169 76911 167287
rect 76633 149329 76751 149447
rect 76793 149329 76911 149447
rect 76633 149169 76751 149287
rect 76793 149169 76911 149287
rect 76633 131329 76751 131447
rect 76793 131329 76911 131447
rect 76633 131169 76751 131287
rect 76793 131169 76911 131287
rect 76633 113329 76751 113447
rect 76793 113329 76911 113447
rect 76633 113169 76751 113287
rect 76793 113169 76911 113287
rect 76633 95329 76751 95447
rect 76793 95329 76911 95447
rect 76633 95169 76751 95287
rect 76793 95169 76911 95287
rect 76633 77329 76751 77447
rect 76793 77329 76911 77447
rect 76633 77169 76751 77287
rect 76793 77169 76911 77287
rect 76633 59329 76751 59447
rect 76793 59329 76911 59447
rect 76633 59169 76751 59287
rect 76793 59169 76911 59287
rect 76633 41329 76751 41447
rect 76793 41329 76911 41447
rect 76633 41169 76751 41287
rect 76793 41169 76911 41287
rect 76633 23329 76751 23447
rect 76793 23329 76911 23447
rect 76633 23169 76751 23287
rect 76793 23169 76911 23287
rect 76633 5329 76751 5447
rect 76793 5329 76911 5447
rect 76633 5169 76751 5287
rect 76793 5169 76911 5287
rect 76633 -2211 76751 -2093
rect 76793 -2211 76911 -2093
rect 76633 -2371 76751 -2253
rect 76793 -2371 76911 -2253
rect 87493 355661 87611 355779
rect 87653 355661 87771 355779
rect 87493 355501 87611 355619
rect 87653 355501 87771 355619
rect 85633 354701 85751 354819
rect 85793 354701 85911 354819
rect 85633 354541 85751 354659
rect 85793 354541 85911 354659
rect 83773 353741 83891 353859
rect 83933 353741 84051 353859
rect 83773 353581 83891 353699
rect 83933 353581 84051 353699
rect 78493 349189 78611 349307
rect 78653 349189 78771 349307
rect 78493 349029 78611 349147
rect 78653 349029 78771 349147
rect 78493 331189 78611 331307
rect 78653 331189 78771 331307
rect 78493 331029 78611 331147
rect 78653 331029 78771 331147
rect 78493 313189 78611 313307
rect 78653 313189 78771 313307
rect 78493 313029 78611 313147
rect 78653 313029 78771 313147
rect 78493 295189 78611 295307
rect 78653 295189 78771 295307
rect 78493 295029 78611 295147
rect 78653 295029 78771 295147
rect 78493 277189 78611 277307
rect 78653 277189 78771 277307
rect 78493 277029 78611 277147
rect 78653 277029 78771 277147
rect 78493 259189 78611 259307
rect 78653 259189 78771 259307
rect 78493 259029 78611 259147
rect 78653 259029 78771 259147
rect 78493 241189 78611 241307
rect 78653 241189 78771 241307
rect 78493 241029 78611 241147
rect 78653 241029 78771 241147
rect 78493 223189 78611 223307
rect 78653 223189 78771 223307
rect 78493 223029 78611 223147
rect 78653 223029 78771 223147
rect 78493 205189 78611 205307
rect 78653 205189 78771 205307
rect 78493 205029 78611 205147
rect 78653 205029 78771 205147
rect 78493 187189 78611 187307
rect 78653 187189 78771 187307
rect 78493 187029 78611 187147
rect 78653 187029 78771 187147
rect 78493 169189 78611 169307
rect 78653 169189 78771 169307
rect 78493 169029 78611 169147
rect 78653 169029 78771 169147
rect 78493 151189 78611 151307
rect 78653 151189 78771 151307
rect 78493 151029 78611 151147
rect 78653 151029 78771 151147
rect 78493 133189 78611 133307
rect 78653 133189 78771 133307
rect 78493 133029 78611 133147
rect 78653 133029 78771 133147
rect 78493 115189 78611 115307
rect 78653 115189 78771 115307
rect 78493 115029 78611 115147
rect 78653 115029 78771 115147
rect 78493 97189 78611 97307
rect 78653 97189 78771 97307
rect 78493 97029 78611 97147
rect 78653 97029 78771 97147
rect 78493 79189 78611 79307
rect 78653 79189 78771 79307
rect 78493 79029 78611 79147
rect 78653 79029 78771 79147
rect 78493 61189 78611 61307
rect 78653 61189 78771 61307
rect 78493 61029 78611 61147
rect 78653 61029 78771 61147
rect 78493 43189 78611 43307
rect 78653 43189 78771 43307
rect 78493 43029 78611 43147
rect 78653 43029 78771 43147
rect 78493 25189 78611 25307
rect 78653 25189 78771 25307
rect 78493 25029 78611 25147
rect 78653 25029 78771 25147
rect 78493 7189 78611 7307
rect 78653 7189 78771 7307
rect 78493 7029 78611 7147
rect 78653 7029 78771 7147
rect 69493 -3651 69611 -3533
rect 69653 -3651 69771 -3533
rect 69493 -3811 69611 -3693
rect 69653 -3811 69771 -3693
rect 81913 352781 82031 352899
rect 82073 352781 82191 352899
rect 81913 352621 82031 352739
rect 82073 352621 82191 352739
rect 81913 334609 82031 334727
rect 82073 334609 82191 334727
rect 81913 334449 82031 334567
rect 82073 334449 82191 334567
rect 81913 316609 82031 316727
rect 82073 316609 82191 316727
rect 81913 316449 82031 316567
rect 82073 316449 82191 316567
rect 81913 298609 82031 298727
rect 82073 298609 82191 298727
rect 81913 298449 82031 298567
rect 82073 298449 82191 298567
rect 81913 280609 82031 280727
rect 82073 280609 82191 280727
rect 81913 280449 82031 280567
rect 82073 280449 82191 280567
rect 81913 262609 82031 262727
rect 82073 262609 82191 262727
rect 81913 262449 82031 262567
rect 82073 262449 82191 262567
rect 81913 244609 82031 244727
rect 82073 244609 82191 244727
rect 81913 244449 82031 244567
rect 82073 244449 82191 244567
rect 81913 226609 82031 226727
rect 82073 226609 82191 226727
rect 81913 226449 82031 226567
rect 82073 226449 82191 226567
rect 81913 208609 82031 208727
rect 82073 208609 82191 208727
rect 81913 208449 82031 208567
rect 82073 208449 82191 208567
rect 81913 190609 82031 190727
rect 82073 190609 82191 190727
rect 81913 190449 82031 190567
rect 82073 190449 82191 190567
rect 81913 172609 82031 172727
rect 82073 172609 82191 172727
rect 81913 172449 82031 172567
rect 82073 172449 82191 172567
rect 81913 154609 82031 154727
rect 82073 154609 82191 154727
rect 81913 154449 82031 154567
rect 82073 154449 82191 154567
rect 81913 136609 82031 136727
rect 82073 136609 82191 136727
rect 81913 136449 82031 136567
rect 82073 136449 82191 136567
rect 81913 118609 82031 118727
rect 82073 118609 82191 118727
rect 81913 118449 82031 118567
rect 82073 118449 82191 118567
rect 81913 100609 82031 100727
rect 82073 100609 82191 100727
rect 81913 100449 82031 100567
rect 82073 100449 82191 100567
rect 81913 82609 82031 82727
rect 82073 82609 82191 82727
rect 81913 82449 82031 82567
rect 82073 82449 82191 82567
rect 81913 64609 82031 64727
rect 82073 64609 82191 64727
rect 81913 64449 82031 64567
rect 82073 64449 82191 64567
rect 81913 46609 82031 46727
rect 82073 46609 82191 46727
rect 81913 46449 82031 46567
rect 82073 46449 82191 46567
rect 81913 28609 82031 28727
rect 82073 28609 82191 28727
rect 81913 28449 82031 28567
rect 82073 28449 82191 28567
rect 81913 10609 82031 10727
rect 82073 10609 82191 10727
rect 81913 10449 82031 10567
rect 82073 10449 82191 10567
rect 81913 -771 82031 -653
rect 82073 -771 82191 -653
rect 81913 -931 82031 -813
rect 82073 -931 82191 -813
rect 83773 336469 83891 336587
rect 83933 336469 84051 336587
rect 83773 336309 83891 336427
rect 83933 336309 84051 336427
rect 83773 318469 83891 318587
rect 83933 318469 84051 318587
rect 83773 318309 83891 318427
rect 83933 318309 84051 318427
rect 83773 300469 83891 300587
rect 83933 300469 84051 300587
rect 83773 300309 83891 300427
rect 83933 300309 84051 300427
rect 83773 282469 83891 282587
rect 83933 282469 84051 282587
rect 83773 282309 83891 282427
rect 83933 282309 84051 282427
rect 83773 264469 83891 264587
rect 83933 264469 84051 264587
rect 83773 264309 83891 264427
rect 83933 264309 84051 264427
rect 83773 246469 83891 246587
rect 83933 246469 84051 246587
rect 83773 246309 83891 246427
rect 83933 246309 84051 246427
rect 83773 228469 83891 228587
rect 83933 228469 84051 228587
rect 83773 228309 83891 228427
rect 83933 228309 84051 228427
rect 83773 210469 83891 210587
rect 83933 210469 84051 210587
rect 83773 210309 83891 210427
rect 83933 210309 84051 210427
rect 83773 192469 83891 192587
rect 83933 192469 84051 192587
rect 83773 192309 83891 192427
rect 83933 192309 84051 192427
rect 83773 174469 83891 174587
rect 83933 174469 84051 174587
rect 83773 174309 83891 174427
rect 83933 174309 84051 174427
rect 83773 156469 83891 156587
rect 83933 156469 84051 156587
rect 83773 156309 83891 156427
rect 83933 156309 84051 156427
rect 83773 138469 83891 138587
rect 83933 138469 84051 138587
rect 83773 138309 83891 138427
rect 83933 138309 84051 138427
rect 83773 120469 83891 120587
rect 83933 120469 84051 120587
rect 83773 120309 83891 120427
rect 83933 120309 84051 120427
rect 83773 102469 83891 102587
rect 83933 102469 84051 102587
rect 83773 102309 83891 102427
rect 83933 102309 84051 102427
rect 83773 84469 83891 84587
rect 83933 84469 84051 84587
rect 83773 84309 83891 84427
rect 83933 84309 84051 84427
rect 83773 66469 83891 66587
rect 83933 66469 84051 66587
rect 83773 66309 83891 66427
rect 83933 66309 84051 66427
rect 83773 48469 83891 48587
rect 83933 48469 84051 48587
rect 83773 48309 83891 48427
rect 83933 48309 84051 48427
rect 83773 30469 83891 30587
rect 83933 30469 84051 30587
rect 83773 30309 83891 30427
rect 83933 30309 84051 30427
rect 83773 12469 83891 12587
rect 83933 12469 84051 12587
rect 83773 12309 83891 12427
rect 83933 12309 84051 12427
rect 83773 -1731 83891 -1613
rect 83933 -1731 84051 -1613
rect 83773 -1891 83891 -1773
rect 83933 -1891 84051 -1773
rect 85633 338329 85751 338447
rect 85793 338329 85911 338447
rect 85633 338169 85751 338287
rect 85793 338169 85911 338287
rect 85633 320329 85751 320447
rect 85793 320329 85911 320447
rect 85633 320169 85751 320287
rect 85793 320169 85911 320287
rect 85633 302329 85751 302447
rect 85793 302329 85911 302447
rect 85633 302169 85751 302287
rect 85793 302169 85911 302287
rect 85633 284329 85751 284447
rect 85793 284329 85911 284447
rect 85633 284169 85751 284287
rect 85793 284169 85911 284287
rect 85633 266329 85751 266447
rect 85793 266329 85911 266447
rect 85633 266169 85751 266287
rect 85793 266169 85911 266287
rect 85633 248329 85751 248447
rect 85793 248329 85911 248447
rect 85633 248169 85751 248287
rect 85793 248169 85911 248287
rect 85633 230329 85751 230447
rect 85793 230329 85911 230447
rect 85633 230169 85751 230287
rect 85793 230169 85911 230287
rect 85633 212329 85751 212447
rect 85793 212329 85911 212447
rect 85633 212169 85751 212287
rect 85793 212169 85911 212287
rect 85633 194329 85751 194447
rect 85793 194329 85911 194447
rect 85633 194169 85751 194287
rect 85793 194169 85911 194287
rect 85633 176329 85751 176447
rect 85793 176329 85911 176447
rect 85633 176169 85751 176287
rect 85793 176169 85911 176287
rect 85633 158329 85751 158447
rect 85793 158329 85911 158447
rect 85633 158169 85751 158287
rect 85793 158169 85911 158287
rect 85633 140329 85751 140447
rect 85793 140329 85911 140447
rect 85633 140169 85751 140287
rect 85793 140169 85911 140287
rect 85633 122329 85751 122447
rect 85793 122329 85911 122447
rect 85633 122169 85751 122287
rect 85793 122169 85911 122287
rect 85633 104329 85751 104447
rect 85793 104329 85911 104447
rect 85633 104169 85751 104287
rect 85793 104169 85911 104287
rect 85633 86329 85751 86447
rect 85793 86329 85911 86447
rect 85633 86169 85751 86287
rect 85793 86169 85911 86287
rect 85633 68329 85751 68447
rect 85793 68329 85911 68447
rect 85633 68169 85751 68287
rect 85793 68169 85911 68287
rect 85633 50329 85751 50447
rect 85793 50329 85911 50447
rect 85633 50169 85751 50287
rect 85793 50169 85911 50287
rect 85633 32329 85751 32447
rect 85793 32329 85911 32447
rect 85633 32169 85751 32287
rect 85793 32169 85911 32287
rect 85633 14329 85751 14447
rect 85793 14329 85911 14447
rect 85633 14169 85751 14287
rect 85793 14169 85911 14287
rect 85633 -2691 85751 -2573
rect 85793 -2691 85911 -2573
rect 85633 -2851 85751 -2733
rect 85793 -2851 85911 -2733
rect 96493 355181 96611 355299
rect 96653 355181 96771 355299
rect 96493 355021 96611 355139
rect 96653 355021 96771 355139
rect 94633 354221 94751 354339
rect 94793 354221 94911 354339
rect 94633 354061 94751 354179
rect 94793 354061 94911 354179
rect 92773 353261 92891 353379
rect 92933 353261 93051 353379
rect 92773 353101 92891 353219
rect 92933 353101 93051 353219
rect 87493 340189 87611 340307
rect 87653 340189 87771 340307
rect 87493 340029 87611 340147
rect 87653 340029 87771 340147
rect 87493 322189 87611 322307
rect 87653 322189 87771 322307
rect 87493 322029 87611 322147
rect 87653 322029 87771 322147
rect 87493 304189 87611 304307
rect 87653 304189 87771 304307
rect 87493 304029 87611 304147
rect 87653 304029 87771 304147
rect 87493 286189 87611 286307
rect 87653 286189 87771 286307
rect 87493 286029 87611 286147
rect 87653 286029 87771 286147
rect 87493 268189 87611 268307
rect 87653 268189 87771 268307
rect 87493 268029 87611 268147
rect 87653 268029 87771 268147
rect 87493 250189 87611 250307
rect 87653 250189 87771 250307
rect 87493 250029 87611 250147
rect 87653 250029 87771 250147
rect 87493 232189 87611 232307
rect 87653 232189 87771 232307
rect 87493 232029 87611 232147
rect 87653 232029 87771 232147
rect 87493 214189 87611 214307
rect 87653 214189 87771 214307
rect 87493 214029 87611 214147
rect 87653 214029 87771 214147
rect 87493 196189 87611 196307
rect 87653 196189 87771 196307
rect 87493 196029 87611 196147
rect 87653 196029 87771 196147
rect 87493 178189 87611 178307
rect 87653 178189 87771 178307
rect 87493 178029 87611 178147
rect 87653 178029 87771 178147
rect 87493 160189 87611 160307
rect 87653 160189 87771 160307
rect 87493 160029 87611 160147
rect 87653 160029 87771 160147
rect 87493 142189 87611 142307
rect 87653 142189 87771 142307
rect 87493 142029 87611 142147
rect 87653 142029 87771 142147
rect 87493 124189 87611 124307
rect 87653 124189 87771 124307
rect 87493 124029 87611 124147
rect 87653 124029 87771 124147
rect 87493 106189 87611 106307
rect 87653 106189 87771 106307
rect 87493 106029 87611 106147
rect 87653 106029 87771 106147
rect 87493 88189 87611 88307
rect 87653 88189 87771 88307
rect 87493 88029 87611 88147
rect 87653 88029 87771 88147
rect 87493 70189 87611 70307
rect 87653 70189 87771 70307
rect 87493 70029 87611 70147
rect 87653 70029 87771 70147
rect 87493 52189 87611 52307
rect 87653 52189 87771 52307
rect 87493 52029 87611 52147
rect 87653 52029 87771 52147
rect 87493 34189 87611 34307
rect 87653 34189 87771 34307
rect 87493 34029 87611 34147
rect 87653 34029 87771 34147
rect 87493 16189 87611 16307
rect 87653 16189 87771 16307
rect 87493 16029 87611 16147
rect 87653 16029 87771 16147
rect 78493 -3171 78611 -3053
rect 78653 -3171 78771 -3053
rect 78493 -3331 78611 -3213
rect 78653 -3331 78771 -3213
rect 90913 352301 91031 352419
rect 91073 352301 91191 352419
rect 90913 352141 91031 352259
rect 91073 352141 91191 352259
rect 90913 343609 91031 343727
rect 91073 343609 91191 343727
rect 90913 343449 91031 343567
rect 91073 343449 91191 343567
rect 90913 325609 91031 325727
rect 91073 325609 91191 325727
rect 90913 325449 91031 325567
rect 91073 325449 91191 325567
rect 90913 307609 91031 307727
rect 91073 307609 91191 307727
rect 90913 307449 91031 307567
rect 91073 307449 91191 307567
rect 90913 289609 91031 289727
rect 91073 289609 91191 289727
rect 90913 289449 91031 289567
rect 91073 289449 91191 289567
rect 90913 271609 91031 271727
rect 91073 271609 91191 271727
rect 90913 271449 91031 271567
rect 91073 271449 91191 271567
rect 90913 253609 91031 253727
rect 91073 253609 91191 253727
rect 90913 253449 91031 253567
rect 91073 253449 91191 253567
rect 90913 235609 91031 235727
rect 91073 235609 91191 235727
rect 90913 235449 91031 235567
rect 91073 235449 91191 235567
rect 90913 217609 91031 217727
rect 91073 217609 91191 217727
rect 90913 217449 91031 217567
rect 91073 217449 91191 217567
rect 90913 199609 91031 199727
rect 91073 199609 91191 199727
rect 90913 199449 91031 199567
rect 91073 199449 91191 199567
rect 90913 181609 91031 181727
rect 91073 181609 91191 181727
rect 90913 181449 91031 181567
rect 91073 181449 91191 181567
rect 90913 163609 91031 163727
rect 91073 163609 91191 163727
rect 90913 163449 91031 163567
rect 91073 163449 91191 163567
rect 90913 145609 91031 145727
rect 91073 145609 91191 145727
rect 90913 145449 91031 145567
rect 91073 145449 91191 145567
rect 90913 127609 91031 127727
rect 91073 127609 91191 127727
rect 90913 127449 91031 127567
rect 91073 127449 91191 127567
rect 90913 109609 91031 109727
rect 91073 109609 91191 109727
rect 90913 109449 91031 109567
rect 91073 109449 91191 109567
rect 90913 91609 91031 91727
rect 91073 91609 91191 91727
rect 90913 91449 91031 91567
rect 91073 91449 91191 91567
rect 90913 73609 91031 73727
rect 91073 73609 91191 73727
rect 90913 73449 91031 73567
rect 91073 73449 91191 73567
rect 90913 55609 91031 55727
rect 91073 55609 91191 55727
rect 90913 55449 91031 55567
rect 91073 55449 91191 55567
rect 90913 37609 91031 37727
rect 91073 37609 91191 37727
rect 90913 37449 91031 37567
rect 91073 37449 91191 37567
rect 90913 19609 91031 19727
rect 91073 19609 91191 19727
rect 90913 19449 91031 19567
rect 91073 19449 91191 19567
rect 90913 1609 91031 1727
rect 91073 1609 91191 1727
rect 90913 1449 91031 1567
rect 91073 1449 91191 1567
rect 90913 -291 91031 -173
rect 91073 -291 91191 -173
rect 90913 -451 91031 -333
rect 91073 -451 91191 -333
rect 92773 345469 92891 345587
rect 92933 345469 93051 345587
rect 92773 345309 92891 345427
rect 92933 345309 93051 345427
rect 92773 327469 92891 327587
rect 92933 327469 93051 327587
rect 92773 327309 92891 327427
rect 92933 327309 93051 327427
rect 92773 309469 92891 309587
rect 92933 309469 93051 309587
rect 92773 309309 92891 309427
rect 92933 309309 93051 309427
rect 92773 291469 92891 291587
rect 92933 291469 93051 291587
rect 92773 291309 92891 291427
rect 92933 291309 93051 291427
rect 92773 273469 92891 273587
rect 92933 273469 93051 273587
rect 92773 273309 92891 273427
rect 92933 273309 93051 273427
rect 92773 255469 92891 255587
rect 92933 255469 93051 255587
rect 92773 255309 92891 255427
rect 92933 255309 93051 255427
rect 92773 237469 92891 237587
rect 92933 237469 93051 237587
rect 92773 237309 92891 237427
rect 92933 237309 93051 237427
rect 92773 219469 92891 219587
rect 92933 219469 93051 219587
rect 92773 219309 92891 219427
rect 92933 219309 93051 219427
rect 92773 201469 92891 201587
rect 92933 201469 93051 201587
rect 92773 201309 92891 201427
rect 92933 201309 93051 201427
rect 92773 183469 92891 183587
rect 92933 183469 93051 183587
rect 92773 183309 92891 183427
rect 92933 183309 93051 183427
rect 92773 165469 92891 165587
rect 92933 165469 93051 165587
rect 92773 165309 92891 165427
rect 92933 165309 93051 165427
rect 92773 147469 92891 147587
rect 92933 147469 93051 147587
rect 92773 147309 92891 147427
rect 92933 147309 93051 147427
rect 92773 129469 92891 129587
rect 92933 129469 93051 129587
rect 92773 129309 92891 129427
rect 92933 129309 93051 129427
rect 92773 111469 92891 111587
rect 92933 111469 93051 111587
rect 92773 111309 92891 111427
rect 92933 111309 93051 111427
rect 92773 93469 92891 93587
rect 92933 93469 93051 93587
rect 92773 93309 92891 93427
rect 92933 93309 93051 93427
rect 92773 75469 92891 75587
rect 92933 75469 93051 75587
rect 92773 75309 92891 75427
rect 92933 75309 93051 75427
rect 92773 57469 92891 57587
rect 92933 57469 93051 57587
rect 92773 57309 92891 57427
rect 92933 57309 93051 57427
rect 92773 39469 92891 39587
rect 92933 39469 93051 39587
rect 92773 39309 92891 39427
rect 92933 39309 93051 39427
rect 92773 21469 92891 21587
rect 92933 21469 93051 21587
rect 92773 21309 92891 21427
rect 92933 21309 93051 21427
rect 92773 3469 92891 3587
rect 92933 3469 93051 3587
rect 92773 3309 92891 3427
rect 92933 3309 93051 3427
rect 92773 -1251 92891 -1133
rect 92933 -1251 93051 -1133
rect 92773 -1411 92891 -1293
rect 92933 -1411 93051 -1293
rect 94633 347329 94751 347447
rect 94793 347329 94911 347447
rect 94633 347169 94751 347287
rect 94793 347169 94911 347287
rect 94633 329329 94751 329447
rect 94793 329329 94911 329447
rect 94633 329169 94751 329287
rect 94793 329169 94911 329287
rect 94633 311329 94751 311447
rect 94793 311329 94911 311447
rect 94633 311169 94751 311287
rect 94793 311169 94911 311287
rect 94633 293329 94751 293447
rect 94793 293329 94911 293447
rect 94633 293169 94751 293287
rect 94793 293169 94911 293287
rect 94633 275329 94751 275447
rect 94793 275329 94911 275447
rect 94633 275169 94751 275287
rect 94793 275169 94911 275287
rect 94633 257329 94751 257447
rect 94793 257329 94911 257447
rect 94633 257169 94751 257287
rect 94793 257169 94911 257287
rect 94633 239329 94751 239447
rect 94793 239329 94911 239447
rect 94633 239169 94751 239287
rect 94793 239169 94911 239287
rect 94633 221329 94751 221447
rect 94793 221329 94911 221447
rect 94633 221169 94751 221287
rect 94793 221169 94911 221287
rect 94633 203329 94751 203447
rect 94793 203329 94911 203447
rect 94633 203169 94751 203287
rect 94793 203169 94911 203287
rect 94633 185329 94751 185447
rect 94793 185329 94911 185447
rect 94633 185169 94751 185287
rect 94793 185169 94911 185287
rect 94633 167329 94751 167447
rect 94793 167329 94911 167447
rect 94633 167169 94751 167287
rect 94793 167169 94911 167287
rect 94633 149329 94751 149447
rect 94793 149329 94911 149447
rect 94633 149169 94751 149287
rect 94793 149169 94911 149287
rect 94633 131329 94751 131447
rect 94793 131329 94911 131447
rect 94633 131169 94751 131287
rect 94793 131169 94911 131287
rect 94633 113329 94751 113447
rect 94793 113329 94911 113447
rect 94633 113169 94751 113287
rect 94793 113169 94911 113287
rect 94633 95329 94751 95447
rect 94793 95329 94911 95447
rect 94633 95169 94751 95287
rect 94793 95169 94911 95287
rect 94633 77329 94751 77447
rect 94793 77329 94911 77447
rect 94633 77169 94751 77287
rect 94793 77169 94911 77287
rect 94633 59329 94751 59447
rect 94793 59329 94911 59447
rect 94633 59169 94751 59287
rect 94793 59169 94911 59287
rect 94633 41329 94751 41447
rect 94793 41329 94911 41447
rect 94633 41169 94751 41287
rect 94793 41169 94911 41287
rect 94633 23329 94751 23447
rect 94793 23329 94911 23447
rect 94633 23169 94751 23287
rect 94793 23169 94911 23287
rect 94633 5329 94751 5447
rect 94793 5329 94911 5447
rect 94633 5169 94751 5287
rect 94793 5169 94911 5287
rect 94633 -2211 94751 -2093
rect 94793 -2211 94911 -2093
rect 94633 -2371 94751 -2253
rect 94793 -2371 94911 -2253
rect 105493 355661 105611 355779
rect 105653 355661 105771 355779
rect 105493 355501 105611 355619
rect 105653 355501 105771 355619
rect 103633 354701 103751 354819
rect 103793 354701 103911 354819
rect 103633 354541 103751 354659
rect 103793 354541 103911 354659
rect 101773 353741 101891 353859
rect 101933 353741 102051 353859
rect 101773 353581 101891 353699
rect 101933 353581 102051 353699
rect 96493 349189 96611 349307
rect 96653 349189 96771 349307
rect 96493 349029 96611 349147
rect 96653 349029 96771 349147
rect 96493 331189 96611 331307
rect 96653 331189 96771 331307
rect 96493 331029 96611 331147
rect 96653 331029 96771 331147
rect 96493 313189 96611 313307
rect 96653 313189 96771 313307
rect 96493 313029 96611 313147
rect 96653 313029 96771 313147
rect 96493 295189 96611 295307
rect 96653 295189 96771 295307
rect 96493 295029 96611 295147
rect 96653 295029 96771 295147
rect 96493 277189 96611 277307
rect 96653 277189 96771 277307
rect 96493 277029 96611 277147
rect 96653 277029 96771 277147
rect 96493 259189 96611 259307
rect 96653 259189 96771 259307
rect 96493 259029 96611 259147
rect 96653 259029 96771 259147
rect 96493 241189 96611 241307
rect 96653 241189 96771 241307
rect 96493 241029 96611 241147
rect 96653 241029 96771 241147
rect 96493 223189 96611 223307
rect 96653 223189 96771 223307
rect 96493 223029 96611 223147
rect 96653 223029 96771 223147
rect 96493 205189 96611 205307
rect 96653 205189 96771 205307
rect 96493 205029 96611 205147
rect 96653 205029 96771 205147
rect 96493 187189 96611 187307
rect 96653 187189 96771 187307
rect 96493 187029 96611 187147
rect 96653 187029 96771 187147
rect 96493 169189 96611 169307
rect 96653 169189 96771 169307
rect 96493 169029 96611 169147
rect 96653 169029 96771 169147
rect 96493 151189 96611 151307
rect 96653 151189 96771 151307
rect 96493 151029 96611 151147
rect 96653 151029 96771 151147
rect 96493 133189 96611 133307
rect 96653 133189 96771 133307
rect 96493 133029 96611 133147
rect 96653 133029 96771 133147
rect 96493 115189 96611 115307
rect 96653 115189 96771 115307
rect 96493 115029 96611 115147
rect 96653 115029 96771 115147
rect 96493 97189 96611 97307
rect 96653 97189 96771 97307
rect 96493 97029 96611 97147
rect 96653 97029 96771 97147
rect 96493 79189 96611 79307
rect 96653 79189 96771 79307
rect 96493 79029 96611 79147
rect 96653 79029 96771 79147
rect 96493 61189 96611 61307
rect 96653 61189 96771 61307
rect 96493 61029 96611 61147
rect 96653 61029 96771 61147
rect 96493 43189 96611 43307
rect 96653 43189 96771 43307
rect 96493 43029 96611 43147
rect 96653 43029 96771 43147
rect 96493 25189 96611 25307
rect 96653 25189 96771 25307
rect 96493 25029 96611 25147
rect 96653 25029 96771 25147
rect 96493 7189 96611 7307
rect 96653 7189 96771 7307
rect 96493 7029 96611 7147
rect 96653 7029 96771 7147
rect 87493 -3651 87611 -3533
rect 87653 -3651 87771 -3533
rect 87493 -3811 87611 -3693
rect 87653 -3811 87771 -3693
rect 99913 352781 100031 352899
rect 100073 352781 100191 352899
rect 99913 352621 100031 352739
rect 100073 352621 100191 352739
rect 99913 334609 100031 334727
rect 100073 334609 100191 334727
rect 99913 334449 100031 334567
rect 100073 334449 100191 334567
rect 99913 316609 100031 316727
rect 100073 316609 100191 316727
rect 99913 316449 100031 316567
rect 100073 316449 100191 316567
rect 99913 298609 100031 298727
rect 100073 298609 100191 298727
rect 99913 298449 100031 298567
rect 100073 298449 100191 298567
rect 99913 280609 100031 280727
rect 100073 280609 100191 280727
rect 99913 280449 100031 280567
rect 100073 280449 100191 280567
rect 99913 262609 100031 262727
rect 100073 262609 100191 262727
rect 99913 262449 100031 262567
rect 100073 262449 100191 262567
rect 99913 244609 100031 244727
rect 100073 244609 100191 244727
rect 99913 244449 100031 244567
rect 100073 244449 100191 244567
rect 99913 226609 100031 226727
rect 100073 226609 100191 226727
rect 99913 226449 100031 226567
rect 100073 226449 100191 226567
rect 99913 208609 100031 208727
rect 100073 208609 100191 208727
rect 99913 208449 100031 208567
rect 100073 208449 100191 208567
rect 99913 190609 100031 190727
rect 100073 190609 100191 190727
rect 99913 190449 100031 190567
rect 100073 190449 100191 190567
rect 99913 172609 100031 172727
rect 100073 172609 100191 172727
rect 99913 172449 100031 172567
rect 100073 172449 100191 172567
rect 99913 154609 100031 154727
rect 100073 154609 100191 154727
rect 99913 154449 100031 154567
rect 100073 154449 100191 154567
rect 99913 136609 100031 136727
rect 100073 136609 100191 136727
rect 99913 136449 100031 136567
rect 100073 136449 100191 136567
rect 99913 118609 100031 118727
rect 100073 118609 100191 118727
rect 99913 118449 100031 118567
rect 100073 118449 100191 118567
rect 99913 100609 100031 100727
rect 100073 100609 100191 100727
rect 99913 100449 100031 100567
rect 100073 100449 100191 100567
rect 99913 82609 100031 82727
rect 100073 82609 100191 82727
rect 99913 82449 100031 82567
rect 100073 82449 100191 82567
rect 99913 64609 100031 64727
rect 100073 64609 100191 64727
rect 99913 64449 100031 64567
rect 100073 64449 100191 64567
rect 99913 46609 100031 46727
rect 100073 46609 100191 46727
rect 99913 46449 100031 46567
rect 100073 46449 100191 46567
rect 99913 28609 100031 28727
rect 100073 28609 100191 28727
rect 99913 28449 100031 28567
rect 100073 28449 100191 28567
rect 99913 10609 100031 10727
rect 100073 10609 100191 10727
rect 99913 10449 100031 10567
rect 100073 10449 100191 10567
rect 99913 -771 100031 -653
rect 100073 -771 100191 -653
rect 99913 -931 100031 -813
rect 100073 -931 100191 -813
rect 101773 336469 101891 336587
rect 101933 336469 102051 336587
rect 101773 336309 101891 336427
rect 101933 336309 102051 336427
rect 101773 318469 101891 318587
rect 101933 318469 102051 318587
rect 101773 318309 101891 318427
rect 101933 318309 102051 318427
rect 101773 300469 101891 300587
rect 101933 300469 102051 300587
rect 101773 300309 101891 300427
rect 101933 300309 102051 300427
rect 101773 282469 101891 282587
rect 101933 282469 102051 282587
rect 101773 282309 101891 282427
rect 101933 282309 102051 282427
rect 101773 264469 101891 264587
rect 101933 264469 102051 264587
rect 101773 264309 101891 264427
rect 101933 264309 102051 264427
rect 101773 246469 101891 246587
rect 101933 246469 102051 246587
rect 101773 246309 101891 246427
rect 101933 246309 102051 246427
rect 101773 228469 101891 228587
rect 101933 228469 102051 228587
rect 101773 228309 101891 228427
rect 101933 228309 102051 228427
rect 101773 210469 101891 210587
rect 101933 210469 102051 210587
rect 101773 210309 101891 210427
rect 101933 210309 102051 210427
rect 101773 192469 101891 192587
rect 101933 192469 102051 192587
rect 101773 192309 101891 192427
rect 101933 192309 102051 192427
rect 101773 174469 101891 174587
rect 101933 174469 102051 174587
rect 101773 174309 101891 174427
rect 101933 174309 102051 174427
rect 101773 156469 101891 156587
rect 101933 156469 102051 156587
rect 101773 156309 101891 156427
rect 101933 156309 102051 156427
rect 101773 138469 101891 138587
rect 101933 138469 102051 138587
rect 101773 138309 101891 138427
rect 101933 138309 102051 138427
rect 101773 120469 101891 120587
rect 101933 120469 102051 120587
rect 101773 120309 101891 120427
rect 101933 120309 102051 120427
rect 101773 102469 101891 102587
rect 101933 102469 102051 102587
rect 101773 102309 101891 102427
rect 101933 102309 102051 102427
rect 101773 84469 101891 84587
rect 101933 84469 102051 84587
rect 101773 84309 101891 84427
rect 101933 84309 102051 84427
rect 101773 66469 101891 66587
rect 101933 66469 102051 66587
rect 101773 66309 101891 66427
rect 101933 66309 102051 66427
rect 101773 48469 101891 48587
rect 101933 48469 102051 48587
rect 101773 48309 101891 48427
rect 101933 48309 102051 48427
rect 101773 30469 101891 30587
rect 101933 30469 102051 30587
rect 101773 30309 101891 30427
rect 101933 30309 102051 30427
rect 101773 12469 101891 12587
rect 101933 12469 102051 12587
rect 101773 12309 101891 12427
rect 101933 12309 102051 12427
rect 101773 -1731 101891 -1613
rect 101933 -1731 102051 -1613
rect 101773 -1891 101891 -1773
rect 101933 -1891 102051 -1773
rect 103633 338329 103751 338447
rect 103793 338329 103911 338447
rect 103633 338169 103751 338287
rect 103793 338169 103911 338287
rect 103633 320329 103751 320447
rect 103793 320329 103911 320447
rect 103633 320169 103751 320287
rect 103793 320169 103911 320287
rect 103633 302329 103751 302447
rect 103793 302329 103911 302447
rect 103633 302169 103751 302287
rect 103793 302169 103911 302287
rect 103633 284329 103751 284447
rect 103793 284329 103911 284447
rect 103633 284169 103751 284287
rect 103793 284169 103911 284287
rect 103633 266329 103751 266447
rect 103793 266329 103911 266447
rect 103633 266169 103751 266287
rect 103793 266169 103911 266287
rect 103633 248329 103751 248447
rect 103793 248329 103911 248447
rect 103633 248169 103751 248287
rect 103793 248169 103911 248287
rect 103633 230329 103751 230447
rect 103793 230329 103911 230447
rect 103633 230169 103751 230287
rect 103793 230169 103911 230287
rect 103633 212329 103751 212447
rect 103793 212329 103911 212447
rect 103633 212169 103751 212287
rect 103793 212169 103911 212287
rect 103633 194329 103751 194447
rect 103793 194329 103911 194447
rect 103633 194169 103751 194287
rect 103793 194169 103911 194287
rect 103633 176329 103751 176447
rect 103793 176329 103911 176447
rect 103633 176169 103751 176287
rect 103793 176169 103911 176287
rect 103633 158329 103751 158447
rect 103793 158329 103911 158447
rect 103633 158169 103751 158287
rect 103793 158169 103911 158287
rect 103633 140329 103751 140447
rect 103793 140329 103911 140447
rect 103633 140169 103751 140287
rect 103793 140169 103911 140287
rect 103633 122329 103751 122447
rect 103793 122329 103911 122447
rect 103633 122169 103751 122287
rect 103793 122169 103911 122287
rect 103633 104329 103751 104447
rect 103793 104329 103911 104447
rect 103633 104169 103751 104287
rect 103793 104169 103911 104287
rect 103633 86329 103751 86447
rect 103793 86329 103911 86447
rect 103633 86169 103751 86287
rect 103793 86169 103911 86287
rect 103633 68329 103751 68447
rect 103793 68329 103911 68447
rect 103633 68169 103751 68287
rect 103793 68169 103911 68287
rect 103633 50329 103751 50447
rect 103793 50329 103911 50447
rect 103633 50169 103751 50287
rect 103793 50169 103911 50287
rect 103633 32329 103751 32447
rect 103793 32329 103911 32447
rect 103633 32169 103751 32287
rect 103793 32169 103911 32287
rect 103633 14329 103751 14447
rect 103793 14329 103911 14447
rect 103633 14169 103751 14287
rect 103793 14169 103911 14287
rect 103633 -2691 103751 -2573
rect 103793 -2691 103911 -2573
rect 103633 -2851 103751 -2733
rect 103793 -2851 103911 -2733
rect 114493 355181 114611 355299
rect 114653 355181 114771 355299
rect 114493 355021 114611 355139
rect 114653 355021 114771 355139
rect 112633 354221 112751 354339
rect 112793 354221 112911 354339
rect 112633 354061 112751 354179
rect 112793 354061 112911 354179
rect 110773 353261 110891 353379
rect 110933 353261 111051 353379
rect 110773 353101 110891 353219
rect 110933 353101 111051 353219
rect 105493 340189 105611 340307
rect 105653 340189 105771 340307
rect 105493 340029 105611 340147
rect 105653 340029 105771 340147
rect 105493 322189 105611 322307
rect 105653 322189 105771 322307
rect 105493 322029 105611 322147
rect 105653 322029 105771 322147
rect 105493 304189 105611 304307
rect 105653 304189 105771 304307
rect 105493 304029 105611 304147
rect 105653 304029 105771 304147
rect 105493 286189 105611 286307
rect 105653 286189 105771 286307
rect 105493 286029 105611 286147
rect 105653 286029 105771 286147
rect 105493 268189 105611 268307
rect 105653 268189 105771 268307
rect 105493 268029 105611 268147
rect 105653 268029 105771 268147
rect 105493 250189 105611 250307
rect 105653 250189 105771 250307
rect 105493 250029 105611 250147
rect 105653 250029 105771 250147
rect 105493 232189 105611 232307
rect 105653 232189 105771 232307
rect 105493 232029 105611 232147
rect 105653 232029 105771 232147
rect 105493 214189 105611 214307
rect 105653 214189 105771 214307
rect 105493 214029 105611 214147
rect 105653 214029 105771 214147
rect 105493 196189 105611 196307
rect 105653 196189 105771 196307
rect 105493 196029 105611 196147
rect 105653 196029 105771 196147
rect 105493 178189 105611 178307
rect 105653 178189 105771 178307
rect 105493 178029 105611 178147
rect 105653 178029 105771 178147
rect 105493 160189 105611 160307
rect 105653 160189 105771 160307
rect 105493 160029 105611 160147
rect 105653 160029 105771 160147
rect 105493 142189 105611 142307
rect 105653 142189 105771 142307
rect 105493 142029 105611 142147
rect 105653 142029 105771 142147
rect 105493 124189 105611 124307
rect 105653 124189 105771 124307
rect 105493 124029 105611 124147
rect 105653 124029 105771 124147
rect 105493 106189 105611 106307
rect 105653 106189 105771 106307
rect 105493 106029 105611 106147
rect 105653 106029 105771 106147
rect 105493 88189 105611 88307
rect 105653 88189 105771 88307
rect 105493 88029 105611 88147
rect 105653 88029 105771 88147
rect 105493 70189 105611 70307
rect 105653 70189 105771 70307
rect 105493 70029 105611 70147
rect 105653 70029 105771 70147
rect 105493 52189 105611 52307
rect 105653 52189 105771 52307
rect 105493 52029 105611 52147
rect 105653 52029 105771 52147
rect 105493 34189 105611 34307
rect 105653 34189 105771 34307
rect 105493 34029 105611 34147
rect 105653 34029 105771 34147
rect 105493 16189 105611 16307
rect 105653 16189 105771 16307
rect 105493 16029 105611 16147
rect 105653 16029 105771 16147
rect 96493 -3171 96611 -3053
rect 96653 -3171 96771 -3053
rect 96493 -3331 96611 -3213
rect 96653 -3331 96771 -3213
rect 108913 352301 109031 352419
rect 109073 352301 109191 352419
rect 108913 352141 109031 352259
rect 109073 352141 109191 352259
rect 108913 343609 109031 343727
rect 109073 343609 109191 343727
rect 108913 343449 109031 343567
rect 109073 343449 109191 343567
rect 108913 325609 109031 325727
rect 109073 325609 109191 325727
rect 108913 325449 109031 325567
rect 109073 325449 109191 325567
rect 108913 307609 109031 307727
rect 109073 307609 109191 307727
rect 108913 307449 109031 307567
rect 109073 307449 109191 307567
rect 108913 289609 109031 289727
rect 109073 289609 109191 289727
rect 108913 289449 109031 289567
rect 109073 289449 109191 289567
rect 108913 271609 109031 271727
rect 109073 271609 109191 271727
rect 108913 271449 109031 271567
rect 109073 271449 109191 271567
rect 108913 253609 109031 253727
rect 109073 253609 109191 253727
rect 108913 253449 109031 253567
rect 109073 253449 109191 253567
rect 108913 235609 109031 235727
rect 109073 235609 109191 235727
rect 108913 235449 109031 235567
rect 109073 235449 109191 235567
rect 108913 217609 109031 217727
rect 109073 217609 109191 217727
rect 108913 217449 109031 217567
rect 109073 217449 109191 217567
rect 108913 199609 109031 199727
rect 109073 199609 109191 199727
rect 108913 199449 109031 199567
rect 109073 199449 109191 199567
rect 108913 181609 109031 181727
rect 109073 181609 109191 181727
rect 108913 181449 109031 181567
rect 109073 181449 109191 181567
rect 108913 163609 109031 163727
rect 109073 163609 109191 163727
rect 108913 163449 109031 163567
rect 109073 163449 109191 163567
rect 108913 145609 109031 145727
rect 109073 145609 109191 145727
rect 108913 145449 109031 145567
rect 109073 145449 109191 145567
rect 108913 127609 109031 127727
rect 109073 127609 109191 127727
rect 108913 127449 109031 127567
rect 109073 127449 109191 127567
rect 108913 109609 109031 109727
rect 109073 109609 109191 109727
rect 108913 109449 109031 109567
rect 109073 109449 109191 109567
rect 108913 91609 109031 91727
rect 109073 91609 109191 91727
rect 108913 91449 109031 91567
rect 109073 91449 109191 91567
rect 108913 73609 109031 73727
rect 109073 73609 109191 73727
rect 108913 73449 109031 73567
rect 109073 73449 109191 73567
rect 108913 55609 109031 55727
rect 109073 55609 109191 55727
rect 108913 55449 109031 55567
rect 109073 55449 109191 55567
rect 108913 37609 109031 37727
rect 109073 37609 109191 37727
rect 108913 37449 109031 37567
rect 109073 37449 109191 37567
rect 108913 19609 109031 19727
rect 109073 19609 109191 19727
rect 108913 19449 109031 19567
rect 109073 19449 109191 19567
rect 108913 1609 109031 1727
rect 109073 1609 109191 1727
rect 108913 1449 109031 1567
rect 109073 1449 109191 1567
rect 108913 -291 109031 -173
rect 109073 -291 109191 -173
rect 108913 -451 109031 -333
rect 109073 -451 109191 -333
rect 110773 345469 110891 345587
rect 110933 345469 111051 345587
rect 110773 345309 110891 345427
rect 110933 345309 111051 345427
rect 110773 327469 110891 327587
rect 110933 327469 111051 327587
rect 110773 327309 110891 327427
rect 110933 327309 111051 327427
rect 110773 309469 110891 309587
rect 110933 309469 111051 309587
rect 110773 309309 110891 309427
rect 110933 309309 111051 309427
rect 110773 291469 110891 291587
rect 110933 291469 111051 291587
rect 110773 291309 110891 291427
rect 110933 291309 111051 291427
rect 110773 273469 110891 273587
rect 110933 273469 111051 273587
rect 110773 273309 110891 273427
rect 110933 273309 111051 273427
rect 110773 255469 110891 255587
rect 110933 255469 111051 255587
rect 110773 255309 110891 255427
rect 110933 255309 111051 255427
rect 110773 237469 110891 237587
rect 110933 237469 111051 237587
rect 110773 237309 110891 237427
rect 110933 237309 111051 237427
rect 110773 219469 110891 219587
rect 110933 219469 111051 219587
rect 110773 219309 110891 219427
rect 110933 219309 111051 219427
rect 110773 201469 110891 201587
rect 110933 201469 111051 201587
rect 110773 201309 110891 201427
rect 110933 201309 111051 201427
rect 110773 183469 110891 183587
rect 110933 183469 111051 183587
rect 110773 183309 110891 183427
rect 110933 183309 111051 183427
rect 110773 165469 110891 165587
rect 110933 165469 111051 165587
rect 110773 165309 110891 165427
rect 110933 165309 111051 165427
rect 110773 147469 110891 147587
rect 110933 147469 111051 147587
rect 110773 147309 110891 147427
rect 110933 147309 111051 147427
rect 110773 129469 110891 129587
rect 110933 129469 111051 129587
rect 110773 129309 110891 129427
rect 110933 129309 111051 129427
rect 110773 111469 110891 111587
rect 110933 111469 111051 111587
rect 110773 111309 110891 111427
rect 110933 111309 111051 111427
rect 110773 93469 110891 93587
rect 110933 93469 111051 93587
rect 110773 93309 110891 93427
rect 110933 93309 111051 93427
rect 110773 75469 110891 75587
rect 110933 75469 111051 75587
rect 110773 75309 110891 75427
rect 110933 75309 111051 75427
rect 110773 57469 110891 57587
rect 110933 57469 111051 57587
rect 110773 57309 110891 57427
rect 110933 57309 111051 57427
rect 110773 39469 110891 39587
rect 110933 39469 111051 39587
rect 110773 39309 110891 39427
rect 110933 39309 111051 39427
rect 110773 21469 110891 21587
rect 110933 21469 111051 21587
rect 110773 21309 110891 21427
rect 110933 21309 111051 21427
rect 110773 3469 110891 3587
rect 110933 3469 111051 3587
rect 110773 3309 110891 3427
rect 110933 3309 111051 3427
rect 110773 -1251 110891 -1133
rect 110933 -1251 111051 -1133
rect 110773 -1411 110891 -1293
rect 110933 -1411 111051 -1293
rect 112633 347329 112751 347447
rect 112793 347329 112911 347447
rect 112633 347169 112751 347287
rect 112793 347169 112911 347287
rect 112633 329329 112751 329447
rect 112793 329329 112911 329447
rect 112633 329169 112751 329287
rect 112793 329169 112911 329287
rect 112633 311329 112751 311447
rect 112793 311329 112911 311447
rect 112633 311169 112751 311287
rect 112793 311169 112911 311287
rect 112633 293329 112751 293447
rect 112793 293329 112911 293447
rect 112633 293169 112751 293287
rect 112793 293169 112911 293287
rect 112633 275329 112751 275447
rect 112793 275329 112911 275447
rect 112633 275169 112751 275287
rect 112793 275169 112911 275287
rect 112633 257329 112751 257447
rect 112793 257329 112911 257447
rect 112633 257169 112751 257287
rect 112793 257169 112911 257287
rect 112633 239329 112751 239447
rect 112793 239329 112911 239447
rect 112633 239169 112751 239287
rect 112793 239169 112911 239287
rect 112633 221329 112751 221447
rect 112793 221329 112911 221447
rect 112633 221169 112751 221287
rect 112793 221169 112911 221287
rect 112633 203329 112751 203447
rect 112793 203329 112911 203447
rect 112633 203169 112751 203287
rect 112793 203169 112911 203287
rect 112633 185329 112751 185447
rect 112793 185329 112911 185447
rect 112633 185169 112751 185287
rect 112793 185169 112911 185287
rect 112633 167329 112751 167447
rect 112793 167329 112911 167447
rect 112633 167169 112751 167287
rect 112793 167169 112911 167287
rect 112633 149329 112751 149447
rect 112793 149329 112911 149447
rect 112633 149169 112751 149287
rect 112793 149169 112911 149287
rect 112633 131329 112751 131447
rect 112793 131329 112911 131447
rect 112633 131169 112751 131287
rect 112793 131169 112911 131287
rect 112633 113329 112751 113447
rect 112793 113329 112911 113447
rect 112633 113169 112751 113287
rect 112793 113169 112911 113287
rect 112633 95329 112751 95447
rect 112793 95329 112911 95447
rect 112633 95169 112751 95287
rect 112793 95169 112911 95287
rect 112633 77329 112751 77447
rect 112793 77329 112911 77447
rect 112633 77169 112751 77287
rect 112793 77169 112911 77287
rect 112633 59329 112751 59447
rect 112793 59329 112911 59447
rect 112633 59169 112751 59287
rect 112793 59169 112911 59287
rect 112633 41329 112751 41447
rect 112793 41329 112911 41447
rect 112633 41169 112751 41287
rect 112793 41169 112911 41287
rect 112633 23329 112751 23447
rect 112793 23329 112911 23447
rect 112633 23169 112751 23287
rect 112793 23169 112911 23287
rect 112633 5329 112751 5447
rect 112793 5329 112911 5447
rect 112633 5169 112751 5287
rect 112793 5169 112911 5287
rect 112633 -2211 112751 -2093
rect 112793 -2211 112911 -2093
rect 112633 -2371 112751 -2253
rect 112793 -2371 112911 -2253
rect 123493 355661 123611 355779
rect 123653 355661 123771 355779
rect 123493 355501 123611 355619
rect 123653 355501 123771 355619
rect 121633 354701 121751 354819
rect 121793 354701 121911 354819
rect 121633 354541 121751 354659
rect 121793 354541 121911 354659
rect 119773 353741 119891 353859
rect 119933 353741 120051 353859
rect 119773 353581 119891 353699
rect 119933 353581 120051 353699
rect 114493 349189 114611 349307
rect 114653 349189 114771 349307
rect 114493 349029 114611 349147
rect 114653 349029 114771 349147
rect 114493 331189 114611 331307
rect 114653 331189 114771 331307
rect 114493 331029 114611 331147
rect 114653 331029 114771 331147
rect 114493 313189 114611 313307
rect 114653 313189 114771 313307
rect 114493 313029 114611 313147
rect 114653 313029 114771 313147
rect 114493 295189 114611 295307
rect 114653 295189 114771 295307
rect 114493 295029 114611 295147
rect 114653 295029 114771 295147
rect 114493 277189 114611 277307
rect 114653 277189 114771 277307
rect 114493 277029 114611 277147
rect 114653 277029 114771 277147
rect 114493 259189 114611 259307
rect 114653 259189 114771 259307
rect 114493 259029 114611 259147
rect 114653 259029 114771 259147
rect 114493 241189 114611 241307
rect 114653 241189 114771 241307
rect 114493 241029 114611 241147
rect 114653 241029 114771 241147
rect 114493 223189 114611 223307
rect 114653 223189 114771 223307
rect 114493 223029 114611 223147
rect 114653 223029 114771 223147
rect 114493 205189 114611 205307
rect 114653 205189 114771 205307
rect 114493 205029 114611 205147
rect 114653 205029 114771 205147
rect 114493 187189 114611 187307
rect 114653 187189 114771 187307
rect 114493 187029 114611 187147
rect 114653 187029 114771 187147
rect 114493 169189 114611 169307
rect 114653 169189 114771 169307
rect 114493 169029 114611 169147
rect 114653 169029 114771 169147
rect 114493 151189 114611 151307
rect 114653 151189 114771 151307
rect 114493 151029 114611 151147
rect 114653 151029 114771 151147
rect 114493 133189 114611 133307
rect 114653 133189 114771 133307
rect 114493 133029 114611 133147
rect 114653 133029 114771 133147
rect 114493 115189 114611 115307
rect 114653 115189 114771 115307
rect 114493 115029 114611 115147
rect 114653 115029 114771 115147
rect 114493 97189 114611 97307
rect 114653 97189 114771 97307
rect 114493 97029 114611 97147
rect 114653 97029 114771 97147
rect 114493 79189 114611 79307
rect 114653 79189 114771 79307
rect 114493 79029 114611 79147
rect 114653 79029 114771 79147
rect 114493 61189 114611 61307
rect 114653 61189 114771 61307
rect 114493 61029 114611 61147
rect 114653 61029 114771 61147
rect 114493 43189 114611 43307
rect 114653 43189 114771 43307
rect 114493 43029 114611 43147
rect 114653 43029 114771 43147
rect 114493 25189 114611 25307
rect 114653 25189 114771 25307
rect 114493 25029 114611 25147
rect 114653 25029 114771 25147
rect 114493 7189 114611 7307
rect 114653 7189 114771 7307
rect 114493 7029 114611 7147
rect 114653 7029 114771 7147
rect 105493 -3651 105611 -3533
rect 105653 -3651 105771 -3533
rect 105493 -3811 105611 -3693
rect 105653 -3811 105771 -3693
rect 117913 352781 118031 352899
rect 118073 352781 118191 352899
rect 117913 352621 118031 352739
rect 118073 352621 118191 352739
rect 117913 334609 118031 334727
rect 118073 334609 118191 334727
rect 117913 334449 118031 334567
rect 118073 334449 118191 334567
rect 117913 316609 118031 316727
rect 118073 316609 118191 316727
rect 117913 316449 118031 316567
rect 118073 316449 118191 316567
rect 117913 298609 118031 298727
rect 118073 298609 118191 298727
rect 117913 298449 118031 298567
rect 118073 298449 118191 298567
rect 117913 280609 118031 280727
rect 118073 280609 118191 280727
rect 117913 280449 118031 280567
rect 118073 280449 118191 280567
rect 117913 262609 118031 262727
rect 118073 262609 118191 262727
rect 117913 262449 118031 262567
rect 118073 262449 118191 262567
rect 117913 244609 118031 244727
rect 118073 244609 118191 244727
rect 117913 244449 118031 244567
rect 118073 244449 118191 244567
rect 117913 226609 118031 226727
rect 118073 226609 118191 226727
rect 117913 226449 118031 226567
rect 118073 226449 118191 226567
rect 117913 208609 118031 208727
rect 118073 208609 118191 208727
rect 117913 208449 118031 208567
rect 118073 208449 118191 208567
rect 117913 190609 118031 190727
rect 118073 190609 118191 190727
rect 117913 190449 118031 190567
rect 118073 190449 118191 190567
rect 117913 172609 118031 172727
rect 118073 172609 118191 172727
rect 117913 172449 118031 172567
rect 118073 172449 118191 172567
rect 117913 154609 118031 154727
rect 118073 154609 118191 154727
rect 117913 154449 118031 154567
rect 118073 154449 118191 154567
rect 117913 136609 118031 136727
rect 118073 136609 118191 136727
rect 117913 136449 118031 136567
rect 118073 136449 118191 136567
rect 117913 118609 118031 118727
rect 118073 118609 118191 118727
rect 117913 118449 118031 118567
rect 118073 118449 118191 118567
rect 117913 100609 118031 100727
rect 118073 100609 118191 100727
rect 117913 100449 118031 100567
rect 118073 100449 118191 100567
rect 117913 82609 118031 82727
rect 118073 82609 118191 82727
rect 117913 82449 118031 82567
rect 118073 82449 118191 82567
rect 117913 64609 118031 64727
rect 118073 64609 118191 64727
rect 117913 64449 118031 64567
rect 118073 64449 118191 64567
rect 117913 46609 118031 46727
rect 118073 46609 118191 46727
rect 117913 46449 118031 46567
rect 118073 46449 118191 46567
rect 117913 28609 118031 28727
rect 118073 28609 118191 28727
rect 117913 28449 118031 28567
rect 118073 28449 118191 28567
rect 117913 10609 118031 10727
rect 118073 10609 118191 10727
rect 117913 10449 118031 10567
rect 118073 10449 118191 10567
rect 117913 -771 118031 -653
rect 118073 -771 118191 -653
rect 117913 -931 118031 -813
rect 118073 -931 118191 -813
rect 119773 336469 119891 336587
rect 119933 336469 120051 336587
rect 119773 336309 119891 336427
rect 119933 336309 120051 336427
rect 119773 318469 119891 318587
rect 119933 318469 120051 318587
rect 119773 318309 119891 318427
rect 119933 318309 120051 318427
rect 119773 300469 119891 300587
rect 119933 300469 120051 300587
rect 119773 300309 119891 300427
rect 119933 300309 120051 300427
rect 119773 282469 119891 282587
rect 119933 282469 120051 282587
rect 119773 282309 119891 282427
rect 119933 282309 120051 282427
rect 119773 264469 119891 264587
rect 119933 264469 120051 264587
rect 119773 264309 119891 264427
rect 119933 264309 120051 264427
rect 119773 246469 119891 246587
rect 119933 246469 120051 246587
rect 119773 246309 119891 246427
rect 119933 246309 120051 246427
rect 119773 228469 119891 228587
rect 119933 228469 120051 228587
rect 119773 228309 119891 228427
rect 119933 228309 120051 228427
rect 119773 210469 119891 210587
rect 119933 210469 120051 210587
rect 119773 210309 119891 210427
rect 119933 210309 120051 210427
rect 119773 192469 119891 192587
rect 119933 192469 120051 192587
rect 119773 192309 119891 192427
rect 119933 192309 120051 192427
rect 119773 174469 119891 174587
rect 119933 174469 120051 174587
rect 119773 174309 119891 174427
rect 119933 174309 120051 174427
rect 119773 156469 119891 156587
rect 119933 156469 120051 156587
rect 119773 156309 119891 156427
rect 119933 156309 120051 156427
rect 119773 138469 119891 138587
rect 119933 138469 120051 138587
rect 119773 138309 119891 138427
rect 119933 138309 120051 138427
rect 119773 120469 119891 120587
rect 119933 120469 120051 120587
rect 119773 120309 119891 120427
rect 119933 120309 120051 120427
rect 119773 102469 119891 102587
rect 119933 102469 120051 102587
rect 119773 102309 119891 102427
rect 119933 102309 120051 102427
rect 119773 84469 119891 84587
rect 119933 84469 120051 84587
rect 119773 84309 119891 84427
rect 119933 84309 120051 84427
rect 119773 66469 119891 66587
rect 119933 66469 120051 66587
rect 119773 66309 119891 66427
rect 119933 66309 120051 66427
rect 119773 48469 119891 48587
rect 119933 48469 120051 48587
rect 119773 48309 119891 48427
rect 119933 48309 120051 48427
rect 119773 30469 119891 30587
rect 119933 30469 120051 30587
rect 119773 30309 119891 30427
rect 119933 30309 120051 30427
rect 119773 12469 119891 12587
rect 119933 12469 120051 12587
rect 119773 12309 119891 12427
rect 119933 12309 120051 12427
rect 119773 -1731 119891 -1613
rect 119933 -1731 120051 -1613
rect 119773 -1891 119891 -1773
rect 119933 -1891 120051 -1773
rect 121633 338329 121751 338447
rect 121793 338329 121911 338447
rect 121633 338169 121751 338287
rect 121793 338169 121911 338287
rect 121633 320329 121751 320447
rect 121793 320329 121911 320447
rect 121633 320169 121751 320287
rect 121793 320169 121911 320287
rect 121633 302329 121751 302447
rect 121793 302329 121911 302447
rect 121633 302169 121751 302287
rect 121793 302169 121911 302287
rect 121633 284329 121751 284447
rect 121793 284329 121911 284447
rect 121633 284169 121751 284287
rect 121793 284169 121911 284287
rect 121633 266329 121751 266447
rect 121793 266329 121911 266447
rect 121633 266169 121751 266287
rect 121793 266169 121911 266287
rect 121633 248329 121751 248447
rect 121793 248329 121911 248447
rect 121633 248169 121751 248287
rect 121793 248169 121911 248287
rect 121633 230329 121751 230447
rect 121793 230329 121911 230447
rect 121633 230169 121751 230287
rect 121793 230169 121911 230287
rect 121633 212329 121751 212447
rect 121793 212329 121911 212447
rect 121633 212169 121751 212287
rect 121793 212169 121911 212287
rect 121633 194329 121751 194447
rect 121793 194329 121911 194447
rect 121633 194169 121751 194287
rect 121793 194169 121911 194287
rect 121633 176329 121751 176447
rect 121793 176329 121911 176447
rect 121633 176169 121751 176287
rect 121793 176169 121911 176287
rect 121633 158329 121751 158447
rect 121793 158329 121911 158447
rect 121633 158169 121751 158287
rect 121793 158169 121911 158287
rect 121633 140329 121751 140447
rect 121793 140329 121911 140447
rect 121633 140169 121751 140287
rect 121793 140169 121911 140287
rect 121633 122329 121751 122447
rect 121793 122329 121911 122447
rect 121633 122169 121751 122287
rect 121793 122169 121911 122287
rect 121633 104329 121751 104447
rect 121793 104329 121911 104447
rect 121633 104169 121751 104287
rect 121793 104169 121911 104287
rect 121633 86329 121751 86447
rect 121793 86329 121911 86447
rect 121633 86169 121751 86287
rect 121793 86169 121911 86287
rect 121633 68329 121751 68447
rect 121793 68329 121911 68447
rect 121633 68169 121751 68287
rect 121793 68169 121911 68287
rect 121633 50329 121751 50447
rect 121793 50329 121911 50447
rect 121633 50169 121751 50287
rect 121793 50169 121911 50287
rect 121633 32329 121751 32447
rect 121793 32329 121911 32447
rect 121633 32169 121751 32287
rect 121793 32169 121911 32287
rect 121633 14329 121751 14447
rect 121793 14329 121911 14447
rect 121633 14169 121751 14287
rect 121793 14169 121911 14287
rect 121633 -2691 121751 -2573
rect 121793 -2691 121911 -2573
rect 121633 -2851 121751 -2733
rect 121793 -2851 121911 -2733
rect 132493 355181 132611 355299
rect 132653 355181 132771 355299
rect 132493 355021 132611 355139
rect 132653 355021 132771 355139
rect 130633 354221 130751 354339
rect 130793 354221 130911 354339
rect 130633 354061 130751 354179
rect 130793 354061 130911 354179
rect 128773 353261 128891 353379
rect 128933 353261 129051 353379
rect 128773 353101 128891 353219
rect 128933 353101 129051 353219
rect 123493 340189 123611 340307
rect 123653 340189 123771 340307
rect 123493 340029 123611 340147
rect 123653 340029 123771 340147
rect 123493 322189 123611 322307
rect 123653 322189 123771 322307
rect 123493 322029 123611 322147
rect 123653 322029 123771 322147
rect 123493 304189 123611 304307
rect 123653 304189 123771 304307
rect 123493 304029 123611 304147
rect 123653 304029 123771 304147
rect 123493 286189 123611 286307
rect 123653 286189 123771 286307
rect 123493 286029 123611 286147
rect 123653 286029 123771 286147
rect 123493 268189 123611 268307
rect 123653 268189 123771 268307
rect 123493 268029 123611 268147
rect 123653 268029 123771 268147
rect 123493 250189 123611 250307
rect 123653 250189 123771 250307
rect 123493 250029 123611 250147
rect 123653 250029 123771 250147
rect 123493 232189 123611 232307
rect 123653 232189 123771 232307
rect 123493 232029 123611 232147
rect 123653 232029 123771 232147
rect 123493 214189 123611 214307
rect 123653 214189 123771 214307
rect 123493 214029 123611 214147
rect 123653 214029 123771 214147
rect 123493 196189 123611 196307
rect 123653 196189 123771 196307
rect 123493 196029 123611 196147
rect 123653 196029 123771 196147
rect 123493 178189 123611 178307
rect 123653 178189 123771 178307
rect 123493 178029 123611 178147
rect 123653 178029 123771 178147
rect 123493 160189 123611 160307
rect 123653 160189 123771 160307
rect 123493 160029 123611 160147
rect 123653 160029 123771 160147
rect 123493 142189 123611 142307
rect 123653 142189 123771 142307
rect 123493 142029 123611 142147
rect 123653 142029 123771 142147
rect 123493 124189 123611 124307
rect 123653 124189 123771 124307
rect 123493 124029 123611 124147
rect 123653 124029 123771 124147
rect 123493 106189 123611 106307
rect 123653 106189 123771 106307
rect 123493 106029 123611 106147
rect 123653 106029 123771 106147
rect 123493 88189 123611 88307
rect 123653 88189 123771 88307
rect 123493 88029 123611 88147
rect 123653 88029 123771 88147
rect 123493 70189 123611 70307
rect 123653 70189 123771 70307
rect 123493 70029 123611 70147
rect 123653 70029 123771 70147
rect 123493 52189 123611 52307
rect 123653 52189 123771 52307
rect 123493 52029 123611 52147
rect 123653 52029 123771 52147
rect 123493 34189 123611 34307
rect 123653 34189 123771 34307
rect 123493 34029 123611 34147
rect 123653 34029 123771 34147
rect 123493 16189 123611 16307
rect 123653 16189 123771 16307
rect 123493 16029 123611 16147
rect 123653 16029 123771 16147
rect 114493 -3171 114611 -3053
rect 114653 -3171 114771 -3053
rect 114493 -3331 114611 -3213
rect 114653 -3331 114771 -3213
rect 126913 352301 127031 352419
rect 127073 352301 127191 352419
rect 126913 352141 127031 352259
rect 127073 352141 127191 352259
rect 126913 343609 127031 343727
rect 127073 343609 127191 343727
rect 126913 343449 127031 343567
rect 127073 343449 127191 343567
rect 126913 325609 127031 325727
rect 127073 325609 127191 325727
rect 126913 325449 127031 325567
rect 127073 325449 127191 325567
rect 126913 307609 127031 307727
rect 127073 307609 127191 307727
rect 126913 307449 127031 307567
rect 127073 307449 127191 307567
rect 126913 289609 127031 289727
rect 127073 289609 127191 289727
rect 126913 289449 127031 289567
rect 127073 289449 127191 289567
rect 126913 271609 127031 271727
rect 127073 271609 127191 271727
rect 126913 271449 127031 271567
rect 127073 271449 127191 271567
rect 126913 253609 127031 253727
rect 127073 253609 127191 253727
rect 126913 253449 127031 253567
rect 127073 253449 127191 253567
rect 126913 235609 127031 235727
rect 127073 235609 127191 235727
rect 126913 235449 127031 235567
rect 127073 235449 127191 235567
rect 126913 217609 127031 217727
rect 127073 217609 127191 217727
rect 126913 217449 127031 217567
rect 127073 217449 127191 217567
rect 126913 199609 127031 199727
rect 127073 199609 127191 199727
rect 126913 199449 127031 199567
rect 127073 199449 127191 199567
rect 126913 181609 127031 181727
rect 127073 181609 127191 181727
rect 126913 181449 127031 181567
rect 127073 181449 127191 181567
rect 126913 163609 127031 163727
rect 127073 163609 127191 163727
rect 126913 163449 127031 163567
rect 127073 163449 127191 163567
rect 126913 145609 127031 145727
rect 127073 145609 127191 145727
rect 126913 145449 127031 145567
rect 127073 145449 127191 145567
rect 126913 127609 127031 127727
rect 127073 127609 127191 127727
rect 126913 127449 127031 127567
rect 127073 127449 127191 127567
rect 126913 109609 127031 109727
rect 127073 109609 127191 109727
rect 126913 109449 127031 109567
rect 127073 109449 127191 109567
rect 126913 91609 127031 91727
rect 127073 91609 127191 91727
rect 126913 91449 127031 91567
rect 127073 91449 127191 91567
rect 126913 73609 127031 73727
rect 127073 73609 127191 73727
rect 126913 73449 127031 73567
rect 127073 73449 127191 73567
rect 126913 55609 127031 55727
rect 127073 55609 127191 55727
rect 126913 55449 127031 55567
rect 127073 55449 127191 55567
rect 126913 37609 127031 37727
rect 127073 37609 127191 37727
rect 126913 37449 127031 37567
rect 127073 37449 127191 37567
rect 126913 19609 127031 19727
rect 127073 19609 127191 19727
rect 126913 19449 127031 19567
rect 127073 19449 127191 19567
rect 126913 1609 127031 1727
rect 127073 1609 127191 1727
rect 126913 1449 127031 1567
rect 127073 1449 127191 1567
rect 126913 -291 127031 -173
rect 127073 -291 127191 -173
rect 126913 -451 127031 -333
rect 127073 -451 127191 -333
rect 128773 345469 128891 345587
rect 128933 345469 129051 345587
rect 128773 345309 128891 345427
rect 128933 345309 129051 345427
rect 128773 327469 128891 327587
rect 128933 327469 129051 327587
rect 128773 327309 128891 327427
rect 128933 327309 129051 327427
rect 128773 309469 128891 309587
rect 128933 309469 129051 309587
rect 128773 309309 128891 309427
rect 128933 309309 129051 309427
rect 128773 291469 128891 291587
rect 128933 291469 129051 291587
rect 128773 291309 128891 291427
rect 128933 291309 129051 291427
rect 128773 273469 128891 273587
rect 128933 273469 129051 273587
rect 128773 273309 128891 273427
rect 128933 273309 129051 273427
rect 128773 255469 128891 255587
rect 128933 255469 129051 255587
rect 128773 255309 128891 255427
rect 128933 255309 129051 255427
rect 128773 237469 128891 237587
rect 128933 237469 129051 237587
rect 128773 237309 128891 237427
rect 128933 237309 129051 237427
rect 128773 219469 128891 219587
rect 128933 219469 129051 219587
rect 128773 219309 128891 219427
rect 128933 219309 129051 219427
rect 128773 201469 128891 201587
rect 128933 201469 129051 201587
rect 128773 201309 128891 201427
rect 128933 201309 129051 201427
rect 128773 183469 128891 183587
rect 128933 183469 129051 183587
rect 128773 183309 128891 183427
rect 128933 183309 129051 183427
rect 128773 165469 128891 165587
rect 128933 165469 129051 165587
rect 128773 165309 128891 165427
rect 128933 165309 129051 165427
rect 128773 147469 128891 147587
rect 128933 147469 129051 147587
rect 128773 147309 128891 147427
rect 128933 147309 129051 147427
rect 128773 129469 128891 129587
rect 128933 129469 129051 129587
rect 128773 129309 128891 129427
rect 128933 129309 129051 129427
rect 128773 111469 128891 111587
rect 128933 111469 129051 111587
rect 128773 111309 128891 111427
rect 128933 111309 129051 111427
rect 128773 93469 128891 93587
rect 128933 93469 129051 93587
rect 128773 93309 128891 93427
rect 128933 93309 129051 93427
rect 128773 75469 128891 75587
rect 128933 75469 129051 75587
rect 128773 75309 128891 75427
rect 128933 75309 129051 75427
rect 128773 57469 128891 57587
rect 128933 57469 129051 57587
rect 128773 57309 128891 57427
rect 128933 57309 129051 57427
rect 128773 39469 128891 39587
rect 128933 39469 129051 39587
rect 128773 39309 128891 39427
rect 128933 39309 129051 39427
rect 128773 21469 128891 21587
rect 128933 21469 129051 21587
rect 128773 21309 128891 21427
rect 128933 21309 129051 21427
rect 128773 3469 128891 3587
rect 128933 3469 129051 3587
rect 128773 3309 128891 3427
rect 128933 3309 129051 3427
rect 128773 -1251 128891 -1133
rect 128933 -1251 129051 -1133
rect 128773 -1411 128891 -1293
rect 128933 -1411 129051 -1293
rect 130633 347329 130751 347447
rect 130793 347329 130911 347447
rect 130633 347169 130751 347287
rect 130793 347169 130911 347287
rect 130633 329329 130751 329447
rect 130793 329329 130911 329447
rect 130633 329169 130751 329287
rect 130793 329169 130911 329287
rect 130633 311329 130751 311447
rect 130793 311329 130911 311447
rect 130633 311169 130751 311287
rect 130793 311169 130911 311287
rect 130633 293329 130751 293447
rect 130793 293329 130911 293447
rect 130633 293169 130751 293287
rect 130793 293169 130911 293287
rect 130633 275329 130751 275447
rect 130793 275329 130911 275447
rect 130633 275169 130751 275287
rect 130793 275169 130911 275287
rect 130633 257329 130751 257447
rect 130793 257329 130911 257447
rect 130633 257169 130751 257287
rect 130793 257169 130911 257287
rect 130633 239329 130751 239447
rect 130793 239329 130911 239447
rect 130633 239169 130751 239287
rect 130793 239169 130911 239287
rect 130633 221329 130751 221447
rect 130793 221329 130911 221447
rect 130633 221169 130751 221287
rect 130793 221169 130911 221287
rect 130633 203329 130751 203447
rect 130793 203329 130911 203447
rect 130633 203169 130751 203287
rect 130793 203169 130911 203287
rect 130633 185329 130751 185447
rect 130793 185329 130911 185447
rect 130633 185169 130751 185287
rect 130793 185169 130911 185287
rect 130633 167329 130751 167447
rect 130793 167329 130911 167447
rect 130633 167169 130751 167287
rect 130793 167169 130911 167287
rect 130633 149329 130751 149447
rect 130793 149329 130911 149447
rect 130633 149169 130751 149287
rect 130793 149169 130911 149287
rect 130633 131329 130751 131447
rect 130793 131329 130911 131447
rect 130633 131169 130751 131287
rect 130793 131169 130911 131287
rect 130633 113329 130751 113447
rect 130793 113329 130911 113447
rect 130633 113169 130751 113287
rect 130793 113169 130911 113287
rect 130633 95329 130751 95447
rect 130793 95329 130911 95447
rect 130633 95169 130751 95287
rect 130793 95169 130911 95287
rect 130633 77329 130751 77447
rect 130793 77329 130911 77447
rect 130633 77169 130751 77287
rect 130793 77169 130911 77287
rect 130633 59329 130751 59447
rect 130793 59329 130911 59447
rect 130633 59169 130751 59287
rect 130793 59169 130911 59287
rect 130633 41329 130751 41447
rect 130793 41329 130911 41447
rect 130633 41169 130751 41287
rect 130793 41169 130911 41287
rect 130633 23329 130751 23447
rect 130793 23329 130911 23447
rect 130633 23169 130751 23287
rect 130793 23169 130911 23287
rect 130633 5329 130751 5447
rect 130793 5329 130911 5447
rect 130633 5169 130751 5287
rect 130793 5169 130911 5287
rect 130633 -2211 130751 -2093
rect 130793 -2211 130911 -2093
rect 130633 -2371 130751 -2253
rect 130793 -2371 130911 -2253
rect 141493 355661 141611 355779
rect 141653 355661 141771 355779
rect 141493 355501 141611 355619
rect 141653 355501 141771 355619
rect 139633 354701 139751 354819
rect 139793 354701 139911 354819
rect 139633 354541 139751 354659
rect 139793 354541 139911 354659
rect 137773 353741 137891 353859
rect 137933 353741 138051 353859
rect 137773 353581 137891 353699
rect 137933 353581 138051 353699
rect 132493 349189 132611 349307
rect 132653 349189 132771 349307
rect 132493 349029 132611 349147
rect 132653 349029 132771 349147
rect 132493 331189 132611 331307
rect 132653 331189 132771 331307
rect 132493 331029 132611 331147
rect 132653 331029 132771 331147
rect 132493 313189 132611 313307
rect 132653 313189 132771 313307
rect 132493 313029 132611 313147
rect 132653 313029 132771 313147
rect 132493 295189 132611 295307
rect 132653 295189 132771 295307
rect 132493 295029 132611 295147
rect 132653 295029 132771 295147
rect 132493 277189 132611 277307
rect 132653 277189 132771 277307
rect 132493 277029 132611 277147
rect 132653 277029 132771 277147
rect 132493 259189 132611 259307
rect 132653 259189 132771 259307
rect 132493 259029 132611 259147
rect 132653 259029 132771 259147
rect 132493 241189 132611 241307
rect 132653 241189 132771 241307
rect 132493 241029 132611 241147
rect 132653 241029 132771 241147
rect 132493 223189 132611 223307
rect 132653 223189 132771 223307
rect 132493 223029 132611 223147
rect 132653 223029 132771 223147
rect 132493 205189 132611 205307
rect 132653 205189 132771 205307
rect 132493 205029 132611 205147
rect 132653 205029 132771 205147
rect 132493 187189 132611 187307
rect 132653 187189 132771 187307
rect 132493 187029 132611 187147
rect 132653 187029 132771 187147
rect 132493 169189 132611 169307
rect 132653 169189 132771 169307
rect 132493 169029 132611 169147
rect 132653 169029 132771 169147
rect 132493 151189 132611 151307
rect 132653 151189 132771 151307
rect 132493 151029 132611 151147
rect 132653 151029 132771 151147
rect 132493 133189 132611 133307
rect 132653 133189 132771 133307
rect 132493 133029 132611 133147
rect 132653 133029 132771 133147
rect 132493 115189 132611 115307
rect 132653 115189 132771 115307
rect 132493 115029 132611 115147
rect 132653 115029 132771 115147
rect 132493 97189 132611 97307
rect 132653 97189 132771 97307
rect 132493 97029 132611 97147
rect 132653 97029 132771 97147
rect 132493 79189 132611 79307
rect 132653 79189 132771 79307
rect 132493 79029 132611 79147
rect 132653 79029 132771 79147
rect 132493 61189 132611 61307
rect 132653 61189 132771 61307
rect 132493 61029 132611 61147
rect 132653 61029 132771 61147
rect 132493 43189 132611 43307
rect 132653 43189 132771 43307
rect 132493 43029 132611 43147
rect 132653 43029 132771 43147
rect 132493 25189 132611 25307
rect 132653 25189 132771 25307
rect 132493 25029 132611 25147
rect 132653 25029 132771 25147
rect 132493 7189 132611 7307
rect 132653 7189 132771 7307
rect 132493 7029 132611 7147
rect 132653 7029 132771 7147
rect 123493 -3651 123611 -3533
rect 123653 -3651 123771 -3533
rect 123493 -3811 123611 -3693
rect 123653 -3811 123771 -3693
rect 135913 352781 136031 352899
rect 136073 352781 136191 352899
rect 135913 352621 136031 352739
rect 136073 352621 136191 352739
rect 135913 334609 136031 334727
rect 136073 334609 136191 334727
rect 135913 334449 136031 334567
rect 136073 334449 136191 334567
rect 135913 316609 136031 316727
rect 136073 316609 136191 316727
rect 135913 316449 136031 316567
rect 136073 316449 136191 316567
rect 135913 298609 136031 298727
rect 136073 298609 136191 298727
rect 135913 298449 136031 298567
rect 136073 298449 136191 298567
rect 135913 280609 136031 280727
rect 136073 280609 136191 280727
rect 135913 280449 136031 280567
rect 136073 280449 136191 280567
rect 135913 262609 136031 262727
rect 136073 262609 136191 262727
rect 135913 262449 136031 262567
rect 136073 262449 136191 262567
rect 135913 244609 136031 244727
rect 136073 244609 136191 244727
rect 135913 244449 136031 244567
rect 136073 244449 136191 244567
rect 135913 226609 136031 226727
rect 136073 226609 136191 226727
rect 135913 226449 136031 226567
rect 136073 226449 136191 226567
rect 135913 208609 136031 208727
rect 136073 208609 136191 208727
rect 135913 208449 136031 208567
rect 136073 208449 136191 208567
rect 135913 190609 136031 190727
rect 136073 190609 136191 190727
rect 135913 190449 136031 190567
rect 136073 190449 136191 190567
rect 135913 172609 136031 172727
rect 136073 172609 136191 172727
rect 135913 172449 136031 172567
rect 136073 172449 136191 172567
rect 135913 154609 136031 154727
rect 136073 154609 136191 154727
rect 135913 154449 136031 154567
rect 136073 154449 136191 154567
rect 135913 136609 136031 136727
rect 136073 136609 136191 136727
rect 135913 136449 136031 136567
rect 136073 136449 136191 136567
rect 135913 118609 136031 118727
rect 136073 118609 136191 118727
rect 135913 118449 136031 118567
rect 136073 118449 136191 118567
rect 135913 100609 136031 100727
rect 136073 100609 136191 100727
rect 135913 100449 136031 100567
rect 136073 100449 136191 100567
rect 135913 82609 136031 82727
rect 136073 82609 136191 82727
rect 135913 82449 136031 82567
rect 136073 82449 136191 82567
rect 135913 64609 136031 64727
rect 136073 64609 136191 64727
rect 135913 64449 136031 64567
rect 136073 64449 136191 64567
rect 135913 46609 136031 46727
rect 136073 46609 136191 46727
rect 135913 46449 136031 46567
rect 136073 46449 136191 46567
rect 135913 28609 136031 28727
rect 136073 28609 136191 28727
rect 135913 28449 136031 28567
rect 136073 28449 136191 28567
rect 135913 10609 136031 10727
rect 136073 10609 136191 10727
rect 135913 10449 136031 10567
rect 136073 10449 136191 10567
rect 135913 -771 136031 -653
rect 136073 -771 136191 -653
rect 135913 -931 136031 -813
rect 136073 -931 136191 -813
rect 137773 336469 137891 336587
rect 137933 336469 138051 336587
rect 137773 336309 137891 336427
rect 137933 336309 138051 336427
rect 137773 318469 137891 318587
rect 137933 318469 138051 318587
rect 137773 318309 137891 318427
rect 137933 318309 138051 318427
rect 137773 300469 137891 300587
rect 137933 300469 138051 300587
rect 137773 300309 137891 300427
rect 137933 300309 138051 300427
rect 137773 282469 137891 282587
rect 137933 282469 138051 282587
rect 137773 282309 137891 282427
rect 137933 282309 138051 282427
rect 137773 264469 137891 264587
rect 137933 264469 138051 264587
rect 137773 264309 137891 264427
rect 137933 264309 138051 264427
rect 137773 246469 137891 246587
rect 137933 246469 138051 246587
rect 137773 246309 137891 246427
rect 137933 246309 138051 246427
rect 137773 228469 137891 228587
rect 137933 228469 138051 228587
rect 137773 228309 137891 228427
rect 137933 228309 138051 228427
rect 137773 210469 137891 210587
rect 137933 210469 138051 210587
rect 137773 210309 137891 210427
rect 137933 210309 138051 210427
rect 137773 192469 137891 192587
rect 137933 192469 138051 192587
rect 137773 192309 137891 192427
rect 137933 192309 138051 192427
rect 137773 174469 137891 174587
rect 137933 174469 138051 174587
rect 137773 174309 137891 174427
rect 137933 174309 138051 174427
rect 137773 156469 137891 156587
rect 137933 156469 138051 156587
rect 137773 156309 137891 156427
rect 137933 156309 138051 156427
rect 137773 138469 137891 138587
rect 137933 138469 138051 138587
rect 137773 138309 137891 138427
rect 137933 138309 138051 138427
rect 137773 120469 137891 120587
rect 137933 120469 138051 120587
rect 137773 120309 137891 120427
rect 137933 120309 138051 120427
rect 137773 102469 137891 102587
rect 137933 102469 138051 102587
rect 137773 102309 137891 102427
rect 137933 102309 138051 102427
rect 137773 84469 137891 84587
rect 137933 84469 138051 84587
rect 137773 84309 137891 84427
rect 137933 84309 138051 84427
rect 137773 66469 137891 66587
rect 137933 66469 138051 66587
rect 137773 66309 137891 66427
rect 137933 66309 138051 66427
rect 137773 48469 137891 48587
rect 137933 48469 138051 48587
rect 137773 48309 137891 48427
rect 137933 48309 138051 48427
rect 137773 30469 137891 30587
rect 137933 30469 138051 30587
rect 137773 30309 137891 30427
rect 137933 30309 138051 30427
rect 137773 12469 137891 12587
rect 137933 12469 138051 12587
rect 137773 12309 137891 12427
rect 137933 12309 138051 12427
rect 137773 -1731 137891 -1613
rect 137933 -1731 138051 -1613
rect 137773 -1891 137891 -1773
rect 137933 -1891 138051 -1773
rect 139633 338329 139751 338447
rect 139793 338329 139911 338447
rect 139633 338169 139751 338287
rect 139793 338169 139911 338287
rect 139633 320329 139751 320447
rect 139793 320329 139911 320447
rect 139633 320169 139751 320287
rect 139793 320169 139911 320287
rect 139633 302329 139751 302447
rect 139793 302329 139911 302447
rect 139633 302169 139751 302287
rect 139793 302169 139911 302287
rect 139633 284329 139751 284447
rect 139793 284329 139911 284447
rect 139633 284169 139751 284287
rect 139793 284169 139911 284287
rect 139633 266329 139751 266447
rect 139793 266329 139911 266447
rect 139633 266169 139751 266287
rect 139793 266169 139911 266287
rect 139633 248329 139751 248447
rect 139793 248329 139911 248447
rect 139633 248169 139751 248287
rect 139793 248169 139911 248287
rect 139633 230329 139751 230447
rect 139793 230329 139911 230447
rect 139633 230169 139751 230287
rect 139793 230169 139911 230287
rect 139633 212329 139751 212447
rect 139793 212329 139911 212447
rect 139633 212169 139751 212287
rect 139793 212169 139911 212287
rect 139633 194329 139751 194447
rect 139793 194329 139911 194447
rect 139633 194169 139751 194287
rect 139793 194169 139911 194287
rect 139633 176329 139751 176447
rect 139793 176329 139911 176447
rect 139633 176169 139751 176287
rect 139793 176169 139911 176287
rect 139633 158329 139751 158447
rect 139793 158329 139911 158447
rect 139633 158169 139751 158287
rect 139793 158169 139911 158287
rect 139633 140329 139751 140447
rect 139793 140329 139911 140447
rect 139633 140169 139751 140287
rect 139793 140169 139911 140287
rect 139633 122329 139751 122447
rect 139793 122329 139911 122447
rect 139633 122169 139751 122287
rect 139793 122169 139911 122287
rect 139633 104329 139751 104447
rect 139793 104329 139911 104447
rect 139633 104169 139751 104287
rect 139793 104169 139911 104287
rect 139633 86329 139751 86447
rect 139793 86329 139911 86447
rect 139633 86169 139751 86287
rect 139793 86169 139911 86287
rect 139633 68329 139751 68447
rect 139793 68329 139911 68447
rect 139633 68169 139751 68287
rect 139793 68169 139911 68287
rect 139633 50329 139751 50447
rect 139793 50329 139911 50447
rect 139633 50169 139751 50287
rect 139793 50169 139911 50287
rect 139633 32329 139751 32447
rect 139793 32329 139911 32447
rect 139633 32169 139751 32287
rect 139793 32169 139911 32287
rect 139633 14329 139751 14447
rect 139793 14329 139911 14447
rect 139633 14169 139751 14287
rect 139793 14169 139911 14287
rect 139633 -2691 139751 -2573
rect 139793 -2691 139911 -2573
rect 139633 -2851 139751 -2733
rect 139793 -2851 139911 -2733
rect 150493 355181 150611 355299
rect 150653 355181 150771 355299
rect 150493 355021 150611 355139
rect 150653 355021 150771 355139
rect 148633 354221 148751 354339
rect 148793 354221 148911 354339
rect 148633 354061 148751 354179
rect 148793 354061 148911 354179
rect 146773 353261 146891 353379
rect 146933 353261 147051 353379
rect 146773 353101 146891 353219
rect 146933 353101 147051 353219
rect 141493 340189 141611 340307
rect 141653 340189 141771 340307
rect 141493 340029 141611 340147
rect 141653 340029 141771 340147
rect 141493 322189 141611 322307
rect 141653 322189 141771 322307
rect 141493 322029 141611 322147
rect 141653 322029 141771 322147
rect 141493 304189 141611 304307
rect 141653 304189 141771 304307
rect 141493 304029 141611 304147
rect 141653 304029 141771 304147
rect 141493 286189 141611 286307
rect 141653 286189 141771 286307
rect 141493 286029 141611 286147
rect 141653 286029 141771 286147
rect 141493 268189 141611 268307
rect 141653 268189 141771 268307
rect 141493 268029 141611 268147
rect 141653 268029 141771 268147
rect 141493 250189 141611 250307
rect 141653 250189 141771 250307
rect 141493 250029 141611 250147
rect 141653 250029 141771 250147
rect 141493 232189 141611 232307
rect 141653 232189 141771 232307
rect 141493 232029 141611 232147
rect 141653 232029 141771 232147
rect 141493 214189 141611 214307
rect 141653 214189 141771 214307
rect 141493 214029 141611 214147
rect 141653 214029 141771 214147
rect 141493 196189 141611 196307
rect 141653 196189 141771 196307
rect 141493 196029 141611 196147
rect 141653 196029 141771 196147
rect 141493 178189 141611 178307
rect 141653 178189 141771 178307
rect 141493 178029 141611 178147
rect 141653 178029 141771 178147
rect 141493 160189 141611 160307
rect 141653 160189 141771 160307
rect 141493 160029 141611 160147
rect 141653 160029 141771 160147
rect 141493 142189 141611 142307
rect 141653 142189 141771 142307
rect 141493 142029 141611 142147
rect 141653 142029 141771 142147
rect 141493 124189 141611 124307
rect 141653 124189 141771 124307
rect 141493 124029 141611 124147
rect 141653 124029 141771 124147
rect 141493 106189 141611 106307
rect 141653 106189 141771 106307
rect 141493 106029 141611 106147
rect 141653 106029 141771 106147
rect 141493 88189 141611 88307
rect 141653 88189 141771 88307
rect 141493 88029 141611 88147
rect 141653 88029 141771 88147
rect 141493 70189 141611 70307
rect 141653 70189 141771 70307
rect 141493 70029 141611 70147
rect 141653 70029 141771 70147
rect 141493 52189 141611 52307
rect 141653 52189 141771 52307
rect 141493 52029 141611 52147
rect 141653 52029 141771 52147
rect 141493 34189 141611 34307
rect 141653 34189 141771 34307
rect 141493 34029 141611 34147
rect 141653 34029 141771 34147
rect 141493 16189 141611 16307
rect 141653 16189 141771 16307
rect 141493 16029 141611 16147
rect 141653 16029 141771 16147
rect 132493 -3171 132611 -3053
rect 132653 -3171 132771 -3053
rect 132493 -3331 132611 -3213
rect 132653 -3331 132771 -3213
rect 144913 352301 145031 352419
rect 145073 352301 145191 352419
rect 144913 352141 145031 352259
rect 145073 352141 145191 352259
rect 144913 343609 145031 343727
rect 145073 343609 145191 343727
rect 144913 343449 145031 343567
rect 145073 343449 145191 343567
rect 144913 325609 145031 325727
rect 145073 325609 145191 325727
rect 144913 325449 145031 325567
rect 145073 325449 145191 325567
rect 144913 307609 145031 307727
rect 145073 307609 145191 307727
rect 144913 307449 145031 307567
rect 145073 307449 145191 307567
rect 144913 289609 145031 289727
rect 145073 289609 145191 289727
rect 144913 289449 145031 289567
rect 145073 289449 145191 289567
rect 144913 271609 145031 271727
rect 145073 271609 145191 271727
rect 144913 271449 145031 271567
rect 145073 271449 145191 271567
rect 144913 253609 145031 253727
rect 145073 253609 145191 253727
rect 144913 253449 145031 253567
rect 145073 253449 145191 253567
rect 144913 235609 145031 235727
rect 145073 235609 145191 235727
rect 144913 235449 145031 235567
rect 145073 235449 145191 235567
rect 144913 217609 145031 217727
rect 145073 217609 145191 217727
rect 144913 217449 145031 217567
rect 145073 217449 145191 217567
rect 144913 199609 145031 199727
rect 145073 199609 145191 199727
rect 144913 199449 145031 199567
rect 145073 199449 145191 199567
rect 144913 181609 145031 181727
rect 145073 181609 145191 181727
rect 144913 181449 145031 181567
rect 145073 181449 145191 181567
rect 144913 163609 145031 163727
rect 145073 163609 145191 163727
rect 144913 163449 145031 163567
rect 145073 163449 145191 163567
rect 144913 145609 145031 145727
rect 145073 145609 145191 145727
rect 144913 145449 145031 145567
rect 145073 145449 145191 145567
rect 144913 127609 145031 127727
rect 145073 127609 145191 127727
rect 144913 127449 145031 127567
rect 145073 127449 145191 127567
rect 144913 109609 145031 109727
rect 145073 109609 145191 109727
rect 144913 109449 145031 109567
rect 145073 109449 145191 109567
rect 144913 91609 145031 91727
rect 145073 91609 145191 91727
rect 144913 91449 145031 91567
rect 145073 91449 145191 91567
rect 144913 73609 145031 73727
rect 145073 73609 145191 73727
rect 144913 73449 145031 73567
rect 145073 73449 145191 73567
rect 144913 55609 145031 55727
rect 145073 55609 145191 55727
rect 144913 55449 145031 55567
rect 145073 55449 145191 55567
rect 144913 37609 145031 37727
rect 145073 37609 145191 37727
rect 144913 37449 145031 37567
rect 145073 37449 145191 37567
rect 144913 19609 145031 19727
rect 145073 19609 145191 19727
rect 144913 19449 145031 19567
rect 145073 19449 145191 19567
rect 144913 1609 145031 1727
rect 145073 1609 145191 1727
rect 144913 1449 145031 1567
rect 145073 1449 145191 1567
rect 144913 -291 145031 -173
rect 145073 -291 145191 -173
rect 144913 -451 145031 -333
rect 145073 -451 145191 -333
rect 146773 345469 146891 345587
rect 146933 345469 147051 345587
rect 146773 345309 146891 345427
rect 146933 345309 147051 345427
rect 146773 327469 146891 327587
rect 146933 327469 147051 327587
rect 146773 327309 146891 327427
rect 146933 327309 147051 327427
rect 146773 309469 146891 309587
rect 146933 309469 147051 309587
rect 146773 309309 146891 309427
rect 146933 309309 147051 309427
rect 146773 291469 146891 291587
rect 146933 291469 147051 291587
rect 146773 291309 146891 291427
rect 146933 291309 147051 291427
rect 146773 273469 146891 273587
rect 146933 273469 147051 273587
rect 146773 273309 146891 273427
rect 146933 273309 147051 273427
rect 146773 255469 146891 255587
rect 146933 255469 147051 255587
rect 146773 255309 146891 255427
rect 146933 255309 147051 255427
rect 146773 237469 146891 237587
rect 146933 237469 147051 237587
rect 146773 237309 146891 237427
rect 146933 237309 147051 237427
rect 146773 219469 146891 219587
rect 146933 219469 147051 219587
rect 146773 219309 146891 219427
rect 146933 219309 147051 219427
rect 146773 201469 146891 201587
rect 146933 201469 147051 201587
rect 146773 201309 146891 201427
rect 146933 201309 147051 201427
rect 146773 183469 146891 183587
rect 146933 183469 147051 183587
rect 146773 183309 146891 183427
rect 146933 183309 147051 183427
rect 146773 165469 146891 165587
rect 146933 165469 147051 165587
rect 146773 165309 146891 165427
rect 146933 165309 147051 165427
rect 146773 147469 146891 147587
rect 146933 147469 147051 147587
rect 146773 147309 146891 147427
rect 146933 147309 147051 147427
rect 146773 129469 146891 129587
rect 146933 129469 147051 129587
rect 146773 129309 146891 129427
rect 146933 129309 147051 129427
rect 146773 111469 146891 111587
rect 146933 111469 147051 111587
rect 146773 111309 146891 111427
rect 146933 111309 147051 111427
rect 146773 93469 146891 93587
rect 146933 93469 147051 93587
rect 146773 93309 146891 93427
rect 146933 93309 147051 93427
rect 146773 75469 146891 75587
rect 146933 75469 147051 75587
rect 146773 75309 146891 75427
rect 146933 75309 147051 75427
rect 146773 57469 146891 57587
rect 146933 57469 147051 57587
rect 146773 57309 146891 57427
rect 146933 57309 147051 57427
rect 146773 39469 146891 39587
rect 146933 39469 147051 39587
rect 146773 39309 146891 39427
rect 146933 39309 147051 39427
rect 146773 21469 146891 21587
rect 146933 21469 147051 21587
rect 146773 21309 146891 21427
rect 146933 21309 147051 21427
rect 146773 3469 146891 3587
rect 146933 3469 147051 3587
rect 146773 3309 146891 3427
rect 146933 3309 147051 3427
rect 146773 -1251 146891 -1133
rect 146933 -1251 147051 -1133
rect 146773 -1411 146891 -1293
rect 146933 -1411 147051 -1293
rect 148633 347329 148751 347447
rect 148793 347329 148911 347447
rect 148633 347169 148751 347287
rect 148793 347169 148911 347287
rect 148633 329329 148751 329447
rect 148793 329329 148911 329447
rect 148633 329169 148751 329287
rect 148793 329169 148911 329287
rect 148633 311329 148751 311447
rect 148793 311329 148911 311447
rect 148633 311169 148751 311287
rect 148793 311169 148911 311287
rect 148633 293329 148751 293447
rect 148793 293329 148911 293447
rect 148633 293169 148751 293287
rect 148793 293169 148911 293287
rect 148633 275329 148751 275447
rect 148793 275329 148911 275447
rect 148633 275169 148751 275287
rect 148793 275169 148911 275287
rect 148633 257329 148751 257447
rect 148793 257329 148911 257447
rect 148633 257169 148751 257287
rect 148793 257169 148911 257287
rect 148633 239329 148751 239447
rect 148793 239329 148911 239447
rect 148633 239169 148751 239287
rect 148793 239169 148911 239287
rect 148633 221329 148751 221447
rect 148793 221329 148911 221447
rect 148633 221169 148751 221287
rect 148793 221169 148911 221287
rect 148633 203329 148751 203447
rect 148793 203329 148911 203447
rect 148633 203169 148751 203287
rect 148793 203169 148911 203287
rect 148633 185329 148751 185447
rect 148793 185329 148911 185447
rect 148633 185169 148751 185287
rect 148793 185169 148911 185287
rect 148633 167329 148751 167447
rect 148793 167329 148911 167447
rect 148633 167169 148751 167287
rect 148793 167169 148911 167287
rect 148633 149329 148751 149447
rect 148793 149329 148911 149447
rect 148633 149169 148751 149287
rect 148793 149169 148911 149287
rect 148633 131329 148751 131447
rect 148793 131329 148911 131447
rect 148633 131169 148751 131287
rect 148793 131169 148911 131287
rect 148633 113329 148751 113447
rect 148793 113329 148911 113447
rect 148633 113169 148751 113287
rect 148793 113169 148911 113287
rect 148633 95329 148751 95447
rect 148793 95329 148911 95447
rect 148633 95169 148751 95287
rect 148793 95169 148911 95287
rect 148633 77329 148751 77447
rect 148793 77329 148911 77447
rect 148633 77169 148751 77287
rect 148793 77169 148911 77287
rect 148633 59329 148751 59447
rect 148793 59329 148911 59447
rect 148633 59169 148751 59287
rect 148793 59169 148911 59287
rect 148633 41329 148751 41447
rect 148793 41329 148911 41447
rect 148633 41169 148751 41287
rect 148793 41169 148911 41287
rect 148633 23329 148751 23447
rect 148793 23329 148911 23447
rect 148633 23169 148751 23287
rect 148793 23169 148911 23287
rect 148633 5329 148751 5447
rect 148793 5329 148911 5447
rect 148633 5169 148751 5287
rect 148793 5169 148911 5287
rect 148633 -2211 148751 -2093
rect 148793 -2211 148911 -2093
rect 148633 -2371 148751 -2253
rect 148793 -2371 148911 -2253
rect 159493 355661 159611 355779
rect 159653 355661 159771 355779
rect 159493 355501 159611 355619
rect 159653 355501 159771 355619
rect 157633 354701 157751 354819
rect 157793 354701 157911 354819
rect 157633 354541 157751 354659
rect 157793 354541 157911 354659
rect 155773 353741 155891 353859
rect 155933 353741 156051 353859
rect 155773 353581 155891 353699
rect 155933 353581 156051 353699
rect 150493 349189 150611 349307
rect 150653 349189 150771 349307
rect 150493 349029 150611 349147
rect 150653 349029 150771 349147
rect 150493 331189 150611 331307
rect 150653 331189 150771 331307
rect 150493 331029 150611 331147
rect 150653 331029 150771 331147
rect 150493 313189 150611 313307
rect 150653 313189 150771 313307
rect 150493 313029 150611 313147
rect 150653 313029 150771 313147
rect 150493 295189 150611 295307
rect 150653 295189 150771 295307
rect 150493 295029 150611 295147
rect 150653 295029 150771 295147
rect 150493 277189 150611 277307
rect 150653 277189 150771 277307
rect 150493 277029 150611 277147
rect 150653 277029 150771 277147
rect 150493 259189 150611 259307
rect 150653 259189 150771 259307
rect 150493 259029 150611 259147
rect 150653 259029 150771 259147
rect 150493 241189 150611 241307
rect 150653 241189 150771 241307
rect 150493 241029 150611 241147
rect 150653 241029 150771 241147
rect 150493 223189 150611 223307
rect 150653 223189 150771 223307
rect 150493 223029 150611 223147
rect 150653 223029 150771 223147
rect 150493 205189 150611 205307
rect 150653 205189 150771 205307
rect 150493 205029 150611 205147
rect 150653 205029 150771 205147
rect 150493 187189 150611 187307
rect 150653 187189 150771 187307
rect 150493 187029 150611 187147
rect 150653 187029 150771 187147
rect 150493 169189 150611 169307
rect 150653 169189 150771 169307
rect 150493 169029 150611 169147
rect 150653 169029 150771 169147
rect 150493 151189 150611 151307
rect 150653 151189 150771 151307
rect 150493 151029 150611 151147
rect 150653 151029 150771 151147
rect 150493 133189 150611 133307
rect 150653 133189 150771 133307
rect 150493 133029 150611 133147
rect 150653 133029 150771 133147
rect 150493 115189 150611 115307
rect 150653 115189 150771 115307
rect 150493 115029 150611 115147
rect 150653 115029 150771 115147
rect 150493 97189 150611 97307
rect 150653 97189 150771 97307
rect 150493 97029 150611 97147
rect 150653 97029 150771 97147
rect 150493 79189 150611 79307
rect 150653 79189 150771 79307
rect 150493 79029 150611 79147
rect 150653 79029 150771 79147
rect 150493 61189 150611 61307
rect 150653 61189 150771 61307
rect 150493 61029 150611 61147
rect 150653 61029 150771 61147
rect 150493 43189 150611 43307
rect 150653 43189 150771 43307
rect 150493 43029 150611 43147
rect 150653 43029 150771 43147
rect 150493 25189 150611 25307
rect 150653 25189 150771 25307
rect 150493 25029 150611 25147
rect 150653 25029 150771 25147
rect 150493 7189 150611 7307
rect 150653 7189 150771 7307
rect 150493 7029 150611 7147
rect 150653 7029 150771 7147
rect 141493 -3651 141611 -3533
rect 141653 -3651 141771 -3533
rect 141493 -3811 141611 -3693
rect 141653 -3811 141771 -3693
rect 153913 352781 154031 352899
rect 154073 352781 154191 352899
rect 153913 352621 154031 352739
rect 154073 352621 154191 352739
rect 153913 334609 154031 334727
rect 154073 334609 154191 334727
rect 153913 334449 154031 334567
rect 154073 334449 154191 334567
rect 153913 316609 154031 316727
rect 154073 316609 154191 316727
rect 153913 316449 154031 316567
rect 154073 316449 154191 316567
rect 153913 298609 154031 298727
rect 154073 298609 154191 298727
rect 153913 298449 154031 298567
rect 154073 298449 154191 298567
rect 153913 280609 154031 280727
rect 154073 280609 154191 280727
rect 153913 280449 154031 280567
rect 154073 280449 154191 280567
rect 153913 262609 154031 262727
rect 154073 262609 154191 262727
rect 153913 262449 154031 262567
rect 154073 262449 154191 262567
rect 153913 244609 154031 244727
rect 154073 244609 154191 244727
rect 153913 244449 154031 244567
rect 154073 244449 154191 244567
rect 153913 226609 154031 226727
rect 154073 226609 154191 226727
rect 153913 226449 154031 226567
rect 154073 226449 154191 226567
rect 153913 208609 154031 208727
rect 154073 208609 154191 208727
rect 153913 208449 154031 208567
rect 154073 208449 154191 208567
rect 153913 190609 154031 190727
rect 154073 190609 154191 190727
rect 153913 190449 154031 190567
rect 154073 190449 154191 190567
rect 153913 172609 154031 172727
rect 154073 172609 154191 172727
rect 153913 172449 154031 172567
rect 154073 172449 154191 172567
rect 153913 154609 154031 154727
rect 154073 154609 154191 154727
rect 153913 154449 154031 154567
rect 154073 154449 154191 154567
rect 153913 136609 154031 136727
rect 154073 136609 154191 136727
rect 153913 136449 154031 136567
rect 154073 136449 154191 136567
rect 153913 118609 154031 118727
rect 154073 118609 154191 118727
rect 153913 118449 154031 118567
rect 154073 118449 154191 118567
rect 153913 100609 154031 100727
rect 154073 100609 154191 100727
rect 153913 100449 154031 100567
rect 154073 100449 154191 100567
rect 153913 82609 154031 82727
rect 154073 82609 154191 82727
rect 153913 82449 154031 82567
rect 154073 82449 154191 82567
rect 153913 64609 154031 64727
rect 154073 64609 154191 64727
rect 153913 64449 154031 64567
rect 154073 64449 154191 64567
rect 153913 46609 154031 46727
rect 154073 46609 154191 46727
rect 153913 46449 154031 46567
rect 154073 46449 154191 46567
rect 153913 28609 154031 28727
rect 154073 28609 154191 28727
rect 153913 28449 154031 28567
rect 154073 28449 154191 28567
rect 153913 10609 154031 10727
rect 154073 10609 154191 10727
rect 153913 10449 154031 10567
rect 154073 10449 154191 10567
rect 153913 -771 154031 -653
rect 154073 -771 154191 -653
rect 153913 -931 154031 -813
rect 154073 -931 154191 -813
rect 155773 336469 155891 336587
rect 155933 336469 156051 336587
rect 155773 336309 155891 336427
rect 155933 336309 156051 336427
rect 155773 318469 155891 318587
rect 155933 318469 156051 318587
rect 155773 318309 155891 318427
rect 155933 318309 156051 318427
rect 155773 300469 155891 300587
rect 155933 300469 156051 300587
rect 155773 300309 155891 300427
rect 155933 300309 156051 300427
rect 155773 282469 155891 282587
rect 155933 282469 156051 282587
rect 155773 282309 155891 282427
rect 155933 282309 156051 282427
rect 155773 264469 155891 264587
rect 155933 264469 156051 264587
rect 155773 264309 155891 264427
rect 155933 264309 156051 264427
rect 155773 246469 155891 246587
rect 155933 246469 156051 246587
rect 155773 246309 155891 246427
rect 155933 246309 156051 246427
rect 155773 228469 155891 228587
rect 155933 228469 156051 228587
rect 155773 228309 155891 228427
rect 155933 228309 156051 228427
rect 155773 210469 155891 210587
rect 155933 210469 156051 210587
rect 155773 210309 155891 210427
rect 155933 210309 156051 210427
rect 155773 192469 155891 192587
rect 155933 192469 156051 192587
rect 155773 192309 155891 192427
rect 155933 192309 156051 192427
rect 155773 174469 155891 174587
rect 155933 174469 156051 174587
rect 155773 174309 155891 174427
rect 155933 174309 156051 174427
rect 155773 156469 155891 156587
rect 155933 156469 156051 156587
rect 155773 156309 155891 156427
rect 155933 156309 156051 156427
rect 155773 138469 155891 138587
rect 155933 138469 156051 138587
rect 155773 138309 155891 138427
rect 155933 138309 156051 138427
rect 155773 120469 155891 120587
rect 155933 120469 156051 120587
rect 155773 120309 155891 120427
rect 155933 120309 156051 120427
rect 155773 102469 155891 102587
rect 155933 102469 156051 102587
rect 155773 102309 155891 102427
rect 155933 102309 156051 102427
rect 155773 84469 155891 84587
rect 155933 84469 156051 84587
rect 155773 84309 155891 84427
rect 155933 84309 156051 84427
rect 155773 66469 155891 66587
rect 155933 66469 156051 66587
rect 155773 66309 155891 66427
rect 155933 66309 156051 66427
rect 155773 48469 155891 48587
rect 155933 48469 156051 48587
rect 155773 48309 155891 48427
rect 155933 48309 156051 48427
rect 155773 30469 155891 30587
rect 155933 30469 156051 30587
rect 155773 30309 155891 30427
rect 155933 30309 156051 30427
rect 155773 12469 155891 12587
rect 155933 12469 156051 12587
rect 155773 12309 155891 12427
rect 155933 12309 156051 12427
rect 155773 -1731 155891 -1613
rect 155933 -1731 156051 -1613
rect 155773 -1891 155891 -1773
rect 155933 -1891 156051 -1773
rect 157633 338329 157751 338447
rect 157793 338329 157911 338447
rect 157633 338169 157751 338287
rect 157793 338169 157911 338287
rect 157633 320329 157751 320447
rect 157793 320329 157911 320447
rect 157633 320169 157751 320287
rect 157793 320169 157911 320287
rect 157633 302329 157751 302447
rect 157793 302329 157911 302447
rect 157633 302169 157751 302287
rect 157793 302169 157911 302287
rect 157633 284329 157751 284447
rect 157793 284329 157911 284447
rect 157633 284169 157751 284287
rect 157793 284169 157911 284287
rect 157633 266329 157751 266447
rect 157793 266329 157911 266447
rect 157633 266169 157751 266287
rect 157793 266169 157911 266287
rect 157633 248329 157751 248447
rect 157793 248329 157911 248447
rect 157633 248169 157751 248287
rect 157793 248169 157911 248287
rect 157633 230329 157751 230447
rect 157793 230329 157911 230447
rect 157633 230169 157751 230287
rect 157793 230169 157911 230287
rect 157633 212329 157751 212447
rect 157793 212329 157911 212447
rect 157633 212169 157751 212287
rect 157793 212169 157911 212287
rect 157633 194329 157751 194447
rect 157793 194329 157911 194447
rect 157633 194169 157751 194287
rect 157793 194169 157911 194287
rect 157633 176329 157751 176447
rect 157793 176329 157911 176447
rect 157633 176169 157751 176287
rect 157793 176169 157911 176287
rect 157633 158329 157751 158447
rect 157793 158329 157911 158447
rect 157633 158169 157751 158287
rect 157793 158169 157911 158287
rect 157633 140329 157751 140447
rect 157793 140329 157911 140447
rect 157633 140169 157751 140287
rect 157793 140169 157911 140287
rect 157633 122329 157751 122447
rect 157793 122329 157911 122447
rect 157633 122169 157751 122287
rect 157793 122169 157911 122287
rect 157633 104329 157751 104447
rect 157793 104329 157911 104447
rect 157633 104169 157751 104287
rect 157793 104169 157911 104287
rect 157633 86329 157751 86447
rect 157793 86329 157911 86447
rect 157633 86169 157751 86287
rect 157793 86169 157911 86287
rect 157633 68329 157751 68447
rect 157793 68329 157911 68447
rect 157633 68169 157751 68287
rect 157793 68169 157911 68287
rect 157633 50329 157751 50447
rect 157793 50329 157911 50447
rect 157633 50169 157751 50287
rect 157793 50169 157911 50287
rect 157633 32329 157751 32447
rect 157793 32329 157911 32447
rect 157633 32169 157751 32287
rect 157793 32169 157911 32287
rect 157633 14329 157751 14447
rect 157793 14329 157911 14447
rect 157633 14169 157751 14287
rect 157793 14169 157911 14287
rect 157633 -2691 157751 -2573
rect 157793 -2691 157911 -2573
rect 157633 -2851 157751 -2733
rect 157793 -2851 157911 -2733
rect 168493 355181 168611 355299
rect 168653 355181 168771 355299
rect 168493 355021 168611 355139
rect 168653 355021 168771 355139
rect 166633 354221 166751 354339
rect 166793 354221 166911 354339
rect 166633 354061 166751 354179
rect 166793 354061 166911 354179
rect 164773 353261 164891 353379
rect 164933 353261 165051 353379
rect 164773 353101 164891 353219
rect 164933 353101 165051 353219
rect 159493 340189 159611 340307
rect 159653 340189 159771 340307
rect 159493 340029 159611 340147
rect 159653 340029 159771 340147
rect 159493 322189 159611 322307
rect 159653 322189 159771 322307
rect 159493 322029 159611 322147
rect 159653 322029 159771 322147
rect 159493 304189 159611 304307
rect 159653 304189 159771 304307
rect 159493 304029 159611 304147
rect 159653 304029 159771 304147
rect 159493 286189 159611 286307
rect 159653 286189 159771 286307
rect 159493 286029 159611 286147
rect 159653 286029 159771 286147
rect 159493 268189 159611 268307
rect 159653 268189 159771 268307
rect 159493 268029 159611 268147
rect 159653 268029 159771 268147
rect 159493 250189 159611 250307
rect 159653 250189 159771 250307
rect 159493 250029 159611 250147
rect 159653 250029 159771 250147
rect 159493 232189 159611 232307
rect 159653 232189 159771 232307
rect 159493 232029 159611 232147
rect 159653 232029 159771 232147
rect 159493 214189 159611 214307
rect 159653 214189 159771 214307
rect 159493 214029 159611 214147
rect 159653 214029 159771 214147
rect 159493 196189 159611 196307
rect 159653 196189 159771 196307
rect 159493 196029 159611 196147
rect 159653 196029 159771 196147
rect 159493 178189 159611 178307
rect 159653 178189 159771 178307
rect 159493 178029 159611 178147
rect 159653 178029 159771 178147
rect 159493 160189 159611 160307
rect 159653 160189 159771 160307
rect 159493 160029 159611 160147
rect 159653 160029 159771 160147
rect 159493 142189 159611 142307
rect 159653 142189 159771 142307
rect 159493 142029 159611 142147
rect 159653 142029 159771 142147
rect 159493 124189 159611 124307
rect 159653 124189 159771 124307
rect 159493 124029 159611 124147
rect 159653 124029 159771 124147
rect 159493 106189 159611 106307
rect 159653 106189 159771 106307
rect 159493 106029 159611 106147
rect 159653 106029 159771 106147
rect 159493 88189 159611 88307
rect 159653 88189 159771 88307
rect 159493 88029 159611 88147
rect 159653 88029 159771 88147
rect 159493 70189 159611 70307
rect 159653 70189 159771 70307
rect 159493 70029 159611 70147
rect 159653 70029 159771 70147
rect 159493 52189 159611 52307
rect 159653 52189 159771 52307
rect 159493 52029 159611 52147
rect 159653 52029 159771 52147
rect 159493 34189 159611 34307
rect 159653 34189 159771 34307
rect 159493 34029 159611 34147
rect 159653 34029 159771 34147
rect 159493 16189 159611 16307
rect 159653 16189 159771 16307
rect 159493 16029 159611 16147
rect 159653 16029 159771 16147
rect 150493 -3171 150611 -3053
rect 150653 -3171 150771 -3053
rect 150493 -3331 150611 -3213
rect 150653 -3331 150771 -3213
rect 162913 352301 163031 352419
rect 163073 352301 163191 352419
rect 162913 352141 163031 352259
rect 163073 352141 163191 352259
rect 162913 343609 163031 343727
rect 163073 343609 163191 343727
rect 162913 343449 163031 343567
rect 163073 343449 163191 343567
rect 162913 325609 163031 325727
rect 163073 325609 163191 325727
rect 162913 325449 163031 325567
rect 163073 325449 163191 325567
rect 162913 307609 163031 307727
rect 163073 307609 163191 307727
rect 162913 307449 163031 307567
rect 163073 307449 163191 307567
rect 162913 289609 163031 289727
rect 163073 289609 163191 289727
rect 162913 289449 163031 289567
rect 163073 289449 163191 289567
rect 162913 271609 163031 271727
rect 163073 271609 163191 271727
rect 162913 271449 163031 271567
rect 163073 271449 163191 271567
rect 162913 253609 163031 253727
rect 163073 253609 163191 253727
rect 162913 253449 163031 253567
rect 163073 253449 163191 253567
rect 162913 235609 163031 235727
rect 163073 235609 163191 235727
rect 162913 235449 163031 235567
rect 163073 235449 163191 235567
rect 162913 217609 163031 217727
rect 163073 217609 163191 217727
rect 162913 217449 163031 217567
rect 163073 217449 163191 217567
rect 162913 199609 163031 199727
rect 163073 199609 163191 199727
rect 162913 199449 163031 199567
rect 163073 199449 163191 199567
rect 162913 181609 163031 181727
rect 163073 181609 163191 181727
rect 162913 181449 163031 181567
rect 163073 181449 163191 181567
rect 162913 163609 163031 163727
rect 163073 163609 163191 163727
rect 162913 163449 163031 163567
rect 163073 163449 163191 163567
rect 162913 145609 163031 145727
rect 163073 145609 163191 145727
rect 162913 145449 163031 145567
rect 163073 145449 163191 145567
rect 162913 127609 163031 127727
rect 163073 127609 163191 127727
rect 162913 127449 163031 127567
rect 163073 127449 163191 127567
rect 162913 109609 163031 109727
rect 163073 109609 163191 109727
rect 162913 109449 163031 109567
rect 163073 109449 163191 109567
rect 162913 91609 163031 91727
rect 163073 91609 163191 91727
rect 162913 91449 163031 91567
rect 163073 91449 163191 91567
rect 162913 73609 163031 73727
rect 163073 73609 163191 73727
rect 162913 73449 163031 73567
rect 163073 73449 163191 73567
rect 162913 55609 163031 55727
rect 163073 55609 163191 55727
rect 162913 55449 163031 55567
rect 163073 55449 163191 55567
rect 162913 37609 163031 37727
rect 163073 37609 163191 37727
rect 162913 37449 163031 37567
rect 163073 37449 163191 37567
rect 162913 19609 163031 19727
rect 163073 19609 163191 19727
rect 162913 19449 163031 19567
rect 163073 19449 163191 19567
rect 162913 1609 163031 1727
rect 163073 1609 163191 1727
rect 162913 1449 163031 1567
rect 163073 1449 163191 1567
rect 162913 -291 163031 -173
rect 163073 -291 163191 -173
rect 162913 -451 163031 -333
rect 163073 -451 163191 -333
rect 164773 345469 164891 345587
rect 164933 345469 165051 345587
rect 164773 345309 164891 345427
rect 164933 345309 165051 345427
rect 164773 327469 164891 327587
rect 164933 327469 165051 327587
rect 164773 327309 164891 327427
rect 164933 327309 165051 327427
rect 164773 309469 164891 309587
rect 164933 309469 165051 309587
rect 164773 309309 164891 309427
rect 164933 309309 165051 309427
rect 164773 291469 164891 291587
rect 164933 291469 165051 291587
rect 164773 291309 164891 291427
rect 164933 291309 165051 291427
rect 164773 273469 164891 273587
rect 164933 273469 165051 273587
rect 164773 273309 164891 273427
rect 164933 273309 165051 273427
rect 164773 255469 164891 255587
rect 164933 255469 165051 255587
rect 164773 255309 164891 255427
rect 164933 255309 165051 255427
rect 164773 237469 164891 237587
rect 164933 237469 165051 237587
rect 164773 237309 164891 237427
rect 164933 237309 165051 237427
rect 164773 219469 164891 219587
rect 164933 219469 165051 219587
rect 164773 219309 164891 219427
rect 164933 219309 165051 219427
rect 164773 201469 164891 201587
rect 164933 201469 165051 201587
rect 164773 201309 164891 201427
rect 164933 201309 165051 201427
rect 164773 183469 164891 183587
rect 164933 183469 165051 183587
rect 164773 183309 164891 183427
rect 164933 183309 165051 183427
rect 164773 165469 164891 165587
rect 164933 165469 165051 165587
rect 164773 165309 164891 165427
rect 164933 165309 165051 165427
rect 164773 147469 164891 147587
rect 164933 147469 165051 147587
rect 164773 147309 164891 147427
rect 164933 147309 165051 147427
rect 164773 129469 164891 129587
rect 164933 129469 165051 129587
rect 164773 129309 164891 129427
rect 164933 129309 165051 129427
rect 164773 111469 164891 111587
rect 164933 111469 165051 111587
rect 164773 111309 164891 111427
rect 164933 111309 165051 111427
rect 164773 93469 164891 93587
rect 164933 93469 165051 93587
rect 164773 93309 164891 93427
rect 164933 93309 165051 93427
rect 164773 75469 164891 75587
rect 164933 75469 165051 75587
rect 164773 75309 164891 75427
rect 164933 75309 165051 75427
rect 164773 57469 164891 57587
rect 164933 57469 165051 57587
rect 164773 57309 164891 57427
rect 164933 57309 165051 57427
rect 164773 39469 164891 39587
rect 164933 39469 165051 39587
rect 164773 39309 164891 39427
rect 164933 39309 165051 39427
rect 164773 21469 164891 21587
rect 164933 21469 165051 21587
rect 164773 21309 164891 21427
rect 164933 21309 165051 21427
rect 164773 3469 164891 3587
rect 164933 3469 165051 3587
rect 164773 3309 164891 3427
rect 164933 3309 165051 3427
rect 164773 -1251 164891 -1133
rect 164933 -1251 165051 -1133
rect 164773 -1411 164891 -1293
rect 164933 -1411 165051 -1293
rect 166633 347329 166751 347447
rect 166793 347329 166911 347447
rect 166633 347169 166751 347287
rect 166793 347169 166911 347287
rect 166633 329329 166751 329447
rect 166793 329329 166911 329447
rect 166633 329169 166751 329287
rect 166793 329169 166911 329287
rect 166633 311329 166751 311447
rect 166793 311329 166911 311447
rect 166633 311169 166751 311287
rect 166793 311169 166911 311287
rect 166633 293329 166751 293447
rect 166793 293329 166911 293447
rect 166633 293169 166751 293287
rect 166793 293169 166911 293287
rect 166633 275329 166751 275447
rect 166793 275329 166911 275447
rect 166633 275169 166751 275287
rect 166793 275169 166911 275287
rect 166633 257329 166751 257447
rect 166793 257329 166911 257447
rect 166633 257169 166751 257287
rect 166793 257169 166911 257287
rect 166633 239329 166751 239447
rect 166793 239329 166911 239447
rect 166633 239169 166751 239287
rect 166793 239169 166911 239287
rect 166633 221329 166751 221447
rect 166793 221329 166911 221447
rect 166633 221169 166751 221287
rect 166793 221169 166911 221287
rect 166633 203329 166751 203447
rect 166793 203329 166911 203447
rect 166633 203169 166751 203287
rect 166793 203169 166911 203287
rect 166633 185329 166751 185447
rect 166793 185329 166911 185447
rect 166633 185169 166751 185287
rect 166793 185169 166911 185287
rect 166633 167329 166751 167447
rect 166793 167329 166911 167447
rect 166633 167169 166751 167287
rect 166793 167169 166911 167287
rect 166633 149329 166751 149447
rect 166793 149329 166911 149447
rect 166633 149169 166751 149287
rect 166793 149169 166911 149287
rect 166633 131329 166751 131447
rect 166793 131329 166911 131447
rect 166633 131169 166751 131287
rect 166793 131169 166911 131287
rect 166633 113329 166751 113447
rect 166793 113329 166911 113447
rect 166633 113169 166751 113287
rect 166793 113169 166911 113287
rect 166633 95329 166751 95447
rect 166793 95329 166911 95447
rect 166633 95169 166751 95287
rect 166793 95169 166911 95287
rect 166633 77329 166751 77447
rect 166793 77329 166911 77447
rect 166633 77169 166751 77287
rect 166793 77169 166911 77287
rect 166633 59329 166751 59447
rect 166793 59329 166911 59447
rect 166633 59169 166751 59287
rect 166793 59169 166911 59287
rect 166633 41329 166751 41447
rect 166793 41329 166911 41447
rect 166633 41169 166751 41287
rect 166793 41169 166911 41287
rect 166633 23329 166751 23447
rect 166793 23329 166911 23447
rect 166633 23169 166751 23287
rect 166793 23169 166911 23287
rect 166633 5329 166751 5447
rect 166793 5329 166911 5447
rect 166633 5169 166751 5287
rect 166793 5169 166911 5287
rect 166633 -2211 166751 -2093
rect 166793 -2211 166911 -2093
rect 166633 -2371 166751 -2253
rect 166793 -2371 166911 -2253
rect 177493 355661 177611 355779
rect 177653 355661 177771 355779
rect 177493 355501 177611 355619
rect 177653 355501 177771 355619
rect 175633 354701 175751 354819
rect 175793 354701 175911 354819
rect 175633 354541 175751 354659
rect 175793 354541 175911 354659
rect 173773 353741 173891 353859
rect 173933 353741 174051 353859
rect 173773 353581 173891 353699
rect 173933 353581 174051 353699
rect 168493 349189 168611 349307
rect 168653 349189 168771 349307
rect 168493 349029 168611 349147
rect 168653 349029 168771 349147
rect 168493 331189 168611 331307
rect 168653 331189 168771 331307
rect 168493 331029 168611 331147
rect 168653 331029 168771 331147
rect 168493 313189 168611 313307
rect 168653 313189 168771 313307
rect 168493 313029 168611 313147
rect 168653 313029 168771 313147
rect 168493 295189 168611 295307
rect 168653 295189 168771 295307
rect 168493 295029 168611 295147
rect 168653 295029 168771 295147
rect 168493 277189 168611 277307
rect 168653 277189 168771 277307
rect 168493 277029 168611 277147
rect 168653 277029 168771 277147
rect 168493 259189 168611 259307
rect 168653 259189 168771 259307
rect 168493 259029 168611 259147
rect 168653 259029 168771 259147
rect 168493 241189 168611 241307
rect 168653 241189 168771 241307
rect 168493 241029 168611 241147
rect 168653 241029 168771 241147
rect 168493 223189 168611 223307
rect 168653 223189 168771 223307
rect 168493 223029 168611 223147
rect 168653 223029 168771 223147
rect 168493 205189 168611 205307
rect 168653 205189 168771 205307
rect 168493 205029 168611 205147
rect 168653 205029 168771 205147
rect 168493 187189 168611 187307
rect 168653 187189 168771 187307
rect 168493 187029 168611 187147
rect 168653 187029 168771 187147
rect 168493 169189 168611 169307
rect 168653 169189 168771 169307
rect 168493 169029 168611 169147
rect 168653 169029 168771 169147
rect 168493 151189 168611 151307
rect 168653 151189 168771 151307
rect 168493 151029 168611 151147
rect 168653 151029 168771 151147
rect 168493 133189 168611 133307
rect 168653 133189 168771 133307
rect 168493 133029 168611 133147
rect 168653 133029 168771 133147
rect 168493 115189 168611 115307
rect 168653 115189 168771 115307
rect 168493 115029 168611 115147
rect 168653 115029 168771 115147
rect 168493 97189 168611 97307
rect 168653 97189 168771 97307
rect 168493 97029 168611 97147
rect 168653 97029 168771 97147
rect 168493 79189 168611 79307
rect 168653 79189 168771 79307
rect 168493 79029 168611 79147
rect 168653 79029 168771 79147
rect 168493 61189 168611 61307
rect 168653 61189 168771 61307
rect 168493 61029 168611 61147
rect 168653 61029 168771 61147
rect 168493 43189 168611 43307
rect 168653 43189 168771 43307
rect 168493 43029 168611 43147
rect 168653 43029 168771 43147
rect 168493 25189 168611 25307
rect 168653 25189 168771 25307
rect 168493 25029 168611 25147
rect 168653 25029 168771 25147
rect 168493 7189 168611 7307
rect 168653 7189 168771 7307
rect 168493 7029 168611 7147
rect 168653 7029 168771 7147
rect 159493 -3651 159611 -3533
rect 159653 -3651 159771 -3533
rect 159493 -3811 159611 -3693
rect 159653 -3811 159771 -3693
rect 171913 352781 172031 352899
rect 172073 352781 172191 352899
rect 171913 352621 172031 352739
rect 172073 352621 172191 352739
rect 171913 334609 172031 334727
rect 172073 334609 172191 334727
rect 171913 334449 172031 334567
rect 172073 334449 172191 334567
rect 171913 316609 172031 316727
rect 172073 316609 172191 316727
rect 171913 316449 172031 316567
rect 172073 316449 172191 316567
rect 171913 298609 172031 298727
rect 172073 298609 172191 298727
rect 171913 298449 172031 298567
rect 172073 298449 172191 298567
rect 171913 280609 172031 280727
rect 172073 280609 172191 280727
rect 171913 280449 172031 280567
rect 172073 280449 172191 280567
rect 171913 262609 172031 262727
rect 172073 262609 172191 262727
rect 171913 262449 172031 262567
rect 172073 262449 172191 262567
rect 171913 244609 172031 244727
rect 172073 244609 172191 244727
rect 171913 244449 172031 244567
rect 172073 244449 172191 244567
rect 171913 226609 172031 226727
rect 172073 226609 172191 226727
rect 171913 226449 172031 226567
rect 172073 226449 172191 226567
rect 171913 208609 172031 208727
rect 172073 208609 172191 208727
rect 171913 208449 172031 208567
rect 172073 208449 172191 208567
rect 171913 190609 172031 190727
rect 172073 190609 172191 190727
rect 171913 190449 172031 190567
rect 172073 190449 172191 190567
rect 171913 172609 172031 172727
rect 172073 172609 172191 172727
rect 171913 172449 172031 172567
rect 172073 172449 172191 172567
rect 171913 154609 172031 154727
rect 172073 154609 172191 154727
rect 171913 154449 172031 154567
rect 172073 154449 172191 154567
rect 171913 136609 172031 136727
rect 172073 136609 172191 136727
rect 171913 136449 172031 136567
rect 172073 136449 172191 136567
rect 171913 118609 172031 118727
rect 172073 118609 172191 118727
rect 171913 118449 172031 118567
rect 172073 118449 172191 118567
rect 171913 100609 172031 100727
rect 172073 100609 172191 100727
rect 171913 100449 172031 100567
rect 172073 100449 172191 100567
rect 171913 82609 172031 82727
rect 172073 82609 172191 82727
rect 171913 82449 172031 82567
rect 172073 82449 172191 82567
rect 171913 64609 172031 64727
rect 172073 64609 172191 64727
rect 171913 64449 172031 64567
rect 172073 64449 172191 64567
rect 171913 46609 172031 46727
rect 172073 46609 172191 46727
rect 171913 46449 172031 46567
rect 172073 46449 172191 46567
rect 171913 28609 172031 28727
rect 172073 28609 172191 28727
rect 171913 28449 172031 28567
rect 172073 28449 172191 28567
rect 171913 10609 172031 10727
rect 172073 10609 172191 10727
rect 171913 10449 172031 10567
rect 172073 10449 172191 10567
rect 171913 -771 172031 -653
rect 172073 -771 172191 -653
rect 171913 -931 172031 -813
rect 172073 -931 172191 -813
rect 173773 336469 173891 336587
rect 173933 336469 174051 336587
rect 173773 336309 173891 336427
rect 173933 336309 174051 336427
rect 173773 318469 173891 318587
rect 173933 318469 174051 318587
rect 173773 318309 173891 318427
rect 173933 318309 174051 318427
rect 173773 300469 173891 300587
rect 173933 300469 174051 300587
rect 173773 300309 173891 300427
rect 173933 300309 174051 300427
rect 173773 282469 173891 282587
rect 173933 282469 174051 282587
rect 173773 282309 173891 282427
rect 173933 282309 174051 282427
rect 173773 264469 173891 264587
rect 173933 264469 174051 264587
rect 173773 264309 173891 264427
rect 173933 264309 174051 264427
rect 173773 246469 173891 246587
rect 173933 246469 174051 246587
rect 173773 246309 173891 246427
rect 173933 246309 174051 246427
rect 173773 228469 173891 228587
rect 173933 228469 174051 228587
rect 173773 228309 173891 228427
rect 173933 228309 174051 228427
rect 173773 210469 173891 210587
rect 173933 210469 174051 210587
rect 173773 210309 173891 210427
rect 173933 210309 174051 210427
rect 173773 192469 173891 192587
rect 173933 192469 174051 192587
rect 173773 192309 173891 192427
rect 173933 192309 174051 192427
rect 173773 174469 173891 174587
rect 173933 174469 174051 174587
rect 173773 174309 173891 174427
rect 173933 174309 174051 174427
rect 173773 156469 173891 156587
rect 173933 156469 174051 156587
rect 173773 156309 173891 156427
rect 173933 156309 174051 156427
rect 173773 138469 173891 138587
rect 173933 138469 174051 138587
rect 173773 138309 173891 138427
rect 173933 138309 174051 138427
rect 173773 120469 173891 120587
rect 173933 120469 174051 120587
rect 173773 120309 173891 120427
rect 173933 120309 174051 120427
rect 173773 102469 173891 102587
rect 173933 102469 174051 102587
rect 173773 102309 173891 102427
rect 173933 102309 174051 102427
rect 173773 84469 173891 84587
rect 173933 84469 174051 84587
rect 173773 84309 173891 84427
rect 173933 84309 174051 84427
rect 173773 66469 173891 66587
rect 173933 66469 174051 66587
rect 173773 66309 173891 66427
rect 173933 66309 174051 66427
rect 173773 48469 173891 48587
rect 173933 48469 174051 48587
rect 173773 48309 173891 48427
rect 173933 48309 174051 48427
rect 173773 30469 173891 30587
rect 173933 30469 174051 30587
rect 173773 30309 173891 30427
rect 173933 30309 174051 30427
rect 173773 12469 173891 12587
rect 173933 12469 174051 12587
rect 173773 12309 173891 12427
rect 173933 12309 174051 12427
rect 173773 -1731 173891 -1613
rect 173933 -1731 174051 -1613
rect 173773 -1891 173891 -1773
rect 173933 -1891 174051 -1773
rect 175633 338329 175751 338447
rect 175793 338329 175911 338447
rect 175633 338169 175751 338287
rect 175793 338169 175911 338287
rect 175633 320329 175751 320447
rect 175793 320329 175911 320447
rect 175633 320169 175751 320287
rect 175793 320169 175911 320287
rect 175633 302329 175751 302447
rect 175793 302329 175911 302447
rect 175633 302169 175751 302287
rect 175793 302169 175911 302287
rect 175633 284329 175751 284447
rect 175793 284329 175911 284447
rect 175633 284169 175751 284287
rect 175793 284169 175911 284287
rect 175633 266329 175751 266447
rect 175793 266329 175911 266447
rect 175633 266169 175751 266287
rect 175793 266169 175911 266287
rect 175633 248329 175751 248447
rect 175793 248329 175911 248447
rect 175633 248169 175751 248287
rect 175793 248169 175911 248287
rect 175633 230329 175751 230447
rect 175793 230329 175911 230447
rect 175633 230169 175751 230287
rect 175793 230169 175911 230287
rect 175633 212329 175751 212447
rect 175793 212329 175911 212447
rect 175633 212169 175751 212287
rect 175793 212169 175911 212287
rect 175633 194329 175751 194447
rect 175793 194329 175911 194447
rect 175633 194169 175751 194287
rect 175793 194169 175911 194287
rect 175633 176329 175751 176447
rect 175793 176329 175911 176447
rect 175633 176169 175751 176287
rect 175793 176169 175911 176287
rect 175633 158329 175751 158447
rect 175793 158329 175911 158447
rect 175633 158169 175751 158287
rect 175793 158169 175911 158287
rect 175633 140329 175751 140447
rect 175793 140329 175911 140447
rect 175633 140169 175751 140287
rect 175793 140169 175911 140287
rect 175633 122329 175751 122447
rect 175793 122329 175911 122447
rect 175633 122169 175751 122287
rect 175793 122169 175911 122287
rect 175633 104329 175751 104447
rect 175793 104329 175911 104447
rect 175633 104169 175751 104287
rect 175793 104169 175911 104287
rect 175633 86329 175751 86447
rect 175793 86329 175911 86447
rect 175633 86169 175751 86287
rect 175793 86169 175911 86287
rect 175633 68329 175751 68447
rect 175793 68329 175911 68447
rect 175633 68169 175751 68287
rect 175793 68169 175911 68287
rect 175633 50329 175751 50447
rect 175793 50329 175911 50447
rect 175633 50169 175751 50287
rect 175793 50169 175911 50287
rect 175633 32329 175751 32447
rect 175793 32329 175911 32447
rect 175633 32169 175751 32287
rect 175793 32169 175911 32287
rect 175633 14329 175751 14447
rect 175793 14329 175911 14447
rect 175633 14169 175751 14287
rect 175793 14169 175911 14287
rect 175633 -2691 175751 -2573
rect 175793 -2691 175911 -2573
rect 175633 -2851 175751 -2733
rect 175793 -2851 175911 -2733
rect 186493 355181 186611 355299
rect 186653 355181 186771 355299
rect 186493 355021 186611 355139
rect 186653 355021 186771 355139
rect 184633 354221 184751 354339
rect 184793 354221 184911 354339
rect 184633 354061 184751 354179
rect 184793 354061 184911 354179
rect 182773 353261 182891 353379
rect 182933 353261 183051 353379
rect 182773 353101 182891 353219
rect 182933 353101 183051 353219
rect 177493 340189 177611 340307
rect 177653 340189 177771 340307
rect 177493 340029 177611 340147
rect 177653 340029 177771 340147
rect 177493 322189 177611 322307
rect 177653 322189 177771 322307
rect 177493 322029 177611 322147
rect 177653 322029 177771 322147
rect 177493 304189 177611 304307
rect 177653 304189 177771 304307
rect 177493 304029 177611 304147
rect 177653 304029 177771 304147
rect 177493 286189 177611 286307
rect 177653 286189 177771 286307
rect 177493 286029 177611 286147
rect 177653 286029 177771 286147
rect 177493 268189 177611 268307
rect 177653 268189 177771 268307
rect 177493 268029 177611 268147
rect 177653 268029 177771 268147
rect 177493 250189 177611 250307
rect 177653 250189 177771 250307
rect 177493 250029 177611 250147
rect 177653 250029 177771 250147
rect 177493 232189 177611 232307
rect 177653 232189 177771 232307
rect 177493 232029 177611 232147
rect 177653 232029 177771 232147
rect 177493 214189 177611 214307
rect 177653 214189 177771 214307
rect 177493 214029 177611 214147
rect 177653 214029 177771 214147
rect 177493 196189 177611 196307
rect 177653 196189 177771 196307
rect 177493 196029 177611 196147
rect 177653 196029 177771 196147
rect 177493 178189 177611 178307
rect 177653 178189 177771 178307
rect 177493 178029 177611 178147
rect 177653 178029 177771 178147
rect 177493 160189 177611 160307
rect 177653 160189 177771 160307
rect 177493 160029 177611 160147
rect 177653 160029 177771 160147
rect 177493 142189 177611 142307
rect 177653 142189 177771 142307
rect 177493 142029 177611 142147
rect 177653 142029 177771 142147
rect 177493 124189 177611 124307
rect 177653 124189 177771 124307
rect 177493 124029 177611 124147
rect 177653 124029 177771 124147
rect 177493 106189 177611 106307
rect 177653 106189 177771 106307
rect 177493 106029 177611 106147
rect 177653 106029 177771 106147
rect 177493 88189 177611 88307
rect 177653 88189 177771 88307
rect 177493 88029 177611 88147
rect 177653 88029 177771 88147
rect 177493 70189 177611 70307
rect 177653 70189 177771 70307
rect 177493 70029 177611 70147
rect 177653 70029 177771 70147
rect 177493 52189 177611 52307
rect 177653 52189 177771 52307
rect 177493 52029 177611 52147
rect 177653 52029 177771 52147
rect 177493 34189 177611 34307
rect 177653 34189 177771 34307
rect 177493 34029 177611 34147
rect 177653 34029 177771 34147
rect 177493 16189 177611 16307
rect 177653 16189 177771 16307
rect 177493 16029 177611 16147
rect 177653 16029 177771 16147
rect 168493 -3171 168611 -3053
rect 168653 -3171 168771 -3053
rect 168493 -3331 168611 -3213
rect 168653 -3331 168771 -3213
rect 180913 352301 181031 352419
rect 181073 352301 181191 352419
rect 180913 352141 181031 352259
rect 181073 352141 181191 352259
rect 180913 343609 181031 343727
rect 181073 343609 181191 343727
rect 180913 343449 181031 343567
rect 181073 343449 181191 343567
rect 180913 325609 181031 325727
rect 181073 325609 181191 325727
rect 180913 325449 181031 325567
rect 181073 325449 181191 325567
rect 180913 307609 181031 307727
rect 181073 307609 181191 307727
rect 180913 307449 181031 307567
rect 181073 307449 181191 307567
rect 180913 289609 181031 289727
rect 181073 289609 181191 289727
rect 180913 289449 181031 289567
rect 181073 289449 181191 289567
rect 180913 271609 181031 271727
rect 181073 271609 181191 271727
rect 180913 271449 181031 271567
rect 181073 271449 181191 271567
rect 180913 253609 181031 253727
rect 181073 253609 181191 253727
rect 180913 253449 181031 253567
rect 181073 253449 181191 253567
rect 180913 235609 181031 235727
rect 181073 235609 181191 235727
rect 180913 235449 181031 235567
rect 181073 235449 181191 235567
rect 180913 217609 181031 217727
rect 181073 217609 181191 217727
rect 180913 217449 181031 217567
rect 181073 217449 181191 217567
rect 180913 199609 181031 199727
rect 181073 199609 181191 199727
rect 180913 199449 181031 199567
rect 181073 199449 181191 199567
rect 180913 181609 181031 181727
rect 181073 181609 181191 181727
rect 180913 181449 181031 181567
rect 181073 181449 181191 181567
rect 180913 163609 181031 163727
rect 181073 163609 181191 163727
rect 180913 163449 181031 163567
rect 181073 163449 181191 163567
rect 180913 145609 181031 145727
rect 181073 145609 181191 145727
rect 180913 145449 181031 145567
rect 181073 145449 181191 145567
rect 180913 127609 181031 127727
rect 181073 127609 181191 127727
rect 180913 127449 181031 127567
rect 181073 127449 181191 127567
rect 180913 109609 181031 109727
rect 181073 109609 181191 109727
rect 180913 109449 181031 109567
rect 181073 109449 181191 109567
rect 180913 91609 181031 91727
rect 181073 91609 181191 91727
rect 180913 91449 181031 91567
rect 181073 91449 181191 91567
rect 180913 73609 181031 73727
rect 181073 73609 181191 73727
rect 180913 73449 181031 73567
rect 181073 73449 181191 73567
rect 180913 55609 181031 55727
rect 181073 55609 181191 55727
rect 180913 55449 181031 55567
rect 181073 55449 181191 55567
rect 180913 37609 181031 37727
rect 181073 37609 181191 37727
rect 180913 37449 181031 37567
rect 181073 37449 181191 37567
rect 180913 19609 181031 19727
rect 181073 19609 181191 19727
rect 180913 19449 181031 19567
rect 181073 19449 181191 19567
rect 180913 1609 181031 1727
rect 181073 1609 181191 1727
rect 180913 1449 181031 1567
rect 181073 1449 181191 1567
rect 180913 -291 181031 -173
rect 181073 -291 181191 -173
rect 180913 -451 181031 -333
rect 181073 -451 181191 -333
rect 182773 345469 182891 345587
rect 182933 345469 183051 345587
rect 182773 345309 182891 345427
rect 182933 345309 183051 345427
rect 182773 327469 182891 327587
rect 182933 327469 183051 327587
rect 182773 327309 182891 327427
rect 182933 327309 183051 327427
rect 182773 309469 182891 309587
rect 182933 309469 183051 309587
rect 182773 309309 182891 309427
rect 182933 309309 183051 309427
rect 182773 291469 182891 291587
rect 182933 291469 183051 291587
rect 182773 291309 182891 291427
rect 182933 291309 183051 291427
rect 182773 273469 182891 273587
rect 182933 273469 183051 273587
rect 182773 273309 182891 273427
rect 182933 273309 183051 273427
rect 182773 255469 182891 255587
rect 182933 255469 183051 255587
rect 182773 255309 182891 255427
rect 182933 255309 183051 255427
rect 182773 237469 182891 237587
rect 182933 237469 183051 237587
rect 182773 237309 182891 237427
rect 182933 237309 183051 237427
rect 182773 219469 182891 219587
rect 182933 219469 183051 219587
rect 182773 219309 182891 219427
rect 182933 219309 183051 219427
rect 182773 201469 182891 201587
rect 182933 201469 183051 201587
rect 182773 201309 182891 201427
rect 182933 201309 183051 201427
rect 182773 183469 182891 183587
rect 182933 183469 183051 183587
rect 182773 183309 182891 183427
rect 182933 183309 183051 183427
rect 182773 165469 182891 165587
rect 182933 165469 183051 165587
rect 182773 165309 182891 165427
rect 182933 165309 183051 165427
rect 182773 147469 182891 147587
rect 182933 147469 183051 147587
rect 182773 147309 182891 147427
rect 182933 147309 183051 147427
rect 182773 129469 182891 129587
rect 182933 129469 183051 129587
rect 182773 129309 182891 129427
rect 182933 129309 183051 129427
rect 182773 111469 182891 111587
rect 182933 111469 183051 111587
rect 182773 111309 182891 111427
rect 182933 111309 183051 111427
rect 182773 93469 182891 93587
rect 182933 93469 183051 93587
rect 182773 93309 182891 93427
rect 182933 93309 183051 93427
rect 182773 75469 182891 75587
rect 182933 75469 183051 75587
rect 182773 75309 182891 75427
rect 182933 75309 183051 75427
rect 182773 57469 182891 57587
rect 182933 57469 183051 57587
rect 182773 57309 182891 57427
rect 182933 57309 183051 57427
rect 182773 39469 182891 39587
rect 182933 39469 183051 39587
rect 182773 39309 182891 39427
rect 182933 39309 183051 39427
rect 182773 21469 182891 21587
rect 182933 21469 183051 21587
rect 182773 21309 182891 21427
rect 182933 21309 183051 21427
rect 182773 3469 182891 3587
rect 182933 3469 183051 3587
rect 182773 3309 182891 3427
rect 182933 3309 183051 3427
rect 182773 -1251 182891 -1133
rect 182933 -1251 183051 -1133
rect 182773 -1411 182891 -1293
rect 182933 -1411 183051 -1293
rect 184633 347329 184751 347447
rect 184793 347329 184911 347447
rect 184633 347169 184751 347287
rect 184793 347169 184911 347287
rect 184633 329329 184751 329447
rect 184793 329329 184911 329447
rect 184633 329169 184751 329287
rect 184793 329169 184911 329287
rect 184633 311329 184751 311447
rect 184793 311329 184911 311447
rect 184633 311169 184751 311287
rect 184793 311169 184911 311287
rect 184633 293329 184751 293447
rect 184793 293329 184911 293447
rect 184633 293169 184751 293287
rect 184793 293169 184911 293287
rect 184633 275329 184751 275447
rect 184793 275329 184911 275447
rect 184633 275169 184751 275287
rect 184793 275169 184911 275287
rect 184633 257329 184751 257447
rect 184793 257329 184911 257447
rect 184633 257169 184751 257287
rect 184793 257169 184911 257287
rect 184633 239329 184751 239447
rect 184793 239329 184911 239447
rect 184633 239169 184751 239287
rect 184793 239169 184911 239287
rect 184633 221329 184751 221447
rect 184793 221329 184911 221447
rect 184633 221169 184751 221287
rect 184793 221169 184911 221287
rect 184633 203329 184751 203447
rect 184793 203329 184911 203447
rect 184633 203169 184751 203287
rect 184793 203169 184911 203287
rect 184633 185329 184751 185447
rect 184793 185329 184911 185447
rect 184633 185169 184751 185287
rect 184793 185169 184911 185287
rect 184633 167329 184751 167447
rect 184793 167329 184911 167447
rect 184633 167169 184751 167287
rect 184793 167169 184911 167287
rect 184633 149329 184751 149447
rect 184793 149329 184911 149447
rect 184633 149169 184751 149287
rect 184793 149169 184911 149287
rect 184633 131329 184751 131447
rect 184793 131329 184911 131447
rect 184633 131169 184751 131287
rect 184793 131169 184911 131287
rect 184633 113329 184751 113447
rect 184793 113329 184911 113447
rect 184633 113169 184751 113287
rect 184793 113169 184911 113287
rect 184633 95329 184751 95447
rect 184793 95329 184911 95447
rect 184633 95169 184751 95287
rect 184793 95169 184911 95287
rect 184633 77329 184751 77447
rect 184793 77329 184911 77447
rect 184633 77169 184751 77287
rect 184793 77169 184911 77287
rect 184633 59329 184751 59447
rect 184793 59329 184911 59447
rect 184633 59169 184751 59287
rect 184793 59169 184911 59287
rect 184633 41329 184751 41447
rect 184793 41329 184911 41447
rect 184633 41169 184751 41287
rect 184793 41169 184911 41287
rect 184633 23329 184751 23447
rect 184793 23329 184911 23447
rect 184633 23169 184751 23287
rect 184793 23169 184911 23287
rect 184633 5329 184751 5447
rect 184793 5329 184911 5447
rect 184633 5169 184751 5287
rect 184793 5169 184911 5287
rect 184633 -2211 184751 -2093
rect 184793 -2211 184911 -2093
rect 184633 -2371 184751 -2253
rect 184793 -2371 184911 -2253
rect 195493 355661 195611 355779
rect 195653 355661 195771 355779
rect 195493 355501 195611 355619
rect 195653 355501 195771 355619
rect 193633 354701 193751 354819
rect 193793 354701 193911 354819
rect 193633 354541 193751 354659
rect 193793 354541 193911 354659
rect 191773 353741 191891 353859
rect 191933 353741 192051 353859
rect 191773 353581 191891 353699
rect 191933 353581 192051 353699
rect 186493 349189 186611 349307
rect 186653 349189 186771 349307
rect 186493 349029 186611 349147
rect 186653 349029 186771 349147
rect 186493 331189 186611 331307
rect 186653 331189 186771 331307
rect 186493 331029 186611 331147
rect 186653 331029 186771 331147
rect 186493 313189 186611 313307
rect 186653 313189 186771 313307
rect 186493 313029 186611 313147
rect 186653 313029 186771 313147
rect 186493 295189 186611 295307
rect 186653 295189 186771 295307
rect 186493 295029 186611 295147
rect 186653 295029 186771 295147
rect 186493 277189 186611 277307
rect 186653 277189 186771 277307
rect 186493 277029 186611 277147
rect 186653 277029 186771 277147
rect 186493 259189 186611 259307
rect 186653 259189 186771 259307
rect 186493 259029 186611 259147
rect 186653 259029 186771 259147
rect 186493 241189 186611 241307
rect 186653 241189 186771 241307
rect 186493 241029 186611 241147
rect 186653 241029 186771 241147
rect 186493 223189 186611 223307
rect 186653 223189 186771 223307
rect 186493 223029 186611 223147
rect 186653 223029 186771 223147
rect 186493 205189 186611 205307
rect 186653 205189 186771 205307
rect 186493 205029 186611 205147
rect 186653 205029 186771 205147
rect 186493 187189 186611 187307
rect 186653 187189 186771 187307
rect 186493 187029 186611 187147
rect 186653 187029 186771 187147
rect 186493 169189 186611 169307
rect 186653 169189 186771 169307
rect 186493 169029 186611 169147
rect 186653 169029 186771 169147
rect 186493 151189 186611 151307
rect 186653 151189 186771 151307
rect 186493 151029 186611 151147
rect 186653 151029 186771 151147
rect 186493 133189 186611 133307
rect 186653 133189 186771 133307
rect 186493 133029 186611 133147
rect 186653 133029 186771 133147
rect 186493 115189 186611 115307
rect 186653 115189 186771 115307
rect 186493 115029 186611 115147
rect 186653 115029 186771 115147
rect 186493 97189 186611 97307
rect 186653 97189 186771 97307
rect 186493 97029 186611 97147
rect 186653 97029 186771 97147
rect 186493 79189 186611 79307
rect 186653 79189 186771 79307
rect 186493 79029 186611 79147
rect 186653 79029 186771 79147
rect 186493 61189 186611 61307
rect 186653 61189 186771 61307
rect 186493 61029 186611 61147
rect 186653 61029 186771 61147
rect 186493 43189 186611 43307
rect 186653 43189 186771 43307
rect 186493 43029 186611 43147
rect 186653 43029 186771 43147
rect 186493 25189 186611 25307
rect 186653 25189 186771 25307
rect 186493 25029 186611 25147
rect 186653 25029 186771 25147
rect 186493 7189 186611 7307
rect 186653 7189 186771 7307
rect 186493 7029 186611 7147
rect 186653 7029 186771 7147
rect 177493 -3651 177611 -3533
rect 177653 -3651 177771 -3533
rect 177493 -3811 177611 -3693
rect 177653 -3811 177771 -3693
rect 189913 352781 190031 352899
rect 190073 352781 190191 352899
rect 189913 352621 190031 352739
rect 190073 352621 190191 352739
rect 189913 334609 190031 334727
rect 190073 334609 190191 334727
rect 189913 334449 190031 334567
rect 190073 334449 190191 334567
rect 189913 316609 190031 316727
rect 190073 316609 190191 316727
rect 189913 316449 190031 316567
rect 190073 316449 190191 316567
rect 189913 298609 190031 298727
rect 190073 298609 190191 298727
rect 189913 298449 190031 298567
rect 190073 298449 190191 298567
rect 189913 280609 190031 280727
rect 190073 280609 190191 280727
rect 189913 280449 190031 280567
rect 190073 280449 190191 280567
rect 189913 262609 190031 262727
rect 190073 262609 190191 262727
rect 189913 262449 190031 262567
rect 190073 262449 190191 262567
rect 189913 244609 190031 244727
rect 190073 244609 190191 244727
rect 189913 244449 190031 244567
rect 190073 244449 190191 244567
rect 189913 226609 190031 226727
rect 190073 226609 190191 226727
rect 189913 226449 190031 226567
rect 190073 226449 190191 226567
rect 189913 208609 190031 208727
rect 190073 208609 190191 208727
rect 189913 208449 190031 208567
rect 190073 208449 190191 208567
rect 189913 190609 190031 190727
rect 190073 190609 190191 190727
rect 189913 190449 190031 190567
rect 190073 190449 190191 190567
rect 189913 172609 190031 172727
rect 190073 172609 190191 172727
rect 189913 172449 190031 172567
rect 190073 172449 190191 172567
rect 189913 154609 190031 154727
rect 190073 154609 190191 154727
rect 189913 154449 190031 154567
rect 190073 154449 190191 154567
rect 189913 136609 190031 136727
rect 190073 136609 190191 136727
rect 189913 136449 190031 136567
rect 190073 136449 190191 136567
rect 189913 118609 190031 118727
rect 190073 118609 190191 118727
rect 189913 118449 190031 118567
rect 190073 118449 190191 118567
rect 189913 100609 190031 100727
rect 190073 100609 190191 100727
rect 189913 100449 190031 100567
rect 190073 100449 190191 100567
rect 189913 82609 190031 82727
rect 190073 82609 190191 82727
rect 189913 82449 190031 82567
rect 190073 82449 190191 82567
rect 189913 64609 190031 64727
rect 190073 64609 190191 64727
rect 189913 64449 190031 64567
rect 190073 64449 190191 64567
rect 189913 46609 190031 46727
rect 190073 46609 190191 46727
rect 189913 46449 190031 46567
rect 190073 46449 190191 46567
rect 189913 28609 190031 28727
rect 190073 28609 190191 28727
rect 189913 28449 190031 28567
rect 190073 28449 190191 28567
rect 189913 10609 190031 10727
rect 190073 10609 190191 10727
rect 189913 10449 190031 10567
rect 190073 10449 190191 10567
rect 189913 -771 190031 -653
rect 190073 -771 190191 -653
rect 189913 -931 190031 -813
rect 190073 -931 190191 -813
rect 191773 336469 191891 336587
rect 191933 336469 192051 336587
rect 191773 336309 191891 336427
rect 191933 336309 192051 336427
rect 191773 318469 191891 318587
rect 191933 318469 192051 318587
rect 191773 318309 191891 318427
rect 191933 318309 192051 318427
rect 191773 300469 191891 300587
rect 191933 300469 192051 300587
rect 191773 300309 191891 300427
rect 191933 300309 192051 300427
rect 191773 282469 191891 282587
rect 191933 282469 192051 282587
rect 191773 282309 191891 282427
rect 191933 282309 192051 282427
rect 191773 264469 191891 264587
rect 191933 264469 192051 264587
rect 191773 264309 191891 264427
rect 191933 264309 192051 264427
rect 191773 246469 191891 246587
rect 191933 246469 192051 246587
rect 191773 246309 191891 246427
rect 191933 246309 192051 246427
rect 191773 228469 191891 228587
rect 191933 228469 192051 228587
rect 191773 228309 191891 228427
rect 191933 228309 192051 228427
rect 191773 210469 191891 210587
rect 191933 210469 192051 210587
rect 191773 210309 191891 210427
rect 191933 210309 192051 210427
rect 191773 192469 191891 192587
rect 191933 192469 192051 192587
rect 191773 192309 191891 192427
rect 191933 192309 192051 192427
rect 191773 174469 191891 174587
rect 191933 174469 192051 174587
rect 191773 174309 191891 174427
rect 191933 174309 192051 174427
rect 191773 156469 191891 156587
rect 191933 156469 192051 156587
rect 191773 156309 191891 156427
rect 191933 156309 192051 156427
rect 191773 138469 191891 138587
rect 191933 138469 192051 138587
rect 191773 138309 191891 138427
rect 191933 138309 192051 138427
rect 191773 120469 191891 120587
rect 191933 120469 192051 120587
rect 191773 120309 191891 120427
rect 191933 120309 192051 120427
rect 191773 102469 191891 102587
rect 191933 102469 192051 102587
rect 191773 102309 191891 102427
rect 191933 102309 192051 102427
rect 191773 84469 191891 84587
rect 191933 84469 192051 84587
rect 191773 84309 191891 84427
rect 191933 84309 192051 84427
rect 191773 66469 191891 66587
rect 191933 66469 192051 66587
rect 191773 66309 191891 66427
rect 191933 66309 192051 66427
rect 191773 48469 191891 48587
rect 191933 48469 192051 48587
rect 191773 48309 191891 48427
rect 191933 48309 192051 48427
rect 191773 30469 191891 30587
rect 191933 30469 192051 30587
rect 191773 30309 191891 30427
rect 191933 30309 192051 30427
rect 191773 12469 191891 12587
rect 191933 12469 192051 12587
rect 191773 12309 191891 12427
rect 191933 12309 192051 12427
rect 191773 -1731 191891 -1613
rect 191933 -1731 192051 -1613
rect 191773 -1891 191891 -1773
rect 191933 -1891 192051 -1773
rect 193633 338329 193751 338447
rect 193793 338329 193911 338447
rect 193633 338169 193751 338287
rect 193793 338169 193911 338287
rect 193633 320329 193751 320447
rect 193793 320329 193911 320447
rect 193633 320169 193751 320287
rect 193793 320169 193911 320287
rect 193633 302329 193751 302447
rect 193793 302329 193911 302447
rect 193633 302169 193751 302287
rect 193793 302169 193911 302287
rect 193633 284329 193751 284447
rect 193793 284329 193911 284447
rect 193633 284169 193751 284287
rect 193793 284169 193911 284287
rect 193633 266329 193751 266447
rect 193793 266329 193911 266447
rect 193633 266169 193751 266287
rect 193793 266169 193911 266287
rect 193633 248329 193751 248447
rect 193793 248329 193911 248447
rect 193633 248169 193751 248287
rect 193793 248169 193911 248287
rect 193633 230329 193751 230447
rect 193793 230329 193911 230447
rect 193633 230169 193751 230287
rect 193793 230169 193911 230287
rect 193633 212329 193751 212447
rect 193793 212329 193911 212447
rect 193633 212169 193751 212287
rect 193793 212169 193911 212287
rect 193633 194329 193751 194447
rect 193793 194329 193911 194447
rect 193633 194169 193751 194287
rect 193793 194169 193911 194287
rect 193633 176329 193751 176447
rect 193793 176329 193911 176447
rect 193633 176169 193751 176287
rect 193793 176169 193911 176287
rect 193633 158329 193751 158447
rect 193793 158329 193911 158447
rect 193633 158169 193751 158287
rect 193793 158169 193911 158287
rect 193633 140329 193751 140447
rect 193793 140329 193911 140447
rect 193633 140169 193751 140287
rect 193793 140169 193911 140287
rect 193633 122329 193751 122447
rect 193793 122329 193911 122447
rect 193633 122169 193751 122287
rect 193793 122169 193911 122287
rect 193633 104329 193751 104447
rect 193793 104329 193911 104447
rect 193633 104169 193751 104287
rect 193793 104169 193911 104287
rect 193633 86329 193751 86447
rect 193793 86329 193911 86447
rect 193633 86169 193751 86287
rect 193793 86169 193911 86287
rect 193633 68329 193751 68447
rect 193793 68329 193911 68447
rect 193633 68169 193751 68287
rect 193793 68169 193911 68287
rect 193633 50329 193751 50447
rect 193793 50329 193911 50447
rect 193633 50169 193751 50287
rect 193793 50169 193911 50287
rect 193633 32329 193751 32447
rect 193793 32329 193911 32447
rect 193633 32169 193751 32287
rect 193793 32169 193911 32287
rect 193633 14329 193751 14447
rect 193793 14329 193911 14447
rect 193633 14169 193751 14287
rect 193793 14169 193911 14287
rect 193633 -2691 193751 -2573
rect 193793 -2691 193911 -2573
rect 193633 -2851 193751 -2733
rect 193793 -2851 193911 -2733
rect 204493 355181 204611 355299
rect 204653 355181 204771 355299
rect 204493 355021 204611 355139
rect 204653 355021 204771 355139
rect 202633 354221 202751 354339
rect 202793 354221 202911 354339
rect 202633 354061 202751 354179
rect 202793 354061 202911 354179
rect 200773 353261 200891 353379
rect 200933 353261 201051 353379
rect 200773 353101 200891 353219
rect 200933 353101 201051 353219
rect 195493 340189 195611 340307
rect 195653 340189 195771 340307
rect 195493 340029 195611 340147
rect 195653 340029 195771 340147
rect 195493 322189 195611 322307
rect 195653 322189 195771 322307
rect 195493 322029 195611 322147
rect 195653 322029 195771 322147
rect 195493 304189 195611 304307
rect 195653 304189 195771 304307
rect 195493 304029 195611 304147
rect 195653 304029 195771 304147
rect 195493 286189 195611 286307
rect 195653 286189 195771 286307
rect 195493 286029 195611 286147
rect 195653 286029 195771 286147
rect 195493 268189 195611 268307
rect 195653 268189 195771 268307
rect 195493 268029 195611 268147
rect 195653 268029 195771 268147
rect 195493 250189 195611 250307
rect 195653 250189 195771 250307
rect 195493 250029 195611 250147
rect 195653 250029 195771 250147
rect 195493 232189 195611 232307
rect 195653 232189 195771 232307
rect 195493 232029 195611 232147
rect 195653 232029 195771 232147
rect 195493 214189 195611 214307
rect 195653 214189 195771 214307
rect 195493 214029 195611 214147
rect 195653 214029 195771 214147
rect 195493 196189 195611 196307
rect 195653 196189 195771 196307
rect 195493 196029 195611 196147
rect 195653 196029 195771 196147
rect 195493 178189 195611 178307
rect 195653 178189 195771 178307
rect 195493 178029 195611 178147
rect 195653 178029 195771 178147
rect 195493 160189 195611 160307
rect 195653 160189 195771 160307
rect 195493 160029 195611 160147
rect 195653 160029 195771 160147
rect 195493 142189 195611 142307
rect 195653 142189 195771 142307
rect 195493 142029 195611 142147
rect 195653 142029 195771 142147
rect 195493 124189 195611 124307
rect 195653 124189 195771 124307
rect 195493 124029 195611 124147
rect 195653 124029 195771 124147
rect 195493 106189 195611 106307
rect 195653 106189 195771 106307
rect 195493 106029 195611 106147
rect 195653 106029 195771 106147
rect 195493 88189 195611 88307
rect 195653 88189 195771 88307
rect 195493 88029 195611 88147
rect 195653 88029 195771 88147
rect 195493 70189 195611 70307
rect 195653 70189 195771 70307
rect 195493 70029 195611 70147
rect 195653 70029 195771 70147
rect 195493 52189 195611 52307
rect 195653 52189 195771 52307
rect 195493 52029 195611 52147
rect 195653 52029 195771 52147
rect 195493 34189 195611 34307
rect 195653 34189 195771 34307
rect 195493 34029 195611 34147
rect 195653 34029 195771 34147
rect 195493 16189 195611 16307
rect 195653 16189 195771 16307
rect 195493 16029 195611 16147
rect 195653 16029 195771 16147
rect 186493 -3171 186611 -3053
rect 186653 -3171 186771 -3053
rect 186493 -3331 186611 -3213
rect 186653 -3331 186771 -3213
rect 198913 352301 199031 352419
rect 199073 352301 199191 352419
rect 198913 352141 199031 352259
rect 199073 352141 199191 352259
rect 198913 343609 199031 343727
rect 199073 343609 199191 343727
rect 198913 343449 199031 343567
rect 199073 343449 199191 343567
rect 198913 325609 199031 325727
rect 199073 325609 199191 325727
rect 198913 325449 199031 325567
rect 199073 325449 199191 325567
rect 198913 307609 199031 307727
rect 199073 307609 199191 307727
rect 198913 307449 199031 307567
rect 199073 307449 199191 307567
rect 198913 289609 199031 289727
rect 199073 289609 199191 289727
rect 198913 289449 199031 289567
rect 199073 289449 199191 289567
rect 198913 271609 199031 271727
rect 199073 271609 199191 271727
rect 198913 271449 199031 271567
rect 199073 271449 199191 271567
rect 198913 253609 199031 253727
rect 199073 253609 199191 253727
rect 198913 253449 199031 253567
rect 199073 253449 199191 253567
rect 198913 235609 199031 235727
rect 199073 235609 199191 235727
rect 198913 235449 199031 235567
rect 199073 235449 199191 235567
rect 198913 217609 199031 217727
rect 199073 217609 199191 217727
rect 198913 217449 199031 217567
rect 199073 217449 199191 217567
rect 198913 199609 199031 199727
rect 199073 199609 199191 199727
rect 198913 199449 199031 199567
rect 199073 199449 199191 199567
rect 198913 181609 199031 181727
rect 199073 181609 199191 181727
rect 198913 181449 199031 181567
rect 199073 181449 199191 181567
rect 198913 163609 199031 163727
rect 199073 163609 199191 163727
rect 198913 163449 199031 163567
rect 199073 163449 199191 163567
rect 198913 145609 199031 145727
rect 199073 145609 199191 145727
rect 198913 145449 199031 145567
rect 199073 145449 199191 145567
rect 198913 127609 199031 127727
rect 199073 127609 199191 127727
rect 198913 127449 199031 127567
rect 199073 127449 199191 127567
rect 198913 109609 199031 109727
rect 199073 109609 199191 109727
rect 198913 109449 199031 109567
rect 199073 109449 199191 109567
rect 198913 91609 199031 91727
rect 199073 91609 199191 91727
rect 198913 91449 199031 91567
rect 199073 91449 199191 91567
rect 198913 73609 199031 73727
rect 199073 73609 199191 73727
rect 198913 73449 199031 73567
rect 199073 73449 199191 73567
rect 198913 55609 199031 55727
rect 199073 55609 199191 55727
rect 198913 55449 199031 55567
rect 199073 55449 199191 55567
rect 198913 37609 199031 37727
rect 199073 37609 199191 37727
rect 198913 37449 199031 37567
rect 199073 37449 199191 37567
rect 198913 19609 199031 19727
rect 199073 19609 199191 19727
rect 198913 19449 199031 19567
rect 199073 19449 199191 19567
rect 198913 1609 199031 1727
rect 199073 1609 199191 1727
rect 198913 1449 199031 1567
rect 199073 1449 199191 1567
rect 198913 -291 199031 -173
rect 199073 -291 199191 -173
rect 198913 -451 199031 -333
rect 199073 -451 199191 -333
rect 200773 345469 200891 345587
rect 200933 345469 201051 345587
rect 200773 345309 200891 345427
rect 200933 345309 201051 345427
rect 200773 327469 200891 327587
rect 200933 327469 201051 327587
rect 200773 327309 200891 327427
rect 200933 327309 201051 327427
rect 200773 309469 200891 309587
rect 200933 309469 201051 309587
rect 200773 309309 200891 309427
rect 200933 309309 201051 309427
rect 200773 291469 200891 291587
rect 200933 291469 201051 291587
rect 200773 291309 200891 291427
rect 200933 291309 201051 291427
rect 200773 273469 200891 273587
rect 200933 273469 201051 273587
rect 200773 273309 200891 273427
rect 200933 273309 201051 273427
rect 200773 255469 200891 255587
rect 200933 255469 201051 255587
rect 200773 255309 200891 255427
rect 200933 255309 201051 255427
rect 200773 237469 200891 237587
rect 200933 237469 201051 237587
rect 200773 237309 200891 237427
rect 200933 237309 201051 237427
rect 200773 219469 200891 219587
rect 200933 219469 201051 219587
rect 200773 219309 200891 219427
rect 200933 219309 201051 219427
rect 200773 201469 200891 201587
rect 200933 201469 201051 201587
rect 200773 201309 200891 201427
rect 200933 201309 201051 201427
rect 200773 183469 200891 183587
rect 200933 183469 201051 183587
rect 200773 183309 200891 183427
rect 200933 183309 201051 183427
rect 200773 165469 200891 165587
rect 200933 165469 201051 165587
rect 200773 165309 200891 165427
rect 200933 165309 201051 165427
rect 200773 147469 200891 147587
rect 200933 147469 201051 147587
rect 200773 147309 200891 147427
rect 200933 147309 201051 147427
rect 200773 129469 200891 129587
rect 200933 129469 201051 129587
rect 200773 129309 200891 129427
rect 200933 129309 201051 129427
rect 200773 111469 200891 111587
rect 200933 111469 201051 111587
rect 200773 111309 200891 111427
rect 200933 111309 201051 111427
rect 200773 93469 200891 93587
rect 200933 93469 201051 93587
rect 200773 93309 200891 93427
rect 200933 93309 201051 93427
rect 200773 75469 200891 75587
rect 200933 75469 201051 75587
rect 200773 75309 200891 75427
rect 200933 75309 201051 75427
rect 200773 57469 200891 57587
rect 200933 57469 201051 57587
rect 200773 57309 200891 57427
rect 200933 57309 201051 57427
rect 200773 39469 200891 39587
rect 200933 39469 201051 39587
rect 200773 39309 200891 39427
rect 200933 39309 201051 39427
rect 200773 21469 200891 21587
rect 200933 21469 201051 21587
rect 200773 21309 200891 21427
rect 200933 21309 201051 21427
rect 200773 3469 200891 3587
rect 200933 3469 201051 3587
rect 200773 3309 200891 3427
rect 200933 3309 201051 3427
rect 200773 -1251 200891 -1133
rect 200933 -1251 201051 -1133
rect 200773 -1411 200891 -1293
rect 200933 -1411 201051 -1293
rect 202633 347329 202751 347447
rect 202793 347329 202911 347447
rect 202633 347169 202751 347287
rect 202793 347169 202911 347287
rect 202633 329329 202751 329447
rect 202793 329329 202911 329447
rect 202633 329169 202751 329287
rect 202793 329169 202911 329287
rect 202633 311329 202751 311447
rect 202793 311329 202911 311447
rect 202633 311169 202751 311287
rect 202793 311169 202911 311287
rect 202633 293329 202751 293447
rect 202793 293329 202911 293447
rect 202633 293169 202751 293287
rect 202793 293169 202911 293287
rect 202633 275329 202751 275447
rect 202793 275329 202911 275447
rect 202633 275169 202751 275287
rect 202793 275169 202911 275287
rect 202633 257329 202751 257447
rect 202793 257329 202911 257447
rect 202633 257169 202751 257287
rect 202793 257169 202911 257287
rect 202633 239329 202751 239447
rect 202793 239329 202911 239447
rect 202633 239169 202751 239287
rect 202793 239169 202911 239287
rect 202633 221329 202751 221447
rect 202793 221329 202911 221447
rect 202633 221169 202751 221287
rect 202793 221169 202911 221287
rect 202633 203329 202751 203447
rect 202793 203329 202911 203447
rect 202633 203169 202751 203287
rect 202793 203169 202911 203287
rect 202633 185329 202751 185447
rect 202793 185329 202911 185447
rect 202633 185169 202751 185287
rect 202793 185169 202911 185287
rect 202633 167329 202751 167447
rect 202793 167329 202911 167447
rect 202633 167169 202751 167287
rect 202793 167169 202911 167287
rect 202633 149329 202751 149447
rect 202793 149329 202911 149447
rect 202633 149169 202751 149287
rect 202793 149169 202911 149287
rect 202633 131329 202751 131447
rect 202793 131329 202911 131447
rect 202633 131169 202751 131287
rect 202793 131169 202911 131287
rect 202633 113329 202751 113447
rect 202793 113329 202911 113447
rect 202633 113169 202751 113287
rect 202793 113169 202911 113287
rect 202633 95329 202751 95447
rect 202793 95329 202911 95447
rect 202633 95169 202751 95287
rect 202793 95169 202911 95287
rect 202633 77329 202751 77447
rect 202793 77329 202911 77447
rect 202633 77169 202751 77287
rect 202793 77169 202911 77287
rect 202633 59329 202751 59447
rect 202793 59329 202911 59447
rect 202633 59169 202751 59287
rect 202793 59169 202911 59287
rect 202633 41329 202751 41447
rect 202793 41329 202911 41447
rect 202633 41169 202751 41287
rect 202793 41169 202911 41287
rect 202633 23329 202751 23447
rect 202793 23329 202911 23447
rect 202633 23169 202751 23287
rect 202793 23169 202911 23287
rect 202633 5329 202751 5447
rect 202793 5329 202911 5447
rect 202633 5169 202751 5287
rect 202793 5169 202911 5287
rect 202633 -2211 202751 -2093
rect 202793 -2211 202911 -2093
rect 202633 -2371 202751 -2253
rect 202793 -2371 202911 -2253
rect 213493 355661 213611 355779
rect 213653 355661 213771 355779
rect 213493 355501 213611 355619
rect 213653 355501 213771 355619
rect 211633 354701 211751 354819
rect 211793 354701 211911 354819
rect 211633 354541 211751 354659
rect 211793 354541 211911 354659
rect 209773 353741 209891 353859
rect 209933 353741 210051 353859
rect 209773 353581 209891 353699
rect 209933 353581 210051 353699
rect 204493 349189 204611 349307
rect 204653 349189 204771 349307
rect 204493 349029 204611 349147
rect 204653 349029 204771 349147
rect 204493 331189 204611 331307
rect 204653 331189 204771 331307
rect 204493 331029 204611 331147
rect 204653 331029 204771 331147
rect 204493 313189 204611 313307
rect 204653 313189 204771 313307
rect 204493 313029 204611 313147
rect 204653 313029 204771 313147
rect 204493 295189 204611 295307
rect 204653 295189 204771 295307
rect 204493 295029 204611 295147
rect 204653 295029 204771 295147
rect 204493 277189 204611 277307
rect 204653 277189 204771 277307
rect 204493 277029 204611 277147
rect 204653 277029 204771 277147
rect 204493 259189 204611 259307
rect 204653 259189 204771 259307
rect 204493 259029 204611 259147
rect 204653 259029 204771 259147
rect 204493 241189 204611 241307
rect 204653 241189 204771 241307
rect 204493 241029 204611 241147
rect 204653 241029 204771 241147
rect 204493 223189 204611 223307
rect 204653 223189 204771 223307
rect 204493 223029 204611 223147
rect 204653 223029 204771 223147
rect 204493 205189 204611 205307
rect 204653 205189 204771 205307
rect 204493 205029 204611 205147
rect 204653 205029 204771 205147
rect 204493 187189 204611 187307
rect 204653 187189 204771 187307
rect 204493 187029 204611 187147
rect 204653 187029 204771 187147
rect 204493 169189 204611 169307
rect 204653 169189 204771 169307
rect 204493 169029 204611 169147
rect 204653 169029 204771 169147
rect 204493 151189 204611 151307
rect 204653 151189 204771 151307
rect 204493 151029 204611 151147
rect 204653 151029 204771 151147
rect 204493 133189 204611 133307
rect 204653 133189 204771 133307
rect 204493 133029 204611 133147
rect 204653 133029 204771 133147
rect 204493 115189 204611 115307
rect 204653 115189 204771 115307
rect 204493 115029 204611 115147
rect 204653 115029 204771 115147
rect 204493 97189 204611 97307
rect 204653 97189 204771 97307
rect 204493 97029 204611 97147
rect 204653 97029 204771 97147
rect 204493 79189 204611 79307
rect 204653 79189 204771 79307
rect 204493 79029 204611 79147
rect 204653 79029 204771 79147
rect 204493 61189 204611 61307
rect 204653 61189 204771 61307
rect 204493 61029 204611 61147
rect 204653 61029 204771 61147
rect 204493 43189 204611 43307
rect 204653 43189 204771 43307
rect 204493 43029 204611 43147
rect 204653 43029 204771 43147
rect 204493 25189 204611 25307
rect 204653 25189 204771 25307
rect 204493 25029 204611 25147
rect 204653 25029 204771 25147
rect 204493 7189 204611 7307
rect 204653 7189 204771 7307
rect 204493 7029 204611 7147
rect 204653 7029 204771 7147
rect 195493 -3651 195611 -3533
rect 195653 -3651 195771 -3533
rect 195493 -3811 195611 -3693
rect 195653 -3811 195771 -3693
rect 207913 352781 208031 352899
rect 208073 352781 208191 352899
rect 207913 352621 208031 352739
rect 208073 352621 208191 352739
rect 207913 334609 208031 334727
rect 208073 334609 208191 334727
rect 207913 334449 208031 334567
rect 208073 334449 208191 334567
rect 207913 316609 208031 316727
rect 208073 316609 208191 316727
rect 207913 316449 208031 316567
rect 208073 316449 208191 316567
rect 207913 298609 208031 298727
rect 208073 298609 208191 298727
rect 207913 298449 208031 298567
rect 208073 298449 208191 298567
rect 207913 280609 208031 280727
rect 208073 280609 208191 280727
rect 207913 280449 208031 280567
rect 208073 280449 208191 280567
rect 207913 262609 208031 262727
rect 208073 262609 208191 262727
rect 207913 262449 208031 262567
rect 208073 262449 208191 262567
rect 207913 244609 208031 244727
rect 208073 244609 208191 244727
rect 207913 244449 208031 244567
rect 208073 244449 208191 244567
rect 207913 226609 208031 226727
rect 208073 226609 208191 226727
rect 207913 226449 208031 226567
rect 208073 226449 208191 226567
rect 207913 208609 208031 208727
rect 208073 208609 208191 208727
rect 207913 208449 208031 208567
rect 208073 208449 208191 208567
rect 207913 190609 208031 190727
rect 208073 190609 208191 190727
rect 207913 190449 208031 190567
rect 208073 190449 208191 190567
rect 207913 172609 208031 172727
rect 208073 172609 208191 172727
rect 207913 172449 208031 172567
rect 208073 172449 208191 172567
rect 207913 154609 208031 154727
rect 208073 154609 208191 154727
rect 207913 154449 208031 154567
rect 208073 154449 208191 154567
rect 207913 136609 208031 136727
rect 208073 136609 208191 136727
rect 207913 136449 208031 136567
rect 208073 136449 208191 136567
rect 207913 118609 208031 118727
rect 208073 118609 208191 118727
rect 207913 118449 208031 118567
rect 208073 118449 208191 118567
rect 207913 100609 208031 100727
rect 208073 100609 208191 100727
rect 207913 100449 208031 100567
rect 208073 100449 208191 100567
rect 207913 82609 208031 82727
rect 208073 82609 208191 82727
rect 207913 82449 208031 82567
rect 208073 82449 208191 82567
rect 207913 64609 208031 64727
rect 208073 64609 208191 64727
rect 207913 64449 208031 64567
rect 208073 64449 208191 64567
rect 207913 46609 208031 46727
rect 208073 46609 208191 46727
rect 207913 46449 208031 46567
rect 208073 46449 208191 46567
rect 207913 28609 208031 28727
rect 208073 28609 208191 28727
rect 207913 28449 208031 28567
rect 208073 28449 208191 28567
rect 207913 10609 208031 10727
rect 208073 10609 208191 10727
rect 207913 10449 208031 10567
rect 208073 10449 208191 10567
rect 207913 -771 208031 -653
rect 208073 -771 208191 -653
rect 207913 -931 208031 -813
rect 208073 -931 208191 -813
rect 209773 336469 209891 336587
rect 209933 336469 210051 336587
rect 209773 336309 209891 336427
rect 209933 336309 210051 336427
rect 209773 318469 209891 318587
rect 209933 318469 210051 318587
rect 209773 318309 209891 318427
rect 209933 318309 210051 318427
rect 209773 300469 209891 300587
rect 209933 300469 210051 300587
rect 209773 300309 209891 300427
rect 209933 300309 210051 300427
rect 209773 282469 209891 282587
rect 209933 282469 210051 282587
rect 209773 282309 209891 282427
rect 209933 282309 210051 282427
rect 209773 264469 209891 264587
rect 209933 264469 210051 264587
rect 209773 264309 209891 264427
rect 209933 264309 210051 264427
rect 209773 246469 209891 246587
rect 209933 246469 210051 246587
rect 209773 246309 209891 246427
rect 209933 246309 210051 246427
rect 209773 228469 209891 228587
rect 209933 228469 210051 228587
rect 209773 228309 209891 228427
rect 209933 228309 210051 228427
rect 209773 210469 209891 210587
rect 209933 210469 210051 210587
rect 209773 210309 209891 210427
rect 209933 210309 210051 210427
rect 209773 192469 209891 192587
rect 209933 192469 210051 192587
rect 209773 192309 209891 192427
rect 209933 192309 210051 192427
rect 209773 174469 209891 174587
rect 209933 174469 210051 174587
rect 209773 174309 209891 174427
rect 209933 174309 210051 174427
rect 209773 156469 209891 156587
rect 209933 156469 210051 156587
rect 209773 156309 209891 156427
rect 209933 156309 210051 156427
rect 209773 138469 209891 138587
rect 209933 138469 210051 138587
rect 209773 138309 209891 138427
rect 209933 138309 210051 138427
rect 209773 120469 209891 120587
rect 209933 120469 210051 120587
rect 209773 120309 209891 120427
rect 209933 120309 210051 120427
rect 209773 102469 209891 102587
rect 209933 102469 210051 102587
rect 209773 102309 209891 102427
rect 209933 102309 210051 102427
rect 209773 84469 209891 84587
rect 209933 84469 210051 84587
rect 209773 84309 209891 84427
rect 209933 84309 210051 84427
rect 209773 66469 209891 66587
rect 209933 66469 210051 66587
rect 209773 66309 209891 66427
rect 209933 66309 210051 66427
rect 209773 48469 209891 48587
rect 209933 48469 210051 48587
rect 209773 48309 209891 48427
rect 209933 48309 210051 48427
rect 209773 30469 209891 30587
rect 209933 30469 210051 30587
rect 209773 30309 209891 30427
rect 209933 30309 210051 30427
rect 209773 12469 209891 12587
rect 209933 12469 210051 12587
rect 209773 12309 209891 12427
rect 209933 12309 210051 12427
rect 209773 -1731 209891 -1613
rect 209933 -1731 210051 -1613
rect 209773 -1891 209891 -1773
rect 209933 -1891 210051 -1773
rect 211633 338329 211751 338447
rect 211793 338329 211911 338447
rect 211633 338169 211751 338287
rect 211793 338169 211911 338287
rect 211633 320329 211751 320447
rect 211793 320329 211911 320447
rect 211633 320169 211751 320287
rect 211793 320169 211911 320287
rect 211633 302329 211751 302447
rect 211793 302329 211911 302447
rect 211633 302169 211751 302287
rect 211793 302169 211911 302287
rect 211633 284329 211751 284447
rect 211793 284329 211911 284447
rect 211633 284169 211751 284287
rect 211793 284169 211911 284287
rect 211633 266329 211751 266447
rect 211793 266329 211911 266447
rect 211633 266169 211751 266287
rect 211793 266169 211911 266287
rect 211633 248329 211751 248447
rect 211793 248329 211911 248447
rect 211633 248169 211751 248287
rect 211793 248169 211911 248287
rect 211633 230329 211751 230447
rect 211793 230329 211911 230447
rect 211633 230169 211751 230287
rect 211793 230169 211911 230287
rect 211633 212329 211751 212447
rect 211793 212329 211911 212447
rect 211633 212169 211751 212287
rect 211793 212169 211911 212287
rect 211633 194329 211751 194447
rect 211793 194329 211911 194447
rect 211633 194169 211751 194287
rect 211793 194169 211911 194287
rect 211633 176329 211751 176447
rect 211793 176329 211911 176447
rect 211633 176169 211751 176287
rect 211793 176169 211911 176287
rect 211633 158329 211751 158447
rect 211793 158329 211911 158447
rect 211633 158169 211751 158287
rect 211793 158169 211911 158287
rect 211633 140329 211751 140447
rect 211793 140329 211911 140447
rect 211633 140169 211751 140287
rect 211793 140169 211911 140287
rect 211633 122329 211751 122447
rect 211793 122329 211911 122447
rect 211633 122169 211751 122287
rect 211793 122169 211911 122287
rect 211633 104329 211751 104447
rect 211793 104329 211911 104447
rect 211633 104169 211751 104287
rect 211793 104169 211911 104287
rect 211633 86329 211751 86447
rect 211793 86329 211911 86447
rect 211633 86169 211751 86287
rect 211793 86169 211911 86287
rect 211633 68329 211751 68447
rect 211793 68329 211911 68447
rect 211633 68169 211751 68287
rect 211793 68169 211911 68287
rect 211633 50329 211751 50447
rect 211793 50329 211911 50447
rect 211633 50169 211751 50287
rect 211793 50169 211911 50287
rect 211633 32329 211751 32447
rect 211793 32329 211911 32447
rect 211633 32169 211751 32287
rect 211793 32169 211911 32287
rect 211633 14329 211751 14447
rect 211793 14329 211911 14447
rect 211633 14169 211751 14287
rect 211793 14169 211911 14287
rect 211633 -2691 211751 -2573
rect 211793 -2691 211911 -2573
rect 211633 -2851 211751 -2733
rect 211793 -2851 211911 -2733
rect 222493 355181 222611 355299
rect 222653 355181 222771 355299
rect 222493 355021 222611 355139
rect 222653 355021 222771 355139
rect 220633 354221 220751 354339
rect 220793 354221 220911 354339
rect 220633 354061 220751 354179
rect 220793 354061 220911 354179
rect 218773 353261 218891 353379
rect 218933 353261 219051 353379
rect 218773 353101 218891 353219
rect 218933 353101 219051 353219
rect 213493 340189 213611 340307
rect 213653 340189 213771 340307
rect 213493 340029 213611 340147
rect 213653 340029 213771 340147
rect 213493 322189 213611 322307
rect 213653 322189 213771 322307
rect 213493 322029 213611 322147
rect 213653 322029 213771 322147
rect 213493 304189 213611 304307
rect 213653 304189 213771 304307
rect 213493 304029 213611 304147
rect 213653 304029 213771 304147
rect 213493 286189 213611 286307
rect 213653 286189 213771 286307
rect 213493 286029 213611 286147
rect 213653 286029 213771 286147
rect 213493 268189 213611 268307
rect 213653 268189 213771 268307
rect 213493 268029 213611 268147
rect 213653 268029 213771 268147
rect 213493 250189 213611 250307
rect 213653 250189 213771 250307
rect 213493 250029 213611 250147
rect 213653 250029 213771 250147
rect 213493 232189 213611 232307
rect 213653 232189 213771 232307
rect 213493 232029 213611 232147
rect 213653 232029 213771 232147
rect 213493 214189 213611 214307
rect 213653 214189 213771 214307
rect 213493 214029 213611 214147
rect 213653 214029 213771 214147
rect 213493 196189 213611 196307
rect 213653 196189 213771 196307
rect 213493 196029 213611 196147
rect 213653 196029 213771 196147
rect 213493 178189 213611 178307
rect 213653 178189 213771 178307
rect 213493 178029 213611 178147
rect 213653 178029 213771 178147
rect 213493 160189 213611 160307
rect 213653 160189 213771 160307
rect 213493 160029 213611 160147
rect 213653 160029 213771 160147
rect 213493 142189 213611 142307
rect 213653 142189 213771 142307
rect 213493 142029 213611 142147
rect 213653 142029 213771 142147
rect 213493 124189 213611 124307
rect 213653 124189 213771 124307
rect 213493 124029 213611 124147
rect 213653 124029 213771 124147
rect 213493 106189 213611 106307
rect 213653 106189 213771 106307
rect 213493 106029 213611 106147
rect 213653 106029 213771 106147
rect 213493 88189 213611 88307
rect 213653 88189 213771 88307
rect 213493 88029 213611 88147
rect 213653 88029 213771 88147
rect 213493 70189 213611 70307
rect 213653 70189 213771 70307
rect 213493 70029 213611 70147
rect 213653 70029 213771 70147
rect 213493 52189 213611 52307
rect 213653 52189 213771 52307
rect 213493 52029 213611 52147
rect 213653 52029 213771 52147
rect 213493 34189 213611 34307
rect 213653 34189 213771 34307
rect 213493 34029 213611 34147
rect 213653 34029 213771 34147
rect 213493 16189 213611 16307
rect 213653 16189 213771 16307
rect 213493 16029 213611 16147
rect 213653 16029 213771 16147
rect 204493 -3171 204611 -3053
rect 204653 -3171 204771 -3053
rect 204493 -3331 204611 -3213
rect 204653 -3331 204771 -3213
rect 216913 352301 217031 352419
rect 217073 352301 217191 352419
rect 216913 352141 217031 352259
rect 217073 352141 217191 352259
rect 216913 343609 217031 343727
rect 217073 343609 217191 343727
rect 216913 343449 217031 343567
rect 217073 343449 217191 343567
rect 216913 325609 217031 325727
rect 217073 325609 217191 325727
rect 216913 325449 217031 325567
rect 217073 325449 217191 325567
rect 216913 307609 217031 307727
rect 217073 307609 217191 307727
rect 216913 307449 217031 307567
rect 217073 307449 217191 307567
rect 216913 289609 217031 289727
rect 217073 289609 217191 289727
rect 216913 289449 217031 289567
rect 217073 289449 217191 289567
rect 216913 271609 217031 271727
rect 217073 271609 217191 271727
rect 216913 271449 217031 271567
rect 217073 271449 217191 271567
rect 216913 253609 217031 253727
rect 217073 253609 217191 253727
rect 216913 253449 217031 253567
rect 217073 253449 217191 253567
rect 216913 235609 217031 235727
rect 217073 235609 217191 235727
rect 216913 235449 217031 235567
rect 217073 235449 217191 235567
rect 216913 217609 217031 217727
rect 217073 217609 217191 217727
rect 216913 217449 217031 217567
rect 217073 217449 217191 217567
rect 216913 199609 217031 199727
rect 217073 199609 217191 199727
rect 216913 199449 217031 199567
rect 217073 199449 217191 199567
rect 216913 181609 217031 181727
rect 217073 181609 217191 181727
rect 216913 181449 217031 181567
rect 217073 181449 217191 181567
rect 216913 163609 217031 163727
rect 217073 163609 217191 163727
rect 216913 163449 217031 163567
rect 217073 163449 217191 163567
rect 216913 145609 217031 145727
rect 217073 145609 217191 145727
rect 216913 145449 217031 145567
rect 217073 145449 217191 145567
rect 216913 127609 217031 127727
rect 217073 127609 217191 127727
rect 216913 127449 217031 127567
rect 217073 127449 217191 127567
rect 216913 109609 217031 109727
rect 217073 109609 217191 109727
rect 216913 109449 217031 109567
rect 217073 109449 217191 109567
rect 216913 91609 217031 91727
rect 217073 91609 217191 91727
rect 216913 91449 217031 91567
rect 217073 91449 217191 91567
rect 216913 73609 217031 73727
rect 217073 73609 217191 73727
rect 216913 73449 217031 73567
rect 217073 73449 217191 73567
rect 216913 55609 217031 55727
rect 217073 55609 217191 55727
rect 216913 55449 217031 55567
rect 217073 55449 217191 55567
rect 216913 37609 217031 37727
rect 217073 37609 217191 37727
rect 216913 37449 217031 37567
rect 217073 37449 217191 37567
rect 216913 19609 217031 19727
rect 217073 19609 217191 19727
rect 216913 19449 217031 19567
rect 217073 19449 217191 19567
rect 216913 1609 217031 1727
rect 217073 1609 217191 1727
rect 216913 1449 217031 1567
rect 217073 1449 217191 1567
rect 216913 -291 217031 -173
rect 217073 -291 217191 -173
rect 216913 -451 217031 -333
rect 217073 -451 217191 -333
rect 218773 345469 218891 345587
rect 218933 345469 219051 345587
rect 218773 345309 218891 345427
rect 218933 345309 219051 345427
rect 218773 327469 218891 327587
rect 218933 327469 219051 327587
rect 218773 327309 218891 327427
rect 218933 327309 219051 327427
rect 218773 309469 218891 309587
rect 218933 309469 219051 309587
rect 218773 309309 218891 309427
rect 218933 309309 219051 309427
rect 218773 291469 218891 291587
rect 218933 291469 219051 291587
rect 218773 291309 218891 291427
rect 218933 291309 219051 291427
rect 218773 273469 218891 273587
rect 218933 273469 219051 273587
rect 218773 273309 218891 273427
rect 218933 273309 219051 273427
rect 218773 255469 218891 255587
rect 218933 255469 219051 255587
rect 218773 255309 218891 255427
rect 218933 255309 219051 255427
rect 218773 237469 218891 237587
rect 218933 237469 219051 237587
rect 218773 237309 218891 237427
rect 218933 237309 219051 237427
rect 218773 219469 218891 219587
rect 218933 219469 219051 219587
rect 218773 219309 218891 219427
rect 218933 219309 219051 219427
rect 218773 201469 218891 201587
rect 218933 201469 219051 201587
rect 218773 201309 218891 201427
rect 218933 201309 219051 201427
rect 218773 183469 218891 183587
rect 218933 183469 219051 183587
rect 218773 183309 218891 183427
rect 218933 183309 219051 183427
rect 218773 165469 218891 165587
rect 218933 165469 219051 165587
rect 218773 165309 218891 165427
rect 218933 165309 219051 165427
rect 218773 147469 218891 147587
rect 218933 147469 219051 147587
rect 218773 147309 218891 147427
rect 218933 147309 219051 147427
rect 218773 129469 218891 129587
rect 218933 129469 219051 129587
rect 218773 129309 218891 129427
rect 218933 129309 219051 129427
rect 218773 111469 218891 111587
rect 218933 111469 219051 111587
rect 218773 111309 218891 111427
rect 218933 111309 219051 111427
rect 218773 93469 218891 93587
rect 218933 93469 219051 93587
rect 218773 93309 218891 93427
rect 218933 93309 219051 93427
rect 218773 75469 218891 75587
rect 218933 75469 219051 75587
rect 218773 75309 218891 75427
rect 218933 75309 219051 75427
rect 218773 57469 218891 57587
rect 218933 57469 219051 57587
rect 218773 57309 218891 57427
rect 218933 57309 219051 57427
rect 218773 39469 218891 39587
rect 218933 39469 219051 39587
rect 218773 39309 218891 39427
rect 218933 39309 219051 39427
rect 218773 21469 218891 21587
rect 218933 21469 219051 21587
rect 218773 21309 218891 21427
rect 218933 21309 219051 21427
rect 218773 3469 218891 3587
rect 218933 3469 219051 3587
rect 218773 3309 218891 3427
rect 218933 3309 219051 3427
rect 218773 -1251 218891 -1133
rect 218933 -1251 219051 -1133
rect 218773 -1411 218891 -1293
rect 218933 -1411 219051 -1293
rect 220633 347329 220751 347447
rect 220793 347329 220911 347447
rect 220633 347169 220751 347287
rect 220793 347169 220911 347287
rect 220633 329329 220751 329447
rect 220793 329329 220911 329447
rect 220633 329169 220751 329287
rect 220793 329169 220911 329287
rect 220633 311329 220751 311447
rect 220793 311329 220911 311447
rect 220633 311169 220751 311287
rect 220793 311169 220911 311287
rect 220633 293329 220751 293447
rect 220793 293329 220911 293447
rect 220633 293169 220751 293287
rect 220793 293169 220911 293287
rect 220633 275329 220751 275447
rect 220793 275329 220911 275447
rect 220633 275169 220751 275287
rect 220793 275169 220911 275287
rect 220633 257329 220751 257447
rect 220793 257329 220911 257447
rect 220633 257169 220751 257287
rect 220793 257169 220911 257287
rect 220633 239329 220751 239447
rect 220793 239329 220911 239447
rect 220633 239169 220751 239287
rect 220793 239169 220911 239287
rect 220633 221329 220751 221447
rect 220793 221329 220911 221447
rect 220633 221169 220751 221287
rect 220793 221169 220911 221287
rect 220633 203329 220751 203447
rect 220793 203329 220911 203447
rect 220633 203169 220751 203287
rect 220793 203169 220911 203287
rect 220633 185329 220751 185447
rect 220793 185329 220911 185447
rect 220633 185169 220751 185287
rect 220793 185169 220911 185287
rect 220633 167329 220751 167447
rect 220793 167329 220911 167447
rect 220633 167169 220751 167287
rect 220793 167169 220911 167287
rect 220633 149329 220751 149447
rect 220793 149329 220911 149447
rect 220633 149169 220751 149287
rect 220793 149169 220911 149287
rect 220633 131329 220751 131447
rect 220793 131329 220911 131447
rect 220633 131169 220751 131287
rect 220793 131169 220911 131287
rect 220633 113329 220751 113447
rect 220793 113329 220911 113447
rect 220633 113169 220751 113287
rect 220793 113169 220911 113287
rect 220633 95329 220751 95447
rect 220793 95329 220911 95447
rect 220633 95169 220751 95287
rect 220793 95169 220911 95287
rect 220633 77329 220751 77447
rect 220793 77329 220911 77447
rect 220633 77169 220751 77287
rect 220793 77169 220911 77287
rect 220633 59329 220751 59447
rect 220793 59329 220911 59447
rect 220633 59169 220751 59287
rect 220793 59169 220911 59287
rect 220633 41329 220751 41447
rect 220793 41329 220911 41447
rect 220633 41169 220751 41287
rect 220793 41169 220911 41287
rect 220633 23329 220751 23447
rect 220793 23329 220911 23447
rect 220633 23169 220751 23287
rect 220793 23169 220911 23287
rect 220633 5329 220751 5447
rect 220793 5329 220911 5447
rect 220633 5169 220751 5287
rect 220793 5169 220911 5287
rect 220633 -2211 220751 -2093
rect 220793 -2211 220911 -2093
rect 220633 -2371 220751 -2253
rect 220793 -2371 220911 -2253
rect 231493 355661 231611 355779
rect 231653 355661 231771 355779
rect 231493 355501 231611 355619
rect 231653 355501 231771 355619
rect 229633 354701 229751 354819
rect 229793 354701 229911 354819
rect 229633 354541 229751 354659
rect 229793 354541 229911 354659
rect 227773 353741 227891 353859
rect 227933 353741 228051 353859
rect 227773 353581 227891 353699
rect 227933 353581 228051 353699
rect 222493 349189 222611 349307
rect 222653 349189 222771 349307
rect 222493 349029 222611 349147
rect 222653 349029 222771 349147
rect 222493 331189 222611 331307
rect 222653 331189 222771 331307
rect 222493 331029 222611 331147
rect 222653 331029 222771 331147
rect 222493 313189 222611 313307
rect 222653 313189 222771 313307
rect 222493 313029 222611 313147
rect 222653 313029 222771 313147
rect 222493 295189 222611 295307
rect 222653 295189 222771 295307
rect 222493 295029 222611 295147
rect 222653 295029 222771 295147
rect 222493 277189 222611 277307
rect 222653 277189 222771 277307
rect 222493 277029 222611 277147
rect 222653 277029 222771 277147
rect 222493 259189 222611 259307
rect 222653 259189 222771 259307
rect 222493 259029 222611 259147
rect 222653 259029 222771 259147
rect 222493 241189 222611 241307
rect 222653 241189 222771 241307
rect 222493 241029 222611 241147
rect 222653 241029 222771 241147
rect 222493 223189 222611 223307
rect 222653 223189 222771 223307
rect 222493 223029 222611 223147
rect 222653 223029 222771 223147
rect 222493 205189 222611 205307
rect 222653 205189 222771 205307
rect 222493 205029 222611 205147
rect 222653 205029 222771 205147
rect 222493 187189 222611 187307
rect 222653 187189 222771 187307
rect 222493 187029 222611 187147
rect 222653 187029 222771 187147
rect 222493 169189 222611 169307
rect 222653 169189 222771 169307
rect 222493 169029 222611 169147
rect 222653 169029 222771 169147
rect 222493 151189 222611 151307
rect 222653 151189 222771 151307
rect 222493 151029 222611 151147
rect 222653 151029 222771 151147
rect 222493 133189 222611 133307
rect 222653 133189 222771 133307
rect 222493 133029 222611 133147
rect 222653 133029 222771 133147
rect 222493 115189 222611 115307
rect 222653 115189 222771 115307
rect 222493 115029 222611 115147
rect 222653 115029 222771 115147
rect 222493 97189 222611 97307
rect 222653 97189 222771 97307
rect 222493 97029 222611 97147
rect 222653 97029 222771 97147
rect 222493 79189 222611 79307
rect 222653 79189 222771 79307
rect 222493 79029 222611 79147
rect 222653 79029 222771 79147
rect 222493 61189 222611 61307
rect 222653 61189 222771 61307
rect 222493 61029 222611 61147
rect 222653 61029 222771 61147
rect 222493 43189 222611 43307
rect 222653 43189 222771 43307
rect 222493 43029 222611 43147
rect 222653 43029 222771 43147
rect 222493 25189 222611 25307
rect 222653 25189 222771 25307
rect 222493 25029 222611 25147
rect 222653 25029 222771 25147
rect 222493 7189 222611 7307
rect 222653 7189 222771 7307
rect 222493 7029 222611 7147
rect 222653 7029 222771 7147
rect 213493 -3651 213611 -3533
rect 213653 -3651 213771 -3533
rect 213493 -3811 213611 -3693
rect 213653 -3811 213771 -3693
rect 225913 352781 226031 352899
rect 226073 352781 226191 352899
rect 225913 352621 226031 352739
rect 226073 352621 226191 352739
rect 225913 334609 226031 334727
rect 226073 334609 226191 334727
rect 225913 334449 226031 334567
rect 226073 334449 226191 334567
rect 225913 316609 226031 316727
rect 226073 316609 226191 316727
rect 225913 316449 226031 316567
rect 226073 316449 226191 316567
rect 225913 298609 226031 298727
rect 226073 298609 226191 298727
rect 225913 298449 226031 298567
rect 226073 298449 226191 298567
rect 225913 280609 226031 280727
rect 226073 280609 226191 280727
rect 225913 280449 226031 280567
rect 226073 280449 226191 280567
rect 225913 262609 226031 262727
rect 226073 262609 226191 262727
rect 225913 262449 226031 262567
rect 226073 262449 226191 262567
rect 225913 244609 226031 244727
rect 226073 244609 226191 244727
rect 225913 244449 226031 244567
rect 226073 244449 226191 244567
rect 225913 226609 226031 226727
rect 226073 226609 226191 226727
rect 225913 226449 226031 226567
rect 226073 226449 226191 226567
rect 225913 208609 226031 208727
rect 226073 208609 226191 208727
rect 225913 208449 226031 208567
rect 226073 208449 226191 208567
rect 225913 190609 226031 190727
rect 226073 190609 226191 190727
rect 225913 190449 226031 190567
rect 226073 190449 226191 190567
rect 225913 172609 226031 172727
rect 226073 172609 226191 172727
rect 225913 172449 226031 172567
rect 226073 172449 226191 172567
rect 225913 154609 226031 154727
rect 226073 154609 226191 154727
rect 225913 154449 226031 154567
rect 226073 154449 226191 154567
rect 225913 136609 226031 136727
rect 226073 136609 226191 136727
rect 225913 136449 226031 136567
rect 226073 136449 226191 136567
rect 225913 118609 226031 118727
rect 226073 118609 226191 118727
rect 225913 118449 226031 118567
rect 226073 118449 226191 118567
rect 225913 100609 226031 100727
rect 226073 100609 226191 100727
rect 225913 100449 226031 100567
rect 226073 100449 226191 100567
rect 225913 82609 226031 82727
rect 226073 82609 226191 82727
rect 225913 82449 226031 82567
rect 226073 82449 226191 82567
rect 225913 64609 226031 64727
rect 226073 64609 226191 64727
rect 225913 64449 226031 64567
rect 226073 64449 226191 64567
rect 225913 46609 226031 46727
rect 226073 46609 226191 46727
rect 225913 46449 226031 46567
rect 226073 46449 226191 46567
rect 225913 28609 226031 28727
rect 226073 28609 226191 28727
rect 225913 28449 226031 28567
rect 226073 28449 226191 28567
rect 225913 10609 226031 10727
rect 226073 10609 226191 10727
rect 225913 10449 226031 10567
rect 226073 10449 226191 10567
rect 225913 -771 226031 -653
rect 226073 -771 226191 -653
rect 225913 -931 226031 -813
rect 226073 -931 226191 -813
rect 227773 336469 227891 336587
rect 227933 336469 228051 336587
rect 227773 336309 227891 336427
rect 227933 336309 228051 336427
rect 227773 318469 227891 318587
rect 227933 318469 228051 318587
rect 227773 318309 227891 318427
rect 227933 318309 228051 318427
rect 227773 300469 227891 300587
rect 227933 300469 228051 300587
rect 227773 300309 227891 300427
rect 227933 300309 228051 300427
rect 227773 282469 227891 282587
rect 227933 282469 228051 282587
rect 227773 282309 227891 282427
rect 227933 282309 228051 282427
rect 227773 264469 227891 264587
rect 227933 264469 228051 264587
rect 227773 264309 227891 264427
rect 227933 264309 228051 264427
rect 227773 246469 227891 246587
rect 227933 246469 228051 246587
rect 227773 246309 227891 246427
rect 227933 246309 228051 246427
rect 227773 228469 227891 228587
rect 227933 228469 228051 228587
rect 227773 228309 227891 228427
rect 227933 228309 228051 228427
rect 227773 210469 227891 210587
rect 227933 210469 228051 210587
rect 227773 210309 227891 210427
rect 227933 210309 228051 210427
rect 227773 192469 227891 192587
rect 227933 192469 228051 192587
rect 227773 192309 227891 192427
rect 227933 192309 228051 192427
rect 227773 174469 227891 174587
rect 227933 174469 228051 174587
rect 227773 174309 227891 174427
rect 227933 174309 228051 174427
rect 227773 156469 227891 156587
rect 227933 156469 228051 156587
rect 227773 156309 227891 156427
rect 227933 156309 228051 156427
rect 227773 138469 227891 138587
rect 227933 138469 228051 138587
rect 227773 138309 227891 138427
rect 227933 138309 228051 138427
rect 227773 120469 227891 120587
rect 227933 120469 228051 120587
rect 227773 120309 227891 120427
rect 227933 120309 228051 120427
rect 227773 102469 227891 102587
rect 227933 102469 228051 102587
rect 227773 102309 227891 102427
rect 227933 102309 228051 102427
rect 227773 84469 227891 84587
rect 227933 84469 228051 84587
rect 227773 84309 227891 84427
rect 227933 84309 228051 84427
rect 227773 66469 227891 66587
rect 227933 66469 228051 66587
rect 227773 66309 227891 66427
rect 227933 66309 228051 66427
rect 227773 48469 227891 48587
rect 227933 48469 228051 48587
rect 227773 48309 227891 48427
rect 227933 48309 228051 48427
rect 227773 30469 227891 30587
rect 227933 30469 228051 30587
rect 227773 30309 227891 30427
rect 227933 30309 228051 30427
rect 227773 12469 227891 12587
rect 227933 12469 228051 12587
rect 227773 12309 227891 12427
rect 227933 12309 228051 12427
rect 227773 -1731 227891 -1613
rect 227933 -1731 228051 -1613
rect 227773 -1891 227891 -1773
rect 227933 -1891 228051 -1773
rect 229633 338329 229751 338447
rect 229793 338329 229911 338447
rect 229633 338169 229751 338287
rect 229793 338169 229911 338287
rect 229633 320329 229751 320447
rect 229793 320329 229911 320447
rect 229633 320169 229751 320287
rect 229793 320169 229911 320287
rect 229633 302329 229751 302447
rect 229793 302329 229911 302447
rect 229633 302169 229751 302287
rect 229793 302169 229911 302287
rect 229633 284329 229751 284447
rect 229793 284329 229911 284447
rect 229633 284169 229751 284287
rect 229793 284169 229911 284287
rect 229633 266329 229751 266447
rect 229793 266329 229911 266447
rect 229633 266169 229751 266287
rect 229793 266169 229911 266287
rect 229633 248329 229751 248447
rect 229793 248329 229911 248447
rect 229633 248169 229751 248287
rect 229793 248169 229911 248287
rect 229633 230329 229751 230447
rect 229793 230329 229911 230447
rect 229633 230169 229751 230287
rect 229793 230169 229911 230287
rect 229633 212329 229751 212447
rect 229793 212329 229911 212447
rect 229633 212169 229751 212287
rect 229793 212169 229911 212287
rect 229633 194329 229751 194447
rect 229793 194329 229911 194447
rect 229633 194169 229751 194287
rect 229793 194169 229911 194287
rect 229633 176329 229751 176447
rect 229793 176329 229911 176447
rect 229633 176169 229751 176287
rect 229793 176169 229911 176287
rect 229633 158329 229751 158447
rect 229793 158329 229911 158447
rect 229633 158169 229751 158287
rect 229793 158169 229911 158287
rect 229633 140329 229751 140447
rect 229793 140329 229911 140447
rect 229633 140169 229751 140287
rect 229793 140169 229911 140287
rect 229633 122329 229751 122447
rect 229793 122329 229911 122447
rect 229633 122169 229751 122287
rect 229793 122169 229911 122287
rect 229633 104329 229751 104447
rect 229793 104329 229911 104447
rect 229633 104169 229751 104287
rect 229793 104169 229911 104287
rect 229633 86329 229751 86447
rect 229793 86329 229911 86447
rect 229633 86169 229751 86287
rect 229793 86169 229911 86287
rect 229633 68329 229751 68447
rect 229793 68329 229911 68447
rect 229633 68169 229751 68287
rect 229793 68169 229911 68287
rect 229633 50329 229751 50447
rect 229793 50329 229911 50447
rect 229633 50169 229751 50287
rect 229793 50169 229911 50287
rect 229633 32329 229751 32447
rect 229793 32329 229911 32447
rect 229633 32169 229751 32287
rect 229793 32169 229911 32287
rect 229633 14329 229751 14447
rect 229793 14329 229911 14447
rect 229633 14169 229751 14287
rect 229793 14169 229911 14287
rect 229633 -2691 229751 -2573
rect 229793 -2691 229911 -2573
rect 229633 -2851 229751 -2733
rect 229793 -2851 229911 -2733
rect 240493 355181 240611 355299
rect 240653 355181 240771 355299
rect 240493 355021 240611 355139
rect 240653 355021 240771 355139
rect 238633 354221 238751 354339
rect 238793 354221 238911 354339
rect 238633 354061 238751 354179
rect 238793 354061 238911 354179
rect 236773 353261 236891 353379
rect 236933 353261 237051 353379
rect 236773 353101 236891 353219
rect 236933 353101 237051 353219
rect 231493 340189 231611 340307
rect 231653 340189 231771 340307
rect 231493 340029 231611 340147
rect 231653 340029 231771 340147
rect 231493 322189 231611 322307
rect 231653 322189 231771 322307
rect 231493 322029 231611 322147
rect 231653 322029 231771 322147
rect 231493 304189 231611 304307
rect 231653 304189 231771 304307
rect 231493 304029 231611 304147
rect 231653 304029 231771 304147
rect 231493 286189 231611 286307
rect 231653 286189 231771 286307
rect 231493 286029 231611 286147
rect 231653 286029 231771 286147
rect 231493 268189 231611 268307
rect 231653 268189 231771 268307
rect 231493 268029 231611 268147
rect 231653 268029 231771 268147
rect 231493 250189 231611 250307
rect 231653 250189 231771 250307
rect 231493 250029 231611 250147
rect 231653 250029 231771 250147
rect 231493 232189 231611 232307
rect 231653 232189 231771 232307
rect 231493 232029 231611 232147
rect 231653 232029 231771 232147
rect 231493 214189 231611 214307
rect 231653 214189 231771 214307
rect 231493 214029 231611 214147
rect 231653 214029 231771 214147
rect 231493 196189 231611 196307
rect 231653 196189 231771 196307
rect 231493 196029 231611 196147
rect 231653 196029 231771 196147
rect 231493 178189 231611 178307
rect 231653 178189 231771 178307
rect 231493 178029 231611 178147
rect 231653 178029 231771 178147
rect 231493 160189 231611 160307
rect 231653 160189 231771 160307
rect 231493 160029 231611 160147
rect 231653 160029 231771 160147
rect 231493 142189 231611 142307
rect 231653 142189 231771 142307
rect 231493 142029 231611 142147
rect 231653 142029 231771 142147
rect 231493 124189 231611 124307
rect 231653 124189 231771 124307
rect 231493 124029 231611 124147
rect 231653 124029 231771 124147
rect 231493 106189 231611 106307
rect 231653 106189 231771 106307
rect 231493 106029 231611 106147
rect 231653 106029 231771 106147
rect 231493 88189 231611 88307
rect 231653 88189 231771 88307
rect 231493 88029 231611 88147
rect 231653 88029 231771 88147
rect 231493 70189 231611 70307
rect 231653 70189 231771 70307
rect 231493 70029 231611 70147
rect 231653 70029 231771 70147
rect 231493 52189 231611 52307
rect 231653 52189 231771 52307
rect 231493 52029 231611 52147
rect 231653 52029 231771 52147
rect 231493 34189 231611 34307
rect 231653 34189 231771 34307
rect 231493 34029 231611 34147
rect 231653 34029 231771 34147
rect 231493 16189 231611 16307
rect 231653 16189 231771 16307
rect 231493 16029 231611 16147
rect 231653 16029 231771 16147
rect 222493 -3171 222611 -3053
rect 222653 -3171 222771 -3053
rect 222493 -3331 222611 -3213
rect 222653 -3331 222771 -3213
rect 234913 352301 235031 352419
rect 235073 352301 235191 352419
rect 234913 352141 235031 352259
rect 235073 352141 235191 352259
rect 234913 343609 235031 343727
rect 235073 343609 235191 343727
rect 234913 343449 235031 343567
rect 235073 343449 235191 343567
rect 234913 325609 235031 325727
rect 235073 325609 235191 325727
rect 234913 325449 235031 325567
rect 235073 325449 235191 325567
rect 234913 307609 235031 307727
rect 235073 307609 235191 307727
rect 234913 307449 235031 307567
rect 235073 307449 235191 307567
rect 234913 289609 235031 289727
rect 235073 289609 235191 289727
rect 234913 289449 235031 289567
rect 235073 289449 235191 289567
rect 234913 271609 235031 271727
rect 235073 271609 235191 271727
rect 234913 271449 235031 271567
rect 235073 271449 235191 271567
rect 234913 253609 235031 253727
rect 235073 253609 235191 253727
rect 234913 253449 235031 253567
rect 235073 253449 235191 253567
rect 234913 235609 235031 235727
rect 235073 235609 235191 235727
rect 234913 235449 235031 235567
rect 235073 235449 235191 235567
rect 234913 217609 235031 217727
rect 235073 217609 235191 217727
rect 234913 217449 235031 217567
rect 235073 217449 235191 217567
rect 234913 199609 235031 199727
rect 235073 199609 235191 199727
rect 234913 199449 235031 199567
rect 235073 199449 235191 199567
rect 234913 181609 235031 181727
rect 235073 181609 235191 181727
rect 234913 181449 235031 181567
rect 235073 181449 235191 181567
rect 234913 163609 235031 163727
rect 235073 163609 235191 163727
rect 234913 163449 235031 163567
rect 235073 163449 235191 163567
rect 234913 145609 235031 145727
rect 235073 145609 235191 145727
rect 234913 145449 235031 145567
rect 235073 145449 235191 145567
rect 234913 127609 235031 127727
rect 235073 127609 235191 127727
rect 234913 127449 235031 127567
rect 235073 127449 235191 127567
rect 234913 109609 235031 109727
rect 235073 109609 235191 109727
rect 234913 109449 235031 109567
rect 235073 109449 235191 109567
rect 234913 91609 235031 91727
rect 235073 91609 235191 91727
rect 234913 91449 235031 91567
rect 235073 91449 235191 91567
rect 234913 73609 235031 73727
rect 235073 73609 235191 73727
rect 234913 73449 235031 73567
rect 235073 73449 235191 73567
rect 234913 55609 235031 55727
rect 235073 55609 235191 55727
rect 234913 55449 235031 55567
rect 235073 55449 235191 55567
rect 234913 37609 235031 37727
rect 235073 37609 235191 37727
rect 234913 37449 235031 37567
rect 235073 37449 235191 37567
rect 234913 19609 235031 19727
rect 235073 19609 235191 19727
rect 234913 19449 235031 19567
rect 235073 19449 235191 19567
rect 234913 1609 235031 1727
rect 235073 1609 235191 1727
rect 234913 1449 235031 1567
rect 235073 1449 235191 1567
rect 234913 -291 235031 -173
rect 235073 -291 235191 -173
rect 234913 -451 235031 -333
rect 235073 -451 235191 -333
rect 236773 345469 236891 345587
rect 236933 345469 237051 345587
rect 236773 345309 236891 345427
rect 236933 345309 237051 345427
rect 236773 327469 236891 327587
rect 236933 327469 237051 327587
rect 236773 327309 236891 327427
rect 236933 327309 237051 327427
rect 236773 309469 236891 309587
rect 236933 309469 237051 309587
rect 236773 309309 236891 309427
rect 236933 309309 237051 309427
rect 236773 291469 236891 291587
rect 236933 291469 237051 291587
rect 236773 291309 236891 291427
rect 236933 291309 237051 291427
rect 236773 273469 236891 273587
rect 236933 273469 237051 273587
rect 236773 273309 236891 273427
rect 236933 273309 237051 273427
rect 236773 255469 236891 255587
rect 236933 255469 237051 255587
rect 236773 255309 236891 255427
rect 236933 255309 237051 255427
rect 236773 237469 236891 237587
rect 236933 237469 237051 237587
rect 236773 237309 236891 237427
rect 236933 237309 237051 237427
rect 236773 219469 236891 219587
rect 236933 219469 237051 219587
rect 236773 219309 236891 219427
rect 236933 219309 237051 219427
rect 236773 201469 236891 201587
rect 236933 201469 237051 201587
rect 236773 201309 236891 201427
rect 236933 201309 237051 201427
rect 236773 183469 236891 183587
rect 236933 183469 237051 183587
rect 236773 183309 236891 183427
rect 236933 183309 237051 183427
rect 236773 165469 236891 165587
rect 236933 165469 237051 165587
rect 236773 165309 236891 165427
rect 236933 165309 237051 165427
rect 236773 147469 236891 147587
rect 236933 147469 237051 147587
rect 236773 147309 236891 147427
rect 236933 147309 237051 147427
rect 236773 129469 236891 129587
rect 236933 129469 237051 129587
rect 236773 129309 236891 129427
rect 236933 129309 237051 129427
rect 236773 111469 236891 111587
rect 236933 111469 237051 111587
rect 236773 111309 236891 111427
rect 236933 111309 237051 111427
rect 236773 93469 236891 93587
rect 236933 93469 237051 93587
rect 236773 93309 236891 93427
rect 236933 93309 237051 93427
rect 236773 75469 236891 75587
rect 236933 75469 237051 75587
rect 236773 75309 236891 75427
rect 236933 75309 237051 75427
rect 236773 57469 236891 57587
rect 236933 57469 237051 57587
rect 236773 57309 236891 57427
rect 236933 57309 237051 57427
rect 236773 39469 236891 39587
rect 236933 39469 237051 39587
rect 236773 39309 236891 39427
rect 236933 39309 237051 39427
rect 236773 21469 236891 21587
rect 236933 21469 237051 21587
rect 236773 21309 236891 21427
rect 236933 21309 237051 21427
rect 236773 3469 236891 3587
rect 236933 3469 237051 3587
rect 236773 3309 236891 3427
rect 236933 3309 237051 3427
rect 236773 -1251 236891 -1133
rect 236933 -1251 237051 -1133
rect 236773 -1411 236891 -1293
rect 236933 -1411 237051 -1293
rect 238633 347329 238751 347447
rect 238793 347329 238911 347447
rect 238633 347169 238751 347287
rect 238793 347169 238911 347287
rect 238633 329329 238751 329447
rect 238793 329329 238911 329447
rect 238633 329169 238751 329287
rect 238793 329169 238911 329287
rect 238633 311329 238751 311447
rect 238793 311329 238911 311447
rect 238633 311169 238751 311287
rect 238793 311169 238911 311287
rect 238633 293329 238751 293447
rect 238793 293329 238911 293447
rect 238633 293169 238751 293287
rect 238793 293169 238911 293287
rect 238633 275329 238751 275447
rect 238793 275329 238911 275447
rect 238633 275169 238751 275287
rect 238793 275169 238911 275287
rect 238633 257329 238751 257447
rect 238793 257329 238911 257447
rect 238633 257169 238751 257287
rect 238793 257169 238911 257287
rect 238633 239329 238751 239447
rect 238793 239329 238911 239447
rect 238633 239169 238751 239287
rect 238793 239169 238911 239287
rect 238633 221329 238751 221447
rect 238793 221329 238911 221447
rect 238633 221169 238751 221287
rect 238793 221169 238911 221287
rect 238633 203329 238751 203447
rect 238793 203329 238911 203447
rect 238633 203169 238751 203287
rect 238793 203169 238911 203287
rect 238633 185329 238751 185447
rect 238793 185329 238911 185447
rect 238633 185169 238751 185287
rect 238793 185169 238911 185287
rect 238633 167329 238751 167447
rect 238793 167329 238911 167447
rect 238633 167169 238751 167287
rect 238793 167169 238911 167287
rect 238633 149329 238751 149447
rect 238793 149329 238911 149447
rect 238633 149169 238751 149287
rect 238793 149169 238911 149287
rect 238633 131329 238751 131447
rect 238793 131329 238911 131447
rect 238633 131169 238751 131287
rect 238793 131169 238911 131287
rect 238633 113329 238751 113447
rect 238793 113329 238911 113447
rect 238633 113169 238751 113287
rect 238793 113169 238911 113287
rect 238633 95329 238751 95447
rect 238793 95329 238911 95447
rect 238633 95169 238751 95287
rect 238793 95169 238911 95287
rect 238633 77329 238751 77447
rect 238793 77329 238911 77447
rect 238633 77169 238751 77287
rect 238793 77169 238911 77287
rect 238633 59329 238751 59447
rect 238793 59329 238911 59447
rect 238633 59169 238751 59287
rect 238793 59169 238911 59287
rect 238633 41329 238751 41447
rect 238793 41329 238911 41447
rect 238633 41169 238751 41287
rect 238793 41169 238911 41287
rect 238633 23329 238751 23447
rect 238793 23329 238911 23447
rect 238633 23169 238751 23287
rect 238793 23169 238911 23287
rect 238633 5329 238751 5447
rect 238793 5329 238911 5447
rect 238633 5169 238751 5287
rect 238793 5169 238911 5287
rect 238633 -2211 238751 -2093
rect 238793 -2211 238911 -2093
rect 238633 -2371 238751 -2253
rect 238793 -2371 238911 -2253
rect 249493 355661 249611 355779
rect 249653 355661 249771 355779
rect 249493 355501 249611 355619
rect 249653 355501 249771 355619
rect 247633 354701 247751 354819
rect 247793 354701 247911 354819
rect 247633 354541 247751 354659
rect 247793 354541 247911 354659
rect 245773 353741 245891 353859
rect 245933 353741 246051 353859
rect 245773 353581 245891 353699
rect 245933 353581 246051 353699
rect 240493 349189 240611 349307
rect 240653 349189 240771 349307
rect 240493 349029 240611 349147
rect 240653 349029 240771 349147
rect 240493 331189 240611 331307
rect 240653 331189 240771 331307
rect 240493 331029 240611 331147
rect 240653 331029 240771 331147
rect 240493 313189 240611 313307
rect 240653 313189 240771 313307
rect 240493 313029 240611 313147
rect 240653 313029 240771 313147
rect 240493 295189 240611 295307
rect 240653 295189 240771 295307
rect 240493 295029 240611 295147
rect 240653 295029 240771 295147
rect 240493 277189 240611 277307
rect 240653 277189 240771 277307
rect 240493 277029 240611 277147
rect 240653 277029 240771 277147
rect 240493 259189 240611 259307
rect 240653 259189 240771 259307
rect 240493 259029 240611 259147
rect 240653 259029 240771 259147
rect 240493 241189 240611 241307
rect 240653 241189 240771 241307
rect 240493 241029 240611 241147
rect 240653 241029 240771 241147
rect 240493 223189 240611 223307
rect 240653 223189 240771 223307
rect 240493 223029 240611 223147
rect 240653 223029 240771 223147
rect 240493 205189 240611 205307
rect 240653 205189 240771 205307
rect 240493 205029 240611 205147
rect 240653 205029 240771 205147
rect 240493 187189 240611 187307
rect 240653 187189 240771 187307
rect 240493 187029 240611 187147
rect 240653 187029 240771 187147
rect 240493 169189 240611 169307
rect 240653 169189 240771 169307
rect 240493 169029 240611 169147
rect 240653 169029 240771 169147
rect 240493 151189 240611 151307
rect 240653 151189 240771 151307
rect 240493 151029 240611 151147
rect 240653 151029 240771 151147
rect 240493 133189 240611 133307
rect 240653 133189 240771 133307
rect 240493 133029 240611 133147
rect 240653 133029 240771 133147
rect 240493 115189 240611 115307
rect 240653 115189 240771 115307
rect 240493 115029 240611 115147
rect 240653 115029 240771 115147
rect 240493 97189 240611 97307
rect 240653 97189 240771 97307
rect 240493 97029 240611 97147
rect 240653 97029 240771 97147
rect 240493 79189 240611 79307
rect 240653 79189 240771 79307
rect 240493 79029 240611 79147
rect 240653 79029 240771 79147
rect 240493 61189 240611 61307
rect 240653 61189 240771 61307
rect 240493 61029 240611 61147
rect 240653 61029 240771 61147
rect 240493 43189 240611 43307
rect 240653 43189 240771 43307
rect 240493 43029 240611 43147
rect 240653 43029 240771 43147
rect 240493 25189 240611 25307
rect 240653 25189 240771 25307
rect 240493 25029 240611 25147
rect 240653 25029 240771 25147
rect 240493 7189 240611 7307
rect 240653 7189 240771 7307
rect 240493 7029 240611 7147
rect 240653 7029 240771 7147
rect 231493 -3651 231611 -3533
rect 231653 -3651 231771 -3533
rect 231493 -3811 231611 -3693
rect 231653 -3811 231771 -3693
rect 243913 352781 244031 352899
rect 244073 352781 244191 352899
rect 243913 352621 244031 352739
rect 244073 352621 244191 352739
rect 243913 334609 244031 334727
rect 244073 334609 244191 334727
rect 243913 334449 244031 334567
rect 244073 334449 244191 334567
rect 243913 316609 244031 316727
rect 244073 316609 244191 316727
rect 243913 316449 244031 316567
rect 244073 316449 244191 316567
rect 243913 298609 244031 298727
rect 244073 298609 244191 298727
rect 243913 298449 244031 298567
rect 244073 298449 244191 298567
rect 243913 280609 244031 280727
rect 244073 280609 244191 280727
rect 243913 280449 244031 280567
rect 244073 280449 244191 280567
rect 243913 262609 244031 262727
rect 244073 262609 244191 262727
rect 243913 262449 244031 262567
rect 244073 262449 244191 262567
rect 243913 244609 244031 244727
rect 244073 244609 244191 244727
rect 243913 244449 244031 244567
rect 244073 244449 244191 244567
rect 243913 226609 244031 226727
rect 244073 226609 244191 226727
rect 243913 226449 244031 226567
rect 244073 226449 244191 226567
rect 243913 208609 244031 208727
rect 244073 208609 244191 208727
rect 243913 208449 244031 208567
rect 244073 208449 244191 208567
rect 243913 190609 244031 190727
rect 244073 190609 244191 190727
rect 243913 190449 244031 190567
rect 244073 190449 244191 190567
rect 243913 172609 244031 172727
rect 244073 172609 244191 172727
rect 243913 172449 244031 172567
rect 244073 172449 244191 172567
rect 243913 154609 244031 154727
rect 244073 154609 244191 154727
rect 243913 154449 244031 154567
rect 244073 154449 244191 154567
rect 243913 136609 244031 136727
rect 244073 136609 244191 136727
rect 243913 136449 244031 136567
rect 244073 136449 244191 136567
rect 243913 118609 244031 118727
rect 244073 118609 244191 118727
rect 243913 118449 244031 118567
rect 244073 118449 244191 118567
rect 243913 100609 244031 100727
rect 244073 100609 244191 100727
rect 243913 100449 244031 100567
rect 244073 100449 244191 100567
rect 243913 82609 244031 82727
rect 244073 82609 244191 82727
rect 243913 82449 244031 82567
rect 244073 82449 244191 82567
rect 243913 64609 244031 64727
rect 244073 64609 244191 64727
rect 243913 64449 244031 64567
rect 244073 64449 244191 64567
rect 243913 46609 244031 46727
rect 244073 46609 244191 46727
rect 243913 46449 244031 46567
rect 244073 46449 244191 46567
rect 243913 28609 244031 28727
rect 244073 28609 244191 28727
rect 243913 28449 244031 28567
rect 244073 28449 244191 28567
rect 243913 10609 244031 10727
rect 244073 10609 244191 10727
rect 243913 10449 244031 10567
rect 244073 10449 244191 10567
rect 243913 -771 244031 -653
rect 244073 -771 244191 -653
rect 243913 -931 244031 -813
rect 244073 -931 244191 -813
rect 245773 336469 245891 336587
rect 245933 336469 246051 336587
rect 245773 336309 245891 336427
rect 245933 336309 246051 336427
rect 245773 318469 245891 318587
rect 245933 318469 246051 318587
rect 245773 318309 245891 318427
rect 245933 318309 246051 318427
rect 245773 300469 245891 300587
rect 245933 300469 246051 300587
rect 245773 300309 245891 300427
rect 245933 300309 246051 300427
rect 245773 282469 245891 282587
rect 245933 282469 246051 282587
rect 245773 282309 245891 282427
rect 245933 282309 246051 282427
rect 245773 264469 245891 264587
rect 245933 264469 246051 264587
rect 245773 264309 245891 264427
rect 245933 264309 246051 264427
rect 245773 246469 245891 246587
rect 245933 246469 246051 246587
rect 245773 246309 245891 246427
rect 245933 246309 246051 246427
rect 245773 228469 245891 228587
rect 245933 228469 246051 228587
rect 245773 228309 245891 228427
rect 245933 228309 246051 228427
rect 245773 210469 245891 210587
rect 245933 210469 246051 210587
rect 245773 210309 245891 210427
rect 245933 210309 246051 210427
rect 245773 192469 245891 192587
rect 245933 192469 246051 192587
rect 245773 192309 245891 192427
rect 245933 192309 246051 192427
rect 245773 174469 245891 174587
rect 245933 174469 246051 174587
rect 245773 174309 245891 174427
rect 245933 174309 246051 174427
rect 245773 156469 245891 156587
rect 245933 156469 246051 156587
rect 245773 156309 245891 156427
rect 245933 156309 246051 156427
rect 245773 138469 245891 138587
rect 245933 138469 246051 138587
rect 245773 138309 245891 138427
rect 245933 138309 246051 138427
rect 245773 120469 245891 120587
rect 245933 120469 246051 120587
rect 245773 120309 245891 120427
rect 245933 120309 246051 120427
rect 245773 102469 245891 102587
rect 245933 102469 246051 102587
rect 245773 102309 245891 102427
rect 245933 102309 246051 102427
rect 245773 84469 245891 84587
rect 245933 84469 246051 84587
rect 245773 84309 245891 84427
rect 245933 84309 246051 84427
rect 245773 66469 245891 66587
rect 245933 66469 246051 66587
rect 245773 66309 245891 66427
rect 245933 66309 246051 66427
rect 245773 48469 245891 48587
rect 245933 48469 246051 48587
rect 245773 48309 245891 48427
rect 245933 48309 246051 48427
rect 245773 30469 245891 30587
rect 245933 30469 246051 30587
rect 245773 30309 245891 30427
rect 245933 30309 246051 30427
rect 245773 12469 245891 12587
rect 245933 12469 246051 12587
rect 245773 12309 245891 12427
rect 245933 12309 246051 12427
rect 245773 -1731 245891 -1613
rect 245933 -1731 246051 -1613
rect 245773 -1891 245891 -1773
rect 245933 -1891 246051 -1773
rect 247633 338329 247751 338447
rect 247793 338329 247911 338447
rect 247633 338169 247751 338287
rect 247793 338169 247911 338287
rect 247633 320329 247751 320447
rect 247793 320329 247911 320447
rect 247633 320169 247751 320287
rect 247793 320169 247911 320287
rect 247633 302329 247751 302447
rect 247793 302329 247911 302447
rect 247633 302169 247751 302287
rect 247793 302169 247911 302287
rect 247633 284329 247751 284447
rect 247793 284329 247911 284447
rect 247633 284169 247751 284287
rect 247793 284169 247911 284287
rect 247633 266329 247751 266447
rect 247793 266329 247911 266447
rect 247633 266169 247751 266287
rect 247793 266169 247911 266287
rect 247633 248329 247751 248447
rect 247793 248329 247911 248447
rect 247633 248169 247751 248287
rect 247793 248169 247911 248287
rect 247633 230329 247751 230447
rect 247793 230329 247911 230447
rect 247633 230169 247751 230287
rect 247793 230169 247911 230287
rect 247633 212329 247751 212447
rect 247793 212329 247911 212447
rect 247633 212169 247751 212287
rect 247793 212169 247911 212287
rect 247633 194329 247751 194447
rect 247793 194329 247911 194447
rect 247633 194169 247751 194287
rect 247793 194169 247911 194287
rect 247633 176329 247751 176447
rect 247793 176329 247911 176447
rect 247633 176169 247751 176287
rect 247793 176169 247911 176287
rect 247633 158329 247751 158447
rect 247793 158329 247911 158447
rect 247633 158169 247751 158287
rect 247793 158169 247911 158287
rect 247633 140329 247751 140447
rect 247793 140329 247911 140447
rect 247633 140169 247751 140287
rect 247793 140169 247911 140287
rect 247633 122329 247751 122447
rect 247793 122329 247911 122447
rect 247633 122169 247751 122287
rect 247793 122169 247911 122287
rect 247633 104329 247751 104447
rect 247793 104329 247911 104447
rect 247633 104169 247751 104287
rect 247793 104169 247911 104287
rect 247633 86329 247751 86447
rect 247793 86329 247911 86447
rect 247633 86169 247751 86287
rect 247793 86169 247911 86287
rect 247633 68329 247751 68447
rect 247793 68329 247911 68447
rect 247633 68169 247751 68287
rect 247793 68169 247911 68287
rect 247633 50329 247751 50447
rect 247793 50329 247911 50447
rect 247633 50169 247751 50287
rect 247793 50169 247911 50287
rect 247633 32329 247751 32447
rect 247793 32329 247911 32447
rect 247633 32169 247751 32287
rect 247793 32169 247911 32287
rect 247633 14329 247751 14447
rect 247793 14329 247911 14447
rect 247633 14169 247751 14287
rect 247793 14169 247911 14287
rect 247633 -2691 247751 -2573
rect 247793 -2691 247911 -2573
rect 247633 -2851 247751 -2733
rect 247793 -2851 247911 -2733
rect 258493 355181 258611 355299
rect 258653 355181 258771 355299
rect 258493 355021 258611 355139
rect 258653 355021 258771 355139
rect 256633 354221 256751 354339
rect 256793 354221 256911 354339
rect 256633 354061 256751 354179
rect 256793 354061 256911 354179
rect 254773 353261 254891 353379
rect 254933 353261 255051 353379
rect 254773 353101 254891 353219
rect 254933 353101 255051 353219
rect 249493 340189 249611 340307
rect 249653 340189 249771 340307
rect 249493 340029 249611 340147
rect 249653 340029 249771 340147
rect 249493 322189 249611 322307
rect 249653 322189 249771 322307
rect 249493 322029 249611 322147
rect 249653 322029 249771 322147
rect 249493 304189 249611 304307
rect 249653 304189 249771 304307
rect 249493 304029 249611 304147
rect 249653 304029 249771 304147
rect 249493 286189 249611 286307
rect 249653 286189 249771 286307
rect 249493 286029 249611 286147
rect 249653 286029 249771 286147
rect 249493 268189 249611 268307
rect 249653 268189 249771 268307
rect 249493 268029 249611 268147
rect 249653 268029 249771 268147
rect 249493 250189 249611 250307
rect 249653 250189 249771 250307
rect 249493 250029 249611 250147
rect 249653 250029 249771 250147
rect 249493 232189 249611 232307
rect 249653 232189 249771 232307
rect 249493 232029 249611 232147
rect 249653 232029 249771 232147
rect 249493 214189 249611 214307
rect 249653 214189 249771 214307
rect 249493 214029 249611 214147
rect 249653 214029 249771 214147
rect 249493 196189 249611 196307
rect 249653 196189 249771 196307
rect 249493 196029 249611 196147
rect 249653 196029 249771 196147
rect 249493 178189 249611 178307
rect 249653 178189 249771 178307
rect 249493 178029 249611 178147
rect 249653 178029 249771 178147
rect 249493 160189 249611 160307
rect 249653 160189 249771 160307
rect 249493 160029 249611 160147
rect 249653 160029 249771 160147
rect 249493 142189 249611 142307
rect 249653 142189 249771 142307
rect 249493 142029 249611 142147
rect 249653 142029 249771 142147
rect 249493 124189 249611 124307
rect 249653 124189 249771 124307
rect 249493 124029 249611 124147
rect 249653 124029 249771 124147
rect 249493 106189 249611 106307
rect 249653 106189 249771 106307
rect 249493 106029 249611 106147
rect 249653 106029 249771 106147
rect 249493 88189 249611 88307
rect 249653 88189 249771 88307
rect 249493 88029 249611 88147
rect 249653 88029 249771 88147
rect 249493 70189 249611 70307
rect 249653 70189 249771 70307
rect 249493 70029 249611 70147
rect 249653 70029 249771 70147
rect 249493 52189 249611 52307
rect 249653 52189 249771 52307
rect 249493 52029 249611 52147
rect 249653 52029 249771 52147
rect 249493 34189 249611 34307
rect 249653 34189 249771 34307
rect 249493 34029 249611 34147
rect 249653 34029 249771 34147
rect 249493 16189 249611 16307
rect 249653 16189 249771 16307
rect 249493 16029 249611 16147
rect 249653 16029 249771 16147
rect 240493 -3171 240611 -3053
rect 240653 -3171 240771 -3053
rect 240493 -3331 240611 -3213
rect 240653 -3331 240771 -3213
rect 252913 352301 253031 352419
rect 253073 352301 253191 352419
rect 252913 352141 253031 352259
rect 253073 352141 253191 352259
rect 252913 343609 253031 343727
rect 253073 343609 253191 343727
rect 252913 343449 253031 343567
rect 253073 343449 253191 343567
rect 252913 325609 253031 325727
rect 253073 325609 253191 325727
rect 252913 325449 253031 325567
rect 253073 325449 253191 325567
rect 252913 307609 253031 307727
rect 253073 307609 253191 307727
rect 252913 307449 253031 307567
rect 253073 307449 253191 307567
rect 252913 289609 253031 289727
rect 253073 289609 253191 289727
rect 252913 289449 253031 289567
rect 253073 289449 253191 289567
rect 252913 271609 253031 271727
rect 253073 271609 253191 271727
rect 252913 271449 253031 271567
rect 253073 271449 253191 271567
rect 252913 253609 253031 253727
rect 253073 253609 253191 253727
rect 252913 253449 253031 253567
rect 253073 253449 253191 253567
rect 252913 235609 253031 235727
rect 253073 235609 253191 235727
rect 252913 235449 253031 235567
rect 253073 235449 253191 235567
rect 252913 217609 253031 217727
rect 253073 217609 253191 217727
rect 252913 217449 253031 217567
rect 253073 217449 253191 217567
rect 252913 199609 253031 199727
rect 253073 199609 253191 199727
rect 252913 199449 253031 199567
rect 253073 199449 253191 199567
rect 252913 181609 253031 181727
rect 253073 181609 253191 181727
rect 252913 181449 253031 181567
rect 253073 181449 253191 181567
rect 252913 163609 253031 163727
rect 253073 163609 253191 163727
rect 252913 163449 253031 163567
rect 253073 163449 253191 163567
rect 252913 145609 253031 145727
rect 253073 145609 253191 145727
rect 252913 145449 253031 145567
rect 253073 145449 253191 145567
rect 252913 127609 253031 127727
rect 253073 127609 253191 127727
rect 252913 127449 253031 127567
rect 253073 127449 253191 127567
rect 252913 109609 253031 109727
rect 253073 109609 253191 109727
rect 252913 109449 253031 109567
rect 253073 109449 253191 109567
rect 252913 91609 253031 91727
rect 253073 91609 253191 91727
rect 252913 91449 253031 91567
rect 253073 91449 253191 91567
rect 252913 73609 253031 73727
rect 253073 73609 253191 73727
rect 252913 73449 253031 73567
rect 253073 73449 253191 73567
rect 252913 55609 253031 55727
rect 253073 55609 253191 55727
rect 252913 55449 253031 55567
rect 253073 55449 253191 55567
rect 252913 37609 253031 37727
rect 253073 37609 253191 37727
rect 252913 37449 253031 37567
rect 253073 37449 253191 37567
rect 252913 19609 253031 19727
rect 253073 19609 253191 19727
rect 252913 19449 253031 19567
rect 253073 19449 253191 19567
rect 252913 1609 253031 1727
rect 253073 1609 253191 1727
rect 252913 1449 253031 1567
rect 253073 1449 253191 1567
rect 252913 -291 253031 -173
rect 253073 -291 253191 -173
rect 252913 -451 253031 -333
rect 253073 -451 253191 -333
rect 254773 345469 254891 345587
rect 254933 345469 255051 345587
rect 254773 345309 254891 345427
rect 254933 345309 255051 345427
rect 254773 327469 254891 327587
rect 254933 327469 255051 327587
rect 254773 327309 254891 327427
rect 254933 327309 255051 327427
rect 254773 309469 254891 309587
rect 254933 309469 255051 309587
rect 254773 309309 254891 309427
rect 254933 309309 255051 309427
rect 254773 291469 254891 291587
rect 254933 291469 255051 291587
rect 254773 291309 254891 291427
rect 254933 291309 255051 291427
rect 254773 273469 254891 273587
rect 254933 273469 255051 273587
rect 254773 273309 254891 273427
rect 254933 273309 255051 273427
rect 254773 255469 254891 255587
rect 254933 255469 255051 255587
rect 254773 255309 254891 255427
rect 254933 255309 255051 255427
rect 254773 237469 254891 237587
rect 254933 237469 255051 237587
rect 254773 237309 254891 237427
rect 254933 237309 255051 237427
rect 254773 219469 254891 219587
rect 254933 219469 255051 219587
rect 254773 219309 254891 219427
rect 254933 219309 255051 219427
rect 254773 201469 254891 201587
rect 254933 201469 255051 201587
rect 254773 201309 254891 201427
rect 254933 201309 255051 201427
rect 254773 183469 254891 183587
rect 254933 183469 255051 183587
rect 254773 183309 254891 183427
rect 254933 183309 255051 183427
rect 254773 165469 254891 165587
rect 254933 165469 255051 165587
rect 254773 165309 254891 165427
rect 254933 165309 255051 165427
rect 254773 147469 254891 147587
rect 254933 147469 255051 147587
rect 254773 147309 254891 147427
rect 254933 147309 255051 147427
rect 254773 129469 254891 129587
rect 254933 129469 255051 129587
rect 254773 129309 254891 129427
rect 254933 129309 255051 129427
rect 254773 111469 254891 111587
rect 254933 111469 255051 111587
rect 254773 111309 254891 111427
rect 254933 111309 255051 111427
rect 254773 93469 254891 93587
rect 254933 93469 255051 93587
rect 254773 93309 254891 93427
rect 254933 93309 255051 93427
rect 254773 75469 254891 75587
rect 254933 75469 255051 75587
rect 254773 75309 254891 75427
rect 254933 75309 255051 75427
rect 254773 57469 254891 57587
rect 254933 57469 255051 57587
rect 254773 57309 254891 57427
rect 254933 57309 255051 57427
rect 254773 39469 254891 39587
rect 254933 39469 255051 39587
rect 254773 39309 254891 39427
rect 254933 39309 255051 39427
rect 254773 21469 254891 21587
rect 254933 21469 255051 21587
rect 254773 21309 254891 21427
rect 254933 21309 255051 21427
rect 254773 3469 254891 3587
rect 254933 3469 255051 3587
rect 254773 3309 254891 3427
rect 254933 3309 255051 3427
rect 254773 -1251 254891 -1133
rect 254933 -1251 255051 -1133
rect 254773 -1411 254891 -1293
rect 254933 -1411 255051 -1293
rect 256633 347329 256751 347447
rect 256793 347329 256911 347447
rect 256633 347169 256751 347287
rect 256793 347169 256911 347287
rect 256633 329329 256751 329447
rect 256793 329329 256911 329447
rect 256633 329169 256751 329287
rect 256793 329169 256911 329287
rect 256633 311329 256751 311447
rect 256793 311329 256911 311447
rect 256633 311169 256751 311287
rect 256793 311169 256911 311287
rect 256633 293329 256751 293447
rect 256793 293329 256911 293447
rect 256633 293169 256751 293287
rect 256793 293169 256911 293287
rect 256633 275329 256751 275447
rect 256793 275329 256911 275447
rect 256633 275169 256751 275287
rect 256793 275169 256911 275287
rect 256633 257329 256751 257447
rect 256793 257329 256911 257447
rect 256633 257169 256751 257287
rect 256793 257169 256911 257287
rect 256633 239329 256751 239447
rect 256793 239329 256911 239447
rect 256633 239169 256751 239287
rect 256793 239169 256911 239287
rect 256633 221329 256751 221447
rect 256793 221329 256911 221447
rect 256633 221169 256751 221287
rect 256793 221169 256911 221287
rect 256633 203329 256751 203447
rect 256793 203329 256911 203447
rect 256633 203169 256751 203287
rect 256793 203169 256911 203287
rect 256633 185329 256751 185447
rect 256793 185329 256911 185447
rect 256633 185169 256751 185287
rect 256793 185169 256911 185287
rect 256633 167329 256751 167447
rect 256793 167329 256911 167447
rect 256633 167169 256751 167287
rect 256793 167169 256911 167287
rect 256633 149329 256751 149447
rect 256793 149329 256911 149447
rect 256633 149169 256751 149287
rect 256793 149169 256911 149287
rect 256633 131329 256751 131447
rect 256793 131329 256911 131447
rect 256633 131169 256751 131287
rect 256793 131169 256911 131287
rect 256633 113329 256751 113447
rect 256793 113329 256911 113447
rect 256633 113169 256751 113287
rect 256793 113169 256911 113287
rect 256633 95329 256751 95447
rect 256793 95329 256911 95447
rect 256633 95169 256751 95287
rect 256793 95169 256911 95287
rect 256633 77329 256751 77447
rect 256793 77329 256911 77447
rect 256633 77169 256751 77287
rect 256793 77169 256911 77287
rect 256633 59329 256751 59447
rect 256793 59329 256911 59447
rect 256633 59169 256751 59287
rect 256793 59169 256911 59287
rect 256633 41329 256751 41447
rect 256793 41329 256911 41447
rect 256633 41169 256751 41287
rect 256793 41169 256911 41287
rect 256633 23329 256751 23447
rect 256793 23329 256911 23447
rect 256633 23169 256751 23287
rect 256793 23169 256911 23287
rect 256633 5329 256751 5447
rect 256793 5329 256911 5447
rect 256633 5169 256751 5287
rect 256793 5169 256911 5287
rect 256633 -2211 256751 -2093
rect 256793 -2211 256911 -2093
rect 256633 -2371 256751 -2253
rect 256793 -2371 256911 -2253
rect 267493 355661 267611 355779
rect 267653 355661 267771 355779
rect 267493 355501 267611 355619
rect 267653 355501 267771 355619
rect 265633 354701 265751 354819
rect 265793 354701 265911 354819
rect 265633 354541 265751 354659
rect 265793 354541 265911 354659
rect 263773 353741 263891 353859
rect 263933 353741 264051 353859
rect 263773 353581 263891 353699
rect 263933 353581 264051 353699
rect 258493 349189 258611 349307
rect 258653 349189 258771 349307
rect 258493 349029 258611 349147
rect 258653 349029 258771 349147
rect 258493 331189 258611 331307
rect 258653 331189 258771 331307
rect 258493 331029 258611 331147
rect 258653 331029 258771 331147
rect 258493 313189 258611 313307
rect 258653 313189 258771 313307
rect 258493 313029 258611 313147
rect 258653 313029 258771 313147
rect 258493 295189 258611 295307
rect 258653 295189 258771 295307
rect 258493 295029 258611 295147
rect 258653 295029 258771 295147
rect 258493 277189 258611 277307
rect 258653 277189 258771 277307
rect 258493 277029 258611 277147
rect 258653 277029 258771 277147
rect 258493 259189 258611 259307
rect 258653 259189 258771 259307
rect 258493 259029 258611 259147
rect 258653 259029 258771 259147
rect 258493 241189 258611 241307
rect 258653 241189 258771 241307
rect 258493 241029 258611 241147
rect 258653 241029 258771 241147
rect 258493 223189 258611 223307
rect 258653 223189 258771 223307
rect 258493 223029 258611 223147
rect 258653 223029 258771 223147
rect 258493 205189 258611 205307
rect 258653 205189 258771 205307
rect 258493 205029 258611 205147
rect 258653 205029 258771 205147
rect 258493 187189 258611 187307
rect 258653 187189 258771 187307
rect 258493 187029 258611 187147
rect 258653 187029 258771 187147
rect 258493 169189 258611 169307
rect 258653 169189 258771 169307
rect 258493 169029 258611 169147
rect 258653 169029 258771 169147
rect 258493 151189 258611 151307
rect 258653 151189 258771 151307
rect 258493 151029 258611 151147
rect 258653 151029 258771 151147
rect 258493 133189 258611 133307
rect 258653 133189 258771 133307
rect 258493 133029 258611 133147
rect 258653 133029 258771 133147
rect 258493 115189 258611 115307
rect 258653 115189 258771 115307
rect 258493 115029 258611 115147
rect 258653 115029 258771 115147
rect 258493 97189 258611 97307
rect 258653 97189 258771 97307
rect 258493 97029 258611 97147
rect 258653 97029 258771 97147
rect 258493 79189 258611 79307
rect 258653 79189 258771 79307
rect 258493 79029 258611 79147
rect 258653 79029 258771 79147
rect 258493 61189 258611 61307
rect 258653 61189 258771 61307
rect 258493 61029 258611 61147
rect 258653 61029 258771 61147
rect 258493 43189 258611 43307
rect 258653 43189 258771 43307
rect 258493 43029 258611 43147
rect 258653 43029 258771 43147
rect 258493 25189 258611 25307
rect 258653 25189 258771 25307
rect 258493 25029 258611 25147
rect 258653 25029 258771 25147
rect 258493 7189 258611 7307
rect 258653 7189 258771 7307
rect 258493 7029 258611 7147
rect 258653 7029 258771 7147
rect 249493 -3651 249611 -3533
rect 249653 -3651 249771 -3533
rect 249493 -3811 249611 -3693
rect 249653 -3811 249771 -3693
rect 261913 352781 262031 352899
rect 262073 352781 262191 352899
rect 261913 352621 262031 352739
rect 262073 352621 262191 352739
rect 261913 334609 262031 334727
rect 262073 334609 262191 334727
rect 261913 334449 262031 334567
rect 262073 334449 262191 334567
rect 261913 316609 262031 316727
rect 262073 316609 262191 316727
rect 261913 316449 262031 316567
rect 262073 316449 262191 316567
rect 261913 298609 262031 298727
rect 262073 298609 262191 298727
rect 261913 298449 262031 298567
rect 262073 298449 262191 298567
rect 261913 280609 262031 280727
rect 262073 280609 262191 280727
rect 261913 280449 262031 280567
rect 262073 280449 262191 280567
rect 261913 262609 262031 262727
rect 262073 262609 262191 262727
rect 261913 262449 262031 262567
rect 262073 262449 262191 262567
rect 261913 244609 262031 244727
rect 262073 244609 262191 244727
rect 261913 244449 262031 244567
rect 262073 244449 262191 244567
rect 261913 226609 262031 226727
rect 262073 226609 262191 226727
rect 261913 226449 262031 226567
rect 262073 226449 262191 226567
rect 261913 208609 262031 208727
rect 262073 208609 262191 208727
rect 261913 208449 262031 208567
rect 262073 208449 262191 208567
rect 261913 190609 262031 190727
rect 262073 190609 262191 190727
rect 261913 190449 262031 190567
rect 262073 190449 262191 190567
rect 261913 172609 262031 172727
rect 262073 172609 262191 172727
rect 261913 172449 262031 172567
rect 262073 172449 262191 172567
rect 261913 154609 262031 154727
rect 262073 154609 262191 154727
rect 261913 154449 262031 154567
rect 262073 154449 262191 154567
rect 261913 136609 262031 136727
rect 262073 136609 262191 136727
rect 261913 136449 262031 136567
rect 262073 136449 262191 136567
rect 261913 118609 262031 118727
rect 262073 118609 262191 118727
rect 261913 118449 262031 118567
rect 262073 118449 262191 118567
rect 261913 100609 262031 100727
rect 262073 100609 262191 100727
rect 261913 100449 262031 100567
rect 262073 100449 262191 100567
rect 261913 82609 262031 82727
rect 262073 82609 262191 82727
rect 261913 82449 262031 82567
rect 262073 82449 262191 82567
rect 261913 64609 262031 64727
rect 262073 64609 262191 64727
rect 261913 64449 262031 64567
rect 262073 64449 262191 64567
rect 261913 46609 262031 46727
rect 262073 46609 262191 46727
rect 261913 46449 262031 46567
rect 262073 46449 262191 46567
rect 261913 28609 262031 28727
rect 262073 28609 262191 28727
rect 261913 28449 262031 28567
rect 262073 28449 262191 28567
rect 261913 10609 262031 10727
rect 262073 10609 262191 10727
rect 261913 10449 262031 10567
rect 262073 10449 262191 10567
rect 261913 -771 262031 -653
rect 262073 -771 262191 -653
rect 261913 -931 262031 -813
rect 262073 -931 262191 -813
rect 263773 336469 263891 336587
rect 263933 336469 264051 336587
rect 263773 336309 263891 336427
rect 263933 336309 264051 336427
rect 263773 318469 263891 318587
rect 263933 318469 264051 318587
rect 263773 318309 263891 318427
rect 263933 318309 264051 318427
rect 263773 300469 263891 300587
rect 263933 300469 264051 300587
rect 263773 300309 263891 300427
rect 263933 300309 264051 300427
rect 263773 282469 263891 282587
rect 263933 282469 264051 282587
rect 263773 282309 263891 282427
rect 263933 282309 264051 282427
rect 263773 264469 263891 264587
rect 263933 264469 264051 264587
rect 263773 264309 263891 264427
rect 263933 264309 264051 264427
rect 263773 246469 263891 246587
rect 263933 246469 264051 246587
rect 263773 246309 263891 246427
rect 263933 246309 264051 246427
rect 263773 228469 263891 228587
rect 263933 228469 264051 228587
rect 263773 228309 263891 228427
rect 263933 228309 264051 228427
rect 263773 210469 263891 210587
rect 263933 210469 264051 210587
rect 263773 210309 263891 210427
rect 263933 210309 264051 210427
rect 263773 192469 263891 192587
rect 263933 192469 264051 192587
rect 263773 192309 263891 192427
rect 263933 192309 264051 192427
rect 263773 174469 263891 174587
rect 263933 174469 264051 174587
rect 263773 174309 263891 174427
rect 263933 174309 264051 174427
rect 263773 156469 263891 156587
rect 263933 156469 264051 156587
rect 263773 156309 263891 156427
rect 263933 156309 264051 156427
rect 263773 138469 263891 138587
rect 263933 138469 264051 138587
rect 263773 138309 263891 138427
rect 263933 138309 264051 138427
rect 263773 120469 263891 120587
rect 263933 120469 264051 120587
rect 263773 120309 263891 120427
rect 263933 120309 264051 120427
rect 263773 102469 263891 102587
rect 263933 102469 264051 102587
rect 263773 102309 263891 102427
rect 263933 102309 264051 102427
rect 263773 84469 263891 84587
rect 263933 84469 264051 84587
rect 263773 84309 263891 84427
rect 263933 84309 264051 84427
rect 263773 66469 263891 66587
rect 263933 66469 264051 66587
rect 263773 66309 263891 66427
rect 263933 66309 264051 66427
rect 263773 48469 263891 48587
rect 263933 48469 264051 48587
rect 263773 48309 263891 48427
rect 263933 48309 264051 48427
rect 263773 30469 263891 30587
rect 263933 30469 264051 30587
rect 263773 30309 263891 30427
rect 263933 30309 264051 30427
rect 263773 12469 263891 12587
rect 263933 12469 264051 12587
rect 263773 12309 263891 12427
rect 263933 12309 264051 12427
rect 263773 -1731 263891 -1613
rect 263933 -1731 264051 -1613
rect 263773 -1891 263891 -1773
rect 263933 -1891 264051 -1773
rect 265633 338329 265751 338447
rect 265793 338329 265911 338447
rect 265633 338169 265751 338287
rect 265793 338169 265911 338287
rect 265633 320329 265751 320447
rect 265793 320329 265911 320447
rect 265633 320169 265751 320287
rect 265793 320169 265911 320287
rect 265633 302329 265751 302447
rect 265793 302329 265911 302447
rect 265633 302169 265751 302287
rect 265793 302169 265911 302287
rect 265633 284329 265751 284447
rect 265793 284329 265911 284447
rect 265633 284169 265751 284287
rect 265793 284169 265911 284287
rect 265633 266329 265751 266447
rect 265793 266329 265911 266447
rect 265633 266169 265751 266287
rect 265793 266169 265911 266287
rect 265633 248329 265751 248447
rect 265793 248329 265911 248447
rect 265633 248169 265751 248287
rect 265793 248169 265911 248287
rect 265633 230329 265751 230447
rect 265793 230329 265911 230447
rect 265633 230169 265751 230287
rect 265793 230169 265911 230287
rect 265633 212329 265751 212447
rect 265793 212329 265911 212447
rect 265633 212169 265751 212287
rect 265793 212169 265911 212287
rect 265633 194329 265751 194447
rect 265793 194329 265911 194447
rect 265633 194169 265751 194287
rect 265793 194169 265911 194287
rect 265633 176329 265751 176447
rect 265793 176329 265911 176447
rect 265633 176169 265751 176287
rect 265793 176169 265911 176287
rect 265633 158329 265751 158447
rect 265793 158329 265911 158447
rect 265633 158169 265751 158287
rect 265793 158169 265911 158287
rect 265633 140329 265751 140447
rect 265793 140329 265911 140447
rect 265633 140169 265751 140287
rect 265793 140169 265911 140287
rect 265633 122329 265751 122447
rect 265793 122329 265911 122447
rect 265633 122169 265751 122287
rect 265793 122169 265911 122287
rect 265633 104329 265751 104447
rect 265793 104329 265911 104447
rect 265633 104169 265751 104287
rect 265793 104169 265911 104287
rect 265633 86329 265751 86447
rect 265793 86329 265911 86447
rect 265633 86169 265751 86287
rect 265793 86169 265911 86287
rect 265633 68329 265751 68447
rect 265793 68329 265911 68447
rect 265633 68169 265751 68287
rect 265793 68169 265911 68287
rect 265633 50329 265751 50447
rect 265793 50329 265911 50447
rect 265633 50169 265751 50287
rect 265793 50169 265911 50287
rect 265633 32329 265751 32447
rect 265793 32329 265911 32447
rect 265633 32169 265751 32287
rect 265793 32169 265911 32287
rect 265633 14329 265751 14447
rect 265793 14329 265911 14447
rect 265633 14169 265751 14287
rect 265793 14169 265911 14287
rect 265633 -2691 265751 -2573
rect 265793 -2691 265911 -2573
rect 265633 -2851 265751 -2733
rect 265793 -2851 265911 -2733
rect 276493 355181 276611 355299
rect 276653 355181 276771 355299
rect 276493 355021 276611 355139
rect 276653 355021 276771 355139
rect 274633 354221 274751 354339
rect 274793 354221 274911 354339
rect 274633 354061 274751 354179
rect 274793 354061 274911 354179
rect 272773 353261 272891 353379
rect 272933 353261 273051 353379
rect 272773 353101 272891 353219
rect 272933 353101 273051 353219
rect 267493 340189 267611 340307
rect 267653 340189 267771 340307
rect 267493 340029 267611 340147
rect 267653 340029 267771 340147
rect 267493 322189 267611 322307
rect 267653 322189 267771 322307
rect 267493 322029 267611 322147
rect 267653 322029 267771 322147
rect 267493 304189 267611 304307
rect 267653 304189 267771 304307
rect 267493 304029 267611 304147
rect 267653 304029 267771 304147
rect 267493 286189 267611 286307
rect 267653 286189 267771 286307
rect 267493 286029 267611 286147
rect 267653 286029 267771 286147
rect 267493 268189 267611 268307
rect 267653 268189 267771 268307
rect 267493 268029 267611 268147
rect 267653 268029 267771 268147
rect 267493 250189 267611 250307
rect 267653 250189 267771 250307
rect 267493 250029 267611 250147
rect 267653 250029 267771 250147
rect 267493 232189 267611 232307
rect 267653 232189 267771 232307
rect 267493 232029 267611 232147
rect 267653 232029 267771 232147
rect 267493 214189 267611 214307
rect 267653 214189 267771 214307
rect 267493 214029 267611 214147
rect 267653 214029 267771 214147
rect 267493 196189 267611 196307
rect 267653 196189 267771 196307
rect 267493 196029 267611 196147
rect 267653 196029 267771 196147
rect 267493 178189 267611 178307
rect 267653 178189 267771 178307
rect 267493 178029 267611 178147
rect 267653 178029 267771 178147
rect 267493 160189 267611 160307
rect 267653 160189 267771 160307
rect 267493 160029 267611 160147
rect 267653 160029 267771 160147
rect 267493 142189 267611 142307
rect 267653 142189 267771 142307
rect 267493 142029 267611 142147
rect 267653 142029 267771 142147
rect 267493 124189 267611 124307
rect 267653 124189 267771 124307
rect 267493 124029 267611 124147
rect 267653 124029 267771 124147
rect 267493 106189 267611 106307
rect 267653 106189 267771 106307
rect 267493 106029 267611 106147
rect 267653 106029 267771 106147
rect 267493 88189 267611 88307
rect 267653 88189 267771 88307
rect 267493 88029 267611 88147
rect 267653 88029 267771 88147
rect 267493 70189 267611 70307
rect 267653 70189 267771 70307
rect 267493 70029 267611 70147
rect 267653 70029 267771 70147
rect 267493 52189 267611 52307
rect 267653 52189 267771 52307
rect 267493 52029 267611 52147
rect 267653 52029 267771 52147
rect 267493 34189 267611 34307
rect 267653 34189 267771 34307
rect 267493 34029 267611 34147
rect 267653 34029 267771 34147
rect 267493 16189 267611 16307
rect 267653 16189 267771 16307
rect 267493 16029 267611 16147
rect 267653 16029 267771 16147
rect 258493 -3171 258611 -3053
rect 258653 -3171 258771 -3053
rect 258493 -3331 258611 -3213
rect 258653 -3331 258771 -3213
rect 270913 352301 271031 352419
rect 271073 352301 271191 352419
rect 270913 352141 271031 352259
rect 271073 352141 271191 352259
rect 270913 343609 271031 343727
rect 271073 343609 271191 343727
rect 270913 343449 271031 343567
rect 271073 343449 271191 343567
rect 270913 325609 271031 325727
rect 271073 325609 271191 325727
rect 270913 325449 271031 325567
rect 271073 325449 271191 325567
rect 270913 307609 271031 307727
rect 271073 307609 271191 307727
rect 270913 307449 271031 307567
rect 271073 307449 271191 307567
rect 270913 289609 271031 289727
rect 271073 289609 271191 289727
rect 270913 289449 271031 289567
rect 271073 289449 271191 289567
rect 270913 271609 271031 271727
rect 271073 271609 271191 271727
rect 270913 271449 271031 271567
rect 271073 271449 271191 271567
rect 270913 253609 271031 253727
rect 271073 253609 271191 253727
rect 270913 253449 271031 253567
rect 271073 253449 271191 253567
rect 270913 235609 271031 235727
rect 271073 235609 271191 235727
rect 270913 235449 271031 235567
rect 271073 235449 271191 235567
rect 270913 217609 271031 217727
rect 271073 217609 271191 217727
rect 270913 217449 271031 217567
rect 271073 217449 271191 217567
rect 270913 199609 271031 199727
rect 271073 199609 271191 199727
rect 270913 199449 271031 199567
rect 271073 199449 271191 199567
rect 270913 181609 271031 181727
rect 271073 181609 271191 181727
rect 270913 181449 271031 181567
rect 271073 181449 271191 181567
rect 270913 163609 271031 163727
rect 271073 163609 271191 163727
rect 270913 163449 271031 163567
rect 271073 163449 271191 163567
rect 270913 145609 271031 145727
rect 271073 145609 271191 145727
rect 270913 145449 271031 145567
rect 271073 145449 271191 145567
rect 270913 127609 271031 127727
rect 271073 127609 271191 127727
rect 270913 127449 271031 127567
rect 271073 127449 271191 127567
rect 270913 109609 271031 109727
rect 271073 109609 271191 109727
rect 270913 109449 271031 109567
rect 271073 109449 271191 109567
rect 270913 91609 271031 91727
rect 271073 91609 271191 91727
rect 270913 91449 271031 91567
rect 271073 91449 271191 91567
rect 270913 73609 271031 73727
rect 271073 73609 271191 73727
rect 270913 73449 271031 73567
rect 271073 73449 271191 73567
rect 270913 55609 271031 55727
rect 271073 55609 271191 55727
rect 270913 55449 271031 55567
rect 271073 55449 271191 55567
rect 270913 37609 271031 37727
rect 271073 37609 271191 37727
rect 270913 37449 271031 37567
rect 271073 37449 271191 37567
rect 270913 19609 271031 19727
rect 271073 19609 271191 19727
rect 270913 19449 271031 19567
rect 271073 19449 271191 19567
rect 270913 1609 271031 1727
rect 271073 1609 271191 1727
rect 270913 1449 271031 1567
rect 271073 1449 271191 1567
rect 270913 -291 271031 -173
rect 271073 -291 271191 -173
rect 270913 -451 271031 -333
rect 271073 -451 271191 -333
rect 272773 345469 272891 345587
rect 272933 345469 273051 345587
rect 272773 345309 272891 345427
rect 272933 345309 273051 345427
rect 272773 327469 272891 327587
rect 272933 327469 273051 327587
rect 272773 327309 272891 327427
rect 272933 327309 273051 327427
rect 272773 309469 272891 309587
rect 272933 309469 273051 309587
rect 272773 309309 272891 309427
rect 272933 309309 273051 309427
rect 272773 291469 272891 291587
rect 272933 291469 273051 291587
rect 272773 291309 272891 291427
rect 272933 291309 273051 291427
rect 272773 273469 272891 273587
rect 272933 273469 273051 273587
rect 272773 273309 272891 273427
rect 272933 273309 273051 273427
rect 272773 255469 272891 255587
rect 272933 255469 273051 255587
rect 272773 255309 272891 255427
rect 272933 255309 273051 255427
rect 272773 237469 272891 237587
rect 272933 237469 273051 237587
rect 272773 237309 272891 237427
rect 272933 237309 273051 237427
rect 272773 219469 272891 219587
rect 272933 219469 273051 219587
rect 272773 219309 272891 219427
rect 272933 219309 273051 219427
rect 272773 201469 272891 201587
rect 272933 201469 273051 201587
rect 272773 201309 272891 201427
rect 272933 201309 273051 201427
rect 272773 183469 272891 183587
rect 272933 183469 273051 183587
rect 272773 183309 272891 183427
rect 272933 183309 273051 183427
rect 272773 165469 272891 165587
rect 272933 165469 273051 165587
rect 272773 165309 272891 165427
rect 272933 165309 273051 165427
rect 272773 147469 272891 147587
rect 272933 147469 273051 147587
rect 272773 147309 272891 147427
rect 272933 147309 273051 147427
rect 272773 129469 272891 129587
rect 272933 129469 273051 129587
rect 272773 129309 272891 129427
rect 272933 129309 273051 129427
rect 272773 111469 272891 111587
rect 272933 111469 273051 111587
rect 272773 111309 272891 111427
rect 272933 111309 273051 111427
rect 272773 93469 272891 93587
rect 272933 93469 273051 93587
rect 272773 93309 272891 93427
rect 272933 93309 273051 93427
rect 272773 75469 272891 75587
rect 272933 75469 273051 75587
rect 272773 75309 272891 75427
rect 272933 75309 273051 75427
rect 272773 57469 272891 57587
rect 272933 57469 273051 57587
rect 272773 57309 272891 57427
rect 272933 57309 273051 57427
rect 272773 39469 272891 39587
rect 272933 39469 273051 39587
rect 272773 39309 272891 39427
rect 272933 39309 273051 39427
rect 272773 21469 272891 21587
rect 272933 21469 273051 21587
rect 272773 21309 272891 21427
rect 272933 21309 273051 21427
rect 272773 3469 272891 3587
rect 272933 3469 273051 3587
rect 272773 3309 272891 3427
rect 272933 3309 273051 3427
rect 272773 -1251 272891 -1133
rect 272933 -1251 273051 -1133
rect 272773 -1411 272891 -1293
rect 272933 -1411 273051 -1293
rect 274633 347329 274751 347447
rect 274793 347329 274911 347447
rect 274633 347169 274751 347287
rect 274793 347169 274911 347287
rect 274633 329329 274751 329447
rect 274793 329329 274911 329447
rect 274633 329169 274751 329287
rect 274793 329169 274911 329287
rect 274633 311329 274751 311447
rect 274793 311329 274911 311447
rect 274633 311169 274751 311287
rect 274793 311169 274911 311287
rect 274633 293329 274751 293447
rect 274793 293329 274911 293447
rect 274633 293169 274751 293287
rect 274793 293169 274911 293287
rect 274633 275329 274751 275447
rect 274793 275329 274911 275447
rect 274633 275169 274751 275287
rect 274793 275169 274911 275287
rect 274633 257329 274751 257447
rect 274793 257329 274911 257447
rect 274633 257169 274751 257287
rect 274793 257169 274911 257287
rect 274633 239329 274751 239447
rect 274793 239329 274911 239447
rect 274633 239169 274751 239287
rect 274793 239169 274911 239287
rect 274633 221329 274751 221447
rect 274793 221329 274911 221447
rect 274633 221169 274751 221287
rect 274793 221169 274911 221287
rect 274633 203329 274751 203447
rect 274793 203329 274911 203447
rect 274633 203169 274751 203287
rect 274793 203169 274911 203287
rect 274633 185329 274751 185447
rect 274793 185329 274911 185447
rect 274633 185169 274751 185287
rect 274793 185169 274911 185287
rect 274633 167329 274751 167447
rect 274793 167329 274911 167447
rect 274633 167169 274751 167287
rect 274793 167169 274911 167287
rect 274633 149329 274751 149447
rect 274793 149329 274911 149447
rect 274633 149169 274751 149287
rect 274793 149169 274911 149287
rect 274633 131329 274751 131447
rect 274793 131329 274911 131447
rect 274633 131169 274751 131287
rect 274793 131169 274911 131287
rect 274633 113329 274751 113447
rect 274793 113329 274911 113447
rect 274633 113169 274751 113287
rect 274793 113169 274911 113287
rect 274633 95329 274751 95447
rect 274793 95329 274911 95447
rect 274633 95169 274751 95287
rect 274793 95169 274911 95287
rect 274633 77329 274751 77447
rect 274793 77329 274911 77447
rect 274633 77169 274751 77287
rect 274793 77169 274911 77287
rect 274633 59329 274751 59447
rect 274793 59329 274911 59447
rect 274633 59169 274751 59287
rect 274793 59169 274911 59287
rect 274633 41329 274751 41447
rect 274793 41329 274911 41447
rect 274633 41169 274751 41287
rect 274793 41169 274911 41287
rect 274633 23329 274751 23447
rect 274793 23329 274911 23447
rect 274633 23169 274751 23287
rect 274793 23169 274911 23287
rect 274633 5329 274751 5447
rect 274793 5329 274911 5447
rect 274633 5169 274751 5287
rect 274793 5169 274911 5287
rect 274633 -2211 274751 -2093
rect 274793 -2211 274911 -2093
rect 274633 -2371 274751 -2253
rect 274793 -2371 274911 -2253
rect 285493 355661 285611 355779
rect 285653 355661 285771 355779
rect 285493 355501 285611 355619
rect 285653 355501 285771 355619
rect 283633 354701 283751 354819
rect 283793 354701 283911 354819
rect 283633 354541 283751 354659
rect 283793 354541 283911 354659
rect 281773 353741 281891 353859
rect 281933 353741 282051 353859
rect 281773 353581 281891 353699
rect 281933 353581 282051 353699
rect 276493 349189 276611 349307
rect 276653 349189 276771 349307
rect 276493 349029 276611 349147
rect 276653 349029 276771 349147
rect 276493 331189 276611 331307
rect 276653 331189 276771 331307
rect 276493 331029 276611 331147
rect 276653 331029 276771 331147
rect 276493 313189 276611 313307
rect 276653 313189 276771 313307
rect 276493 313029 276611 313147
rect 276653 313029 276771 313147
rect 276493 295189 276611 295307
rect 276653 295189 276771 295307
rect 276493 295029 276611 295147
rect 276653 295029 276771 295147
rect 276493 277189 276611 277307
rect 276653 277189 276771 277307
rect 276493 277029 276611 277147
rect 276653 277029 276771 277147
rect 276493 259189 276611 259307
rect 276653 259189 276771 259307
rect 276493 259029 276611 259147
rect 276653 259029 276771 259147
rect 276493 241189 276611 241307
rect 276653 241189 276771 241307
rect 276493 241029 276611 241147
rect 276653 241029 276771 241147
rect 276493 223189 276611 223307
rect 276653 223189 276771 223307
rect 276493 223029 276611 223147
rect 276653 223029 276771 223147
rect 276493 205189 276611 205307
rect 276653 205189 276771 205307
rect 276493 205029 276611 205147
rect 276653 205029 276771 205147
rect 276493 187189 276611 187307
rect 276653 187189 276771 187307
rect 276493 187029 276611 187147
rect 276653 187029 276771 187147
rect 276493 169189 276611 169307
rect 276653 169189 276771 169307
rect 276493 169029 276611 169147
rect 276653 169029 276771 169147
rect 276493 151189 276611 151307
rect 276653 151189 276771 151307
rect 276493 151029 276611 151147
rect 276653 151029 276771 151147
rect 276493 133189 276611 133307
rect 276653 133189 276771 133307
rect 276493 133029 276611 133147
rect 276653 133029 276771 133147
rect 276493 115189 276611 115307
rect 276653 115189 276771 115307
rect 276493 115029 276611 115147
rect 276653 115029 276771 115147
rect 276493 97189 276611 97307
rect 276653 97189 276771 97307
rect 276493 97029 276611 97147
rect 276653 97029 276771 97147
rect 276493 79189 276611 79307
rect 276653 79189 276771 79307
rect 276493 79029 276611 79147
rect 276653 79029 276771 79147
rect 276493 61189 276611 61307
rect 276653 61189 276771 61307
rect 276493 61029 276611 61147
rect 276653 61029 276771 61147
rect 276493 43189 276611 43307
rect 276653 43189 276771 43307
rect 276493 43029 276611 43147
rect 276653 43029 276771 43147
rect 276493 25189 276611 25307
rect 276653 25189 276771 25307
rect 276493 25029 276611 25147
rect 276653 25029 276771 25147
rect 276493 7189 276611 7307
rect 276653 7189 276771 7307
rect 276493 7029 276611 7147
rect 276653 7029 276771 7147
rect 267493 -3651 267611 -3533
rect 267653 -3651 267771 -3533
rect 267493 -3811 267611 -3693
rect 267653 -3811 267771 -3693
rect 279913 352781 280031 352899
rect 280073 352781 280191 352899
rect 279913 352621 280031 352739
rect 280073 352621 280191 352739
rect 279913 334609 280031 334727
rect 280073 334609 280191 334727
rect 279913 334449 280031 334567
rect 280073 334449 280191 334567
rect 279913 316609 280031 316727
rect 280073 316609 280191 316727
rect 279913 316449 280031 316567
rect 280073 316449 280191 316567
rect 279913 298609 280031 298727
rect 280073 298609 280191 298727
rect 279913 298449 280031 298567
rect 280073 298449 280191 298567
rect 279913 280609 280031 280727
rect 280073 280609 280191 280727
rect 279913 280449 280031 280567
rect 280073 280449 280191 280567
rect 279913 262609 280031 262727
rect 280073 262609 280191 262727
rect 279913 262449 280031 262567
rect 280073 262449 280191 262567
rect 279913 244609 280031 244727
rect 280073 244609 280191 244727
rect 279913 244449 280031 244567
rect 280073 244449 280191 244567
rect 279913 226609 280031 226727
rect 280073 226609 280191 226727
rect 279913 226449 280031 226567
rect 280073 226449 280191 226567
rect 279913 208609 280031 208727
rect 280073 208609 280191 208727
rect 279913 208449 280031 208567
rect 280073 208449 280191 208567
rect 279913 190609 280031 190727
rect 280073 190609 280191 190727
rect 279913 190449 280031 190567
rect 280073 190449 280191 190567
rect 279913 172609 280031 172727
rect 280073 172609 280191 172727
rect 279913 172449 280031 172567
rect 280073 172449 280191 172567
rect 279913 154609 280031 154727
rect 280073 154609 280191 154727
rect 279913 154449 280031 154567
rect 280073 154449 280191 154567
rect 279913 136609 280031 136727
rect 280073 136609 280191 136727
rect 279913 136449 280031 136567
rect 280073 136449 280191 136567
rect 279913 118609 280031 118727
rect 280073 118609 280191 118727
rect 279913 118449 280031 118567
rect 280073 118449 280191 118567
rect 279913 100609 280031 100727
rect 280073 100609 280191 100727
rect 279913 100449 280031 100567
rect 280073 100449 280191 100567
rect 279913 82609 280031 82727
rect 280073 82609 280191 82727
rect 279913 82449 280031 82567
rect 280073 82449 280191 82567
rect 279913 64609 280031 64727
rect 280073 64609 280191 64727
rect 279913 64449 280031 64567
rect 280073 64449 280191 64567
rect 279913 46609 280031 46727
rect 280073 46609 280191 46727
rect 279913 46449 280031 46567
rect 280073 46449 280191 46567
rect 279913 28609 280031 28727
rect 280073 28609 280191 28727
rect 279913 28449 280031 28567
rect 280073 28449 280191 28567
rect 279913 10609 280031 10727
rect 280073 10609 280191 10727
rect 279913 10449 280031 10567
rect 280073 10449 280191 10567
rect 279913 -771 280031 -653
rect 280073 -771 280191 -653
rect 279913 -931 280031 -813
rect 280073 -931 280191 -813
rect 281773 336469 281891 336587
rect 281933 336469 282051 336587
rect 281773 336309 281891 336427
rect 281933 336309 282051 336427
rect 281773 318469 281891 318587
rect 281933 318469 282051 318587
rect 281773 318309 281891 318427
rect 281933 318309 282051 318427
rect 281773 300469 281891 300587
rect 281933 300469 282051 300587
rect 281773 300309 281891 300427
rect 281933 300309 282051 300427
rect 281773 282469 281891 282587
rect 281933 282469 282051 282587
rect 281773 282309 281891 282427
rect 281933 282309 282051 282427
rect 281773 264469 281891 264587
rect 281933 264469 282051 264587
rect 281773 264309 281891 264427
rect 281933 264309 282051 264427
rect 281773 246469 281891 246587
rect 281933 246469 282051 246587
rect 281773 246309 281891 246427
rect 281933 246309 282051 246427
rect 281773 228469 281891 228587
rect 281933 228469 282051 228587
rect 281773 228309 281891 228427
rect 281933 228309 282051 228427
rect 281773 210469 281891 210587
rect 281933 210469 282051 210587
rect 281773 210309 281891 210427
rect 281933 210309 282051 210427
rect 281773 192469 281891 192587
rect 281933 192469 282051 192587
rect 281773 192309 281891 192427
rect 281933 192309 282051 192427
rect 281773 174469 281891 174587
rect 281933 174469 282051 174587
rect 281773 174309 281891 174427
rect 281933 174309 282051 174427
rect 281773 156469 281891 156587
rect 281933 156469 282051 156587
rect 281773 156309 281891 156427
rect 281933 156309 282051 156427
rect 281773 138469 281891 138587
rect 281933 138469 282051 138587
rect 281773 138309 281891 138427
rect 281933 138309 282051 138427
rect 281773 120469 281891 120587
rect 281933 120469 282051 120587
rect 281773 120309 281891 120427
rect 281933 120309 282051 120427
rect 281773 102469 281891 102587
rect 281933 102469 282051 102587
rect 281773 102309 281891 102427
rect 281933 102309 282051 102427
rect 281773 84469 281891 84587
rect 281933 84469 282051 84587
rect 281773 84309 281891 84427
rect 281933 84309 282051 84427
rect 281773 66469 281891 66587
rect 281933 66469 282051 66587
rect 281773 66309 281891 66427
rect 281933 66309 282051 66427
rect 281773 48469 281891 48587
rect 281933 48469 282051 48587
rect 281773 48309 281891 48427
rect 281933 48309 282051 48427
rect 281773 30469 281891 30587
rect 281933 30469 282051 30587
rect 281773 30309 281891 30427
rect 281933 30309 282051 30427
rect 281773 12469 281891 12587
rect 281933 12469 282051 12587
rect 281773 12309 281891 12427
rect 281933 12309 282051 12427
rect 281773 -1731 281891 -1613
rect 281933 -1731 282051 -1613
rect 281773 -1891 281891 -1773
rect 281933 -1891 282051 -1773
rect 283633 338329 283751 338447
rect 283793 338329 283911 338447
rect 283633 338169 283751 338287
rect 283793 338169 283911 338287
rect 283633 320329 283751 320447
rect 283793 320329 283911 320447
rect 283633 320169 283751 320287
rect 283793 320169 283911 320287
rect 283633 302329 283751 302447
rect 283793 302329 283911 302447
rect 283633 302169 283751 302287
rect 283793 302169 283911 302287
rect 283633 284329 283751 284447
rect 283793 284329 283911 284447
rect 283633 284169 283751 284287
rect 283793 284169 283911 284287
rect 283633 266329 283751 266447
rect 283793 266329 283911 266447
rect 283633 266169 283751 266287
rect 283793 266169 283911 266287
rect 283633 248329 283751 248447
rect 283793 248329 283911 248447
rect 283633 248169 283751 248287
rect 283793 248169 283911 248287
rect 283633 230329 283751 230447
rect 283793 230329 283911 230447
rect 283633 230169 283751 230287
rect 283793 230169 283911 230287
rect 283633 212329 283751 212447
rect 283793 212329 283911 212447
rect 283633 212169 283751 212287
rect 283793 212169 283911 212287
rect 283633 194329 283751 194447
rect 283793 194329 283911 194447
rect 283633 194169 283751 194287
rect 283793 194169 283911 194287
rect 283633 176329 283751 176447
rect 283793 176329 283911 176447
rect 283633 176169 283751 176287
rect 283793 176169 283911 176287
rect 283633 158329 283751 158447
rect 283793 158329 283911 158447
rect 283633 158169 283751 158287
rect 283793 158169 283911 158287
rect 283633 140329 283751 140447
rect 283793 140329 283911 140447
rect 283633 140169 283751 140287
rect 283793 140169 283911 140287
rect 283633 122329 283751 122447
rect 283793 122329 283911 122447
rect 283633 122169 283751 122287
rect 283793 122169 283911 122287
rect 283633 104329 283751 104447
rect 283793 104329 283911 104447
rect 283633 104169 283751 104287
rect 283793 104169 283911 104287
rect 283633 86329 283751 86447
rect 283793 86329 283911 86447
rect 283633 86169 283751 86287
rect 283793 86169 283911 86287
rect 283633 68329 283751 68447
rect 283793 68329 283911 68447
rect 283633 68169 283751 68287
rect 283793 68169 283911 68287
rect 283633 50329 283751 50447
rect 283793 50329 283911 50447
rect 283633 50169 283751 50287
rect 283793 50169 283911 50287
rect 283633 32329 283751 32447
rect 283793 32329 283911 32447
rect 283633 32169 283751 32287
rect 283793 32169 283911 32287
rect 283633 14329 283751 14447
rect 283793 14329 283911 14447
rect 283633 14169 283751 14287
rect 283793 14169 283911 14287
rect 283633 -2691 283751 -2573
rect 283793 -2691 283911 -2573
rect 283633 -2851 283751 -2733
rect 283793 -2851 283911 -2733
rect 296031 355661 296149 355779
rect 296191 355661 296309 355779
rect 296031 355501 296149 355619
rect 296191 355501 296309 355619
rect 295551 355181 295669 355299
rect 295711 355181 295829 355299
rect 295551 355021 295669 355139
rect 295711 355021 295829 355139
rect 295071 354701 295189 354819
rect 295231 354701 295349 354819
rect 295071 354541 295189 354659
rect 295231 354541 295349 354659
rect 294591 354221 294709 354339
rect 294751 354221 294869 354339
rect 294591 354061 294709 354179
rect 294751 354061 294869 354179
rect 294111 353741 294229 353859
rect 294271 353741 294389 353859
rect 294111 353581 294229 353699
rect 294271 353581 294389 353699
rect 290773 353261 290891 353379
rect 290933 353261 291051 353379
rect 290773 353101 290891 353219
rect 290933 353101 291051 353219
rect 285493 340189 285611 340307
rect 285653 340189 285771 340307
rect 285493 340029 285611 340147
rect 285653 340029 285771 340147
rect 285493 322189 285611 322307
rect 285653 322189 285771 322307
rect 285493 322029 285611 322147
rect 285653 322029 285771 322147
rect 285493 304189 285611 304307
rect 285653 304189 285771 304307
rect 285493 304029 285611 304147
rect 285653 304029 285771 304147
rect 285493 286189 285611 286307
rect 285653 286189 285771 286307
rect 285493 286029 285611 286147
rect 285653 286029 285771 286147
rect 285493 268189 285611 268307
rect 285653 268189 285771 268307
rect 285493 268029 285611 268147
rect 285653 268029 285771 268147
rect 285493 250189 285611 250307
rect 285653 250189 285771 250307
rect 285493 250029 285611 250147
rect 285653 250029 285771 250147
rect 285493 232189 285611 232307
rect 285653 232189 285771 232307
rect 285493 232029 285611 232147
rect 285653 232029 285771 232147
rect 285493 214189 285611 214307
rect 285653 214189 285771 214307
rect 285493 214029 285611 214147
rect 285653 214029 285771 214147
rect 285493 196189 285611 196307
rect 285653 196189 285771 196307
rect 285493 196029 285611 196147
rect 285653 196029 285771 196147
rect 285493 178189 285611 178307
rect 285653 178189 285771 178307
rect 285493 178029 285611 178147
rect 285653 178029 285771 178147
rect 285493 160189 285611 160307
rect 285653 160189 285771 160307
rect 285493 160029 285611 160147
rect 285653 160029 285771 160147
rect 285493 142189 285611 142307
rect 285653 142189 285771 142307
rect 285493 142029 285611 142147
rect 285653 142029 285771 142147
rect 285493 124189 285611 124307
rect 285653 124189 285771 124307
rect 285493 124029 285611 124147
rect 285653 124029 285771 124147
rect 285493 106189 285611 106307
rect 285653 106189 285771 106307
rect 285493 106029 285611 106147
rect 285653 106029 285771 106147
rect 285493 88189 285611 88307
rect 285653 88189 285771 88307
rect 285493 88029 285611 88147
rect 285653 88029 285771 88147
rect 285493 70189 285611 70307
rect 285653 70189 285771 70307
rect 285493 70029 285611 70147
rect 285653 70029 285771 70147
rect 285493 52189 285611 52307
rect 285653 52189 285771 52307
rect 285493 52029 285611 52147
rect 285653 52029 285771 52147
rect 285493 34189 285611 34307
rect 285653 34189 285771 34307
rect 285493 34029 285611 34147
rect 285653 34029 285771 34147
rect 285493 16189 285611 16307
rect 285653 16189 285771 16307
rect 285493 16029 285611 16147
rect 285653 16029 285771 16147
rect 276493 -3171 276611 -3053
rect 276653 -3171 276771 -3053
rect 276493 -3331 276611 -3213
rect 276653 -3331 276771 -3213
rect 288913 352301 289031 352419
rect 289073 352301 289191 352419
rect 288913 352141 289031 352259
rect 289073 352141 289191 352259
rect 288913 343609 289031 343727
rect 289073 343609 289191 343727
rect 288913 343449 289031 343567
rect 289073 343449 289191 343567
rect 288913 325609 289031 325727
rect 289073 325609 289191 325727
rect 288913 325449 289031 325567
rect 289073 325449 289191 325567
rect 288913 307609 289031 307727
rect 289073 307609 289191 307727
rect 288913 307449 289031 307567
rect 289073 307449 289191 307567
rect 288913 289609 289031 289727
rect 289073 289609 289191 289727
rect 288913 289449 289031 289567
rect 289073 289449 289191 289567
rect 288913 271609 289031 271727
rect 289073 271609 289191 271727
rect 288913 271449 289031 271567
rect 289073 271449 289191 271567
rect 288913 253609 289031 253727
rect 289073 253609 289191 253727
rect 288913 253449 289031 253567
rect 289073 253449 289191 253567
rect 288913 235609 289031 235727
rect 289073 235609 289191 235727
rect 288913 235449 289031 235567
rect 289073 235449 289191 235567
rect 288913 217609 289031 217727
rect 289073 217609 289191 217727
rect 288913 217449 289031 217567
rect 289073 217449 289191 217567
rect 288913 199609 289031 199727
rect 289073 199609 289191 199727
rect 288913 199449 289031 199567
rect 289073 199449 289191 199567
rect 288913 181609 289031 181727
rect 289073 181609 289191 181727
rect 288913 181449 289031 181567
rect 289073 181449 289191 181567
rect 288913 163609 289031 163727
rect 289073 163609 289191 163727
rect 288913 163449 289031 163567
rect 289073 163449 289191 163567
rect 288913 145609 289031 145727
rect 289073 145609 289191 145727
rect 288913 145449 289031 145567
rect 289073 145449 289191 145567
rect 288913 127609 289031 127727
rect 289073 127609 289191 127727
rect 288913 127449 289031 127567
rect 289073 127449 289191 127567
rect 288913 109609 289031 109727
rect 289073 109609 289191 109727
rect 288913 109449 289031 109567
rect 289073 109449 289191 109567
rect 288913 91609 289031 91727
rect 289073 91609 289191 91727
rect 288913 91449 289031 91567
rect 289073 91449 289191 91567
rect 288913 73609 289031 73727
rect 289073 73609 289191 73727
rect 288913 73449 289031 73567
rect 289073 73449 289191 73567
rect 288913 55609 289031 55727
rect 289073 55609 289191 55727
rect 288913 55449 289031 55567
rect 289073 55449 289191 55567
rect 288913 37609 289031 37727
rect 289073 37609 289191 37727
rect 288913 37449 289031 37567
rect 289073 37449 289191 37567
rect 288913 19609 289031 19727
rect 289073 19609 289191 19727
rect 288913 19449 289031 19567
rect 289073 19449 289191 19567
rect 288913 1609 289031 1727
rect 289073 1609 289191 1727
rect 288913 1449 289031 1567
rect 289073 1449 289191 1567
rect 288913 -291 289031 -173
rect 289073 -291 289191 -173
rect 288913 -451 289031 -333
rect 289073 -451 289191 -333
rect 293631 353261 293749 353379
rect 293791 353261 293909 353379
rect 293631 353101 293749 353219
rect 293791 353101 293909 353219
rect 293151 352781 293269 352899
rect 293311 352781 293429 352899
rect 293151 352621 293269 352739
rect 293311 352621 293429 352739
rect 290773 345469 290891 345587
rect 290933 345469 291051 345587
rect 290773 345309 290891 345427
rect 290933 345309 291051 345427
rect 290773 327469 290891 327587
rect 290933 327469 291051 327587
rect 290773 327309 290891 327427
rect 290933 327309 291051 327427
rect 290773 309469 290891 309587
rect 290933 309469 291051 309587
rect 290773 309309 290891 309427
rect 290933 309309 291051 309427
rect 290773 291469 290891 291587
rect 290933 291469 291051 291587
rect 290773 291309 290891 291427
rect 290933 291309 291051 291427
rect 290773 273469 290891 273587
rect 290933 273469 291051 273587
rect 290773 273309 290891 273427
rect 290933 273309 291051 273427
rect 290773 255469 290891 255587
rect 290933 255469 291051 255587
rect 290773 255309 290891 255427
rect 290933 255309 291051 255427
rect 290773 237469 290891 237587
rect 290933 237469 291051 237587
rect 290773 237309 290891 237427
rect 290933 237309 291051 237427
rect 290773 219469 290891 219587
rect 290933 219469 291051 219587
rect 290773 219309 290891 219427
rect 290933 219309 291051 219427
rect 290773 201469 290891 201587
rect 290933 201469 291051 201587
rect 290773 201309 290891 201427
rect 290933 201309 291051 201427
rect 290773 183469 290891 183587
rect 290933 183469 291051 183587
rect 290773 183309 290891 183427
rect 290933 183309 291051 183427
rect 290773 165469 290891 165587
rect 290933 165469 291051 165587
rect 290773 165309 290891 165427
rect 290933 165309 291051 165427
rect 290773 147469 290891 147587
rect 290933 147469 291051 147587
rect 290773 147309 290891 147427
rect 290933 147309 291051 147427
rect 290773 129469 290891 129587
rect 290933 129469 291051 129587
rect 290773 129309 290891 129427
rect 290933 129309 291051 129427
rect 290773 111469 290891 111587
rect 290933 111469 291051 111587
rect 290773 111309 290891 111427
rect 290933 111309 291051 111427
rect 290773 93469 290891 93587
rect 290933 93469 291051 93587
rect 290773 93309 290891 93427
rect 290933 93309 291051 93427
rect 290773 75469 290891 75587
rect 290933 75469 291051 75587
rect 290773 75309 290891 75427
rect 290933 75309 291051 75427
rect 290773 57469 290891 57587
rect 290933 57469 291051 57587
rect 290773 57309 290891 57427
rect 290933 57309 291051 57427
rect 290773 39469 290891 39587
rect 290933 39469 291051 39587
rect 290773 39309 290891 39427
rect 290933 39309 291051 39427
rect 290773 21469 290891 21587
rect 290933 21469 291051 21587
rect 290773 21309 290891 21427
rect 290933 21309 291051 21427
rect 290773 3469 290891 3587
rect 290933 3469 291051 3587
rect 290773 3309 290891 3427
rect 290933 3309 291051 3427
rect 292671 352301 292789 352419
rect 292831 352301 292949 352419
rect 292671 352141 292789 352259
rect 292831 352141 292949 352259
rect 292671 343609 292789 343727
rect 292831 343609 292949 343727
rect 292671 343449 292789 343567
rect 292831 343449 292949 343567
rect 292671 325609 292789 325727
rect 292831 325609 292949 325727
rect 292671 325449 292789 325567
rect 292831 325449 292949 325567
rect 292671 307609 292789 307727
rect 292831 307609 292949 307727
rect 292671 307449 292789 307567
rect 292831 307449 292949 307567
rect 292671 289609 292789 289727
rect 292831 289609 292949 289727
rect 292671 289449 292789 289567
rect 292831 289449 292949 289567
rect 292671 271609 292789 271727
rect 292831 271609 292949 271727
rect 292671 271449 292789 271567
rect 292831 271449 292949 271567
rect 292671 253609 292789 253727
rect 292831 253609 292949 253727
rect 292671 253449 292789 253567
rect 292831 253449 292949 253567
rect 292671 235609 292789 235727
rect 292831 235609 292949 235727
rect 292671 235449 292789 235567
rect 292831 235449 292949 235567
rect 292671 217609 292789 217727
rect 292831 217609 292949 217727
rect 292671 217449 292789 217567
rect 292831 217449 292949 217567
rect 292671 199609 292789 199727
rect 292831 199609 292949 199727
rect 292671 199449 292789 199567
rect 292831 199449 292949 199567
rect 292671 181609 292789 181727
rect 292831 181609 292949 181727
rect 292671 181449 292789 181567
rect 292831 181449 292949 181567
rect 292671 163609 292789 163727
rect 292831 163609 292949 163727
rect 292671 163449 292789 163567
rect 292831 163449 292949 163567
rect 292671 145609 292789 145727
rect 292831 145609 292949 145727
rect 292671 145449 292789 145567
rect 292831 145449 292949 145567
rect 292671 127609 292789 127727
rect 292831 127609 292949 127727
rect 292671 127449 292789 127567
rect 292831 127449 292949 127567
rect 292671 109609 292789 109727
rect 292831 109609 292949 109727
rect 292671 109449 292789 109567
rect 292831 109449 292949 109567
rect 292671 91609 292789 91727
rect 292831 91609 292949 91727
rect 292671 91449 292789 91567
rect 292831 91449 292949 91567
rect 292671 73609 292789 73727
rect 292831 73609 292949 73727
rect 292671 73449 292789 73567
rect 292831 73449 292949 73567
rect 292671 55609 292789 55727
rect 292831 55609 292949 55727
rect 292671 55449 292789 55567
rect 292831 55449 292949 55567
rect 292671 37609 292789 37727
rect 292831 37609 292949 37727
rect 292671 37449 292789 37567
rect 292831 37449 292949 37567
rect 292671 19609 292789 19727
rect 292831 19609 292949 19727
rect 292671 19449 292789 19567
rect 292831 19449 292949 19567
rect 292671 1609 292789 1727
rect 292831 1609 292949 1727
rect 292671 1449 292789 1567
rect 292831 1449 292949 1567
rect 292671 -291 292789 -173
rect 292831 -291 292949 -173
rect 292671 -451 292789 -333
rect 292831 -451 292949 -333
rect 293151 334609 293269 334727
rect 293311 334609 293429 334727
rect 293151 334449 293269 334567
rect 293311 334449 293429 334567
rect 293151 316609 293269 316727
rect 293311 316609 293429 316727
rect 293151 316449 293269 316567
rect 293311 316449 293429 316567
rect 293151 298609 293269 298727
rect 293311 298609 293429 298727
rect 293151 298449 293269 298567
rect 293311 298449 293429 298567
rect 293151 280609 293269 280727
rect 293311 280609 293429 280727
rect 293151 280449 293269 280567
rect 293311 280449 293429 280567
rect 293151 262609 293269 262727
rect 293311 262609 293429 262727
rect 293151 262449 293269 262567
rect 293311 262449 293429 262567
rect 293151 244609 293269 244727
rect 293311 244609 293429 244727
rect 293151 244449 293269 244567
rect 293311 244449 293429 244567
rect 293151 226609 293269 226727
rect 293311 226609 293429 226727
rect 293151 226449 293269 226567
rect 293311 226449 293429 226567
rect 293151 208609 293269 208727
rect 293311 208609 293429 208727
rect 293151 208449 293269 208567
rect 293311 208449 293429 208567
rect 293151 190609 293269 190727
rect 293311 190609 293429 190727
rect 293151 190449 293269 190567
rect 293311 190449 293429 190567
rect 293151 172609 293269 172727
rect 293311 172609 293429 172727
rect 293151 172449 293269 172567
rect 293311 172449 293429 172567
rect 293151 154609 293269 154727
rect 293311 154609 293429 154727
rect 293151 154449 293269 154567
rect 293311 154449 293429 154567
rect 293151 136609 293269 136727
rect 293311 136609 293429 136727
rect 293151 136449 293269 136567
rect 293311 136449 293429 136567
rect 293151 118609 293269 118727
rect 293311 118609 293429 118727
rect 293151 118449 293269 118567
rect 293311 118449 293429 118567
rect 293151 100609 293269 100727
rect 293311 100609 293429 100727
rect 293151 100449 293269 100567
rect 293311 100449 293429 100567
rect 293151 82609 293269 82727
rect 293311 82609 293429 82727
rect 293151 82449 293269 82567
rect 293311 82449 293429 82567
rect 293151 64609 293269 64727
rect 293311 64609 293429 64727
rect 293151 64449 293269 64567
rect 293311 64449 293429 64567
rect 293151 46609 293269 46727
rect 293311 46609 293429 46727
rect 293151 46449 293269 46567
rect 293311 46449 293429 46567
rect 293151 28609 293269 28727
rect 293311 28609 293429 28727
rect 293151 28449 293269 28567
rect 293311 28449 293429 28567
rect 293151 10609 293269 10727
rect 293311 10609 293429 10727
rect 293151 10449 293269 10567
rect 293311 10449 293429 10567
rect 293151 -771 293269 -653
rect 293311 -771 293429 -653
rect 293151 -931 293269 -813
rect 293311 -931 293429 -813
rect 293631 345469 293749 345587
rect 293791 345469 293909 345587
rect 293631 345309 293749 345427
rect 293791 345309 293909 345427
rect 293631 327469 293749 327587
rect 293791 327469 293909 327587
rect 293631 327309 293749 327427
rect 293791 327309 293909 327427
rect 293631 309469 293749 309587
rect 293791 309469 293909 309587
rect 293631 309309 293749 309427
rect 293791 309309 293909 309427
rect 293631 291469 293749 291587
rect 293791 291469 293909 291587
rect 293631 291309 293749 291427
rect 293791 291309 293909 291427
rect 293631 273469 293749 273587
rect 293791 273469 293909 273587
rect 293631 273309 293749 273427
rect 293791 273309 293909 273427
rect 293631 255469 293749 255587
rect 293791 255469 293909 255587
rect 293631 255309 293749 255427
rect 293791 255309 293909 255427
rect 293631 237469 293749 237587
rect 293791 237469 293909 237587
rect 293631 237309 293749 237427
rect 293791 237309 293909 237427
rect 293631 219469 293749 219587
rect 293791 219469 293909 219587
rect 293631 219309 293749 219427
rect 293791 219309 293909 219427
rect 293631 201469 293749 201587
rect 293791 201469 293909 201587
rect 293631 201309 293749 201427
rect 293791 201309 293909 201427
rect 293631 183469 293749 183587
rect 293791 183469 293909 183587
rect 293631 183309 293749 183427
rect 293791 183309 293909 183427
rect 293631 165469 293749 165587
rect 293791 165469 293909 165587
rect 293631 165309 293749 165427
rect 293791 165309 293909 165427
rect 293631 147469 293749 147587
rect 293791 147469 293909 147587
rect 293631 147309 293749 147427
rect 293791 147309 293909 147427
rect 293631 129469 293749 129587
rect 293791 129469 293909 129587
rect 293631 129309 293749 129427
rect 293791 129309 293909 129427
rect 293631 111469 293749 111587
rect 293791 111469 293909 111587
rect 293631 111309 293749 111427
rect 293791 111309 293909 111427
rect 293631 93469 293749 93587
rect 293791 93469 293909 93587
rect 293631 93309 293749 93427
rect 293791 93309 293909 93427
rect 293631 75469 293749 75587
rect 293791 75469 293909 75587
rect 293631 75309 293749 75427
rect 293791 75309 293909 75427
rect 293631 57469 293749 57587
rect 293791 57469 293909 57587
rect 293631 57309 293749 57427
rect 293791 57309 293909 57427
rect 293631 39469 293749 39587
rect 293791 39469 293909 39587
rect 293631 39309 293749 39427
rect 293791 39309 293909 39427
rect 293631 21469 293749 21587
rect 293791 21469 293909 21587
rect 293631 21309 293749 21427
rect 293791 21309 293909 21427
rect 293631 3469 293749 3587
rect 293791 3469 293909 3587
rect 293631 3309 293749 3427
rect 293791 3309 293909 3427
rect 290773 -1251 290891 -1133
rect 290933 -1251 291051 -1133
rect 290773 -1411 290891 -1293
rect 290933 -1411 291051 -1293
rect 293631 -1251 293749 -1133
rect 293791 -1251 293909 -1133
rect 293631 -1411 293749 -1293
rect 293791 -1411 293909 -1293
rect 294111 336469 294229 336587
rect 294271 336469 294389 336587
rect 294111 336309 294229 336427
rect 294271 336309 294389 336427
rect 294111 318469 294229 318587
rect 294271 318469 294389 318587
rect 294111 318309 294229 318427
rect 294271 318309 294389 318427
rect 294111 300469 294229 300587
rect 294271 300469 294389 300587
rect 294111 300309 294229 300427
rect 294271 300309 294389 300427
rect 294111 282469 294229 282587
rect 294271 282469 294389 282587
rect 294111 282309 294229 282427
rect 294271 282309 294389 282427
rect 294111 264469 294229 264587
rect 294271 264469 294389 264587
rect 294111 264309 294229 264427
rect 294271 264309 294389 264427
rect 294111 246469 294229 246587
rect 294271 246469 294389 246587
rect 294111 246309 294229 246427
rect 294271 246309 294389 246427
rect 294111 228469 294229 228587
rect 294271 228469 294389 228587
rect 294111 228309 294229 228427
rect 294271 228309 294389 228427
rect 294111 210469 294229 210587
rect 294271 210469 294389 210587
rect 294111 210309 294229 210427
rect 294271 210309 294389 210427
rect 294111 192469 294229 192587
rect 294271 192469 294389 192587
rect 294111 192309 294229 192427
rect 294271 192309 294389 192427
rect 294111 174469 294229 174587
rect 294271 174469 294389 174587
rect 294111 174309 294229 174427
rect 294271 174309 294389 174427
rect 294111 156469 294229 156587
rect 294271 156469 294389 156587
rect 294111 156309 294229 156427
rect 294271 156309 294389 156427
rect 294111 138469 294229 138587
rect 294271 138469 294389 138587
rect 294111 138309 294229 138427
rect 294271 138309 294389 138427
rect 294111 120469 294229 120587
rect 294271 120469 294389 120587
rect 294111 120309 294229 120427
rect 294271 120309 294389 120427
rect 294111 102469 294229 102587
rect 294271 102469 294389 102587
rect 294111 102309 294229 102427
rect 294271 102309 294389 102427
rect 294111 84469 294229 84587
rect 294271 84469 294389 84587
rect 294111 84309 294229 84427
rect 294271 84309 294389 84427
rect 294111 66469 294229 66587
rect 294271 66469 294389 66587
rect 294111 66309 294229 66427
rect 294271 66309 294389 66427
rect 294111 48469 294229 48587
rect 294271 48469 294389 48587
rect 294111 48309 294229 48427
rect 294271 48309 294389 48427
rect 294111 30469 294229 30587
rect 294271 30469 294389 30587
rect 294111 30309 294229 30427
rect 294271 30309 294389 30427
rect 294111 12469 294229 12587
rect 294271 12469 294389 12587
rect 294111 12309 294229 12427
rect 294271 12309 294389 12427
rect 294111 -1731 294229 -1613
rect 294271 -1731 294389 -1613
rect 294111 -1891 294229 -1773
rect 294271 -1891 294389 -1773
rect 294591 347329 294709 347447
rect 294751 347329 294869 347447
rect 294591 347169 294709 347287
rect 294751 347169 294869 347287
rect 294591 329329 294709 329447
rect 294751 329329 294869 329447
rect 294591 329169 294709 329287
rect 294751 329169 294869 329287
rect 294591 311329 294709 311447
rect 294751 311329 294869 311447
rect 294591 311169 294709 311287
rect 294751 311169 294869 311287
rect 294591 293329 294709 293447
rect 294751 293329 294869 293447
rect 294591 293169 294709 293287
rect 294751 293169 294869 293287
rect 294591 275329 294709 275447
rect 294751 275329 294869 275447
rect 294591 275169 294709 275287
rect 294751 275169 294869 275287
rect 294591 257329 294709 257447
rect 294751 257329 294869 257447
rect 294591 257169 294709 257287
rect 294751 257169 294869 257287
rect 294591 239329 294709 239447
rect 294751 239329 294869 239447
rect 294591 239169 294709 239287
rect 294751 239169 294869 239287
rect 294591 221329 294709 221447
rect 294751 221329 294869 221447
rect 294591 221169 294709 221287
rect 294751 221169 294869 221287
rect 294591 203329 294709 203447
rect 294751 203329 294869 203447
rect 294591 203169 294709 203287
rect 294751 203169 294869 203287
rect 294591 185329 294709 185447
rect 294751 185329 294869 185447
rect 294591 185169 294709 185287
rect 294751 185169 294869 185287
rect 294591 167329 294709 167447
rect 294751 167329 294869 167447
rect 294591 167169 294709 167287
rect 294751 167169 294869 167287
rect 294591 149329 294709 149447
rect 294751 149329 294869 149447
rect 294591 149169 294709 149287
rect 294751 149169 294869 149287
rect 294591 131329 294709 131447
rect 294751 131329 294869 131447
rect 294591 131169 294709 131287
rect 294751 131169 294869 131287
rect 294591 113329 294709 113447
rect 294751 113329 294869 113447
rect 294591 113169 294709 113287
rect 294751 113169 294869 113287
rect 294591 95329 294709 95447
rect 294751 95329 294869 95447
rect 294591 95169 294709 95287
rect 294751 95169 294869 95287
rect 294591 77329 294709 77447
rect 294751 77329 294869 77447
rect 294591 77169 294709 77287
rect 294751 77169 294869 77287
rect 294591 59329 294709 59447
rect 294751 59329 294869 59447
rect 294591 59169 294709 59287
rect 294751 59169 294869 59287
rect 294591 41329 294709 41447
rect 294751 41329 294869 41447
rect 294591 41169 294709 41287
rect 294751 41169 294869 41287
rect 294591 23329 294709 23447
rect 294751 23329 294869 23447
rect 294591 23169 294709 23287
rect 294751 23169 294869 23287
rect 294591 5329 294709 5447
rect 294751 5329 294869 5447
rect 294591 5169 294709 5287
rect 294751 5169 294869 5287
rect 294591 -2211 294709 -2093
rect 294751 -2211 294869 -2093
rect 294591 -2371 294709 -2253
rect 294751 -2371 294869 -2253
rect 295071 338329 295189 338447
rect 295231 338329 295349 338447
rect 295071 338169 295189 338287
rect 295231 338169 295349 338287
rect 295071 320329 295189 320447
rect 295231 320329 295349 320447
rect 295071 320169 295189 320287
rect 295231 320169 295349 320287
rect 295071 302329 295189 302447
rect 295231 302329 295349 302447
rect 295071 302169 295189 302287
rect 295231 302169 295349 302287
rect 295071 284329 295189 284447
rect 295231 284329 295349 284447
rect 295071 284169 295189 284287
rect 295231 284169 295349 284287
rect 295071 266329 295189 266447
rect 295231 266329 295349 266447
rect 295071 266169 295189 266287
rect 295231 266169 295349 266287
rect 295071 248329 295189 248447
rect 295231 248329 295349 248447
rect 295071 248169 295189 248287
rect 295231 248169 295349 248287
rect 295071 230329 295189 230447
rect 295231 230329 295349 230447
rect 295071 230169 295189 230287
rect 295231 230169 295349 230287
rect 295071 212329 295189 212447
rect 295231 212329 295349 212447
rect 295071 212169 295189 212287
rect 295231 212169 295349 212287
rect 295071 194329 295189 194447
rect 295231 194329 295349 194447
rect 295071 194169 295189 194287
rect 295231 194169 295349 194287
rect 295071 176329 295189 176447
rect 295231 176329 295349 176447
rect 295071 176169 295189 176287
rect 295231 176169 295349 176287
rect 295071 158329 295189 158447
rect 295231 158329 295349 158447
rect 295071 158169 295189 158287
rect 295231 158169 295349 158287
rect 295071 140329 295189 140447
rect 295231 140329 295349 140447
rect 295071 140169 295189 140287
rect 295231 140169 295349 140287
rect 295071 122329 295189 122447
rect 295231 122329 295349 122447
rect 295071 122169 295189 122287
rect 295231 122169 295349 122287
rect 295071 104329 295189 104447
rect 295231 104329 295349 104447
rect 295071 104169 295189 104287
rect 295231 104169 295349 104287
rect 295071 86329 295189 86447
rect 295231 86329 295349 86447
rect 295071 86169 295189 86287
rect 295231 86169 295349 86287
rect 295071 68329 295189 68447
rect 295231 68329 295349 68447
rect 295071 68169 295189 68287
rect 295231 68169 295349 68287
rect 295071 50329 295189 50447
rect 295231 50329 295349 50447
rect 295071 50169 295189 50287
rect 295231 50169 295349 50287
rect 295071 32329 295189 32447
rect 295231 32329 295349 32447
rect 295071 32169 295189 32287
rect 295231 32169 295349 32287
rect 295071 14329 295189 14447
rect 295231 14329 295349 14447
rect 295071 14169 295189 14287
rect 295231 14169 295349 14287
rect 295071 -2691 295189 -2573
rect 295231 -2691 295349 -2573
rect 295071 -2851 295189 -2733
rect 295231 -2851 295349 -2733
rect 295551 349189 295669 349307
rect 295711 349189 295829 349307
rect 295551 349029 295669 349147
rect 295711 349029 295829 349147
rect 295551 331189 295669 331307
rect 295711 331189 295829 331307
rect 295551 331029 295669 331147
rect 295711 331029 295829 331147
rect 295551 313189 295669 313307
rect 295711 313189 295829 313307
rect 295551 313029 295669 313147
rect 295711 313029 295829 313147
rect 295551 295189 295669 295307
rect 295711 295189 295829 295307
rect 295551 295029 295669 295147
rect 295711 295029 295829 295147
rect 295551 277189 295669 277307
rect 295711 277189 295829 277307
rect 295551 277029 295669 277147
rect 295711 277029 295829 277147
rect 295551 259189 295669 259307
rect 295711 259189 295829 259307
rect 295551 259029 295669 259147
rect 295711 259029 295829 259147
rect 295551 241189 295669 241307
rect 295711 241189 295829 241307
rect 295551 241029 295669 241147
rect 295711 241029 295829 241147
rect 295551 223189 295669 223307
rect 295711 223189 295829 223307
rect 295551 223029 295669 223147
rect 295711 223029 295829 223147
rect 295551 205189 295669 205307
rect 295711 205189 295829 205307
rect 295551 205029 295669 205147
rect 295711 205029 295829 205147
rect 295551 187189 295669 187307
rect 295711 187189 295829 187307
rect 295551 187029 295669 187147
rect 295711 187029 295829 187147
rect 295551 169189 295669 169307
rect 295711 169189 295829 169307
rect 295551 169029 295669 169147
rect 295711 169029 295829 169147
rect 295551 151189 295669 151307
rect 295711 151189 295829 151307
rect 295551 151029 295669 151147
rect 295711 151029 295829 151147
rect 295551 133189 295669 133307
rect 295711 133189 295829 133307
rect 295551 133029 295669 133147
rect 295711 133029 295829 133147
rect 295551 115189 295669 115307
rect 295711 115189 295829 115307
rect 295551 115029 295669 115147
rect 295711 115029 295829 115147
rect 295551 97189 295669 97307
rect 295711 97189 295829 97307
rect 295551 97029 295669 97147
rect 295711 97029 295829 97147
rect 295551 79189 295669 79307
rect 295711 79189 295829 79307
rect 295551 79029 295669 79147
rect 295711 79029 295829 79147
rect 295551 61189 295669 61307
rect 295711 61189 295829 61307
rect 295551 61029 295669 61147
rect 295711 61029 295829 61147
rect 295551 43189 295669 43307
rect 295711 43189 295829 43307
rect 295551 43029 295669 43147
rect 295711 43029 295829 43147
rect 295551 25189 295669 25307
rect 295711 25189 295829 25307
rect 295551 25029 295669 25147
rect 295711 25029 295829 25147
rect 295551 7189 295669 7307
rect 295711 7189 295829 7307
rect 295551 7029 295669 7147
rect 295711 7029 295829 7147
rect 295551 -3171 295669 -3053
rect 295711 -3171 295829 -3053
rect 295551 -3331 295669 -3213
rect 295711 -3331 295829 -3213
rect 296031 340189 296149 340307
rect 296191 340189 296309 340307
rect 296031 340029 296149 340147
rect 296191 340029 296309 340147
rect 296031 322189 296149 322307
rect 296191 322189 296309 322307
rect 296031 322029 296149 322147
rect 296191 322029 296309 322147
rect 296031 304189 296149 304307
rect 296191 304189 296309 304307
rect 296031 304029 296149 304147
rect 296191 304029 296309 304147
rect 296031 286189 296149 286307
rect 296191 286189 296309 286307
rect 296031 286029 296149 286147
rect 296191 286029 296309 286147
rect 296031 268189 296149 268307
rect 296191 268189 296309 268307
rect 296031 268029 296149 268147
rect 296191 268029 296309 268147
rect 296031 250189 296149 250307
rect 296191 250189 296309 250307
rect 296031 250029 296149 250147
rect 296191 250029 296309 250147
rect 296031 232189 296149 232307
rect 296191 232189 296309 232307
rect 296031 232029 296149 232147
rect 296191 232029 296309 232147
rect 296031 214189 296149 214307
rect 296191 214189 296309 214307
rect 296031 214029 296149 214147
rect 296191 214029 296309 214147
rect 296031 196189 296149 196307
rect 296191 196189 296309 196307
rect 296031 196029 296149 196147
rect 296191 196029 296309 196147
rect 296031 178189 296149 178307
rect 296191 178189 296309 178307
rect 296031 178029 296149 178147
rect 296191 178029 296309 178147
rect 296031 160189 296149 160307
rect 296191 160189 296309 160307
rect 296031 160029 296149 160147
rect 296191 160029 296309 160147
rect 296031 142189 296149 142307
rect 296191 142189 296309 142307
rect 296031 142029 296149 142147
rect 296191 142029 296309 142147
rect 296031 124189 296149 124307
rect 296191 124189 296309 124307
rect 296031 124029 296149 124147
rect 296191 124029 296309 124147
rect 296031 106189 296149 106307
rect 296191 106189 296309 106307
rect 296031 106029 296149 106147
rect 296191 106029 296309 106147
rect 296031 88189 296149 88307
rect 296191 88189 296309 88307
rect 296031 88029 296149 88147
rect 296191 88029 296309 88147
rect 296031 70189 296149 70307
rect 296191 70189 296309 70307
rect 296031 70029 296149 70147
rect 296191 70029 296309 70147
rect 296031 52189 296149 52307
rect 296191 52189 296309 52307
rect 296031 52029 296149 52147
rect 296191 52029 296309 52147
rect 296031 34189 296149 34307
rect 296191 34189 296309 34307
rect 296031 34029 296149 34147
rect 296191 34029 296309 34147
rect 296031 16189 296149 16307
rect 296191 16189 296309 16307
rect 296031 16029 296149 16147
rect 296191 16029 296309 16147
rect 285493 -3651 285611 -3533
rect 285653 -3651 285771 -3533
rect 285493 -3811 285611 -3693
rect 285653 -3811 285771 -3693
rect 296031 -3651 296149 -3533
rect 296191 -3651 296309 -3533
rect 296031 -3811 296149 -3693
rect 296191 -3811 296309 -3693
<< metal5 >>
rect -4363 355779 296325 355795
rect -4363 355661 -4347 355779
rect -4229 355661 -4187 355779
rect -4069 355661 15493 355779
rect 15611 355661 15653 355779
rect 15771 355661 33493 355779
rect 33611 355661 33653 355779
rect 33771 355661 51493 355779
rect 51611 355661 51653 355779
rect 51771 355661 69493 355779
rect 69611 355661 69653 355779
rect 69771 355661 87493 355779
rect 87611 355661 87653 355779
rect 87771 355661 105493 355779
rect 105611 355661 105653 355779
rect 105771 355661 123493 355779
rect 123611 355661 123653 355779
rect 123771 355661 141493 355779
rect 141611 355661 141653 355779
rect 141771 355661 159493 355779
rect 159611 355661 159653 355779
rect 159771 355661 177493 355779
rect 177611 355661 177653 355779
rect 177771 355661 195493 355779
rect 195611 355661 195653 355779
rect 195771 355661 213493 355779
rect 213611 355661 213653 355779
rect 213771 355661 231493 355779
rect 231611 355661 231653 355779
rect 231771 355661 249493 355779
rect 249611 355661 249653 355779
rect 249771 355661 267493 355779
rect 267611 355661 267653 355779
rect 267771 355661 285493 355779
rect 285611 355661 285653 355779
rect 285771 355661 296031 355779
rect 296149 355661 296191 355779
rect 296309 355661 296325 355779
rect -4363 355619 296325 355661
rect -4363 355501 -4347 355619
rect -4229 355501 -4187 355619
rect -4069 355501 15493 355619
rect 15611 355501 15653 355619
rect 15771 355501 33493 355619
rect 33611 355501 33653 355619
rect 33771 355501 51493 355619
rect 51611 355501 51653 355619
rect 51771 355501 69493 355619
rect 69611 355501 69653 355619
rect 69771 355501 87493 355619
rect 87611 355501 87653 355619
rect 87771 355501 105493 355619
rect 105611 355501 105653 355619
rect 105771 355501 123493 355619
rect 123611 355501 123653 355619
rect 123771 355501 141493 355619
rect 141611 355501 141653 355619
rect 141771 355501 159493 355619
rect 159611 355501 159653 355619
rect 159771 355501 177493 355619
rect 177611 355501 177653 355619
rect 177771 355501 195493 355619
rect 195611 355501 195653 355619
rect 195771 355501 213493 355619
rect 213611 355501 213653 355619
rect 213771 355501 231493 355619
rect 231611 355501 231653 355619
rect 231771 355501 249493 355619
rect 249611 355501 249653 355619
rect 249771 355501 267493 355619
rect 267611 355501 267653 355619
rect 267771 355501 285493 355619
rect 285611 355501 285653 355619
rect 285771 355501 296031 355619
rect 296149 355501 296191 355619
rect 296309 355501 296325 355619
rect -4363 355485 296325 355501
rect -3883 355299 295845 355315
rect -3883 355181 -3867 355299
rect -3749 355181 -3707 355299
rect -3589 355181 6493 355299
rect 6611 355181 6653 355299
rect 6771 355181 24493 355299
rect 24611 355181 24653 355299
rect 24771 355181 42493 355299
rect 42611 355181 42653 355299
rect 42771 355181 60493 355299
rect 60611 355181 60653 355299
rect 60771 355181 78493 355299
rect 78611 355181 78653 355299
rect 78771 355181 96493 355299
rect 96611 355181 96653 355299
rect 96771 355181 114493 355299
rect 114611 355181 114653 355299
rect 114771 355181 132493 355299
rect 132611 355181 132653 355299
rect 132771 355181 150493 355299
rect 150611 355181 150653 355299
rect 150771 355181 168493 355299
rect 168611 355181 168653 355299
rect 168771 355181 186493 355299
rect 186611 355181 186653 355299
rect 186771 355181 204493 355299
rect 204611 355181 204653 355299
rect 204771 355181 222493 355299
rect 222611 355181 222653 355299
rect 222771 355181 240493 355299
rect 240611 355181 240653 355299
rect 240771 355181 258493 355299
rect 258611 355181 258653 355299
rect 258771 355181 276493 355299
rect 276611 355181 276653 355299
rect 276771 355181 295551 355299
rect 295669 355181 295711 355299
rect 295829 355181 295845 355299
rect -3883 355139 295845 355181
rect -3883 355021 -3867 355139
rect -3749 355021 -3707 355139
rect -3589 355021 6493 355139
rect 6611 355021 6653 355139
rect 6771 355021 24493 355139
rect 24611 355021 24653 355139
rect 24771 355021 42493 355139
rect 42611 355021 42653 355139
rect 42771 355021 60493 355139
rect 60611 355021 60653 355139
rect 60771 355021 78493 355139
rect 78611 355021 78653 355139
rect 78771 355021 96493 355139
rect 96611 355021 96653 355139
rect 96771 355021 114493 355139
rect 114611 355021 114653 355139
rect 114771 355021 132493 355139
rect 132611 355021 132653 355139
rect 132771 355021 150493 355139
rect 150611 355021 150653 355139
rect 150771 355021 168493 355139
rect 168611 355021 168653 355139
rect 168771 355021 186493 355139
rect 186611 355021 186653 355139
rect 186771 355021 204493 355139
rect 204611 355021 204653 355139
rect 204771 355021 222493 355139
rect 222611 355021 222653 355139
rect 222771 355021 240493 355139
rect 240611 355021 240653 355139
rect 240771 355021 258493 355139
rect 258611 355021 258653 355139
rect 258771 355021 276493 355139
rect 276611 355021 276653 355139
rect 276771 355021 295551 355139
rect 295669 355021 295711 355139
rect 295829 355021 295845 355139
rect -3883 355005 295845 355021
rect -3403 354819 295365 354835
rect -3403 354701 -3387 354819
rect -3269 354701 -3227 354819
rect -3109 354701 13633 354819
rect 13751 354701 13793 354819
rect 13911 354701 31633 354819
rect 31751 354701 31793 354819
rect 31911 354701 49633 354819
rect 49751 354701 49793 354819
rect 49911 354701 67633 354819
rect 67751 354701 67793 354819
rect 67911 354701 85633 354819
rect 85751 354701 85793 354819
rect 85911 354701 103633 354819
rect 103751 354701 103793 354819
rect 103911 354701 121633 354819
rect 121751 354701 121793 354819
rect 121911 354701 139633 354819
rect 139751 354701 139793 354819
rect 139911 354701 157633 354819
rect 157751 354701 157793 354819
rect 157911 354701 175633 354819
rect 175751 354701 175793 354819
rect 175911 354701 193633 354819
rect 193751 354701 193793 354819
rect 193911 354701 211633 354819
rect 211751 354701 211793 354819
rect 211911 354701 229633 354819
rect 229751 354701 229793 354819
rect 229911 354701 247633 354819
rect 247751 354701 247793 354819
rect 247911 354701 265633 354819
rect 265751 354701 265793 354819
rect 265911 354701 283633 354819
rect 283751 354701 283793 354819
rect 283911 354701 295071 354819
rect 295189 354701 295231 354819
rect 295349 354701 295365 354819
rect -3403 354659 295365 354701
rect -3403 354541 -3387 354659
rect -3269 354541 -3227 354659
rect -3109 354541 13633 354659
rect 13751 354541 13793 354659
rect 13911 354541 31633 354659
rect 31751 354541 31793 354659
rect 31911 354541 49633 354659
rect 49751 354541 49793 354659
rect 49911 354541 67633 354659
rect 67751 354541 67793 354659
rect 67911 354541 85633 354659
rect 85751 354541 85793 354659
rect 85911 354541 103633 354659
rect 103751 354541 103793 354659
rect 103911 354541 121633 354659
rect 121751 354541 121793 354659
rect 121911 354541 139633 354659
rect 139751 354541 139793 354659
rect 139911 354541 157633 354659
rect 157751 354541 157793 354659
rect 157911 354541 175633 354659
rect 175751 354541 175793 354659
rect 175911 354541 193633 354659
rect 193751 354541 193793 354659
rect 193911 354541 211633 354659
rect 211751 354541 211793 354659
rect 211911 354541 229633 354659
rect 229751 354541 229793 354659
rect 229911 354541 247633 354659
rect 247751 354541 247793 354659
rect 247911 354541 265633 354659
rect 265751 354541 265793 354659
rect 265911 354541 283633 354659
rect 283751 354541 283793 354659
rect 283911 354541 295071 354659
rect 295189 354541 295231 354659
rect 295349 354541 295365 354659
rect -3403 354525 295365 354541
rect -2923 354339 294885 354355
rect -2923 354221 -2907 354339
rect -2789 354221 -2747 354339
rect -2629 354221 4633 354339
rect 4751 354221 4793 354339
rect 4911 354221 22633 354339
rect 22751 354221 22793 354339
rect 22911 354221 40633 354339
rect 40751 354221 40793 354339
rect 40911 354221 58633 354339
rect 58751 354221 58793 354339
rect 58911 354221 76633 354339
rect 76751 354221 76793 354339
rect 76911 354221 94633 354339
rect 94751 354221 94793 354339
rect 94911 354221 112633 354339
rect 112751 354221 112793 354339
rect 112911 354221 130633 354339
rect 130751 354221 130793 354339
rect 130911 354221 148633 354339
rect 148751 354221 148793 354339
rect 148911 354221 166633 354339
rect 166751 354221 166793 354339
rect 166911 354221 184633 354339
rect 184751 354221 184793 354339
rect 184911 354221 202633 354339
rect 202751 354221 202793 354339
rect 202911 354221 220633 354339
rect 220751 354221 220793 354339
rect 220911 354221 238633 354339
rect 238751 354221 238793 354339
rect 238911 354221 256633 354339
rect 256751 354221 256793 354339
rect 256911 354221 274633 354339
rect 274751 354221 274793 354339
rect 274911 354221 294591 354339
rect 294709 354221 294751 354339
rect 294869 354221 294885 354339
rect -2923 354179 294885 354221
rect -2923 354061 -2907 354179
rect -2789 354061 -2747 354179
rect -2629 354061 4633 354179
rect 4751 354061 4793 354179
rect 4911 354061 22633 354179
rect 22751 354061 22793 354179
rect 22911 354061 40633 354179
rect 40751 354061 40793 354179
rect 40911 354061 58633 354179
rect 58751 354061 58793 354179
rect 58911 354061 76633 354179
rect 76751 354061 76793 354179
rect 76911 354061 94633 354179
rect 94751 354061 94793 354179
rect 94911 354061 112633 354179
rect 112751 354061 112793 354179
rect 112911 354061 130633 354179
rect 130751 354061 130793 354179
rect 130911 354061 148633 354179
rect 148751 354061 148793 354179
rect 148911 354061 166633 354179
rect 166751 354061 166793 354179
rect 166911 354061 184633 354179
rect 184751 354061 184793 354179
rect 184911 354061 202633 354179
rect 202751 354061 202793 354179
rect 202911 354061 220633 354179
rect 220751 354061 220793 354179
rect 220911 354061 238633 354179
rect 238751 354061 238793 354179
rect 238911 354061 256633 354179
rect 256751 354061 256793 354179
rect 256911 354061 274633 354179
rect 274751 354061 274793 354179
rect 274911 354061 294591 354179
rect 294709 354061 294751 354179
rect 294869 354061 294885 354179
rect -2923 354045 294885 354061
rect -2443 353859 294405 353875
rect -2443 353741 -2427 353859
rect -2309 353741 -2267 353859
rect -2149 353741 11773 353859
rect 11891 353741 11933 353859
rect 12051 353741 29773 353859
rect 29891 353741 29933 353859
rect 30051 353741 47773 353859
rect 47891 353741 47933 353859
rect 48051 353741 65773 353859
rect 65891 353741 65933 353859
rect 66051 353741 83773 353859
rect 83891 353741 83933 353859
rect 84051 353741 101773 353859
rect 101891 353741 101933 353859
rect 102051 353741 119773 353859
rect 119891 353741 119933 353859
rect 120051 353741 137773 353859
rect 137891 353741 137933 353859
rect 138051 353741 155773 353859
rect 155891 353741 155933 353859
rect 156051 353741 173773 353859
rect 173891 353741 173933 353859
rect 174051 353741 191773 353859
rect 191891 353741 191933 353859
rect 192051 353741 209773 353859
rect 209891 353741 209933 353859
rect 210051 353741 227773 353859
rect 227891 353741 227933 353859
rect 228051 353741 245773 353859
rect 245891 353741 245933 353859
rect 246051 353741 263773 353859
rect 263891 353741 263933 353859
rect 264051 353741 281773 353859
rect 281891 353741 281933 353859
rect 282051 353741 294111 353859
rect 294229 353741 294271 353859
rect 294389 353741 294405 353859
rect -2443 353699 294405 353741
rect -2443 353581 -2427 353699
rect -2309 353581 -2267 353699
rect -2149 353581 11773 353699
rect 11891 353581 11933 353699
rect 12051 353581 29773 353699
rect 29891 353581 29933 353699
rect 30051 353581 47773 353699
rect 47891 353581 47933 353699
rect 48051 353581 65773 353699
rect 65891 353581 65933 353699
rect 66051 353581 83773 353699
rect 83891 353581 83933 353699
rect 84051 353581 101773 353699
rect 101891 353581 101933 353699
rect 102051 353581 119773 353699
rect 119891 353581 119933 353699
rect 120051 353581 137773 353699
rect 137891 353581 137933 353699
rect 138051 353581 155773 353699
rect 155891 353581 155933 353699
rect 156051 353581 173773 353699
rect 173891 353581 173933 353699
rect 174051 353581 191773 353699
rect 191891 353581 191933 353699
rect 192051 353581 209773 353699
rect 209891 353581 209933 353699
rect 210051 353581 227773 353699
rect 227891 353581 227933 353699
rect 228051 353581 245773 353699
rect 245891 353581 245933 353699
rect 246051 353581 263773 353699
rect 263891 353581 263933 353699
rect 264051 353581 281773 353699
rect 281891 353581 281933 353699
rect 282051 353581 294111 353699
rect 294229 353581 294271 353699
rect 294389 353581 294405 353699
rect -2443 353565 294405 353581
rect -1963 353379 293925 353395
rect -1963 353261 -1947 353379
rect -1829 353261 -1787 353379
rect -1669 353261 2773 353379
rect 2891 353261 2933 353379
rect 3051 353261 20773 353379
rect 20891 353261 20933 353379
rect 21051 353261 38773 353379
rect 38891 353261 38933 353379
rect 39051 353261 56773 353379
rect 56891 353261 56933 353379
rect 57051 353261 74773 353379
rect 74891 353261 74933 353379
rect 75051 353261 92773 353379
rect 92891 353261 92933 353379
rect 93051 353261 110773 353379
rect 110891 353261 110933 353379
rect 111051 353261 128773 353379
rect 128891 353261 128933 353379
rect 129051 353261 146773 353379
rect 146891 353261 146933 353379
rect 147051 353261 164773 353379
rect 164891 353261 164933 353379
rect 165051 353261 182773 353379
rect 182891 353261 182933 353379
rect 183051 353261 200773 353379
rect 200891 353261 200933 353379
rect 201051 353261 218773 353379
rect 218891 353261 218933 353379
rect 219051 353261 236773 353379
rect 236891 353261 236933 353379
rect 237051 353261 254773 353379
rect 254891 353261 254933 353379
rect 255051 353261 272773 353379
rect 272891 353261 272933 353379
rect 273051 353261 290773 353379
rect 290891 353261 290933 353379
rect 291051 353261 293631 353379
rect 293749 353261 293791 353379
rect 293909 353261 293925 353379
rect -1963 353219 293925 353261
rect -1963 353101 -1947 353219
rect -1829 353101 -1787 353219
rect -1669 353101 2773 353219
rect 2891 353101 2933 353219
rect 3051 353101 20773 353219
rect 20891 353101 20933 353219
rect 21051 353101 38773 353219
rect 38891 353101 38933 353219
rect 39051 353101 56773 353219
rect 56891 353101 56933 353219
rect 57051 353101 74773 353219
rect 74891 353101 74933 353219
rect 75051 353101 92773 353219
rect 92891 353101 92933 353219
rect 93051 353101 110773 353219
rect 110891 353101 110933 353219
rect 111051 353101 128773 353219
rect 128891 353101 128933 353219
rect 129051 353101 146773 353219
rect 146891 353101 146933 353219
rect 147051 353101 164773 353219
rect 164891 353101 164933 353219
rect 165051 353101 182773 353219
rect 182891 353101 182933 353219
rect 183051 353101 200773 353219
rect 200891 353101 200933 353219
rect 201051 353101 218773 353219
rect 218891 353101 218933 353219
rect 219051 353101 236773 353219
rect 236891 353101 236933 353219
rect 237051 353101 254773 353219
rect 254891 353101 254933 353219
rect 255051 353101 272773 353219
rect 272891 353101 272933 353219
rect 273051 353101 290773 353219
rect 290891 353101 290933 353219
rect 291051 353101 293631 353219
rect 293749 353101 293791 353219
rect 293909 353101 293925 353219
rect -1963 353085 293925 353101
rect -1483 352899 293445 352915
rect -1483 352781 -1467 352899
rect -1349 352781 -1307 352899
rect -1189 352781 9913 352899
rect 10031 352781 10073 352899
rect 10191 352781 27913 352899
rect 28031 352781 28073 352899
rect 28191 352781 45913 352899
rect 46031 352781 46073 352899
rect 46191 352781 63913 352899
rect 64031 352781 64073 352899
rect 64191 352781 81913 352899
rect 82031 352781 82073 352899
rect 82191 352781 99913 352899
rect 100031 352781 100073 352899
rect 100191 352781 117913 352899
rect 118031 352781 118073 352899
rect 118191 352781 135913 352899
rect 136031 352781 136073 352899
rect 136191 352781 153913 352899
rect 154031 352781 154073 352899
rect 154191 352781 171913 352899
rect 172031 352781 172073 352899
rect 172191 352781 189913 352899
rect 190031 352781 190073 352899
rect 190191 352781 207913 352899
rect 208031 352781 208073 352899
rect 208191 352781 225913 352899
rect 226031 352781 226073 352899
rect 226191 352781 243913 352899
rect 244031 352781 244073 352899
rect 244191 352781 261913 352899
rect 262031 352781 262073 352899
rect 262191 352781 279913 352899
rect 280031 352781 280073 352899
rect 280191 352781 293151 352899
rect 293269 352781 293311 352899
rect 293429 352781 293445 352899
rect -1483 352739 293445 352781
rect -1483 352621 -1467 352739
rect -1349 352621 -1307 352739
rect -1189 352621 9913 352739
rect 10031 352621 10073 352739
rect 10191 352621 27913 352739
rect 28031 352621 28073 352739
rect 28191 352621 45913 352739
rect 46031 352621 46073 352739
rect 46191 352621 63913 352739
rect 64031 352621 64073 352739
rect 64191 352621 81913 352739
rect 82031 352621 82073 352739
rect 82191 352621 99913 352739
rect 100031 352621 100073 352739
rect 100191 352621 117913 352739
rect 118031 352621 118073 352739
rect 118191 352621 135913 352739
rect 136031 352621 136073 352739
rect 136191 352621 153913 352739
rect 154031 352621 154073 352739
rect 154191 352621 171913 352739
rect 172031 352621 172073 352739
rect 172191 352621 189913 352739
rect 190031 352621 190073 352739
rect 190191 352621 207913 352739
rect 208031 352621 208073 352739
rect 208191 352621 225913 352739
rect 226031 352621 226073 352739
rect 226191 352621 243913 352739
rect 244031 352621 244073 352739
rect 244191 352621 261913 352739
rect 262031 352621 262073 352739
rect 262191 352621 279913 352739
rect 280031 352621 280073 352739
rect 280191 352621 293151 352739
rect 293269 352621 293311 352739
rect 293429 352621 293445 352739
rect -1483 352605 293445 352621
rect -1003 352419 292965 352435
rect -1003 352301 -987 352419
rect -869 352301 -827 352419
rect -709 352301 913 352419
rect 1031 352301 1073 352419
rect 1191 352301 18913 352419
rect 19031 352301 19073 352419
rect 19191 352301 36913 352419
rect 37031 352301 37073 352419
rect 37191 352301 54913 352419
rect 55031 352301 55073 352419
rect 55191 352301 72913 352419
rect 73031 352301 73073 352419
rect 73191 352301 90913 352419
rect 91031 352301 91073 352419
rect 91191 352301 108913 352419
rect 109031 352301 109073 352419
rect 109191 352301 126913 352419
rect 127031 352301 127073 352419
rect 127191 352301 144913 352419
rect 145031 352301 145073 352419
rect 145191 352301 162913 352419
rect 163031 352301 163073 352419
rect 163191 352301 180913 352419
rect 181031 352301 181073 352419
rect 181191 352301 198913 352419
rect 199031 352301 199073 352419
rect 199191 352301 216913 352419
rect 217031 352301 217073 352419
rect 217191 352301 234913 352419
rect 235031 352301 235073 352419
rect 235191 352301 252913 352419
rect 253031 352301 253073 352419
rect 253191 352301 270913 352419
rect 271031 352301 271073 352419
rect 271191 352301 288913 352419
rect 289031 352301 289073 352419
rect 289191 352301 292671 352419
rect 292789 352301 292831 352419
rect 292949 352301 292965 352419
rect -1003 352259 292965 352301
rect -1003 352141 -987 352259
rect -869 352141 -827 352259
rect -709 352141 913 352259
rect 1031 352141 1073 352259
rect 1191 352141 18913 352259
rect 19031 352141 19073 352259
rect 19191 352141 36913 352259
rect 37031 352141 37073 352259
rect 37191 352141 54913 352259
rect 55031 352141 55073 352259
rect 55191 352141 72913 352259
rect 73031 352141 73073 352259
rect 73191 352141 90913 352259
rect 91031 352141 91073 352259
rect 91191 352141 108913 352259
rect 109031 352141 109073 352259
rect 109191 352141 126913 352259
rect 127031 352141 127073 352259
rect 127191 352141 144913 352259
rect 145031 352141 145073 352259
rect 145191 352141 162913 352259
rect 163031 352141 163073 352259
rect 163191 352141 180913 352259
rect 181031 352141 181073 352259
rect 181191 352141 198913 352259
rect 199031 352141 199073 352259
rect 199191 352141 216913 352259
rect 217031 352141 217073 352259
rect 217191 352141 234913 352259
rect 235031 352141 235073 352259
rect 235191 352141 252913 352259
rect 253031 352141 253073 352259
rect 253191 352141 270913 352259
rect 271031 352141 271073 352259
rect 271191 352141 288913 352259
rect 289031 352141 289073 352259
rect 289191 352141 292671 352259
rect 292789 352141 292831 352259
rect 292949 352141 292965 352259
rect -1003 352125 292965 352141
rect -4363 349307 296325 349323
rect -4363 349189 -3867 349307
rect -3749 349189 -3707 349307
rect -3589 349189 6493 349307
rect 6611 349189 6653 349307
rect 6771 349189 24493 349307
rect 24611 349189 24653 349307
rect 24771 349189 42493 349307
rect 42611 349189 42653 349307
rect 42771 349189 60493 349307
rect 60611 349189 60653 349307
rect 60771 349189 78493 349307
rect 78611 349189 78653 349307
rect 78771 349189 96493 349307
rect 96611 349189 96653 349307
rect 96771 349189 114493 349307
rect 114611 349189 114653 349307
rect 114771 349189 132493 349307
rect 132611 349189 132653 349307
rect 132771 349189 150493 349307
rect 150611 349189 150653 349307
rect 150771 349189 168493 349307
rect 168611 349189 168653 349307
rect 168771 349189 186493 349307
rect 186611 349189 186653 349307
rect 186771 349189 204493 349307
rect 204611 349189 204653 349307
rect 204771 349189 222493 349307
rect 222611 349189 222653 349307
rect 222771 349189 240493 349307
rect 240611 349189 240653 349307
rect 240771 349189 258493 349307
rect 258611 349189 258653 349307
rect 258771 349189 276493 349307
rect 276611 349189 276653 349307
rect 276771 349189 295551 349307
rect 295669 349189 295711 349307
rect 295829 349189 296325 349307
rect -4363 349147 296325 349189
rect -4363 349029 -3867 349147
rect -3749 349029 -3707 349147
rect -3589 349029 6493 349147
rect 6611 349029 6653 349147
rect 6771 349029 24493 349147
rect 24611 349029 24653 349147
rect 24771 349029 42493 349147
rect 42611 349029 42653 349147
rect 42771 349029 60493 349147
rect 60611 349029 60653 349147
rect 60771 349029 78493 349147
rect 78611 349029 78653 349147
rect 78771 349029 96493 349147
rect 96611 349029 96653 349147
rect 96771 349029 114493 349147
rect 114611 349029 114653 349147
rect 114771 349029 132493 349147
rect 132611 349029 132653 349147
rect 132771 349029 150493 349147
rect 150611 349029 150653 349147
rect 150771 349029 168493 349147
rect 168611 349029 168653 349147
rect 168771 349029 186493 349147
rect 186611 349029 186653 349147
rect 186771 349029 204493 349147
rect 204611 349029 204653 349147
rect 204771 349029 222493 349147
rect 222611 349029 222653 349147
rect 222771 349029 240493 349147
rect 240611 349029 240653 349147
rect 240771 349029 258493 349147
rect 258611 349029 258653 349147
rect 258771 349029 276493 349147
rect 276611 349029 276653 349147
rect 276771 349029 295551 349147
rect 295669 349029 295711 349147
rect 295829 349029 296325 349147
rect -4363 349013 296325 349029
rect -3403 347447 295365 347463
rect -3403 347329 -2907 347447
rect -2789 347329 -2747 347447
rect -2629 347329 4633 347447
rect 4751 347329 4793 347447
rect 4911 347329 22633 347447
rect 22751 347329 22793 347447
rect 22911 347329 40633 347447
rect 40751 347329 40793 347447
rect 40911 347329 58633 347447
rect 58751 347329 58793 347447
rect 58911 347329 76633 347447
rect 76751 347329 76793 347447
rect 76911 347329 94633 347447
rect 94751 347329 94793 347447
rect 94911 347329 112633 347447
rect 112751 347329 112793 347447
rect 112911 347329 130633 347447
rect 130751 347329 130793 347447
rect 130911 347329 148633 347447
rect 148751 347329 148793 347447
rect 148911 347329 166633 347447
rect 166751 347329 166793 347447
rect 166911 347329 184633 347447
rect 184751 347329 184793 347447
rect 184911 347329 202633 347447
rect 202751 347329 202793 347447
rect 202911 347329 220633 347447
rect 220751 347329 220793 347447
rect 220911 347329 238633 347447
rect 238751 347329 238793 347447
rect 238911 347329 256633 347447
rect 256751 347329 256793 347447
rect 256911 347329 274633 347447
rect 274751 347329 274793 347447
rect 274911 347329 294591 347447
rect 294709 347329 294751 347447
rect 294869 347329 295365 347447
rect -3403 347287 295365 347329
rect -3403 347169 -2907 347287
rect -2789 347169 -2747 347287
rect -2629 347169 4633 347287
rect 4751 347169 4793 347287
rect 4911 347169 22633 347287
rect 22751 347169 22793 347287
rect 22911 347169 40633 347287
rect 40751 347169 40793 347287
rect 40911 347169 58633 347287
rect 58751 347169 58793 347287
rect 58911 347169 76633 347287
rect 76751 347169 76793 347287
rect 76911 347169 94633 347287
rect 94751 347169 94793 347287
rect 94911 347169 112633 347287
rect 112751 347169 112793 347287
rect 112911 347169 130633 347287
rect 130751 347169 130793 347287
rect 130911 347169 148633 347287
rect 148751 347169 148793 347287
rect 148911 347169 166633 347287
rect 166751 347169 166793 347287
rect 166911 347169 184633 347287
rect 184751 347169 184793 347287
rect 184911 347169 202633 347287
rect 202751 347169 202793 347287
rect 202911 347169 220633 347287
rect 220751 347169 220793 347287
rect 220911 347169 238633 347287
rect 238751 347169 238793 347287
rect 238911 347169 256633 347287
rect 256751 347169 256793 347287
rect 256911 347169 274633 347287
rect 274751 347169 274793 347287
rect 274911 347169 294591 347287
rect 294709 347169 294751 347287
rect 294869 347169 295365 347287
rect -3403 347153 295365 347169
rect -2443 345587 294405 345603
rect -2443 345469 -1947 345587
rect -1829 345469 -1787 345587
rect -1669 345469 2773 345587
rect 2891 345469 2933 345587
rect 3051 345469 20773 345587
rect 20891 345469 20933 345587
rect 21051 345469 38773 345587
rect 38891 345469 38933 345587
rect 39051 345469 56773 345587
rect 56891 345469 56933 345587
rect 57051 345469 74773 345587
rect 74891 345469 74933 345587
rect 75051 345469 92773 345587
rect 92891 345469 92933 345587
rect 93051 345469 110773 345587
rect 110891 345469 110933 345587
rect 111051 345469 128773 345587
rect 128891 345469 128933 345587
rect 129051 345469 146773 345587
rect 146891 345469 146933 345587
rect 147051 345469 164773 345587
rect 164891 345469 164933 345587
rect 165051 345469 182773 345587
rect 182891 345469 182933 345587
rect 183051 345469 200773 345587
rect 200891 345469 200933 345587
rect 201051 345469 218773 345587
rect 218891 345469 218933 345587
rect 219051 345469 236773 345587
rect 236891 345469 236933 345587
rect 237051 345469 254773 345587
rect 254891 345469 254933 345587
rect 255051 345469 272773 345587
rect 272891 345469 272933 345587
rect 273051 345469 290773 345587
rect 290891 345469 290933 345587
rect 291051 345469 293631 345587
rect 293749 345469 293791 345587
rect 293909 345469 294405 345587
rect -2443 345427 294405 345469
rect -2443 345309 -1947 345427
rect -1829 345309 -1787 345427
rect -1669 345309 2773 345427
rect 2891 345309 2933 345427
rect 3051 345309 20773 345427
rect 20891 345309 20933 345427
rect 21051 345309 38773 345427
rect 38891 345309 38933 345427
rect 39051 345309 56773 345427
rect 56891 345309 56933 345427
rect 57051 345309 74773 345427
rect 74891 345309 74933 345427
rect 75051 345309 92773 345427
rect 92891 345309 92933 345427
rect 93051 345309 110773 345427
rect 110891 345309 110933 345427
rect 111051 345309 128773 345427
rect 128891 345309 128933 345427
rect 129051 345309 146773 345427
rect 146891 345309 146933 345427
rect 147051 345309 164773 345427
rect 164891 345309 164933 345427
rect 165051 345309 182773 345427
rect 182891 345309 182933 345427
rect 183051 345309 200773 345427
rect 200891 345309 200933 345427
rect 201051 345309 218773 345427
rect 218891 345309 218933 345427
rect 219051 345309 236773 345427
rect 236891 345309 236933 345427
rect 237051 345309 254773 345427
rect 254891 345309 254933 345427
rect 255051 345309 272773 345427
rect 272891 345309 272933 345427
rect 273051 345309 290773 345427
rect 290891 345309 290933 345427
rect 291051 345309 293631 345427
rect 293749 345309 293791 345427
rect 293909 345309 294405 345427
rect -2443 345293 294405 345309
rect -1483 343727 293445 343743
rect -1483 343609 -987 343727
rect -869 343609 -827 343727
rect -709 343609 913 343727
rect 1031 343609 1073 343727
rect 1191 343609 18913 343727
rect 19031 343609 19073 343727
rect 19191 343609 36913 343727
rect 37031 343609 37073 343727
rect 37191 343609 54913 343727
rect 55031 343609 55073 343727
rect 55191 343609 72913 343727
rect 73031 343609 73073 343727
rect 73191 343609 90913 343727
rect 91031 343609 91073 343727
rect 91191 343609 108913 343727
rect 109031 343609 109073 343727
rect 109191 343609 126913 343727
rect 127031 343609 127073 343727
rect 127191 343609 144913 343727
rect 145031 343609 145073 343727
rect 145191 343609 162913 343727
rect 163031 343609 163073 343727
rect 163191 343609 180913 343727
rect 181031 343609 181073 343727
rect 181191 343609 198913 343727
rect 199031 343609 199073 343727
rect 199191 343609 216913 343727
rect 217031 343609 217073 343727
rect 217191 343609 234913 343727
rect 235031 343609 235073 343727
rect 235191 343609 252913 343727
rect 253031 343609 253073 343727
rect 253191 343609 270913 343727
rect 271031 343609 271073 343727
rect 271191 343609 288913 343727
rect 289031 343609 289073 343727
rect 289191 343609 292671 343727
rect 292789 343609 292831 343727
rect 292949 343609 293445 343727
rect -1483 343567 293445 343609
rect -1483 343449 -987 343567
rect -869 343449 -827 343567
rect -709 343449 913 343567
rect 1031 343449 1073 343567
rect 1191 343449 18913 343567
rect 19031 343449 19073 343567
rect 19191 343449 36913 343567
rect 37031 343449 37073 343567
rect 37191 343449 54913 343567
rect 55031 343449 55073 343567
rect 55191 343449 72913 343567
rect 73031 343449 73073 343567
rect 73191 343449 90913 343567
rect 91031 343449 91073 343567
rect 91191 343449 108913 343567
rect 109031 343449 109073 343567
rect 109191 343449 126913 343567
rect 127031 343449 127073 343567
rect 127191 343449 144913 343567
rect 145031 343449 145073 343567
rect 145191 343449 162913 343567
rect 163031 343449 163073 343567
rect 163191 343449 180913 343567
rect 181031 343449 181073 343567
rect 181191 343449 198913 343567
rect 199031 343449 199073 343567
rect 199191 343449 216913 343567
rect 217031 343449 217073 343567
rect 217191 343449 234913 343567
rect 235031 343449 235073 343567
rect 235191 343449 252913 343567
rect 253031 343449 253073 343567
rect 253191 343449 270913 343567
rect 271031 343449 271073 343567
rect 271191 343449 288913 343567
rect 289031 343449 289073 343567
rect 289191 343449 292671 343567
rect 292789 343449 292831 343567
rect 292949 343449 293445 343567
rect -1483 343433 293445 343449
rect -4363 340307 296325 340323
rect -4363 340189 -4347 340307
rect -4229 340189 -4187 340307
rect -4069 340189 15493 340307
rect 15611 340189 15653 340307
rect 15771 340189 33493 340307
rect 33611 340189 33653 340307
rect 33771 340189 51493 340307
rect 51611 340189 51653 340307
rect 51771 340189 69493 340307
rect 69611 340189 69653 340307
rect 69771 340189 87493 340307
rect 87611 340189 87653 340307
rect 87771 340189 105493 340307
rect 105611 340189 105653 340307
rect 105771 340189 123493 340307
rect 123611 340189 123653 340307
rect 123771 340189 141493 340307
rect 141611 340189 141653 340307
rect 141771 340189 159493 340307
rect 159611 340189 159653 340307
rect 159771 340189 177493 340307
rect 177611 340189 177653 340307
rect 177771 340189 195493 340307
rect 195611 340189 195653 340307
rect 195771 340189 213493 340307
rect 213611 340189 213653 340307
rect 213771 340189 231493 340307
rect 231611 340189 231653 340307
rect 231771 340189 249493 340307
rect 249611 340189 249653 340307
rect 249771 340189 267493 340307
rect 267611 340189 267653 340307
rect 267771 340189 285493 340307
rect 285611 340189 285653 340307
rect 285771 340189 296031 340307
rect 296149 340189 296191 340307
rect 296309 340189 296325 340307
rect -4363 340147 296325 340189
rect -4363 340029 -4347 340147
rect -4229 340029 -4187 340147
rect -4069 340029 15493 340147
rect 15611 340029 15653 340147
rect 15771 340029 33493 340147
rect 33611 340029 33653 340147
rect 33771 340029 51493 340147
rect 51611 340029 51653 340147
rect 51771 340029 69493 340147
rect 69611 340029 69653 340147
rect 69771 340029 87493 340147
rect 87611 340029 87653 340147
rect 87771 340029 105493 340147
rect 105611 340029 105653 340147
rect 105771 340029 123493 340147
rect 123611 340029 123653 340147
rect 123771 340029 141493 340147
rect 141611 340029 141653 340147
rect 141771 340029 159493 340147
rect 159611 340029 159653 340147
rect 159771 340029 177493 340147
rect 177611 340029 177653 340147
rect 177771 340029 195493 340147
rect 195611 340029 195653 340147
rect 195771 340029 213493 340147
rect 213611 340029 213653 340147
rect 213771 340029 231493 340147
rect 231611 340029 231653 340147
rect 231771 340029 249493 340147
rect 249611 340029 249653 340147
rect 249771 340029 267493 340147
rect 267611 340029 267653 340147
rect 267771 340029 285493 340147
rect 285611 340029 285653 340147
rect 285771 340029 296031 340147
rect 296149 340029 296191 340147
rect 296309 340029 296325 340147
rect -4363 340013 296325 340029
rect -3403 338447 295365 338463
rect -3403 338329 -3387 338447
rect -3269 338329 -3227 338447
rect -3109 338329 13633 338447
rect 13751 338329 13793 338447
rect 13911 338329 31633 338447
rect 31751 338329 31793 338447
rect 31911 338329 49633 338447
rect 49751 338329 49793 338447
rect 49911 338329 67633 338447
rect 67751 338329 67793 338447
rect 67911 338329 85633 338447
rect 85751 338329 85793 338447
rect 85911 338329 103633 338447
rect 103751 338329 103793 338447
rect 103911 338329 121633 338447
rect 121751 338329 121793 338447
rect 121911 338329 139633 338447
rect 139751 338329 139793 338447
rect 139911 338329 157633 338447
rect 157751 338329 157793 338447
rect 157911 338329 175633 338447
rect 175751 338329 175793 338447
rect 175911 338329 193633 338447
rect 193751 338329 193793 338447
rect 193911 338329 211633 338447
rect 211751 338329 211793 338447
rect 211911 338329 229633 338447
rect 229751 338329 229793 338447
rect 229911 338329 247633 338447
rect 247751 338329 247793 338447
rect 247911 338329 265633 338447
rect 265751 338329 265793 338447
rect 265911 338329 283633 338447
rect 283751 338329 283793 338447
rect 283911 338329 295071 338447
rect 295189 338329 295231 338447
rect 295349 338329 295365 338447
rect -3403 338287 295365 338329
rect -3403 338169 -3387 338287
rect -3269 338169 -3227 338287
rect -3109 338169 13633 338287
rect 13751 338169 13793 338287
rect 13911 338169 31633 338287
rect 31751 338169 31793 338287
rect 31911 338169 49633 338287
rect 49751 338169 49793 338287
rect 49911 338169 67633 338287
rect 67751 338169 67793 338287
rect 67911 338169 85633 338287
rect 85751 338169 85793 338287
rect 85911 338169 103633 338287
rect 103751 338169 103793 338287
rect 103911 338169 121633 338287
rect 121751 338169 121793 338287
rect 121911 338169 139633 338287
rect 139751 338169 139793 338287
rect 139911 338169 157633 338287
rect 157751 338169 157793 338287
rect 157911 338169 175633 338287
rect 175751 338169 175793 338287
rect 175911 338169 193633 338287
rect 193751 338169 193793 338287
rect 193911 338169 211633 338287
rect 211751 338169 211793 338287
rect 211911 338169 229633 338287
rect 229751 338169 229793 338287
rect 229911 338169 247633 338287
rect 247751 338169 247793 338287
rect 247911 338169 265633 338287
rect 265751 338169 265793 338287
rect 265911 338169 283633 338287
rect 283751 338169 283793 338287
rect 283911 338169 295071 338287
rect 295189 338169 295231 338287
rect 295349 338169 295365 338287
rect -3403 338153 295365 338169
rect -2443 336587 294405 336603
rect -2443 336469 -2427 336587
rect -2309 336469 -2267 336587
rect -2149 336469 11773 336587
rect 11891 336469 11933 336587
rect 12051 336469 29773 336587
rect 29891 336469 29933 336587
rect 30051 336469 47773 336587
rect 47891 336469 47933 336587
rect 48051 336469 65773 336587
rect 65891 336469 65933 336587
rect 66051 336469 83773 336587
rect 83891 336469 83933 336587
rect 84051 336469 101773 336587
rect 101891 336469 101933 336587
rect 102051 336469 119773 336587
rect 119891 336469 119933 336587
rect 120051 336469 137773 336587
rect 137891 336469 137933 336587
rect 138051 336469 155773 336587
rect 155891 336469 155933 336587
rect 156051 336469 173773 336587
rect 173891 336469 173933 336587
rect 174051 336469 191773 336587
rect 191891 336469 191933 336587
rect 192051 336469 209773 336587
rect 209891 336469 209933 336587
rect 210051 336469 227773 336587
rect 227891 336469 227933 336587
rect 228051 336469 245773 336587
rect 245891 336469 245933 336587
rect 246051 336469 263773 336587
rect 263891 336469 263933 336587
rect 264051 336469 281773 336587
rect 281891 336469 281933 336587
rect 282051 336469 294111 336587
rect 294229 336469 294271 336587
rect 294389 336469 294405 336587
rect -2443 336427 294405 336469
rect -2443 336309 -2427 336427
rect -2309 336309 -2267 336427
rect -2149 336309 11773 336427
rect 11891 336309 11933 336427
rect 12051 336309 29773 336427
rect 29891 336309 29933 336427
rect 30051 336309 47773 336427
rect 47891 336309 47933 336427
rect 48051 336309 65773 336427
rect 65891 336309 65933 336427
rect 66051 336309 83773 336427
rect 83891 336309 83933 336427
rect 84051 336309 101773 336427
rect 101891 336309 101933 336427
rect 102051 336309 119773 336427
rect 119891 336309 119933 336427
rect 120051 336309 137773 336427
rect 137891 336309 137933 336427
rect 138051 336309 155773 336427
rect 155891 336309 155933 336427
rect 156051 336309 173773 336427
rect 173891 336309 173933 336427
rect 174051 336309 191773 336427
rect 191891 336309 191933 336427
rect 192051 336309 209773 336427
rect 209891 336309 209933 336427
rect 210051 336309 227773 336427
rect 227891 336309 227933 336427
rect 228051 336309 245773 336427
rect 245891 336309 245933 336427
rect 246051 336309 263773 336427
rect 263891 336309 263933 336427
rect 264051 336309 281773 336427
rect 281891 336309 281933 336427
rect 282051 336309 294111 336427
rect 294229 336309 294271 336427
rect 294389 336309 294405 336427
rect -2443 336293 294405 336309
rect -1483 334727 293445 334743
rect -1483 334609 -1467 334727
rect -1349 334609 -1307 334727
rect -1189 334609 9913 334727
rect 10031 334609 10073 334727
rect 10191 334609 27913 334727
rect 28031 334609 28073 334727
rect 28191 334609 45913 334727
rect 46031 334609 46073 334727
rect 46191 334609 63913 334727
rect 64031 334609 64073 334727
rect 64191 334609 81913 334727
rect 82031 334609 82073 334727
rect 82191 334609 99913 334727
rect 100031 334609 100073 334727
rect 100191 334609 117913 334727
rect 118031 334609 118073 334727
rect 118191 334609 135913 334727
rect 136031 334609 136073 334727
rect 136191 334609 153913 334727
rect 154031 334609 154073 334727
rect 154191 334609 171913 334727
rect 172031 334609 172073 334727
rect 172191 334609 189913 334727
rect 190031 334609 190073 334727
rect 190191 334609 207913 334727
rect 208031 334609 208073 334727
rect 208191 334609 225913 334727
rect 226031 334609 226073 334727
rect 226191 334609 243913 334727
rect 244031 334609 244073 334727
rect 244191 334609 261913 334727
rect 262031 334609 262073 334727
rect 262191 334609 279913 334727
rect 280031 334609 280073 334727
rect 280191 334609 293151 334727
rect 293269 334609 293311 334727
rect 293429 334609 293445 334727
rect -1483 334567 293445 334609
rect -1483 334449 -1467 334567
rect -1349 334449 -1307 334567
rect -1189 334449 9913 334567
rect 10031 334449 10073 334567
rect 10191 334449 27913 334567
rect 28031 334449 28073 334567
rect 28191 334449 45913 334567
rect 46031 334449 46073 334567
rect 46191 334449 63913 334567
rect 64031 334449 64073 334567
rect 64191 334449 81913 334567
rect 82031 334449 82073 334567
rect 82191 334449 99913 334567
rect 100031 334449 100073 334567
rect 100191 334449 117913 334567
rect 118031 334449 118073 334567
rect 118191 334449 135913 334567
rect 136031 334449 136073 334567
rect 136191 334449 153913 334567
rect 154031 334449 154073 334567
rect 154191 334449 171913 334567
rect 172031 334449 172073 334567
rect 172191 334449 189913 334567
rect 190031 334449 190073 334567
rect 190191 334449 207913 334567
rect 208031 334449 208073 334567
rect 208191 334449 225913 334567
rect 226031 334449 226073 334567
rect 226191 334449 243913 334567
rect 244031 334449 244073 334567
rect 244191 334449 261913 334567
rect 262031 334449 262073 334567
rect 262191 334449 279913 334567
rect 280031 334449 280073 334567
rect 280191 334449 293151 334567
rect 293269 334449 293311 334567
rect 293429 334449 293445 334567
rect -1483 334433 293445 334449
rect -4363 331307 296325 331323
rect -4363 331189 -3867 331307
rect -3749 331189 -3707 331307
rect -3589 331189 6493 331307
rect 6611 331189 6653 331307
rect 6771 331189 24493 331307
rect 24611 331189 24653 331307
rect 24771 331189 42493 331307
rect 42611 331189 42653 331307
rect 42771 331189 60493 331307
rect 60611 331189 60653 331307
rect 60771 331189 78493 331307
rect 78611 331189 78653 331307
rect 78771 331189 96493 331307
rect 96611 331189 96653 331307
rect 96771 331189 114493 331307
rect 114611 331189 114653 331307
rect 114771 331189 132493 331307
rect 132611 331189 132653 331307
rect 132771 331189 150493 331307
rect 150611 331189 150653 331307
rect 150771 331189 168493 331307
rect 168611 331189 168653 331307
rect 168771 331189 186493 331307
rect 186611 331189 186653 331307
rect 186771 331189 204493 331307
rect 204611 331189 204653 331307
rect 204771 331189 222493 331307
rect 222611 331189 222653 331307
rect 222771 331189 240493 331307
rect 240611 331189 240653 331307
rect 240771 331189 258493 331307
rect 258611 331189 258653 331307
rect 258771 331189 276493 331307
rect 276611 331189 276653 331307
rect 276771 331189 295551 331307
rect 295669 331189 295711 331307
rect 295829 331189 296325 331307
rect -4363 331147 296325 331189
rect -4363 331029 -3867 331147
rect -3749 331029 -3707 331147
rect -3589 331029 6493 331147
rect 6611 331029 6653 331147
rect 6771 331029 24493 331147
rect 24611 331029 24653 331147
rect 24771 331029 42493 331147
rect 42611 331029 42653 331147
rect 42771 331029 60493 331147
rect 60611 331029 60653 331147
rect 60771 331029 78493 331147
rect 78611 331029 78653 331147
rect 78771 331029 96493 331147
rect 96611 331029 96653 331147
rect 96771 331029 114493 331147
rect 114611 331029 114653 331147
rect 114771 331029 132493 331147
rect 132611 331029 132653 331147
rect 132771 331029 150493 331147
rect 150611 331029 150653 331147
rect 150771 331029 168493 331147
rect 168611 331029 168653 331147
rect 168771 331029 186493 331147
rect 186611 331029 186653 331147
rect 186771 331029 204493 331147
rect 204611 331029 204653 331147
rect 204771 331029 222493 331147
rect 222611 331029 222653 331147
rect 222771 331029 240493 331147
rect 240611 331029 240653 331147
rect 240771 331029 258493 331147
rect 258611 331029 258653 331147
rect 258771 331029 276493 331147
rect 276611 331029 276653 331147
rect 276771 331029 295551 331147
rect 295669 331029 295711 331147
rect 295829 331029 296325 331147
rect -4363 331013 296325 331029
rect -3403 329447 295365 329463
rect -3403 329329 -2907 329447
rect -2789 329329 -2747 329447
rect -2629 329329 4633 329447
rect 4751 329329 4793 329447
rect 4911 329329 22633 329447
rect 22751 329329 22793 329447
rect 22911 329329 40633 329447
rect 40751 329329 40793 329447
rect 40911 329329 58633 329447
rect 58751 329329 58793 329447
rect 58911 329329 76633 329447
rect 76751 329329 76793 329447
rect 76911 329329 94633 329447
rect 94751 329329 94793 329447
rect 94911 329329 112633 329447
rect 112751 329329 112793 329447
rect 112911 329329 130633 329447
rect 130751 329329 130793 329447
rect 130911 329329 148633 329447
rect 148751 329329 148793 329447
rect 148911 329329 166633 329447
rect 166751 329329 166793 329447
rect 166911 329329 184633 329447
rect 184751 329329 184793 329447
rect 184911 329329 202633 329447
rect 202751 329329 202793 329447
rect 202911 329329 220633 329447
rect 220751 329329 220793 329447
rect 220911 329329 238633 329447
rect 238751 329329 238793 329447
rect 238911 329329 256633 329447
rect 256751 329329 256793 329447
rect 256911 329329 274633 329447
rect 274751 329329 274793 329447
rect 274911 329329 294591 329447
rect 294709 329329 294751 329447
rect 294869 329329 295365 329447
rect -3403 329287 295365 329329
rect -3403 329169 -2907 329287
rect -2789 329169 -2747 329287
rect -2629 329169 4633 329287
rect 4751 329169 4793 329287
rect 4911 329169 22633 329287
rect 22751 329169 22793 329287
rect 22911 329169 40633 329287
rect 40751 329169 40793 329287
rect 40911 329169 58633 329287
rect 58751 329169 58793 329287
rect 58911 329169 76633 329287
rect 76751 329169 76793 329287
rect 76911 329169 94633 329287
rect 94751 329169 94793 329287
rect 94911 329169 112633 329287
rect 112751 329169 112793 329287
rect 112911 329169 130633 329287
rect 130751 329169 130793 329287
rect 130911 329169 148633 329287
rect 148751 329169 148793 329287
rect 148911 329169 166633 329287
rect 166751 329169 166793 329287
rect 166911 329169 184633 329287
rect 184751 329169 184793 329287
rect 184911 329169 202633 329287
rect 202751 329169 202793 329287
rect 202911 329169 220633 329287
rect 220751 329169 220793 329287
rect 220911 329169 238633 329287
rect 238751 329169 238793 329287
rect 238911 329169 256633 329287
rect 256751 329169 256793 329287
rect 256911 329169 274633 329287
rect 274751 329169 274793 329287
rect 274911 329169 294591 329287
rect 294709 329169 294751 329287
rect 294869 329169 295365 329287
rect -3403 329153 295365 329169
rect -2443 327587 294405 327603
rect -2443 327469 -1947 327587
rect -1829 327469 -1787 327587
rect -1669 327469 2773 327587
rect 2891 327469 2933 327587
rect 3051 327469 20773 327587
rect 20891 327469 20933 327587
rect 21051 327469 38773 327587
rect 38891 327469 38933 327587
rect 39051 327469 56773 327587
rect 56891 327469 56933 327587
rect 57051 327469 74773 327587
rect 74891 327469 74933 327587
rect 75051 327469 92773 327587
rect 92891 327469 92933 327587
rect 93051 327469 110773 327587
rect 110891 327469 110933 327587
rect 111051 327469 128773 327587
rect 128891 327469 128933 327587
rect 129051 327469 146773 327587
rect 146891 327469 146933 327587
rect 147051 327469 164773 327587
rect 164891 327469 164933 327587
rect 165051 327469 182773 327587
rect 182891 327469 182933 327587
rect 183051 327469 200773 327587
rect 200891 327469 200933 327587
rect 201051 327469 218773 327587
rect 218891 327469 218933 327587
rect 219051 327469 236773 327587
rect 236891 327469 236933 327587
rect 237051 327469 254773 327587
rect 254891 327469 254933 327587
rect 255051 327469 272773 327587
rect 272891 327469 272933 327587
rect 273051 327469 290773 327587
rect 290891 327469 290933 327587
rect 291051 327469 293631 327587
rect 293749 327469 293791 327587
rect 293909 327469 294405 327587
rect -2443 327427 294405 327469
rect -2443 327309 -1947 327427
rect -1829 327309 -1787 327427
rect -1669 327309 2773 327427
rect 2891 327309 2933 327427
rect 3051 327309 20773 327427
rect 20891 327309 20933 327427
rect 21051 327309 38773 327427
rect 38891 327309 38933 327427
rect 39051 327309 56773 327427
rect 56891 327309 56933 327427
rect 57051 327309 74773 327427
rect 74891 327309 74933 327427
rect 75051 327309 92773 327427
rect 92891 327309 92933 327427
rect 93051 327309 110773 327427
rect 110891 327309 110933 327427
rect 111051 327309 128773 327427
rect 128891 327309 128933 327427
rect 129051 327309 146773 327427
rect 146891 327309 146933 327427
rect 147051 327309 164773 327427
rect 164891 327309 164933 327427
rect 165051 327309 182773 327427
rect 182891 327309 182933 327427
rect 183051 327309 200773 327427
rect 200891 327309 200933 327427
rect 201051 327309 218773 327427
rect 218891 327309 218933 327427
rect 219051 327309 236773 327427
rect 236891 327309 236933 327427
rect 237051 327309 254773 327427
rect 254891 327309 254933 327427
rect 255051 327309 272773 327427
rect 272891 327309 272933 327427
rect 273051 327309 290773 327427
rect 290891 327309 290933 327427
rect 291051 327309 293631 327427
rect 293749 327309 293791 327427
rect 293909 327309 294405 327427
rect -2443 327293 294405 327309
rect -1483 325727 293445 325743
rect -1483 325609 -987 325727
rect -869 325609 -827 325727
rect -709 325609 913 325727
rect 1031 325609 1073 325727
rect 1191 325609 18913 325727
rect 19031 325609 19073 325727
rect 19191 325609 36913 325727
rect 37031 325609 37073 325727
rect 37191 325609 54913 325727
rect 55031 325609 55073 325727
rect 55191 325609 72913 325727
rect 73031 325609 73073 325727
rect 73191 325609 90913 325727
rect 91031 325609 91073 325727
rect 91191 325609 108913 325727
rect 109031 325609 109073 325727
rect 109191 325609 126913 325727
rect 127031 325609 127073 325727
rect 127191 325609 144913 325727
rect 145031 325609 145073 325727
rect 145191 325609 162913 325727
rect 163031 325609 163073 325727
rect 163191 325609 180913 325727
rect 181031 325609 181073 325727
rect 181191 325609 198913 325727
rect 199031 325609 199073 325727
rect 199191 325609 216913 325727
rect 217031 325609 217073 325727
rect 217191 325609 234913 325727
rect 235031 325609 235073 325727
rect 235191 325609 252913 325727
rect 253031 325609 253073 325727
rect 253191 325609 270913 325727
rect 271031 325609 271073 325727
rect 271191 325609 288913 325727
rect 289031 325609 289073 325727
rect 289191 325609 292671 325727
rect 292789 325609 292831 325727
rect 292949 325609 293445 325727
rect -1483 325567 293445 325609
rect -1483 325449 -987 325567
rect -869 325449 -827 325567
rect -709 325449 913 325567
rect 1031 325449 1073 325567
rect 1191 325449 18913 325567
rect 19031 325449 19073 325567
rect 19191 325449 36913 325567
rect 37031 325449 37073 325567
rect 37191 325449 54913 325567
rect 55031 325449 55073 325567
rect 55191 325449 72913 325567
rect 73031 325449 73073 325567
rect 73191 325449 90913 325567
rect 91031 325449 91073 325567
rect 91191 325449 108913 325567
rect 109031 325449 109073 325567
rect 109191 325449 126913 325567
rect 127031 325449 127073 325567
rect 127191 325449 144913 325567
rect 145031 325449 145073 325567
rect 145191 325449 162913 325567
rect 163031 325449 163073 325567
rect 163191 325449 180913 325567
rect 181031 325449 181073 325567
rect 181191 325449 198913 325567
rect 199031 325449 199073 325567
rect 199191 325449 216913 325567
rect 217031 325449 217073 325567
rect 217191 325449 234913 325567
rect 235031 325449 235073 325567
rect 235191 325449 252913 325567
rect 253031 325449 253073 325567
rect 253191 325449 270913 325567
rect 271031 325449 271073 325567
rect 271191 325449 288913 325567
rect 289031 325449 289073 325567
rect 289191 325449 292671 325567
rect 292789 325449 292831 325567
rect 292949 325449 293445 325567
rect -1483 325433 293445 325449
rect -4363 322307 296325 322323
rect -4363 322189 -4347 322307
rect -4229 322189 -4187 322307
rect -4069 322189 15493 322307
rect 15611 322189 15653 322307
rect 15771 322189 33493 322307
rect 33611 322189 33653 322307
rect 33771 322189 51493 322307
rect 51611 322189 51653 322307
rect 51771 322189 69493 322307
rect 69611 322189 69653 322307
rect 69771 322189 87493 322307
rect 87611 322189 87653 322307
rect 87771 322189 105493 322307
rect 105611 322189 105653 322307
rect 105771 322189 123493 322307
rect 123611 322189 123653 322307
rect 123771 322189 141493 322307
rect 141611 322189 141653 322307
rect 141771 322189 159493 322307
rect 159611 322189 159653 322307
rect 159771 322189 177493 322307
rect 177611 322189 177653 322307
rect 177771 322189 195493 322307
rect 195611 322189 195653 322307
rect 195771 322189 213493 322307
rect 213611 322189 213653 322307
rect 213771 322189 231493 322307
rect 231611 322189 231653 322307
rect 231771 322189 249493 322307
rect 249611 322189 249653 322307
rect 249771 322189 267493 322307
rect 267611 322189 267653 322307
rect 267771 322189 285493 322307
rect 285611 322189 285653 322307
rect 285771 322189 296031 322307
rect 296149 322189 296191 322307
rect 296309 322189 296325 322307
rect -4363 322147 296325 322189
rect -4363 322029 -4347 322147
rect -4229 322029 -4187 322147
rect -4069 322029 15493 322147
rect 15611 322029 15653 322147
rect 15771 322029 33493 322147
rect 33611 322029 33653 322147
rect 33771 322029 51493 322147
rect 51611 322029 51653 322147
rect 51771 322029 69493 322147
rect 69611 322029 69653 322147
rect 69771 322029 87493 322147
rect 87611 322029 87653 322147
rect 87771 322029 105493 322147
rect 105611 322029 105653 322147
rect 105771 322029 123493 322147
rect 123611 322029 123653 322147
rect 123771 322029 141493 322147
rect 141611 322029 141653 322147
rect 141771 322029 159493 322147
rect 159611 322029 159653 322147
rect 159771 322029 177493 322147
rect 177611 322029 177653 322147
rect 177771 322029 195493 322147
rect 195611 322029 195653 322147
rect 195771 322029 213493 322147
rect 213611 322029 213653 322147
rect 213771 322029 231493 322147
rect 231611 322029 231653 322147
rect 231771 322029 249493 322147
rect 249611 322029 249653 322147
rect 249771 322029 267493 322147
rect 267611 322029 267653 322147
rect 267771 322029 285493 322147
rect 285611 322029 285653 322147
rect 285771 322029 296031 322147
rect 296149 322029 296191 322147
rect 296309 322029 296325 322147
rect -4363 322013 296325 322029
rect -3403 320447 295365 320463
rect -3403 320329 -3387 320447
rect -3269 320329 -3227 320447
rect -3109 320329 13633 320447
rect 13751 320329 13793 320447
rect 13911 320329 31633 320447
rect 31751 320329 31793 320447
rect 31911 320329 49633 320447
rect 49751 320329 49793 320447
rect 49911 320329 67633 320447
rect 67751 320329 67793 320447
rect 67911 320329 85633 320447
rect 85751 320329 85793 320447
rect 85911 320329 103633 320447
rect 103751 320329 103793 320447
rect 103911 320329 121633 320447
rect 121751 320329 121793 320447
rect 121911 320329 139633 320447
rect 139751 320329 139793 320447
rect 139911 320329 157633 320447
rect 157751 320329 157793 320447
rect 157911 320329 175633 320447
rect 175751 320329 175793 320447
rect 175911 320329 193633 320447
rect 193751 320329 193793 320447
rect 193911 320329 211633 320447
rect 211751 320329 211793 320447
rect 211911 320329 229633 320447
rect 229751 320329 229793 320447
rect 229911 320329 247633 320447
rect 247751 320329 247793 320447
rect 247911 320329 265633 320447
rect 265751 320329 265793 320447
rect 265911 320329 283633 320447
rect 283751 320329 283793 320447
rect 283911 320329 295071 320447
rect 295189 320329 295231 320447
rect 295349 320329 295365 320447
rect -3403 320287 295365 320329
rect -3403 320169 -3387 320287
rect -3269 320169 -3227 320287
rect -3109 320169 13633 320287
rect 13751 320169 13793 320287
rect 13911 320169 31633 320287
rect 31751 320169 31793 320287
rect 31911 320169 49633 320287
rect 49751 320169 49793 320287
rect 49911 320169 67633 320287
rect 67751 320169 67793 320287
rect 67911 320169 85633 320287
rect 85751 320169 85793 320287
rect 85911 320169 103633 320287
rect 103751 320169 103793 320287
rect 103911 320169 121633 320287
rect 121751 320169 121793 320287
rect 121911 320169 139633 320287
rect 139751 320169 139793 320287
rect 139911 320169 157633 320287
rect 157751 320169 157793 320287
rect 157911 320169 175633 320287
rect 175751 320169 175793 320287
rect 175911 320169 193633 320287
rect 193751 320169 193793 320287
rect 193911 320169 211633 320287
rect 211751 320169 211793 320287
rect 211911 320169 229633 320287
rect 229751 320169 229793 320287
rect 229911 320169 247633 320287
rect 247751 320169 247793 320287
rect 247911 320169 265633 320287
rect 265751 320169 265793 320287
rect 265911 320169 283633 320287
rect 283751 320169 283793 320287
rect 283911 320169 295071 320287
rect 295189 320169 295231 320287
rect 295349 320169 295365 320287
rect -3403 320153 295365 320169
rect -2443 318587 294405 318603
rect -2443 318469 -2427 318587
rect -2309 318469 -2267 318587
rect -2149 318469 11773 318587
rect 11891 318469 11933 318587
rect 12051 318469 29773 318587
rect 29891 318469 29933 318587
rect 30051 318469 47773 318587
rect 47891 318469 47933 318587
rect 48051 318469 65773 318587
rect 65891 318469 65933 318587
rect 66051 318469 83773 318587
rect 83891 318469 83933 318587
rect 84051 318469 101773 318587
rect 101891 318469 101933 318587
rect 102051 318469 119773 318587
rect 119891 318469 119933 318587
rect 120051 318469 137773 318587
rect 137891 318469 137933 318587
rect 138051 318469 155773 318587
rect 155891 318469 155933 318587
rect 156051 318469 173773 318587
rect 173891 318469 173933 318587
rect 174051 318469 191773 318587
rect 191891 318469 191933 318587
rect 192051 318469 209773 318587
rect 209891 318469 209933 318587
rect 210051 318469 227773 318587
rect 227891 318469 227933 318587
rect 228051 318469 245773 318587
rect 245891 318469 245933 318587
rect 246051 318469 263773 318587
rect 263891 318469 263933 318587
rect 264051 318469 281773 318587
rect 281891 318469 281933 318587
rect 282051 318469 294111 318587
rect 294229 318469 294271 318587
rect 294389 318469 294405 318587
rect -2443 318427 294405 318469
rect -2443 318309 -2427 318427
rect -2309 318309 -2267 318427
rect -2149 318309 11773 318427
rect 11891 318309 11933 318427
rect 12051 318309 29773 318427
rect 29891 318309 29933 318427
rect 30051 318309 47773 318427
rect 47891 318309 47933 318427
rect 48051 318309 65773 318427
rect 65891 318309 65933 318427
rect 66051 318309 83773 318427
rect 83891 318309 83933 318427
rect 84051 318309 101773 318427
rect 101891 318309 101933 318427
rect 102051 318309 119773 318427
rect 119891 318309 119933 318427
rect 120051 318309 137773 318427
rect 137891 318309 137933 318427
rect 138051 318309 155773 318427
rect 155891 318309 155933 318427
rect 156051 318309 173773 318427
rect 173891 318309 173933 318427
rect 174051 318309 191773 318427
rect 191891 318309 191933 318427
rect 192051 318309 209773 318427
rect 209891 318309 209933 318427
rect 210051 318309 227773 318427
rect 227891 318309 227933 318427
rect 228051 318309 245773 318427
rect 245891 318309 245933 318427
rect 246051 318309 263773 318427
rect 263891 318309 263933 318427
rect 264051 318309 281773 318427
rect 281891 318309 281933 318427
rect 282051 318309 294111 318427
rect 294229 318309 294271 318427
rect 294389 318309 294405 318427
rect -2443 318293 294405 318309
rect -1483 316727 293445 316743
rect -1483 316609 -1467 316727
rect -1349 316609 -1307 316727
rect -1189 316609 9913 316727
rect 10031 316609 10073 316727
rect 10191 316609 27913 316727
rect 28031 316609 28073 316727
rect 28191 316609 45913 316727
rect 46031 316609 46073 316727
rect 46191 316609 63913 316727
rect 64031 316609 64073 316727
rect 64191 316609 81913 316727
rect 82031 316609 82073 316727
rect 82191 316609 99913 316727
rect 100031 316609 100073 316727
rect 100191 316609 117913 316727
rect 118031 316609 118073 316727
rect 118191 316609 135913 316727
rect 136031 316609 136073 316727
rect 136191 316609 153913 316727
rect 154031 316609 154073 316727
rect 154191 316609 171913 316727
rect 172031 316609 172073 316727
rect 172191 316609 189913 316727
rect 190031 316609 190073 316727
rect 190191 316609 207913 316727
rect 208031 316609 208073 316727
rect 208191 316609 225913 316727
rect 226031 316609 226073 316727
rect 226191 316609 243913 316727
rect 244031 316609 244073 316727
rect 244191 316609 261913 316727
rect 262031 316609 262073 316727
rect 262191 316609 279913 316727
rect 280031 316609 280073 316727
rect 280191 316609 293151 316727
rect 293269 316609 293311 316727
rect 293429 316609 293445 316727
rect -1483 316567 293445 316609
rect -1483 316449 -1467 316567
rect -1349 316449 -1307 316567
rect -1189 316449 9913 316567
rect 10031 316449 10073 316567
rect 10191 316449 27913 316567
rect 28031 316449 28073 316567
rect 28191 316449 45913 316567
rect 46031 316449 46073 316567
rect 46191 316449 63913 316567
rect 64031 316449 64073 316567
rect 64191 316449 81913 316567
rect 82031 316449 82073 316567
rect 82191 316449 99913 316567
rect 100031 316449 100073 316567
rect 100191 316449 117913 316567
rect 118031 316449 118073 316567
rect 118191 316449 135913 316567
rect 136031 316449 136073 316567
rect 136191 316449 153913 316567
rect 154031 316449 154073 316567
rect 154191 316449 171913 316567
rect 172031 316449 172073 316567
rect 172191 316449 189913 316567
rect 190031 316449 190073 316567
rect 190191 316449 207913 316567
rect 208031 316449 208073 316567
rect 208191 316449 225913 316567
rect 226031 316449 226073 316567
rect 226191 316449 243913 316567
rect 244031 316449 244073 316567
rect 244191 316449 261913 316567
rect 262031 316449 262073 316567
rect 262191 316449 279913 316567
rect 280031 316449 280073 316567
rect 280191 316449 293151 316567
rect 293269 316449 293311 316567
rect 293429 316449 293445 316567
rect -1483 316433 293445 316449
rect -4363 313307 296325 313323
rect -4363 313189 -3867 313307
rect -3749 313189 -3707 313307
rect -3589 313189 6493 313307
rect 6611 313189 6653 313307
rect 6771 313189 24493 313307
rect 24611 313189 24653 313307
rect 24771 313189 42493 313307
rect 42611 313189 42653 313307
rect 42771 313189 60493 313307
rect 60611 313189 60653 313307
rect 60771 313189 78493 313307
rect 78611 313189 78653 313307
rect 78771 313189 96493 313307
rect 96611 313189 96653 313307
rect 96771 313189 114493 313307
rect 114611 313189 114653 313307
rect 114771 313189 132493 313307
rect 132611 313189 132653 313307
rect 132771 313189 150493 313307
rect 150611 313189 150653 313307
rect 150771 313189 168493 313307
rect 168611 313189 168653 313307
rect 168771 313189 186493 313307
rect 186611 313189 186653 313307
rect 186771 313189 204493 313307
rect 204611 313189 204653 313307
rect 204771 313189 222493 313307
rect 222611 313189 222653 313307
rect 222771 313189 240493 313307
rect 240611 313189 240653 313307
rect 240771 313189 258493 313307
rect 258611 313189 258653 313307
rect 258771 313189 276493 313307
rect 276611 313189 276653 313307
rect 276771 313189 295551 313307
rect 295669 313189 295711 313307
rect 295829 313189 296325 313307
rect -4363 313147 296325 313189
rect -4363 313029 -3867 313147
rect -3749 313029 -3707 313147
rect -3589 313029 6493 313147
rect 6611 313029 6653 313147
rect 6771 313029 24493 313147
rect 24611 313029 24653 313147
rect 24771 313029 42493 313147
rect 42611 313029 42653 313147
rect 42771 313029 60493 313147
rect 60611 313029 60653 313147
rect 60771 313029 78493 313147
rect 78611 313029 78653 313147
rect 78771 313029 96493 313147
rect 96611 313029 96653 313147
rect 96771 313029 114493 313147
rect 114611 313029 114653 313147
rect 114771 313029 132493 313147
rect 132611 313029 132653 313147
rect 132771 313029 150493 313147
rect 150611 313029 150653 313147
rect 150771 313029 168493 313147
rect 168611 313029 168653 313147
rect 168771 313029 186493 313147
rect 186611 313029 186653 313147
rect 186771 313029 204493 313147
rect 204611 313029 204653 313147
rect 204771 313029 222493 313147
rect 222611 313029 222653 313147
rect 222771 313029 240493 313147
rect 240611 313029 240653 313147
rect 240771 313029 258493 313147
rect 258611 313029 258653 313147
rect 258771 313029 276493 313147
rect 276611 313029 276653 313147
rect 276771 313029 295551 313147
rect 295669 313029 295711 313147
rect 295829 313029 296325 313147
rect -4363 313013 296325 313029
rect -3403 311447 295365 311463
rect -3403 311329 -2907 311447
rect -2789 311329 -2747 311447
rect -2629 311329 4633 311447
rect 4751 311329 4793 311447
rect 4911 311329 22633 311447
rect 22751 311329 22793 311447
rect 22911 311329 40633 311447
rect 40751 311329 40793 311447
rect 40911 311329 58633 311447
rect 58751 311329 58793 311447
rect 58911 311329 76633 311447
rect 76751 311329 76793 311447
rect 76911 311329 94633 311447
rect 94751 311329 94793 311447
rect 94911 311329 112633 311447
rect 112751 311329 112793 311447
rect 112911 311329 130633 311447
rect 130751 311329 130793 311447
rect 130911 311329 148633 311447
rect 148751 311329 148793 311447
rect 148911 311329 166633 311447
rect 166751 311329 166793 311447
rect 166911 311329 184633 311447
rect 184751 311329 184793 311447
rect 184911 311329 202633 311447
rect 202751 311329 202793 311447
rect 202911 311329 220633 311447
rect 220751 311329 220793 311447
rect 220911 311329 238633 311447
rect 238751 311329 238793 311447
rect 238911 311329 256633 311447
rect 256751 311329 256793 311447
rect 256911 311329 274633 311447
rect 274751 311329 274793 311447
rect 274911 311329 294591 311447
rect 294709 311329 294751 311447
rect 294869 311329 295365 311447
rect -3403 311287 295365 311329
rect -3403 311169 -2907 311287
rect -2789 311169 -2747 311287
rect -2629 311169 4633 311287
rect 4751 311169 4793 311287
rect 4911 311169 22633 311287
rect 22751 311169 22793 311287
rect 22911 311169 40633 311287
rect 40751 311169 40793 311287
rect 40911 311169 58633 311287
rect 58751 311169 58793 311287
rect 58911 311169 76633 311287
rect 76751 311169 76793 311287
rect 76911 311169 94633 311287
rect 94751 311169 94793 311287
rect 94911 311169 112633 311287
rect 112751 311169 112793 311287
rect 112911 311169 130633 311287
rect 130751 311169 130793 311287
rect 130911 311169 148633 311287
rect 148751 311169 148793 311287
rect 148911 311169 166633 311287
rect 166751 311169 166793 311287
rect 166911 311169 184633 311287
rect 184751 311169 184793 311287
rect 184911 311169 202633 311287
rect 202751 311169 202793 311287
rect 202911 311169 220633 311287
rect 220751 311169 220793 311287
rect 220911 311169 238633 311287
rect 238751 311169 238793 311287
rect 238911 311169 256633 311287
rect 256751 311169 256793 311287
rect 256911 311169 274633 311287
rect 274751 311169 274793 311287
rect 274911 311169 294591 311287
rect 294709 311169 294751 311287
rect 294869 311169 295365 311287
rect -3403 311153 295365 311169
rect -2443 309587 294405 309603
rect -2443 309469 -1947 309587
rect -1829 309469 -1787 309587
rect -1669 309469 2773 309587
rect 2891 309469 2933 309587
rect 3051 309469 20773 309587
rect 20891 309469 20933 309587
rect 21051 309469 38773 309587
rect 38891 309469 38933 309587
rect 39051 309469 56773 309587
rect 56891 309469 56933 309587
rect 57051 309469 74773 309587
rect 74891 309469 74933 309587
rect 75051 309469 92773 309587
rect 92891 309469 92933 309587
rect 93051 309469 110773 309587
rect 110891 309469 110933 309587
rect 111051 309469 128773 309587
rect 128891 309469 128933 309587
rect 129051 309469 146773 309587
rect 146891 309469 146933 309587
rect 147051 309469 164773 309587
rect 164891 309469 164933 309587
rect 165051 309469 182773 309587
rect 182891 309469 182933 309587
rect 183051 309469 200773 309587
rect 200891 309469 200933 309587
rect 201051 309469 218773 309587
rect 218891 309469 218933 309587
rect 219051 309469 236773 309587
rect 236891 309469 236933 309587
rect 237051 309469 254773 309587
rect 254891 309469 254933 309587
rect 255051 309469 272773 309587
rect 272891 309469 272933 309587
rect 273051 309469 290773 309587
rect 290891 309469 290933 309587
rect 291051 309469 293631 309587
rect 293749 309469 293791 309587
rect 293909 309469 294405 309587
rect -2443 309427 294405 309469
rect -2443 309309 -1947 309427
rect -1829 309309 -1787 309427
rect -1669 309309 2773 309427
rect 2891 309309 2933 309427
rect 3051 309309 20773 309427
rect 20891 309309 20933 309427
rect 21051 309309 38773 309427
rect 38891 309309 38933 309427
rect 39051 309309 56773 309427
rect 56891 309309 56933 309427
rect 57051 309309 74773 309427
rect 74891 309309 74933 309427
rect 75051 309309 92773 309427
rect 92891 309309 92933 309427
rect 93051 309309 110773 309427
rect 110891 309309 110933 309427
rect 111051 309309 128773 309427
rect 128891 309309 128933 309427
rect 129051 309309 146773 309427
rect 146891 309309 146933 309427
rect 147051 309309 164773 309427
rect 164891 309309 164933 309427
rect 165051 309309 182773 309427
rect 182891 309309 182933 309427
rect 183051 309309 200773 309427
rect 200891 309309 200933 309427
rect 201051 309309 218773 309427
rect 218891 309309 218933 309427
rect 219051 309309 236773 309427
rect 236891 309309 236933 309427
rect 237051 309309 254773 309427
rect 254891 309309 254933 309427
rect 255051 309309 272773 309427
rect 272891 309309 272933 309427
rect 273051 309309 290773 309427
rect 290891 309309 290933 309427
rect 291051 309309 293631 309427
rect 293749 309309 293791 309427
rect 293909 309309 294405 309427
rect -2443 309293 294405 309309
rect -1483 307727 293445 307743
rect -1483 307609 -987 307727
rect -869 307609 -827 307727
rect -709 307609 913 307727
rect 1031 307609 1073 307727
rect 1191 307609 18913 307727
rect 19031 307609 19073 307727
rect 19191 307609 36913 307727
rect 37031 307609 37073 307727
rect 37191 307609 54913 307727
rect 55031 307609 55073 307727
rect 55191 307609 72913 307727
rect 73031 307609 73073 307727
rect 73191 307609 90913 307727
rect 91031 307609 91073 307727
rect 91191 307609 108913 307727
rect 109031 307609 109073 307727
rect 109191 307609 126913 307727
rect 127031 307609 127073 307727
rect 127191 307609 144913 307727
rect 145031 307609 145073 307727
rect 145191 307609 162913 307727
rect 163031 307609 163073 307727
rect 163191 307609 180913 307727
rect 181031 307609 181073 307727
rect 181191 307609 198913 307727
rect 199031 307609 199073 307727
rect 199191 307609 216913 307727
rect 217031 307609 217073 307727
rect 217191 307609 234913 307727
rect 235031 307609 235073 307727
rect 235191 307609 252913 307727
rect 253031 307609 253073 307727
rect 253191 307609 270913 307727
rect 271031 307609 271073 307727
rect 271191 307609 288913 307727
rect 289031 307609 289073 307727
rect 289191 307609 292671 307727
rect 292789 307609 292831 307727
rect 292949 307609 293445 307727
rect -1483 307567 293445 307609
rect -1483 307449 -987 307567
rect -869 307449 -827 307567
rect -709 307449 913 307567
rect 1031 307449 1073 307567
rect 1191 307449 18913 307567
rect 19031 307449 19073 307567
rect 19191 307449 36913 307567
rect 37031 307449 37073 307567
rect 37191 307449 54913 307567
rect 55031 307449 55073 307567
rect 55191 307449 72913 307567
rect 73031 307449 73073 307567
rect 73191 307449 90913 307567
rect 91031 307449 91073 307567
rect 91191 307449 108913 307567
rect 109031 307449 109073 307567
rect 109191 307449 126913 307567
rect 127031 307449 127073 307567
rect 127191 307449 144913 307567
rect 145031 307449 145073 307567
rect 145191 307449 162913 307567
rect 163031 307449 163073 307567
rect 163191 307449 180913 307567
rect 181031 307449 181073 307567
rect 181191 307449 198913 307567
rect 199031 307449 199073 307567
rect 199191 307449 216913 307567
rect 217031 307449 217073 307567
rect 217191 307449 234913 307567
rect 235031 307449 235073 307567
rect 235191 307449 252913 307567
rect 253031 307449 253073 307567
rect 253191 307449 270913 307567
rect 271031 307449 271073 307567
rect 271191 307449 288913 307567
rect 289031 307449 289073 307567
rect 289191 307449 292671 307567
rect 292789 307449 292831 307567
rect 292949 307449 293445 307567
rect -1483 307433 293445 307449
rect -4363 304307 296325 304323
rect -4363 304189 -4347 304307
rect -4229 304189 -4187 304307
rect -4069 304189 15493 304307
rect 15611 304189 15653 304307
rect 15771 304189 33493 304307
rect 33611 304189 33653 304307
rect 33771 304189 51493 304307
rect 51611 304189 51653 304307
rect 51771 304189 69493 304307
rect 69611 304189 69653 304307
rect 69771 304189 87493 304307
rect 87611 304189 87653 304307
rect 87771 304189 105493 304307
rect 105611 304189 105653 304307
rect 105771 304189 123493 304307
rect 123611 304189 123653 304307
rect 123771 304189 141493 304307
rect 141611 304189 141653 304307
rect 141771 304189 159493 304307
rect 159611 304189 159653 304307
rect 159771 304189 177493 304307
rect 177611 304189 177653 304307
rect 177771 304189 195493 304307
rect 195611 304189 195653 304307
rect 195771 304189 213493 304307
rect 213611 304189 213653 304307
rect 213771 304189 231493 304307
rect 231611 304189 231653 304307
rect 231771 304189 249493 304307
rect 249611 304189 249653 304307
rect 249771 304189 267493 304307
rect 267611 304189 267653 304307
rect 267771 304189 285493 304307
rect 285611 304189 285653 304307
rect 285771 304189 296031 304307
rect 296149 304189 296191 304307
rect 296309 304189 296325 304307
rect -4363 304147 296325 304189
rect -4363 304029 -4347 304147
rect -4229 304029 -4187 304147
rect -4069 304029 15493 304147
rect 15611 304029 15653 304147
rect 15771 304029 33493 304147
rect 33611 304029 33653 304147
rect 33771 304029 51493 304147
rect 51611 304029 51653 304147
rect 51771 304029 69493 304147
rect 69611 304029 69653 304147
rect 69771 304029 87493 304147
rect 87611 304029 87653 304147
rect 87771 304029 105493 304147
rect 105611 304029 105653 304147
rect 105771 304029 123493 304147
rect 123611 304029 123653 304147
rect 123771 304029 141493 304147
rect 141611 304029 141653 304147
rect 141771 304029 159493 304147
rect 159611 304029 159653 304147
rect 159771 304029 177493 304147
rect 177611 304029 177653 304147
rect 177771 304029 195493 304147
rect 195611 304029 195653 304147
rect 195771 304029 213493 304147
rect 213611 304029 213653 304147
rect 213771 304029 231493 304147
rect 231611 304029 231653 304147
rect 231771 304029 249493 304147
rect 249611 304029 249653 304147
rect 249771 304029 267493 304147
rect 267611 304029 267653 304147
rect 267771 304029 285493 304147
rect 285611 304029 285653 304147
rect 285771 304029 296031 304147
rect 296149 304029 296191 304147
rect 296309 304029 296325 304147
rect -4363 304013 296325 304029
rect -3403 302447 295365 302463
rect -3403 302329 -3387 302447
rect -3269 302329 -3227 302447
rect -3109 302329 13633 302447
rect 13751 302329 13793 302447
rect 13911 302329 31633 302447
rect 31751 302329 31793 302447
rect 31911 302329 49633 302447
rect 49751 302329 49793 302447
rect 49911 302329 67633 302447
rect 67751 302329 67793 302447
rect 67911 302329 85633 302447
rect 85751 302329 85793 302447
rect 85911 302329 103633 302447
rect 103751 302329 103793 302447
rect 103911 302329 121633 302447
rect 121751 302329 121793 302447
rect 121911 302329 139633 302447
rect 139751 302329 139793 302447
rect 139911 302329 157633 302447
rect 157751 302329 157793 302447
rect 157911 302329 175633 302447
rect 175751 302329 175793 302447
rect 175911 302329 193633 302447
rect 193751 302329 193793 302447
rect 193911 302329 211633 302447
rect 211751 302329 211793 302447
rect 211911 302329 229633 302447
rect 229751 302329 229793 302447
rect 229911 302329 247633 302447
rect 247751 302329 247793 302447
rect 247911 302329 265633 302447
rect 265751 302329 265793 302447
rect 265911 302329 283633 302447
rect 283751 302329 283793 302447
rect 283911 302329 295071 302447
rect 295189 302329 295231 302447
rect 295349 302329 295365 302447
rect -3403 302287 295365 302329
rect -3403 302169 -3387 302287
rect -3269 302169 -3227 302287
rect -3109 302169 13633 302287
rect 13751 302169 13793 302287
rect 13911 302169 31633 302287
rect 31751 302169 31793 302287
rect 31911 302169 49633 302287
rect 49751 302169 49793 302287
rect 49911 302169 67633 302287
rect 67751 302169 67793 302287
rect 67911 302169 85633 302287
rect 85751 302169 85793 302287
rect 85911 302169 103633 302287
rect 103751 302169 103793 302287
rect 103911 302169 121633 302287
rect 121751 302169 121793 302287
rect 121911 302169 139633 302287
rect 139751 302169 139793 302287
rect 139911 302169 157633 302287
rect 157751 302169 157793 302287
rect 157911 302169 175633 302287
rect 175751 302169 175793 302287
rect 175911 302169 193633 302287
rect 193751 302169 193793 302287
rect 193911 302169 211633 302287
rect 211751 302169 211793 302287
rect 211911 302169 229633 302287
rect 229751 302169 229793 302287
rect 229911 302169 247633 302287
rect 247751 302169 247793 302287
rect 247911 302169 265633 302287
rect 265751 302169 265793 302287
rect 265911 302169 283633 302287
rect 283751 302169 283793 302287
rect 283911 302169 295071 302287
rect 295189 302169 295231 302287
rect 295349 302169 295365 302287
rect -3403 302153 295365 302169
rect -2443 300587 294405 300603
rect -2443 300469 -2427 300587
rect -2309 300469 -2267 300587
rect -2149 300469 11773 300587
rect 11891 300469 11933 300587
rect 12051 300469 29773 300587
rect 29891 300469 29933 300587
rect 30051 300469 47773 300587
rect 47891 300469 47933 300587
rect 48051 300469 65773 300587
rect 65891 300469 65933 300587
rect 66051 300469 83773 300587
rect 83891 300469 83933 300587
rect 84051 300469 101773 300587
rect 101891 300469 101933 300587
rect 102051 300469 119773 300587
rect 119891 300469 119933 300587
rect 120051 300469 137773 300587
rect 137891 300469 137933 300587
rect 138051 300469 155773 300587
rect 155891 300469 155933 300587
rect 156051 300469 173773 300587
rect 173891 300469 173933 300587
rect 174051 300469 191773 300587
rect 191891 300469 191933 300587
rect 192051 300469 209773 300587
rect 209891 300469 209933 300587
rect 210051 300469 227773 300587
rect 227891 300469 227933 300587
rect 228051 300469 245773 300587
rect 245891 300469 245933 300587
rect 246051 300469 263773 300587
rect 263891 300469 263933 300587
rect 264051 300469 281773 300587
rect 281891 300469 281933 300587
rect 282051 300469 294111 300587
rect 294229 300469 294271 300587
rect 294389 300469 294405 300587
rect -2443 300427 294405 300469
rect -2443 300309 -2427 300427
rect -2309 300309 -2267 300427
rect -2149 300309 11773 300427
rect 11891 300309 11933 300427
rect 12051 300309 29773 300427
rect 29891 300309 29933 300427
rect 30051 300309 47773 300427
rect 47891 300309 47933 300427
rect 48051 300309 65773 300427
rect 65891 300309 65933 300427
rect 66051 300309 83773 300427
rect 83891 300309 83933 300427
rect 84051 300309 101773 300427
rect 101891 300309 101933 300427
rect 102051 300309 119773 300427
rect 119891 300309 119933 300427
rect 120051 300309 137773 300427
rect 137891 300309 137933 300427
rect 138051 300309 155773 300427
rect 155891 300309 155933 300427
rect 156051 300309 173773 300427
rect 173891 300309 173933 300427
rect 174051 300309 191773 300427
rect 191891 300309 191933 300427
rect 192051 300309 209773 300427
rect 209891 300309 209933 300427
rect 210051 300309 227773 300427
rect 227891 300309 227933 300427
rect 228051 300309 245773 300427
rect 245891 300309 245933 300427
rect 246051 300309 263773 300427
rect 263891 300309 263933 300427
rect 264051 300309 281773 300427
rect 281891 300309 281933 300427
rect 282051 300309 294111 300427
rect 294229 300309 294271 300427
rect 294389 300309 294405 300427
rect -2443 300293 294405 300309
rect -1483 298727 293445 298743
rect -1483 298609 -1467 298727
rect -1349 298609 -1307 298727
rect -1189 298609 9913 298727
rect 10031 298609 10073 298727
rect 10191 298609 27913 298727
rect 28031 298609 28073 298727
rect 28191 298609 45913 298727
rect 46031 298609 46073 298727
rect 46191 298609 63913 298727
rect 64031 298609 64073 298727
rect 64191 298609 81913 298727
rect 82031 298609 82073 298727
rect 82191 298609 99913 298727
rect 100031 298609 100073 298727
rect 100191 298609 117913 298727
rect 118031 298609 118073 298727
rect 118191 298609 135913 298727
rect 136031 298609 136073 298727
rect 136191 298609 153913 298727
rect 154031 298609 154073 298727
rect 154191 298609 171913 298727
rect 172031 298609 172073 298727
rect 172191 298609 189913 298727
rect 190031 298609 190073 298727
rect 190191 298609 207913 298727
rect 208031 298609 208073 298727
rect 208191 298609 225913 298727
rect 226031 298609 226073 298727
rect 226191 298609 243913 298727
rect 244031 298609 244073 298727
rect 244191 298609 261913 298727
rect 262031 298609 262073 298727
rect 262191 298609 279913 298727
rect 280031 298609 280073 298727
rect 280191 298609 293151 298727
rect 293269 298609 293311 298727
rect 293429 298609 293445 298727
rect -1483 298567 293445 298609
rect -1483 298449 -1467 298567
rect -1349 298449 -1307 298567
rect -1189 298449 9913 298567
rect 10031 298449 10073 298567
rect 10191 298449 27913 298567
rect 28031 298449 28073 298567
rect 28191 298449 45913 298567
rect 46031 298449 46073 298567
rect 46191 298449 63913 298567
rect 64031 298449 64073 298567
rect 64191 298449 81913 298567
rect 82031 298449 82073 298567
rect 82191 298449 99913 298567
rect 100031 298449 100073 298567
rect 100191 298449 117913 298567
rect 118031 298449 118073 298567
rect 118191 298449 135913 298567
rect 136031 298449 136073 298567
rect 136191 298449 153913 298567
rect 154031 298449 154073 298567
rect 154191 298449 171913 298567
rect 172031 298449 172073 298567
rect 172191 298449 189913 298567
rect 190031 298449 190073 298567
rect 190191 298449 207913 298567
rect 208031 298449 208073 298567
rect 208191 298449 225913 298567
rect 226031 298449 226073 298567
rect 226191 298449 243913 298567
rect 244031 298449 244073 298567
rect 244191 298449 261913 298567
rect 262031 298449 262073 298567
rect 262191 298449 279913 298567
rect 280031 298449 280073 298567
rect 280191 298449 293151 298567
rect 293269 298449 293311 298567
rect 293429 298449 293445 298567
rect -1483 298433 293445 298449
rect -4363 295307 296325 295323
rect -4363 295189 -3867 295307
rect -3749 295189 -3707 295307
rect -3589 295189 6493 295307
rect 6611 295189 6653 295307
rect 6771 295189 24493 295307
rect 24611 295189 24653 295307
rect 24771 295189 42493 295307
rect 42611 295189 42653 295307
rect 42771 295189 60493 295307
rect 60611 295189 60653 295307
rect 60771 295189 78493 295307
rect 78611 295189 78653 295307
rect 78771 295189 96493 295307
rect 96611 295189 96653 295307
rect 96771 295189 114493 295307
rect 114611 295189 114653 295307
rect 114771 295189 132493 295307
rect 132611 295189 132653 295307
rect 132771 295189 150493 295307
rect 150611 295189 150653 295307
rect 150771 295189 168493 295307
rect 168611 295189 168653 295307
rect 168771 295189 186493 295307
rect 186611 295189 186653 295307
rect 186771 295189 204493 295307
rect 204611 295189 204653 295307
rect 204771 295189 222493 295307
rect 222611 295189 222653 295307
rect 222771 295189 240493 295307
rect 240611 295189 240653 295307
rect 240771 295189 258493 295307
rect 258611 295189 258653 295307
rect 258771 295189 276493 295307
rect 276611 295189 276653 295307
rect 276771 295189 295551 295307
rect 295669 295189 295711 295307
rect 295829 295189 296325 295307
rect -4363 295147 296325 295189
rect -4363 295029 -3867 295147
rect -3749 295029 -3707 295147
rect -3589 295029 6493 295147
rect 6611 295029 6653 295147
rect 6771 295029 24493 295147
rect 24611 295029 24653 295147
rect 24771 295029 42493 295147
rect 42611 295029 42653 295147
rect 42771 295029 60493 295147
rect 60611 295029 60653 295147
rect 60771 295029 78493 295147
rect 78611 295029 78653 295147
rect 78771 295029 96493 295147
rect 96611 295029 96653 295147
rect 96771 295029 114493 295147
rect 114611 295029 114653 295147
rect 114771 295029 132493 295147
rect 132611 295029 132653 295147
rect 132771 295029 150493 295147
rect 150611 295029 150653 295147
rect 150771 295029 168493 295147
rect 168611 295029 168653 295147
rect 168771 295029 186493 295147
rect 186611 295029 186653 295147
rect 186771 295029 204493 295147
rect 204611 295029 204653 295147
rect 204771 295029 222493 295147
rect 222611 295029 222653 295147
rect 222771 295029 240493 295147
rect 240611 295029 240653 295147
rect 240771 295029 258493 295147
rect 258611 295029 258653 295147
rect 258771 295029 276493 295147
rect 276611 295029 276653 295147
rect 276771 295029 295551 295147
rect 295669 295029 295711 295147
rect 295829 295029 296325 295147
rect -4363 295013 296325 295029
rect -3403 293447 295365 293463
rect -3403 293329 -2907 293447
rect -2789 293329 -2747 293447
rect -2629 293329 4633 293447
rect 4751 293329 4793 293447
rect 4911 293329 22633 293447
rect 22751 293329 22793 293447
rect 22911 293329 40633 293447
rect 40751 293329 40793 293447
rect 40911 293329 58633 293447
rect 58751 293329 58793 293447
rect 58911 293329 76633 293447
rect 76751 293329 76793 293447
rect 76911 293329 94633 293447
rect 94751 293329 94793 293447
rect 94911 293329 112633 293447
rect 112751 293329 112793 293447
rect 112911 293329 130633 293447
rect 130751 293329 130793 293447
rect 130911 293329 148633 293447
rect 148751 293329 148793 293447
rect 148911 293329 166633 293447
rect 166751 293329 166793 293447
rect 166911 293329 184633 293447
rect 184751 293329 184793 293447
rect 184911 293329 202633 293447
rect 202751 293329 202793 293447
rect 202911 293329 220633 293447
rect 220751 293329 220793 293447
rect 220911 293329 238633 293447
rect 238751 293329 238793 293447
rect 238911 293329 256633 293447
rect 256751 293329 256793 293447
rect 256911 293329 274633 293447
rect 274751 293329 274793 293447
rect 274911 293329 294591 293447
rect 294709 293329 294751 293447
rect 294869 293329 295365 293447
rect -3403 293287 295365 293329
rect -3403 293169 -2907 293287
rect -2789 293169 -2747 293287
rect -2629 293169 4633 293287
rect 4751 293169 4793 293287
rect 4911 293169 22633 293287
rect 22751 293169 22793 293287
rect 22911 293169 40633 293287
rect 40751 293169 40793 293287
rect 40911 293169 58633 293287
rect 58751 293169 58793 293287
rect 58911 293169 76633 293287
rect 76751 293169 76793 293287
rect 76911 293169 94633 293287
rect 94751 293169 94793 293287
rect 94911 293169 112633 293287
rect 112751 293169 112793 293287
rect 112911 293169 130633 293287
rect 130751 293169 130793 293287
rect 130911 293169 148633 293287
rect 148751 293169 148793 293287
rect 148911 293169 166633 293287
rect 166751 293169 166793 293287
rect 166911 293169 184633 293287
rect 184751 293169 184793 293287
rect 184911 293169 202633 293287
rect 202751 293169 202793 293287
rect 202911 293169 220633 293287
rect 220751 293169 220793 293287
rect 220911 293169 238633 293287
rect 238751 293169 238793 293287
rect 238911 293169 256633 293287
rect 256751 293169 256793 293287
rect 256911 293169 274633 293287
rect 274751 293169 274793 293287
rect 274911 293169 294591 293287
rect 294709 293169 294751 293287
rect 294869 293169 295365 293287
rect -3403 293153 295365 293169
rect -2443 291587 294405 291603
rect -2443 291469 -1947 291587
rect -1829 291469 -1787 291587
rect -1669 291469 2773 291587
rect 2891 291469 2933 291587
rect 3051 291469 20773 291587
rect 20891 291469 20933 291587
rect 21051 291469 38773 291587
rect 38891 291469 38933 291587
rect 39051 291469 56773 291587
rect 56891 291469 56933 291587
rect 57051 291469 74773 291587
rect 74891 291469 74933 291587
rect 75051 291469 92773 291587
rect 92891 291469 92933 291587
rect 93051 291469 110773 291587
rect 110891 291469 110933 291587
rect 111051 291469 128773 291587
rect 128891 291469 128933 291587
rect 129051 291469 146773 291587
rect 146891 291469 146933 291587
rect 147051 291469 164773 291587
rect 164891 291469 164933 291587
rect 165051 291469 182773 291587
rect 182891 291469 182933 291587
rect 183051 291469 200773 291587
rect 200891 291469 200933 291587
rect 201051 291469 218773 291587
rect 218891 291469 218933 291587
rect 219051 291469 236773 291587
rect 236891 291469 236933 291587
rect 237051 291469 254773 291587
rect 254891 291469 254933 291587
rect 255051 291469 272773 291587
rect 272891 291469 272933 291587
rect 273051 291469 290773 291587
rect 290891 291469 290933 291587
rect 291051 291469 293631 291587
rect 293749 291469 293791 291587
rect 293909 291469 294405 291587
rect -2443 291427 294405 291469
rect -2443 291309 -1947 291427
rect -1829 291309 -1787 291427
rect -1669 291309 2773 291427
rect 2891 291309 2933 291427
rect 3051 291309 20773 291427
rect 20891 291309 20933 291427
rect 21051 291309 38773 291427
rect 38891 291309 38933 291427
rect 39051 291309 56773 291427
rect 56891 291309 56933 291427
rect 57051 291309 74773 291427
rect 74891 291309 74933 291427
rect 75051 291309 92773 291427
rect 92891 291309 92933 291427
rect 93051 291309 110773 291427
rect 110891 291309 110933 291427
rect 111051 291309 128773 291427
rect 128891 291309 128933 291427
rect 129051 291309 146773 291427
rect 146891 291309 146933 291427
rect 147051 291309 164773 291427
rect 164891 291309 164933 291427
rect 165051 291309 182773 291427
rect 182891 291309 182933 291427
rect 183051 291309 200773 291427
rect 200891 291309 200933 291427
rect 201051 291309 218773 291427
rect 218891 291309 218933 291427
rect 219051 291309 236773 291427
rect 236891 291309 236933 291427
rect 237051 291309 254773 291427
rect 254891 291309 254933 291427
rect 255051 291309 272773 291427
rect 272891 291309 272933 291427
rect 273051 291309 290773 291427
rect 290891 291309 290933 291427
rect 291051 291309 293631 291427
rect 293749 291309 293791 291427
rect 293909 291309 294405 291427
rect -2443 291293 294405 291309
rect -1483 289727 293445 289743
rect -1483 289609 -987 289727
rect -869 289609 -827 289727
rect -709 289609 913 289727
rect 1031 289609 1073 289727
rect 1191 289609 18913 289727
rect 19031 289609 19073 289727
rect 19191 289609 36913 289727
rect 37031 289609 37073 289727
rect 37191 289609 54913 289727
rect 55031 289609 55073 289727
rect 55191 289609 72913 289727
rect 73031 289609 73073 289727
rect 73191 289609 90913 289727
rect 91031 289609 91073 289727
rect 91191 289609 108913 289727
rect 109031 289609 109073 289727
rect 109191 289609 126913 289727
rect 127031 289609 127073 289727
rect 127191 289609 144913 289727
rect 145031 289609 145073 289727
rect 145191 289609 162913 289727
rect 163031 289609 163073 289727
rect 163191 289609 180913 289727
rect 181031 289609 181073 289727
rect 181191 289609 198913 289727
rect 199031 289609 199073 289727
rect 199191 289609 216913 289727
rect 217031 289609 217073 289727
rect 217191 289609 234913 289727
rect 235031 289609 235073 289727
rect 235191 289609 252913 289727
rect 253031 289609 253073 289727
rect 253191 289609 270913 289727
rect 271031 289609 271073 289727
rect 271191 289609 288913 289727
rect 289031 289609 289073 289727
rect 289191 289609 292671 289727
rect 292789 289609 292831 289727
rect 292949 289609 293445 289727
rect -1483 289567 293445 289609
rect -1483 289449 -987 289567
rect -869 289449 -827 289567
rect -709 289449 913 289567
rect 1031 289449 1073 289567
rect 1191 289449 18913 289567
rect 19031 289449 19073 289567
rect 19191 289449 36913 289567
rect 37031 289449 37073 289567
rect 37191 289449 54913 289567
rect 55031 289449 55073 289567
rect 55191 289449 72913 289567
rect 73031 289449 73073 289567
rect 73191 289449 90913 289567
rect 91031 289449 91073 289567
rect 91191 289449 108913 289567
rect 109031 289449 109073 289567
rect 109191 289449 126913 289567
rect 127031 289449 127073 289567
rect 127191 289449 144913 289567
rect 145031 289449 145073 289567
rect 145191 289449 162913 289567
rect 163031 289449 163073 289567
rect 163191 289449 180913 289567
rect 181031 289449 181073 289567
rect 181191 289449 198913 289567
rect 199031 289449 199073 289567
rect 199191 289449 216913 289567
rect 217031 289449 217073 289567
rect 217191 289449 234913 289567
rect 235031 289449 235073 289567
rect 235191 289449 252913 289567
rect 253031 289449 253073 289567
rect 253191 289449 270913 289567
rect 271031 289449 271073 289567
rect 271191 289449 288913 289567
rect 289031 289449 289073 289567
rect 289191 289449 292671 289567
rect 292789 289449 292831 289567
rect 292949 289449 293445 289567
rect -1483 289433 293445 289449
rect -4363 286307 296325 286323
rect -4363 286189 -4347 286307
rect -4229 286189 -4187 286307
rect -4069 286189 15493 286307
rect 15611 286189 15653 286307
rect 15771 286189 33493 286307
rect 33611 286189 33653 286307
rect 33771 286189 51493 286307
rect 51611 286189 51653 286307
rect 51771 286189 69493 286307
rect 69611 286189 69653 286307
rect 69771 286189 87493 286307
rect 87611 286189 87653 286307
rect 87771 286189 105493 286307
rect 105611 286189 105653 286307
rect 105771 286189 123493 286307
rect 123611 286189 123653 286307
rect 123771 286189 141493 286307
rect 141611 286189 141653 286307
rect 141771 286189 159493 286307
rect 159611 286189 159653 286307
rect 159771 286189 177493 286307
rect 177611 286189 177653 286307
rect 177771 286189 195493 286307
rect 195611 286189 195653 286307
rect 195771 286189 213493 286307
rect 213611 286189 213653 286307
rect 213771 286189 231493 286307
rect 231611 286189 231653 286307
rect 231771 286189 249493 286307
rect 249611 286189 249653 286307
rect 249771 286189 267493 286307
rect 267611 286189 267653 286307
rect 267771 286189 285493 286307
rect 285611 286189 285653 286307
rect 285771 286189 296031 286307
rect 296149 286189 296191 286307
rect 296309 286189 296325 286307
rect -4363 286147 296325 286189
rect -4363 286029 -4347 286147
rect -4229 286029 -4187 286147
rect -4069 286029 15493 286147
rect 15611 286029 15653 286147
rect 15771 286029 33493 286147
rect 33611 286029 33653 286147
rect 33771 286029 51493 286147
rect 51611 286029 51653 286147
rect 51771 286029 69493 286147
rect 69611 286029 69653 286147
rect 69771 286029 87493 286147
rect 87611 286029 87653 286147
rect 87771 286029 105493 286147
rect 105611 286029 105653 286147
rect 105771 286029 123493 286147
rect 123611 286029 123653 286147
rect 123771 286029 141493 286147
rect 141611 286029 141653 286147
rect 141771 286029 159493 286147
rect 159611 286029 159653 286147
rect 159771 286029 177493 286147
rect 177611 286029 177653 286147
rect 177771 286029 195493 286147
rect 195611 286029 195653 286147
rect 195771 286029 213493 286147
rect 213611 286029 213653 286147
rect 213771 286029 231493 286147
rect 231611 286029 231653 286147
rect 231771 286029 249493 286147
rect 249611 286029 249653 286147
rect 249771 286029 267493 286147
rect 267611 286029 267653 286147
rect 267771 286029 285493 286147
rect 285611 286029 285653 286147
rect 285771 286029 296031 286147
rect 296149 286029 296191 286147
rect 296309 286029 296325 286147
rect -4363 286013 296325 286029
rect -3403 284447 295365 284463
rect -3403 284329 -3387 284447
rect -3269 284329 -3227 284447
rect -3109 284329 13633 284447
rect 13751 284329 13793 284447
rect 13911 284329 31633 284447
rect 31751 284329 31793 284447
rect 31911 284329 49633 284447
rect 49751 284329 49793 284447
rect 49911 284329 67633 284447
rect 67751 284329 67793 284447
rect 67911 284329 85633 284447
rect 85751 284329 85793 284447
rect 85911 284329 103633 284447
rect 103751 284329 103793 284447
rect 103911 284329 121633 284447
rect 121751 284329 121793 284447
rect 121911 284329 139633 284447
rect 139751 284329 139793 284447
rect 139911 284329 157633 284447
rect 157751 284329 157793 284447
rect 157911 284329 175633 284447
rect 175751 284329 175793 284447
rect 175911 284329 193633 284447
rect 193751 284329 193793 284447
rect 193911 284329 211633 284447
rect 211751 284329 211793 284447
rect 211911 284329 229633 284447
rect 229751 284329 229793 284447
rect 229911 284329 247633 284447
rect 247751 284329 247793 284447
rect 247911 284329 265633 284447
rect 265751 284329 265793 284447
rect 265911 284329 283633 284447
rect 283751 284329 283793 284447
rect 283911 284329 295071 284447
rect 295189 284329 295231 284447
rect 295349 284329 295365 284447
rect -3403 284287 295365 284329
rect -3403 284169 -3387 284287
rect -3269 284169 -3227 284287
rect -3109 284169 13633 284287
rect 13751 284169 13793 284287
rect 13911 284169 31633 284287
rect 31751 284169 31793 284287
rect 31911 284169 49633 284287
rect 49751 284169 49793 284287
rect 49911 284169 67633 284287
rect 67751 284169 67793 284287
rect 67911 284169 85633 284287
rect 85751 284169 85793 284287
rect 85911 284169 103633 284287
rect 103751 284169 103793 284287
rect 103911 284169 121633 284287
rect 121751 284169 121793 284287
rect 121911 284169 139633 284287
rect 139751 284169 139793 284287
rect 139911 284169 157633 284287
rect 157751 284169 157793 284287
rect 157911 284169 175633 284287
rect 175751 284169 175793 284287
rect 175911 284169 193633 284287
rect 193751 284169 193793 284287
rect 193911 284169 211633 284287
rect 211751 284169 211793 284287
rect 211911 284169 229633 284287
rect 229751 284169 229793 284287
rect 229911 284169 247633 284287
rect 247751 284169 247793 284287
rect 247911 284169 265633 284287
rect 265751 284169 265793 284287
rect 265911 284169 283633 284287
rect 283751 284169 283793 284287
rect 283911 284169 295071 284287
rect 295189 284169 295231 284287
rect 295349 284169 295365 284287
rect -3403 284153 295365 284169
rect -2443 282587 294405 282603
rect -2443 282469 -2427 282587
rect -2309 282469 -2267 282587
rect -2149 282469 11773 282587
rect 11891 282469 11933 282587
rect 12051 282469 29773 282587
rect 29891 282469 29933 282587
rect 30051 282469 47773 282587
rect 47891 282469 47933 282587
rect 48051 282469 65773 282587
rect 65891 282469 65933 282587
rect 66051 282469 83773 282587
rect 83891 282469 83933 282587
rect 84051 282469 101773 282587
rect 101891 282469 101933 282587
rect 102051 282469 119773 282587
rect 119891 282469 119933 282587
rect 120051 282469 137773 282587
rect 137891 282469 137933 282587
rect 138051 282469 155773 282587
rect 155891 282469 155933 282587
rect 156051 282469 173773 282587
rect 173891 282469 173933 282587
rect 174051 282469 191773 282587
rect 191891 282469 191933 282587
rect 192051 282469 209773 282587
rect 209891 282469 209933 282587
rect 210051 282469 227773 282587
rect 227891 282469 227933 282587
rect 228051 282469 245773 282587
rect 245891 282469 245933 282587
rect 246051 282469 263773 282587
rect 263891 282469 263933 282587
rect 264051 282469 281773 282587
rect 281891 282469 281933 282587
rect 282051 282469 294111 282587
rect 294229 282469 294271 282587
rect 294389 282469 294405 282587
rect -2443 282427 294405 282469
rect -2443 282309 -2427 282427
rect -2309 282309 -2267 282427
rect -2149 282309 11773 282427
rect 11891 282309 11933 282427
rect 12051 282309 29773 282427
rect 29891 282309 29933 282427
rect 30051 282309 47773 282427
rect 47891 282309 47933 282427
rect 48051 282309 65773 282427
rect 65891 282309 65933 282427
rect 66051 282309 83773 282427
rect 83891 282309 83933 282427
rect 84051 282309 101773 282427
rect 101891 282309 101933 282427
rect 102051 282309 119773 282427
rect 119891 282309 119933 282427
rect 120051 282309 137773 282427
rect 137891 282309 137933 282427
rect 138051 282309 155773 282427
rect 155891 282309 155933 282427
rect 156051 282309 173773 282427
rect 173891 282309 173933 282427
rect 174051 282309 191773 282427
rect 191891 282309 191933 282427
rect 192051 282309 209773 282427
rect 209891 282309 209933 282427
rect 210051 282309 227773 282427
rect 227891 282309 227933 282427
rect 228051 282309 245773 282427
rect 245891 282309 245933 282427
rect 246051 282309 263773 282427
rect 263891 282309 263933 282427
rect 264051 282309 281773 282427
rect 281891 282309 281933 282427
rect 282051 282309 294111 282427
rect 294229 282309 294271 282427
rect 294389 282309 294405 282427
rect -2443 282293 294405 282309
rect -1483 280727 293445 280743
rect -1483 280609 -1467 280727
rect -1349 280609 -1307 280727
rect -1189 280609 9913 280727
rect 10031 280609 10073 280727
rect 10191 280609 27913 280727
rect 28031 280609 28073 280727
rect 28191 280609 45913 280727
rect 46031 280609 46073 280727
rect 46191 280609 63913 280727
rect 64031 280609 64073 280727
rect 64191 280609 81913 280727
rect 82031 280609 82073 280727
rect 82191 280609 99913 280727
rect 100031 280609 100073 280727
rect 100191 280609 117913 280727
rect 118031 280609 118073 280727
rect 118191 280609 135913 280727
rect 136031 280609 136073 280727
rect 136191 280609 153913 280727
rect 154031 280609 154073 280727
rect 154191 280609 171913 280727
rect 172031 280609 172073 280727
rect 172191 280609 189913 280727
rect 190031 280609 190073 280727
rect 190191 280609 207913 280727
rect 208031 280609 208073 280727
rect 208191 280609 225913 280727
rect 226031 280609 226073 280727
rect 226191 280609 243913 280727
rect 244031 280609 244073 280727
rect 244191 280609 261913 280727
rect 262031 280609 262073 280727
rect 262191 280609 279913 280727
rect 280031 280609 280073 280727
rect 280191 280609 293151 280727
rect 293269 280609 293311 280727
rect 293429 280609 293445 280727
rect -1483 280567 293445 280609
rect -1483 280449 -1467 280567
rect -1349 280449 -1307 280567
rect -1189 280449 9913 280567
rect 10031 280449 10073 280567
rect 10191 280449 27913 280567
rect 28031 280449 28073 280567
rect 28191 280449 45913 280567
rect 46031 280449 46073 280567
rect 46191 280449 63913 280567
rect 64031 280449 64073 280567
rect 64191 280449 81913 280567
rect 82031 280449 82073 280567
rect 82191 280449 99913 280567
rect 100031 280449 100073 280567
rect 100191 280449 117913 280567
rect 118031 280449 118073 280567
rect 118191 280449 135913 280567
rect 136031 280449 136073 280567
rect 136191 280449 153913 280567
rect 154031 280449 154073 280567
rect 154191 280449 171913 280567
rect 172031 280449 172073 280567
rect 172191 280449 189913 280567
rect 190031 280449 190073 280567
rect 190191 280449 207913 280567
rect 208031 280449 208073 280567
rect 208191 280449 225913 280567
rect 226031 280449 226073 280567
rect 226191 280449 243913 280567
rect 244031 280449 244073 280567
rect 244191 280449 261913 280567
rect 262031 280449 262073 280567
rect 262191 280449 279913 280567
rect 280031 280449 280073 280567
rect 280191 280449 293151 280567
rect 293269 280449 293311 280567
rect 293429 280449 293445 280567
rect -1483 280433 293445 280449
rect -4363 277307 296325 277323
rect -4363 277189 -3867 277307
rect -3749 277189 -3707 277307
rect -3589 277189 6493 277307
rect 6611 277189 6653 277307
rect 6771 277189 24493 277307
rect 24611 277189 24653 277307
rect 24771 277189 42493 277307
rect 42611 277189 42653 277307
rect 42771 277189 60493 277307
rect 60611 277189 60653 277307
rect 60771 277189 78493 277307
rect 78611 277189 78653 277307
rect 78771 277189 96493 277307
rect 96611 277189 96653 277307
rect 96771 277189 114493 277307
rect 114611 277189 114653 277307
rect 114771 277189 132493 277307
rect 132611 277189 132653 277307
rect 132771 277189 150493 277307
rect 150611 277189 150653 277307
rect 150771 277189 168493 277307
rect 168611 277189 168653 277307
rect 168771 277189 186493 277307
rect 186611 277189 186653 277307
rect 186771 277189 204493 277307
rect 204611 277189 204653 277307
rect 204771 277189 222493 277307
rect 222611 277189 222653 277307
rect 222771 277189 240493 277307
rect 240611 277189 240653 277307
rect 240771 277189 258493 277307
rect 258611 277189 258653 277307
rect 258771 277189 276493 277307
rect 276611 277189 276653 277307
rect 276771 277189 295551 277307
rect 295669 277189 295711 277307
rect 295829 277189 296325 277307
rect -4363 277147 296325 277189
rect -4363 277029 -3867 277147
rect -3749 277029 -3707 277147
rect -3589 277029 6493 277147
rect 6611 277029 6653 277147
rect 6771 277029 24493 277147
rect 24611 277029 24653 277147
rect 24771 277029 42493 277147
rect 42611 277029 42653 277147
rect 42771 277029 60493 277147
rect 60611 277029 60653 277147
rect 60771 277029 78493 277147
rect 78611 277029 78653 277147
rect 78771 277029 96493 277147
rect 96611 277029 96653 277147
rect 96771 277029 114493 277147
rect 114611 277029 114653 277147
rect 114771 277029 132493 277147
rect 132611 277029 132653 277147
rect 132771 277029 150493 277147
rect 150611 277029 150653 277147
rect 150771 277029 168493 277147
rect 168611 277029 168653 277147
rect 168771 277029 186493 277147
rect 186611 277029 186653 277147
rect 186771 277029 204493 277147
rect 204611 277029 204653 277147
rect 204771 277029 222493 277147
rect 222611 277029 222653 277147
rect 222771 277029 240493 277147
rect 240611 277029 240653 277147
rect 240771 277029 258493 277147
rect 258611 277029 258653 277147
rect 258771 277029 276493 277147
rect 276611 277029 276653 277147
rect 276771 277029 295551 277147
rect 295669 277029 295711 277147
rect 295829 277029 296325 277147
rect -4363 277013 296325 277029
rect -3403 275447 295365 275463
rect -3403 275329 -2907 275447
rect -2789 275329 -2747 275447
rect -2629 275329 4633 275447
rect 4751 275329 4793 275447
rect 4911 275329 22633 275447
rect 22751 275329 22793 275447
rect 22911 275329 40633 275447
rect 40751 275329 40793 275447
rect 40911 275329 58633 275447
rect 58751 275329 58793 275447
rect 58911 275329 76633 275447
rect 76751 275329 76793 275447
rect 76911 275329 94633 275447
rect 94751 275329 94793 275447
rect 94911 275329 112633 275447
rect 112751 275329 112793 275447
rect 112911 275329 130633 275447
rect 130751 275329 130793 275447
rect 130911 275329 148633 275447
rect 148751 275329 148793 275447
rect 148911 275329 166633 275447
rect 166751 275329 166793 275447
rect 166911 275329 184633 275447
rect 184751 275329 184793 275447
rect 184911 275329 202633 275447
rect 202751 275329 202793 275447
rect 202911 275329 220633 275447
rect 220751 275329 220793 275447
rect 220911 275329 238633 275447
rect 238751 275329 238793 275447
rect 238911 275329 256633 275447
rect 256751 275329 256793 275447
rect 256911 275329 274633 275447
rect 274751 275329 274793 275447
rect 274911 275329 294591 275447
rect 294709 275329 294751 275447
rect 294869 275329 295365 275447
rect -3403 275287 295365 275329
rect -3403 275169 -2907 275287
rect -2789 275169 -2747 275287
rect -2629 275169 4633 275287
rect 4751 275169 4793 275287
rect 4911 275169 22633 275287
rect 22751 275169 22793 275287
rect 22911 275169 40633 275287
rect 40751 275169 40793 275287
rect 40911 275169 58633 275287
rect 58751 275169 58793 275287
rect 58911 275169 76633 275287
rect 76751 275169 76793 275287
rect 76911 275169 94633 275287
rect 94751 275169 94793 275287
rect 94911 275169 112633 275287
rect 112751 275169 112793 275287
rect 112911 275169 130633 275287
rect 130751 275169 130793 275287
rect 130911 275169 148633 275287
rect 148751 275169 148793 275287
rect 148911 275169 166633 275287
rect 166751 275169 166793 275287
rect 166911 275169 184633 275287
rect 184751 275169 184793 275287
rect 184911 275169 202633 275287
rect 202751 275169 202793 275287
rect 202911 275169 220633 275287
rect 220751 275169 220793 275287
rect 220911 275169 238633 275287
rect 238751 275169 238793 275287
rect 238911 275169 256633 275287
rect 256751 275169 256793 275287
rect 256911 275169 274633 275287
rect 274751 275169 274793 275287
rect 274911 275169 294591 275287
rect 294709 275169 294751 275287
rect 294869 275169 295365 275287
rect -3403 275153 295365 275169
rect -2443 273587 294405 273603
rect -2443 273469 -1947 273587
rect -1829 273469 -1787 273587
rect -1669 273469 2773 273587
rect 2891 273469 2933 273587
rect 3051 273469 20773 273587
rect 20891 273469 20933 273587
rect 21051 273469 38773 273587
rect 38891 273469 38933 273587
rect 39051 273469 56773 273587
rect 56891 273469 56933 273587
rect 57051 273469 74773 273587
rect 74891 273469 74933 273587
rect 75051 273469 92773 273587
rect 92891 273469 92933 273587
rect 93051 273469 110773 273587
rect 110891 273469 110933 273587
rect 111051 273469 128773 273587
rect 128891 273469 128933 273587
rect 129051 273469 146773 273587
rect 146891 273469 146933 273587
rect 147051 273469 164773 273587
rect 164891 273469 164933 273587
rect 165051 273469 182773 273587
rect 182891 273469 182933 273587
rect 183051 273469 200773 273587
rect 200891 273469 200933 273587
rect 201051 273469 218773 273587
rect 218891 273469 218933 273587
rect 219051 273469 236773 273587
rect 236891 273469 236933 273587
rect 237051 273469 254773 273587
rect 254891 273469 254933 273587
rect 255051 273469 272773 273587
rect 272891 273469 272933 273587
rect 273051 273469 290773 273587
rect 290891 273469 290933 273587
rect 291051 273469 293631 273587
rect 293749 273469 293791 273587
rect 293909 273469 294405 273587
rect -2443 273427 294405 273469
rect -2443 273309 -1947 273427
rect -1829 273309 -1787 273427
rect -1669 273309 2773 273427
rect 2891 273309 2933 273427
rect 3051 273309 20773 273427
rect 20891 273309 20933 273427
rect 21051 273309 38773 273427
rect 38891 273309 38933 273427
rect 39051 273309 56773 273427
rect 56891 273309 56933 273427
rect 57051 273309 74773 273427
rect 74891 273309 74933 273427
rect 75051 273309 92773 273427
rect 92891 273309 92933 273427
rect 93051 273309 110773 273427
rect 110891 273309 110933 273427
rect 111051 273309 128773 273427
rect 128891 273309 128933 273427
rect 129051 273309 146773 273427
rect 146891 273309 146933 273427
rect 147051 273309 164773 273427
rect 164891 273309 164933 273427
rect 165051 273309 182773 273427
rect 182891 273309 182933 273427
rect 183051 273309 200773 273427
rect 200891 273309 200933 273427
rect 201051 273309 218773 273427
rect 218891 273309 218933 273427
rect 219051 273309 236773 273427
rect 236891 273309 236933 273427
rect 237051 273309 254773 273427
rect 254891 273309 254933 273427
rect 255051 273309 272773 273427
rect 272891 273309 272933 273427
rect 273051 273309 290773 273427
rect 290891 273309 290933 273427
rect 291051 273309 293631 273427
rect 293749 273309 293791 273427
rect 293909 273309 294405 273427
rect -2443 273293 294405 273309
rect -1483 271727 293445 271743
rect -1483 271609 -987 271727
rect -869 271609 -827 271727
rect -709 271609 913 271727
rect 1031 271609 1073 271727
rect 1191 271609 18913 271727
rect 19031 271609 19073 271727
rect 19191 271609 36913 271727
rect 37031 271609 37073 271727
rect 37191 271609 54913 271727
rect 55031 271609 55073 271727
rect 55191 271609 72913 271727
rect 73031 271609 73073 271727
rect 73191 271609 90913 271727
rect 91031 271609 91073 271727
rect 91191 271609 108913 271727
rect 109031 271609 109073 271727
rect 109191 271609 126913 271727
rect 127031 271609 127073 271727
rect 127191 271609 144913 271727
rect 145031 271609 145073 271727
rect 145191 271609 162913 271727
rect 163031 271609 163073 271727
rect 163191 271609 180913 271727
rect 181031 271609 181073 271727
rect 181191 271609 198913 271727
rect 199031 271609 199073 271727
rect 199191 271609 216913 271727
rect 217031 271609 217073 271727
rect 217191 271609 234913 271727
rect 235031 271609 235073 271727
rect 235191 271609 252913 271727
rect 253031 271609 253073 271727
rect 253191 271609 270913 271727
rect 271031 271609 271073 271727
rect 271191 271609 288913 271727
rect 289031 271609 289073 271727
rect 289191 271609 292671 271727
rect 292789 271609 292831 271727
rect 292949 271609 293445 271727
rect -1483 271567 293445 271609
rect -1483 271449 -987 271567
rect -869 271449 -827 271567
rect -709 271449 913 271567
rect 1031 271449 1073 271567
rect 1191 271449 18913 271567
rect 19031 271449 19073 271567
rect 19191 271449 36913 271567
rect 37031 271449 37073 271567
rect 37191 271449 54913 271567
rect 55031 271449 55073 271567
rect 55191 271449 72913 271567
rect 73031 271449 73073 271567
rect 73191 271449 90913 271567
rect 91031 271449 91073 271567
rect 91191 271449 108913 271567
rect 109031 271449 109073 271567
rect 109191 271449 126913 271567
rect 127031 271449 127073 271567
rect 127191 271449 144913 271567
rect 145031 271449 145073 271567
rect 145191 271449 162913 271567
rect 163031 271449 163073 271567
rect 163191 271449 180913 271567
rect 181031 271449 181073 271567
rect 181191 271449 198913 271567
rect 199031 271449 199073 271567
rect 199191 271449 216913 271567
rect 217031 271449 217073 271567
rect 217191 271449 234913 271567
rect 235031 271449 235073 271567
rect 235191 271449 252913 271567
rect 253031 271449 253073 271567
rect 253191 271449 270913 271567
rect 271031 271449 271073 271567
rect 271191 271449 288913 271567
rect 289031 271449 289073 271567
rect 289191 271449 292671 271567
rect 292789 271449 292831 271567
rect 292949 271449 293445 271567
rect -1483 271433 293445 271449
rect -4363 268307 296325 268323
rect -4363 268189 -4347 268307
rect -4229 268189 -4187 268307
rect -4069 268189 15493 268307
rect 15611 268189 15653 268307
rect 15771 268189 33493 268307
rect 33611 268189 33653 268307
rect 33771 268189 51493 268307
rect 51611 268189 51653 268307
rect 51771 268189 69493 268307
rect 69611 268189 69653 268307
rect 69771 268189 87493 268307
rect 87611 268189 87653 268307
rect 87771 268189 105493 268307
rect 105611 268189 105653 268307
rect 105771 268189 123493 268307
rect 123611 268189 123653 268307
rect 123771 268189 141493 268307
rect 141611 268189 141653 268307
rect 141771 268189 159493 268307
rect 159611 268189 159653 268307
rect 159771 268189 177493 268307
rect 177611 268189 177653 268307
rect 177771 268189 195493 268307
rect 195611 268189 195653 268307
rect 195771 268189 213493 268307
rect 213611 268189 213653 268307
rect 213771 268189 231493 268307
rect 231611 268189 231653 268307
rect 231771 268189 249493 268307
rect 249611 268189 249653 268307
rect 249771 268189 267493 268307
rect 267611 268189 267653 268307
rect 267771 268189 285493 268307
rect 285611 268189 285653 268307
rect 285771 268189 296031 268307
rect 296149 268189 296191 268307
rect 296309 268189 296325 268307
rect -4363 268147 296325 268189
rect -4363 268029 -4347 268147
rect -4229 268029 -4187 268147
rect -4069 268029 15493 268147
rect 15611 268029 15653 268147
rect 15771 268029 33493 268147
rect 33611 268029 33653 268147
rect 33771 268029 51493 268147
rect 51611 268029 51653 268147
rect 51771 268029 69493 268147
rect 69611 268029 69653 268147
rect 69771 268029 87493 268147
rect 87611 268029 87653 268147
rect 87771 268029 105493 268147
rect 105611 268029 105653 268147
rect 105771 268029 123493 268147
rect 123611 268029 123653 268147
rect 123771 268029 141493 268147
rect 141611 268029 141653 268147
rect 141771 268029 159493 268147
rect 159611 268029 159653 268147
rect 159771 268029 177493 268147
rect 177611 268029 177653 268147
rect 177771 268029 195493 268147
rect 195611 268029 195653 268147
rect 195771 268029 213493 268147
rect 213611 268029 213653 268147
rect 213771 268029 231493 268147
rect 231611 268029 231653 268147
rect 231771 268029 249493 268147
rect 249611 268029 249653 268147
rect 249771 268029 267493 268147
rect 267611 268029 267653 268147
rect 267771 268029 285493 268147
rect 285611 268029 285653 268147
rect 285771 268029 296031 268147
rect 296149 268029 296191 268147
rect 296309 268029 296325 268147
rect -4363 268013 296325 268029
rect -3403 266447 295365 266463
rect -3403 266329 -3387 266447
rect -3269 266329 -3227 266447
rect -3109 266329 13633 266447
rect 13751 266329 13793 266447
rect 13911 266329 31633 266447
rect 31751 266329 31793 266447
rect 31911 266329 49633 266447
rect 49751 266329 49793 266447
rect 49911 266329 67633 266447
rect 67751 266329 67793 266447
rect 67911 266329 85633 266447
rect 85751 266329 85793 266447
rect 85911 266329 103633 266447
rect 103751 266329 103793 266447
rect 103911 266329 121633 266447
rect 121751 266329 121793 266447
rect 121911 266329 139633 266447
rect 139751 266329 139793 266447
rect 139911 266329 157633 266447
rect 157751 266329 157793 266447
rect 157911 266329 175633 266447
rect 175751 266329 175793 266447
rect 175911 266329 193633 266447
rect 193751 266329 193793 266447
rect 193911 266329 211633 266447
rect 211751 266329 211793 266447
rect 211911 266329 229633 266447
rect 229751 266329 229793 266447
rect 229911 266329 247633 266447
rect 247751 266329 247793 266447
rect 247911 266329 265633 266447
rect 265751 266329 265793 266447
rect 265911 266329 283633 266447
rect 283751 266329 283793 266447
rect 283911 266329 295071 266447
rect 295189 266329 295231 266447
rect 295349 266329 295365 266447
rect -3403 266287 295365 266329
rect -3403 266169 -3387 266287
rect -3269 266169 -3227 266287
rect -3109 266169 13633 266287
rect 13751 266169 13793 266287
rect 13911 266169 31633 266287
rect 31751 266169 31793 266287
rect 31911 266169 49633 266287
rect 49751 266169 49793 266287
rect 49911 266169 67633 266287
rect 67751 266169 67793 266287
rect 67911 266169 85633 266287
rect 85751 266169 85793 266287
rect 85911 266169 103633 266287
rect 103751 266169 103793 266287
rect 103911 266169 121633 266287
rect 121751 266169 121793 266287
rect 121911 266169 139633 266287
rect 139751 266169 139793 266287
rect 139911 266169 157633 266287
rect 157751 266169 157793 266287
rect 157911 266169 175633 266287
rect 175751 266169 175793 266287
rect 175911 266169 193633 266287
rect 193751 266169 193793 266287
rect 193911 266169 211633 266287
rect 211751 266169 211793 266287
rect 211911 266169 229633 266287
rect 229751 266169 229793 266287
rect 229911 266169 247633 266287
rect 247751 266169 247793 266287
rect 247911 266169 265633 266287
rect 265751 266169 265793 266287
rect 265911 266169 283633 266287
rect 283751 266169 283793 266287
rect 283911 266169 295071 266287
rect 295189 266169 295231 266287
rect 295349 266169 295365 266287
rect -3403 266153 295365 266169
rect -2443 264587 294405 264603
rect -2443 264469 -2427 264587
rect -2309 264469 -2267 264587
rect -2149 264469 11773 264587
rect 11891 264469 11933 264587
rect 12051 264469 29773 264587
rect 29891 264469 29933 264587
rect 30051 264469 47773 264587
rect 47891 264469 47933 264587
rect 48051 264469 65773 264587
rect 65891 264469 65933 264587
rect 66051 264469 83773 264587
rect 83891 264469 83933 264587
rect 84051 264469 101773 264587
rect 101891 264469 101933 264587
rect 102051 264469 119773 264587
rect 119891 264469 119933 264587
rect 120051 264469 137773 264587
rect 137891 264469 137933 264587
rect 138051 264469 155773 264587
rect 155891 264469 155933 264587
rect 156051 264469 173773 264587
rect 173891 264469 173933 264587
rect 174051 264469 191773 264587
rect 191891 264469 191933 264587
rect 192051 264469 209773 264587
rect 209891 264469 209933 264587
rect 210051 264469 227773 264587
rect 227891 264469 227933 264587
rect 228051 264469 245773 264587
rect 245891 264469 245933 264587
rect 246051 264469 263773 264587
rect 263891 264469 263933 264587
rect 264051 264469 281773 264587
rect 281891 264469 281933 264587
rect 282051 264469 294111 264587
rect 294229 264469 294271 264587
rect 294389 264469 294405 264587
rect -2443 264427 294405 264469
rect -2443 264309 -2427 264427
rect -2309 264309 -2267 264427
rect -2149 264309 11773 264427
rect 11891 264309 11933 264427
rect 12051 264309 29773 264427
rect 29891 264309 29933 264427
rect 30051 264309 47773 264427
rect 47891 264309 47933 264427
rect 48051 264309 65773 264427
rect 65891 264309 65933 264427
rect 66051 264309 83773 264427
rect 83891 264309 83933 264427
rect 84051 264309 101773 264427
rect 101891 264309 101933 264427
rect 102051 264309 119773 264427
rect 119891 264309 119933 264427
rect 120051 264309 137773 264427
rect 137891 264309 137933 264427
rect 138051 264309 155773 264427
rect 155891 264309 155933 264427
rect 156051 264309 173773 264427
rect 173891 264309 173933 264427
rect 174051 264309 191773 264427
rect 191891 264309 191933 264427
rect 192051 264309 209773 264427
rect 209891 264309 209933 264427
rect 210051 264309 227773 264427
rect 227891 264309 227933 264427
rect 228051 264309 245773 264427
rect 245891 264309 245933 264427
rect 246051 264309 263773 264427
rect 263891 264309 263933 264427
rect 264051 264309 281773 264427
rect 281891 264309 281933 264427
rect 282051 264309 294111 264427
rect 294229 264309 294271 264427
rect 294389 264309 294405 264427
rect -2443 264293 294405 264309
rect -1483 262727 293445 262743
rect -1483 262609 -1467 262727
rect -1349 262609 -1307 262727
rect -1189 262609 9913 262727
rect 10031 262609 10073 262727
rect 10191 262609 27913 262727
rect 28031 262609 28073 262727
rect 28191 262609 45913 262727
rect 46031 262609 46073 262727
rect 46191 262609 63913 262727
rect 64031 262609 64073 262727
rect 64191 262609 81913 262727
rect 82031 262609 82073 262727
rect 82191 262609 99913 262727
rect 100031 262609 100073 262727
rect 100191 262609 117913 262727
rect 118031 262609 118073 262727
rect 118191 262609 135913 262727
rect 136031 262609 136073 262727
rect 136191 262609 153913 262727
rect 154031 262609 154073 262727
rect 154191 262609 171913 262727
rect 172031 262609 172073 262727
rect 172191 262609 189913 262727
rect 190031 262609 190073 262727
rect 190191 262609 207913 262727
rect 208031 262609 208073 262727
rect 208191 262609 225913 262727
rect 226031 262609 226073 262727
rect 226191 262609 243913 262727
rect 244031 262609 244073 262727
rect 244191 262609 261913 262727
rect 262031 262609 262073 262727
rect 262191 262609 279913 262727
rect 280031 262609 280073 262727
rect 280191 262609 293151 262727
rect 293269 262609 293311 262727
rect 293429 262609 293445 262727
rect -1483 262567 293445 262609
rect -1483 262449 -1467 262567
rect -1349 262449 -1307 262567
rect -1189 262449 9913 262567
rect 10031 262449 10073 262567
rect 10191 262449 27913 262567
rect 28031 262449 28073 262567
rect 28191 262449 45913 262567
rect 46031 262449 46073 262567
rect 46191 262449 63913 262567
rect 64031 262449 64073 262567
rect 64191 262449 81913 262567
rect 82031 262449 82073 262567
rect 82191 262449 99913 262567
rect 100031 262449 100073 262567
rect 100191 262449 117913 262567
rect 118031 262449 118073 262567
rect 118191 262449 135913 262567
rect 136031 262449 136073 262567
rect 136191 262449 153913 262567
rect 154031 262449 154073 262567
rect 154191 262449 171913 262567
rect 172031 262449 172073 262567
rect 172191 262449 189913 262567
rect 190031 262449 190073 262567
rect 190191 262449 207913 262567
rect 208031 262449 208073 262567
rect 208191 262449 225913 262567
rect 226031 262449 226073 262567
rect 226191 262449 243913 262567
rect 244031 262449 244073 262567
rect 244191 262449 261913 262567
rect 262031 262449 262073 262567
rect 262191 262449 279913 262567
rect 280031 262449 280073 262567
rect 280191 262449 293151 262567
rect 293269 262449 293311 262567
rect 293429 262449 293445 262567
rect -1483 262433 293445 262449
rect -4363 259307 296325 259323
rect -4363 259189 -3867 259307
rect -3749 259189 -3707 259307
rect -3589 259189 6493 259307
rect 6611 259189 6653 259307
rect 6771 259189 24493 259307
rect 24611 259189 24653 259307
rect 24771 259189 42493 259307
rect 42611 259189 42653 259307
rect 42771 259189 60493 259307
rect 60611 259189 60653 259307
rect 60771 259189 78493 259307
rect 78611 259189 78653 259307
rect 78771 259189 96493 259307
rect 96611 259189 96653 259307
rect 96771 259189 114493 259307
rect 114611 259189 114653 259307
rect 114771 259189 132493 259307
rect 132611 259189 132653 259307
rect 132771 259189 150493 259307
rect 150611 259189 150653 259307
rect 150771 259189 168493 259307
rect 168611 259189 168653 259307
rect 168771 259189 186493 259307
rect 186611 259189 186653 259307
rect 186771 259189 204493 259307
rect 204611 259189 204653 259307
rect 204771 259189 222493 259307
rect 222611 259189 222653 259307
rect 222771 259189 240493 259307
rect 240611 259189 240653 259307
rect 240771 259189 258493 259307
rect 258611 259189 258653 259307
rect 258771 259189 276493 259307
rect 276611 259189 276653 259307
rect 276771 259189 295551 259307
rect 295669 259189 295711 259307
rect 295829 259189 296325 259307
rect -4363 259147 296325 259189
rect -4363 259029 -3867 259147
rect -3749 259029 -3707 259147
rect -3589 259029 6493 259147
rect 6611 259029 6653 259147
rect 6771 259029 24493 259147
rect 24611 259029 24653 259147
rect 24771 259029 42493 259147
rect 42611 259029 42653 259147
rect 42771 259029 60493 259147
rect 60611 259029 60653 259147
rect 60771 259029 78493 259147
rect 78611 259029 78653 259147
rect 78771 259029 96493 259147
rect 96611 259029 96653 259147
rect 96771 259029 114493 259147
rect 114611 259029 114653 259147
rect 114771 259029 132493 259147
rect 132611 259029 132653 259147
rect 132771 259029 150493 259147
rect 150611 259029 150653 259147
rect 150771 259029 168493 259147
rect 168611 259029 168653 259147
rect 168771 259029 186493 259147
rect 186611 259029 186653 259147
rect 186771 259029 204493 259147
rect 204611 259029 204653 259147
rect 204771 259029 222493 259147
rect 222611 259029 222653 259147
rect 222771 259029 240493 259147
rect 240611 259029 240653 259147
rect 240771 259029 258493 259147
rect 258611 259029 258653 259147
rect 258771 259029 276493 259147
rect 276611 259029 276653 259147
rect 276771 259029 295551 259147
rect 295669 259029 295711 259147
rect 295829 259029 296325 259147
rect -4363 259013 296325 259029
rect -3403 257447 295365 257463
rect -3403 257329 -2907 257447
rect -2789 257329 -2747 257447
rect -2629 257329 4633 257447
rect 4751 257329 4793 257447
rect 4911 257329 22633 257447
rect 22751 257329 22793 257447
rect 22911 257329 40633 257447
rect 40751 257329 40793 257447
rect 40911 257329 58633 257447
rect 58751 257329 58793 257447
rect 58911 257329 76633 257447
rect 76751 257329 76793 257447
rect 76911 257329 94633 257447
rect 94751 257329 94793 257447
rect 94911 257329 112633 257447
rect 112751 257329 112793 257447
rect 112911 257329 130633 257447
rect 130751 257329 130793 257447
rect 130911 257329 148633 257447
rect 148751 257329 148793 257447
rect 148911 257329 166633 257447
rect 166751 257329 166793 257447
rect 166911 257329 184633 257447
rect 184751 257329 184793 257447
rect 184911 257329 202633 257447
rect 202751 257329 202793 257447
rect 202911 257329 220633 257447
rect 220751 257329 220793 257447
rect 220911 257329 238633 257447
rect 238751 257329 238793 257447
rect 238911 257329 256633 257447
rect 256751 257329 256793 257447
rect 256911 257329 274633 257447
rect 274751 257329 274793 257447
rect 274911 257329 294591 257447
rect 294709 257329 294751 257447
rect 294869 257329 295365 257447
rect -3403 257287 295365 257329
rect -3403 257169 -2907 257287
rect -2789 257169 -2747 257287
rect -2629 257169 4633 257287
rect 4751 257169 4793 257287
rect 4911 257169 22633 257287
rect 22751 257169 22793 257287
rect 22911 257169 40633 257287
rect 40751 257169 40793 257287
rect 40911 257169 58633 257287
rect 58751 257169 58793 257287
rect 58911 257169 76633 257287
rect 76751 257169 76793 257287
rect 76911 257169 94633 257287
rect 94751 257169 94793 257287
rect 94911 257169 112633 257287
rect 112751 257169 112793 257287
rect 112911 257169 130633 257287
rect 130751 257169 130793 257287
rect 130911 257169 148633 257287
rect 148751 257169 148793 257287
rect 148911 257169 166633 257287
rect 166751 257169 166793 257287
rect 166911 257169 184633 257287
rect 184751 257169 184793 257287
rect 184911 257169 202633 257287
rect 202751 257169 202793 257287
rect 202911 257169 220633 257287
rect 220751 257169 220793 257287
rect 220911 257169 238633 257287
rect 238751 257169 238793 257287
rect 238911 257169 256633 257287
rect 256751 257169 256793 257287
rect 256911 257169 274633 257287
rect 274751 257169 274793 257287
rect 274911 257169 294591 257287
rect 294709 257169 294751 257287
rect 294869 257169 295365 257287
rect -3403 257153 295365 257169
rect -2443 255587 294405 255603
rect -2443 255469 -1947 255587
rect -1829 255469 -1787 255587
rect -1669 255469 2773 255587
rect 2891 255469 2933 255587
rect 3051 255469 20773 255587
rect 20891 255469 20933 255587
rect 21051 255469 38773 255587
rect 38891 255469 38933 255587
rect 39051 255469 56773 255587
rect 56891 255469 56933 255587
rect 57051 255469 74773 255587
rect 74891 255469 74933 255587
rect 75051 255469 92773 255587
rect 92891 255469 92933 255587
rect 93051 255469 110773 255587
rect 110891 255469 110933 255587
rect 111051 255469 128773 255587
rect 128891 255469 128933 255587
rect 129051 255469 146773 255587
rect 146891 255469 146933 255587
rect 147051 255469 164773 255587
rect 164891 255469 164933 255587
rect 165051 255469 182773 255587
rect 182891 255469 182933 255587
rect 183051 255469 200773 255587
rect 200891 255469 200933 255587
rect 201051 255469 218773 255587
rect 218891 255469 218933 255587
rect 219051 255469 236773 255587
rect 236891 255469 236933 255587
rect 237051 255469 254773 255587
rect 254891 255469 254933 255587
rect 255051 255469 272773 255587
rect 272891 255469 272933 255587
rect 273051 255469 290773 255587
rect 290891 255469 290933 255587
rect 291051 255469 293631 255587
rect 293749 255469 293791 255587
rect 293909 255469 294405 255587
rect -2443 255427 294405 255469
rect -2443 255309 -1947 255427
rect -1829 255309 -1787 255427
rect -1669 255309 2773 255427
rect 2891 255309 2933 255427
rect 3051 255309 20773 255427
rect 20891 255309 20933 255427
rect 21051 255309 38773 255427
rect 38891 255309 38933 255427
rect 39051 255309 56773 255427
rect 56891 255309 56933 255427
rect 57051 255309 74773 255427
rect 74891 255309 74933 255427
rect 75051 255309 92773 255427
rect 92891 255309 92933 255427
rect 93051 255309 110773 255427
rect 110891 255309 110933 255427
rect 111051 255309 128773 255427
rect 128891 255309 128933 255427
rect 129051 255309 146773 255427
rect 146891 255309 146933 255427
rect 147051 255309 164773 255427
rect 164891 255309 164933 255427
rect 165051 255309 182773 255427
rect 182891 255309 182933 255427
rect 183051 255309 200773 255427
rect 200891 255309 200933 255427
rect 201051 255309 218773 255427
rect 218891 255309 218933 255427
rect 219051 255309 236773 255427
rect 236891 255309 236933 255427
rect 237051 255309 254773 255427
rect 254891 255309 254933 255427
rect 255051 255309 272773 255427
rect 272891 255309 272933 255427
rect 273051 255309 290773 255427
rect 290891 255309 290933 255427
rect 291051 255309 293631 255427
rect 293749 255309 293791 255427
rect 293909 255309 294405 255427
rect -2443 255293 294405 255309
rect -1483 253727 293445 253743
rect -1483 253609 -987 253727
rect -869 253609 -827 253727
rect -709 253609 913 253727
rect 1031 253609 1073 253727
rect 1191 253609 18913 253727
rect 19031 253609 19073 253727
rect 19191 253609 36913 253727
rect 37031 253609 37073 253727
rect 37191 253609 54913 253727
rect 55031 253609 55073 253727
rect 55191 253609 72913 253727
rect 73031 253609 73073 253727
rect 73191 253609 90913 253727
rect 91031 253609 91073 253727
rect 91191 253609 108913 253727
rect 109031 253609 109073 253727
rect 109191 253609 126913 253727
rect 127031 253609 127073 253727
rect 127191 253609 144913 253727
rect 145031 253609 145073 253727
rect 145191 253609 162913 253727
rect 163031 253609 163073 253727
rect 163191 253609 180913 253727
rect 181031 253609 181073 253727
rect 181191 253609 198913 253727
rect 199031 253609 199073 253727
rect 199191 253609 216913 253727
rect 217031 253609 217073 253727
rect 217191 253609 234913 253727
rect 235031 253609 235073 253727
rect 235191 253609 252913 253727
rect 253031 253609 253073 253727
rect 253191 253609 270913 253727
rect 271031 253609 271073 253727
rect 271191 253609 288913 253727
rect 289031 253609 289073 253727
rect 289191 253609 292671 253727
rect 292789 253609 292831 253727
rect 292949 253609 293445 253727
rect -1483 253567 293445 253609
rect -1483 253449 -987 253567
rect -869 253449 -827 253567
rect -709 253449 913 253567
rect 1031 253449 1073 253567
rect 1191 253449 18913 253567
rect 19031 253449 19073 253567
rect 19191 253449 36913 253567
rect 37031 253449 37073 253567
rect 37191 253449 54913 253567
rect 55031 253449 55073 253567
rect 55191 253449 72913 253567
rect 73031 253449 73073 253567
rect 73191 253449 90913 253567
rect 91031 253449 91073 253567
rect 91191 253449 108913 253567
rect 109031 253449 109073 253567
rect 109191 253449 126913 253567
rect 127031 253449 127073 253567
rect 127191 253449 144913 253567
rect 145031 253449 145073 253567
rect 145191 253449 162913 253567
rect 163031 253449 163073 253567
rect 163191 253449 180913 253567
rect 181031 253449 181073 253567
rect 181191 253449 198913 253567
rect 199031 253449 199073 253567
rect 199191 253449 216913 253567
rect 217031 253449 217073 253567
rect 217191 253449 234913 253567
rect 235031 253449 235073 253567
rect 235191 253449 252913 253567
rect 253031 253449 253073 253567
rect 253191 253449 270913 253567
rect 271031 253449 271073 253567
rect 271191 253449 288913 253567
rect 289031 253449 289073 253567
rect 289191 253449 292671 253567
rect 292789 253449 292831 253567
rect 292949 253449 293445 253567
rect -1483 253433 293445 253449
rect -4363 250307 296325 250323
rect -4363 250189 -4347 250307
rect -4229 250189 -4187 250307
rect -4069 250189 15493 250307
rect 15611 250189 15653 250307
rect 15771 250189 33493 250307
rect 33611 250189 33653 250307
rect 33771 250189 51493 250307
rect 51611 250189 51653 250307
rect 51771 250189 69493 250307
rect 69611 250189 69653 250307
rect 69771 250189 87493 250307
rect 87611 250189 87653 250307
rect 87771 250189 105493 250307
rect 105611 250189 105653 250307
rect 105771 250189 123493 250307
rect 123611 250189 123653 250307
rect 123771 250189 141493 250307
rect 141611 250189 141653 250307
rect 141771 250189 159493 250307
rect 159611 250189 159653 250307
rect 159771 250189 177493 250307
rect 177611 250189 177653 250307
rect 177771 250189 195493 250307
rect 195611 250189 195653 250307
rect 195771 250189 213493 250307
rect 213611 250189 213653 250307
rect 213771 250189 231493 250307
rect 231611 250189 231653 250307
rect 231771 250189 249493 250307
rect 249611 250189 249653 250307
rect 249771 250189 267493 250307
rect 267611 250189 267653 250307
rect 267771 250189 285493 250307
rect 285611 250189 285653 250307
rect 285771 250189 296031 250307
rect 296149 250189 296191 250307
rect 296309 250189 296325 250307
rect -4363 250147 296325 250189
rect -4363 250029 -4347 250147
rect -4229 250029 -4187 250147
rect -4069 250029 15493 250147
rect 15611 250029 15653 250147
rect 15771 250029 33493 250147
rect 33611 250029 33653 250147
rect 33771 250029 51493 250147
rect 51611 250029 51653 250147
rect 51771 250029 69493 250147
rect 69611 250029 69653 250147
rect 69771 250029 87493 250147
rect 87611 250029 87653 250147
rect 87771 250029 105493 250147
rect 105611 250029 105653 250147
rect 105771 250029 123493 250147
rect 123611 250029 123653 250147
rect 123771 250029 141493 250147
rect 141611 250029 141653 250147
rect 141771 250029 159493 250147
rect 159611 250029 159653 250147
rect 159771 250029 177493 250147
rect 177611 250029 177653 250147
rect 177771 250029 195493 250147
rect 195611 250029 195653 250147
rect 195771 250029 213493 250147
rect 213611 250029 213653 250147
rect 213771 250029 231493 250147
rect 231611 250029 231653 250147
rect 231771 250029 249493 250147
rect 249611 250029 249653 250147
rect 249771 250029 267493 250147
rect 267611 250029 267653 250147
rect 267771 250029 285493 250147
rect 285611 250029 285653 250147
rect 285771 250029 296031 250147
rect 296149 250029 296191 250147
rect 296309 250029 296325 250147
rect -4363 250013 296325 250029
rect -3403 248447 295365 248463
rect -3403 248329 -3387 248447
rect -3269 248329 -3227 248447
rect -3109 248329 13633 248447
rect 13751 248329 13793 248447
rect 13911 248329 31633 248447
rect 31751 248329 31793 248447
rect 31911 248329 49633 248447
rect 49751 248329 49793 248447
rect 49911 248329 67633 248447
rect 67751 248329 67793 248447
rect 67911 248329 85633 248447
rect 85751 248329 85793 248447
rect 85911 248329 103633 248447
rect 103751 248329 103793 248447
rect 103911 248329 121633 248447
rect 121751 248329 121793 248447
rect 121911 248329 139633 248447
rect 139751 248329 139793 248447
rect 139911 248329 157633 248447
rect 157751 248329 157793 248447
rect 157911 248329 175633 248447
rect 175751 248329 175793 248447
rect 175911 248329 193633 248447
rect 193751 248329 193793 248447
rect 193911 248329 211633 248447
rect 211751 248329 211793 248447
rect 211911 248329 229633 248447
rect 229751 248329 229793 248447
rect 229911 248329 247633 248447
rect 247751 248329 247793 248447
rect 247911 248329 265633 248447
rect 265751 248329 265793 248447
rect 265911 248329 283633 248447
rect 283751 248329 283793 248447
rect 283911 248329 295071 248447
rect 295189 248329 295231 248447
rect 295349 248329 295365 248447
rect -3403 248287 295365 248329
rect -3403 248169 -3387 248287
rect -3269 248169 -3227 248287
rect -3109 248169 13633 248287
rect 13751 248169 13793 248287
rect 13911 248169 31633 248287
rect 31751 248169 31793 248287
rect 31911 248169 49633 248287
rect 49751 248169 49793 248287
rect 49911 248169 67633 248287
rect 67751 248169 67793 248287
rect 67911 248169 85633 248287
rect 85751 248169 85793 248287
rect 85911 248169 103633 248287
rect 103751 248169 103793 248287
rect 103911 248169 121633 248287
rect 121751 248169 121793 248287
rect 121911 248169 139633 248287
rect 139751 248169 139793 248287
rect 139911 248169 157633 248287
rect 157751 248169 157793 248287
rect 157911 248169 175633 248287
rect 175751 248169 175793 248287
rect 175911 248169 193633 248287
rect 193751 248169 193793 248287
rect 193911 248169 211633 248287
rect 211751 248169 211793 248287
rect 211911 248169 229633 248287
rect 229751 248169 229793 248287
rect 229911 248169 247633 248287
rect 247751 248169 247793 248287
rect 247911 248169 265633 248287
rect 265751 248169 265793 248287
rect 265911 248169 283633 248287
rect 283751 248169 283793 248287
rect 283911 248169 295071 248287
rect 295189 248169 295231 248287
rect 295349 248169 295365 248287
rect -3403 248153 295365 248169
rect -2443 246587 294405 246603
rect -2443 246469 -2427 246587
rect -2309 246469 -2267 246587
rect -2149 246469 11773 246587
rect 11891 246469 11933 246587
rect 12051 246469 29773 246587
rect 29891 246469 29933 246587
rect 30051 246469 47773 246587
rect 47891 246469 47933 246587
rect 48051 246469 65773 246587
rect 65891 246469 65933 246587
rect 66051 246469 83773 246587
rect 83891 246469 83933 246587
rect 84051 246469 101773 246587
rect 101891 246469 101933 246587
rect 102051 246469 119773 246587
rect 119891 246469 119933 246587
rect 120051 246469 137773 246587
rect 137891 246469 137933 246587
rect 138051 246469 155773 246587
rect 155891 246469 155933 246587
rect 156051 246469 173773 246587
rect 173891 246469 173933 246587
rect 174051 246469 191773 246587
rect 191891 246469 191933 246587
rect 192051 246469 209773 246587
rect 209891 246469 209933 246587
rect 210051 246469 227773 246587
rect 227891 246469 227933 246587
rect 228051 246469 245773 246587
rect 245891 246469 245933 246587
rect 246051 246469 263773 246587
rect 263891 246469 263933 246587
rect 264051 246469 281773 246587
rect 281891 246469 281933 246587
rect 282051 246469 294111 246587
rect 294229 246469 294271 246587
rect 294389 246469 294405 246587
rect -2443 246427 294405 246469
rect -2443 246309 -2427 246427
rect -2309 246309 -2267 246427
rect -2149 246309 11773 246427
rect 11891 246309 11933 246427
rect 12051 246309 29773 246427
rect 29891 246309 29933 246427
rect 30051 246309 47773 246427
rect 47891 246309 47933 246427
rect 48051 246309 65773 246427
rect 65891 246309 65933 246427
rect 66051 246309 83773 246427
rect 83891 246309 83933 246427
rect 84051 246309 101773 246427
rect 101891 246309 101933 246427
rect 102051 246309 119773 246427
rect 119891 246309 119933 246427
rect 120051 246309 137773 246427
rect 137891 246309 137933 246427
rect 138051 246309 155773 246427
rect 155891 246309 155933 246427
rect 156051 246309 173773 246427
rect 173891 246309 173933 246427
rect 174051 246309 191773 246427
rect 191891 246309 191933 246427
rect 192051 246309 209773 246427
rect 209891 246309 209933 246427
rect 210051 246309 227773 246427
rect 227891 246309 227933 246427
rect 228051 246309 245773 246427
rect 245891 246309 245933 246427
rect 246051 246309 263773 246427
rect 263891 246309 263933 246427
rect 264051 246309 281773 246427
rect 281891 246309 281933 246427
rect 282051 246309 294111 246427
rect 294229 246309 294271 246427
rect 294389 246309 294405 246427
rect -2443 246293 294405 246309
rect -1483 244727 293445 244743
rect -1483 244609 -1467 244727
rect -1349 244609 -1307 244727
rect -1189 244609 9913 244727
rect 10031 244609 10073 244727
rect 10191 244609 27913 244727
rect 28031 244609 28073 244727
rect 28191 244609 45913 244727
rect 46031 244609 46073 244727
rect 46191 244609 63913 244727
rect 64031 244609 64073 244727
rect 64191 244609 81913 244727
rect 82031 244609 82073 244727
rect 82191 244609 99913 244727
rect 100031 244609 100073 244727
rect 100191 244609 117913 244727
rect 118031 244609 118073 244727
rect 118191 244609 135913 244727
rect 136031 244609 136073 244727
rect 136191 244609 153913 244727
rect 154031 244609 154073 244727
rect 154191 244609 171913 244727
rect 172031 244609 172073 244727
rect 172191 244609 189913 244727
rect 190031 244609 190073 244727
rect 190191 244609 207913 244727
rect 208031 244609 208073 244727
rect 208191 244609 225913 244727
rect 226031 244609 226073 244727
rect 226191 244609 243913 244727
rect 244031 244609 244073 244727
rect 244191 244609 261913 244727
rect 262031 244609 262073 244727
rect 262191 244609 279913 244727
rect 280031 244609 280073 244727
rect 280191 244609 293151 244727
rect 293269 244609 293311 244727
rect 293429 244609 293445 244727
rect -1483 244567 293445 244609
rect -1483 244449 -1467 244567
rect -1349 244449 -1307 244567
rect -1189 244449 9913 244567
rect 10031 244449 10073 244567
rect 10191 244449 27913 244567
rect 28031 244449 28073 244567
rect 28191 244449 45913 244567
rect 46031 244449 46073 244567
rect 46191 244449 63913 244567
rect 64031 244449 64073 244567
rect 64191 244449 81913 244567
rect 82031 244449 82073 244567
rect 82191 244449 99913 244567
rect 100031 244449 100073 244567
rect 100191 244449 117913 244567
rect 118031 244449 118073 244567
rect 118191 244449 135913 244567
rect 136031 244449 136073 244567
rect 136191 244449 153913 244567
rect 154031 244449 154073 244567
rect 154191 244449 171913 244567
rect 172031 244449 172073 244567
rect 172191 244449 189913 244567
rect 190031 244449 190073 244567
rect 190191 244449 207913 244567
rect 208031 244449 208073 244567
rect 208191 244449 225913 244567
rect 226031 244449 226073 244567
rect 226191 244449 243913 244567
rect 244031 244449 244073 244567
rect 244191 244449 261913 244567
rect 262031 244449 262073 244567
rect 262191 244449 279913 244567
rect 280031 244449 280073 244567
rect 280191 244449 293151 244567
rect 293269 244449 293311 244567
rect 293429 244449 293445 244567
rect -1483 244433 293445 244449
rect -4363 241307 296325 241323
rect -4363 241189 -3867 241307
rect -3749 241189 -3707 241307
rect -3589 241189 6493 241307
rect 6611 241189 6653 241307
rect 6771 241189 24493 241307
rect 24611 241189 24653 241307
rect 24771 241189 42493 241307
rect 42611 241189 42653 241307
rect 42771 241189 60493 241307
rect 60611 241189 60653 241307
rect 60771 241189 78493 241307
rect 78611 241189 78653 241307
rect 78771 241189 96493 241307
rect 96611 241189 96653 241307
rect 96771 241189 114493 241307
rect 114611 241189 114653 241307
rect 114771 241189 132493 241307
rect 132611 241189 132653 241307
rect 132771 241189 150493 241307
rect 150611 241189 150653 241307
rect 150771 241189 168493 241307
rect 168611 241189 168653 241307
rect 168771 241189 186493 241307
rect 186611 241189 186653 241307
rect 186771 241189 204493 241307
rect 204611 241189 204653 241307
rect 204771 241189 222493 241307
rect 222611 241189 222653 241307
rect 222771 241189 240493 241307
rect 240611 241189 240653 241307
rect 240771 241189 258493 241307
rect 258611 241189 258653 241307
rect 258771 241189 276493 241307
rect 276611 241189 276653 241307
rect 276771 241189 295551 241307
rect 295669 241189 295711 241307
rect 295829 241189 296325 241307
rect -4363 241147 296325 241189
rect -4363 241029 -3867 241147
rect -3749 241029 -3707 241147
rect -3589 241029 6493 241147
rect 6611 241029 6653 241147
rect 6771 241029 24493 241147
rect 24611 241029 24653 241147
rect 24771 241029 42493 241147
rect 42611 241029 42653 241147
rect 42771 241029 60493 241147
rect 60611 241029 60653 241147
rect 60771 241029 78493 241147
rect 78611 241029 78653 241147
rect 78771 241029 96493 241147
rect 96611 241029 96653 241147
rect 96771 241029 114493 241147
rect 114611 241029 114653 241147
rect 114771 241029 132493 241147
rect 132611 241029 132653 241147
rect 132771 241029 150493 241147
rect 150611 241029 150653 241147
rect 150771 241029 168493 241147
rect 168611 241029 168653 241147
rect 168771 241029 186493 241147
rect 186611 241029 186653 241147
rect 186771 241029 204493 241147
rect 204611 241029 204653 241147
rect 204771 241029 222493 241147
rect 222611 241029 222653 241147
rect 222771 241029 240493 241147
rect 240611 241029 240653 241147
rect 240771 241029 258493 241147
rect 258611 241029 258653 241147
rect 258771 241029 276493 241147
rect 276611 241029 276653 241147
rect 276771 241029 295551 241147
rect 295669 241029 295711 241147
rect 295829 241029 296325 241147
rect -4363 241013 296325 241029
rect -3403 239447 295365 239463
rect -3403 239329 -2907 239447
rect -2789 239329 -2747 239447
rect -2629 239329 4633 239447
rect 4751 239329 4793 239447
rect 4911 239329 22633 239447
rect 22751 239329 22793 239447
rect 22911 239329 40633 239447
rect 40751 239329 40793 239447
rect 40911 239329 58633 239447
rect 58751 239329 58793 239447
rect 58911 239329 76633 239447
rect 76751 239329 76793 239447
rect 76911 239329 94633 239447
rect 94751 239329 94793 239447
rect 94911 239329 112633 239447
rect 112751 239329 112793 239447
rect 112911 239329 130633 239447
rect 130751 239329 130793 239447
rect 130911 239329 148633 239447
rect 148751 239329 148793 239447
rect 148911 239329 166633 239447
rect 166751 239329 166793 239447
rect 166911 239329 184633 239447
rect 184751 239329 184793 239447
rect 184911 239329 202633 239447
rect 202751 239329 202793 239447
rect 202911 239329 220633 239447
rect 220751 239329 220793 239447
rect 220911 239329 238633 239447
rect 238751 239329 238793 239447
rect 238911 239329 256633 239447
rect 256751 239329 256793 239447
rect 256911 239329 274633 239447
rect 274751 239329 274793 239447
rect 274911 239329 294591 239447
rect 294709 239329 294751 239447
rect 294869 239329 295365 239447
rect -3403 239287 295365 239329
rect -3403 239169 -2907 239287
rect -2789 239169 -2747 239287
rect -2629 239169 4633 239287
rect 4751 239169 4793 239287
rect 4911 239169 22633 239287
rect 22751 239169 22793 239287
rect 22911 239169 40633 239287
rect 40751 239169 40793 239287
rect 40911 239169 58633 239287
rect 58751 239169 58793 239287
rect 58911 239169 76633 239287
rect 76751 239169 76793 239287
rect 76911 239169 94633 239287
rect 94751 239169 94793 239287
rect 94911 239169 112633 239287
rect 112751 239169 112793 239287
rect 112911 239169 130633 239287
rect 130751 239169 130793 239287
rect 130911 239169 148633 239287
rect 148751 239169 148793 239287
rect 148911 239169 166633 239287
rect 166751 239169 166793 239287
rect 166911 239169 184633 239287
rect 184751 239169 184793 239287
rect 184911 239169 202633 239287
rect 202751 239169 202793 239287
rect 202911 239169 220633 239287
rect 220751 239169 220793 239287
rect 220911 239169 238633 239287
rect 238751 239169 238793 239287
rect 238911 239169 256633 239287
rect 256751 239169 256793 239287
rect 256911 239169 274633 239287
rect 274751 239169 274793 239287
rect 274911 239169 294591 239287
rect 294709 239169 294751 239287
rect 294869 239169 295365 239287
rect -3403 239153 295365 239169
rect -2443 237587 294405 237603
rect -2443 237469 -1947 237587
rect -1829 237469 -1787 237587
rect -1669 237469 2773 237587
rect 2891 237469 2933 237587
rect 3051 237469 20773 237587
rect 20891 237469 20933 237587
rect 21051 237469 38773 237587
rect 38891 237469 38933 237587
rect 39051 237469 56773 237587
rect 56891 237469 56933 237587
rect 57051 237469 74773 237587
rect 74891 237469 74933 237587
rect 75051 237469 92773 237587
rect 92891 237469 92933 237587
rect 93051 237469 110773 237587
rect 110891 237469 110933 237587
rect 111051 237469 128773 237587
rect 128891 237469 128933 237587
rect 129051 237469 146773 237587
rect 146891 237469 146933 237587
rect 147051 237469 164773 237587
rect 164891 237469 164933 237587
rect 165051 237469 182773 237587
rect 182891 237469 182933 237587
rect 183051 237469 200773 237587
rect 200891 237469 200933 237587
rect 201051 237469 218773 237587
rect 218891 237469 218933 237587
rect 219051 237469 236773 237587
rect 236891 237469 236933 237587
rect 237051 237469 254773 237587
rect 254891 237469 254933 237587
rect 255051 237469 272773 237587
rect 272891 237469 272933 237587
rect 273051 237469 290773 237587
rect 290891 237469 290933 237587
rect 291051 237469 293631 237587
rect 293749 237469 293791 237587
rect 293909 237469 294405 237587
rect -2443 237427 294405 237469
rect -2443 237309 -1947 237427
rect -1829 237309 -1787 237427
rect -1669 237309 2773 237427
rect 2891 237309 2933 237427
rect 3051 237309 20773 237427
rect 20891 237309 20933 237427
rect 21051 237309 38773 237427
rect 38891 237309 38933 237427
rect 39051 237309 56773 237427
rect 56891 237309 56933 237427
rect 57051 237309 74773 237427
rect 74891 237309 74933 237427
rect 75051 237309 92773 237427
rect 92891 237309 92933 237427
rect 93051 237309 110773 237427
rect 110891 237309 110933 237427
rect 111051 237309 128773 237427
rect 128891 237309 128933 237427
rect 129051 237309 146773 237427
rect 146891 237309 146933 237427
rect 147051 237309 164773 237427
rect 164891 237309 164933 237427
rect 165051 237309 182773 237427
rect 182891 237309 182933 237427
rect 183051 237309 200773 237427
rect 200891 237309 200933 237427
rect 201051 237309 218773 237427
rect 218891 237309 218933 237427
rect 219051 237309 236773 237427
rect 236891 237309 236933 237427
rect 237051 237309 254773 237427
rect 254891 237309 254933 237427
rect 255051 237309 272773 237427
rect 272891 237309 272933 237427
rect 273051 237309 290773 237427
rect 290891 237309 290933 237427
rect 291051 237309 293631 237427
rect 293749 237309 293791 237427
rect 293909 237309 294405 237427
rect -2443 237293 294405 237309
rect -1483 235727 293445 235743
rect -1483 235609 -987 235727
rect -869 235609 -827 235727
rect -709 235609 913 235727
rect 1031 235609 1073 235727
rect 1191 235609 18913 235727
rect 19031 235609 19073 235727
rect 19191 235609 36913 235727
rect 37031 235609 37073 235727
rect 37191 235609 54913 235727
rect 55031 235609 55073 235727
rect 55191 235609 72913 235727
rect 73031 235609 73073 235727
rect 73191 235609 90913 235727
rect 91031 235609 91073 235727
rect 91191 235609 108913 235727
rect 109031 235609 109073 235727
rect 109191 235609 126913 235727
rect 127031 235609 127073 235727
rect 127191 235609 144913 235727
rect 145031 235609 145073 235727
rect 145191 235609 162913 235727
rect 163031 235609 163073 235727
rect 163191 235609 180913 235727
rect 181031 235609 181073 235727
rect 181191 235609 198913 235727
rect 199031 235609 199073 235727
rect 199191 235609 216913 235727
rect 217031 235609 217073 235727
rect 217191 235609 234913 235727
rect 235031 235609 235073 235727
rect 235191 235609 252913 235727
rect 253031 235609 253073 235727
rect 253191 235609 270913 235727
rect 271031 235609 271073 235727
rect 271191 235609 288913 235727
rect 289031 235609 289073 235727
rect 289191 235609 292671 235727
rect 292789 235609 292831 235727
rect 292949 235609 293445 235727
rect -1483 235567 293445 235609
rect -1483 235449 -987 235567
rect -869 235449 -827 235567
rect -709 235449 913 235567
rect 1031 235449 1073 235567
rect 1191 235449 18913 235567
rect 19031 235449 19073 235567
rect 19191 235449 36913 235567
rect 37031 235449 37073 235567
rect 37191 235449 54913 235567
rect 55031 235449 55073 235567
rect 55191 235449 72913 235567
rect 73031 235449 73073 235567
rect 73191 235449 90913 235567
rect 91031 235449 91073 235567
rect 91191 235449 108913 235567
rect 109031 235449 109073 235567
rect 109191 235449 126913 235567
rect 127031 235449 127073 235567
rect 127191 235449 144913 235567
rect 145031 235449 145073 235567
rect 145191 235449 162913 235567
rect 163031 235449 163073 235567
rect 163191 235449 180913 235567
rect 181031 235449 181073 235567
rect 181191 235449 198913 235567
rect 199031 235449 199073 235567
rect 199191 235449 216913 235567
rect 217031 235449 217073 235567
rect 217191 235449 234913 235567
rect 235031 235449 235073 235567
rect 235191 235449 252913 235567
rect 253031 235449 253073 235567
rect 253191 235449 270913 235567
rect 271031 235449 271073 235567
rect 271191 235449 288913 235567
rect 289031 235449 289073 235567
rect 289191 235449 292671 235567
rect 292789 235449 292831 235567
rect 292949 235449 293445 235567
rect -1483 235433 293445 235449
rect -4363 232307 296325 232323
rect -4363 232189 -4347 232307
rect -4229 232189 -4187 232307
rect -4069 232189 15493 232307
rect 15611 232189 15653 232307
rect 15771 232189 33493 232307
rect 33611 232189 33653 232307
rect 33771 232189 51493 232307
rect 51611 232189 51653 232307
rect 51771 232189 69493 232307
rect 69611 232189 69653 232307
rect 69771 232189 87493 232307
rect 87611 232189 87653 232307
rect 87771 232189 105493 232307
rect 105611 232189 105653 232307
rect 105771 232189 123493 232307
rect 123611 232189 123653 232307
rect 123771 232189 141493 232307
rect 141611 232189 141653 232307
rect 141771 232189 159493 232307
rect 159611 232189 159653 232307
rect 159771 232189 177493 232307
rect 177611 232189 177653 232307
rect 177771 232189 195493 232307
rect 195611 232189 195653 232307
rect 195771 232189 213493 232307
rect 213611 232189 213653 232307
rect 213771 232189 231493 232307
rect 231611 232189 231653 232307
rect 231771 232189 249493 232307
rect 249611 232189 249653 232307
rect 249771 232189 267493 232307
rect 267611 232189 267653 232307
rect 267771 232189 285493 232307
rect 285611 232189 285653 232307
rect 285771 232189 296031 232307
rect 296149 232189 296191 232307
rect 296309 232189 296325 232307
rect -4363 232147 296325 232189
rect -4363 232029 -4347 232147
rect -4229 232029 -4187 232147
rect -4069 232029 15493 232147
rect 15611 232029 15653 232147
rect 15771 232029 33493 232147
rect 33611 232029 33653 232147
rect 33771 232029 51493 232147
rect 51611 232029 51653 232147
rect 51771 232029 69493 232147
rect 69611 232029 69653 232147
rect 69771 232029 87493 232147
rect 87611 232029 87653 232147
rect 87771 232029 105493 232147
rect 105611 232029 105653 232147
rect 105771 232029 123493 232147
rect 123611 232029 123653 232147
rect 123771 232029 141493 232147
rect 141611 232029 141653 232147
rect 141771 232029 159493 232147
rect 159611 232029 159653 232147
rect 159771 232029 177493 232147
rect 177611 232029 177653 232147
rect 177771 232029 195493 232147
rect 195611 232029 195653 232147
rect 195771 232029 213493 232147
rect 213611 232029 213653 232147
rect 213771 232029 231493 232147
rect 231611 232029 231653 232147
rect 231771 232029 249493 232147
rect 249611 232029 249653 232147
rect 249771 232029 267493 232147
rect 267611 232029 267653 232147
rect 267771 232029 285493 232147
rect 285611 232029 285653 232147
rect 285771 232029 296031 232147
rect 296149 232029 296191 232147
rect 296309 232029 296325 232147
rect -4363 232013 296325 232029
rect -3403 230447 295365 230463
rect -3403 230329 -3387 230447
rect -3269 230329 -3227 230447
rect -3109 230329 13633 230447
rect 13751 230329 13793 230447
rect 13911 230329 31633 230447
rect 31751 230329 31793 230447
rect 31911 230329 49633 230447
rect 49751 230329 49793 230447
rect 49911 230329 67633 230447
rect 67751 230329 67793 230447
rect 67911 230329 85633 230447
rect 85751 230329 85793 230447
rect 85911 230329 103633 230447
rect 103751 230329 103793 230447
rect 103911 230329 121633 230447
rect 121751 230329 121793 230447
rect 121911 230329 139633 230447
rect 139751 230329 139793 230447
rect 139911 230329 157633 230447
rect 157751 230329 157793 230447
rect 157911 230329 175633 230447
rect 175751 230329 175793 230447
rect 175911 230329 193633 230447
rect 193751 230329 193793 230447
rect 193911 230329 211633 230447
rect 211751 230329 211793 230447
rect 211911 230329 229633 230447
rect 229751 230329 229793 230447
rect 229911 230329 247633 230447
rect 247751 230329 247793 230447
rect 247911 230329 265633 230447
rect 265751 230329 265793 230447
rect 265911 230329 283633 230447
rect 283751 230329 283793 230447
rect 283911 230329 295071 230447
rect 295189 230329 295231 230447
rect 295349 230329 295365 230447
rect -3403 230287 295365 230329
rect -3403 230169 -3387 230287
rect -3269 230169 -3227 230287
rect -3109 230169 13633 230287
rect 13751 230169 13793 230287
rect 13911 230169 31633 230287
rect 31751 230169 31793 230287
rect 31911 230169 49633 230287
rect 49751 230169 49793 230287
rect 49911 230169 67633 230287
rect 67751 230169 67793 230287
rect 67911 230169 85633 230287
rect 85751 230169 85793 230287
rect 85911 230169 103633 230287
rect 103751 230169 103793 230287
rect 103911 230169 121633 230287
rect 121751 230169 121793 230287
rect 121911 230169 139633 230287
rect 139751 230169 139793 230287
rect 139911 230169 157633 230287
rect 157751 230169 157793 230287
rect 157911 230169 175633 230287
rect 175751 230169 175793 230287
rect 175911 230169 193633 230287
rect 193751 230169 193793 230287
rect 193911 230169 211633 230287
rect 211751 230169 211793 230287
rect 211911 230169 229633 230287
rect 229751 230169 229793 230287
rect 229911 230169 247633 230287
rect 247751 230169 247793 230287
rect 247911 230169 265633 230287
rect 265751 230169 265793 230287
rect 265911 230169 283633 230287
rect 283751 230169 283793 230287
rect 283911 230169 295071 230287
rect 295189 230169 295231 230287
rect 295349 230169 295365 230287
rect -3403 230153 295365 230169
rect -2443 228587 294405 228603
rect -2443 228469 -2427 228587
rect -2309 228469 -2267 228587
rect -2149 228469 11773 228587
rect 11891 228469 11933 228587
rect 12051 228469 29773 228587
rect 29891 228469 29933 228587
rect 30051 228469 47773 228587
rect 47891 228469 47933 228587
rect 48051 228469 65773 228587
rect 65891 228469 65933 228587
rect 66051 228469 83773 228587
rect 83891 228469 83933 228587
rect 84051 228469 101773 228587
rect 101891 228469 101933 228587
rect 102051 228469 119773 228587
rect 119891 228469 119933 228587
rect 120051 228469 137773 228587
rect 137891 228469 137933 228587
rect 138051 228469 155773 228587
rect 155891 228469 155933 228587
rect 156051 228469 173773 228587
rect 173891 228469 173933 228587
rect 174051 228469 191773 228587
rect 191891 228469 191933 228587
rect 192051 228469 209773 228587
rect 209891 228469 209933 228587
rect 210051 228469 227773 228587
rect 227891 228469 227933 228587
rect 228051 228469 245773 228587
rect 245891 228469 245933 228587
rect 246051 228469 263773 228587
rect 263891 228469 263933 228587
rect 264051 228469 281773 228587
rect 281891 228469 281933 228587
rect 282051 228469 294111 228587
rect 294229 228469 294271 228587
rect 294389 228469 294405 228587
rect -2443 228427 294405 228469
rect -2443 228309 -2427 228427
rect -2309 228309 -2267 228427
rect -2149 228309 11773 228427
rect 11891 228309 11933 228427
rect 12051 228309 29773 228427
rect 29891 228309 29933 228427
rect 30051 228309 47773 228427
rect 47891 228309 47933 228427
rect 48051 228309 65773 228427
rect 65891 228309 65933 228427
rect 66051 228309 83773 228427
rect 83891 228309 83933 228427
rect 84051 228309 101773 228427
rect 101891 228309 101933 228427
rect 102051 228309 119773 228427
rect 119891 228309 119933 228427
rect 120051 228309 137773 228427
rect 137891 228309 137933 228427
rect 138051 228309 155773 228427
rect 155891 228309 155933 228427
rect 156051 228309 173773 228427
rect 173891 228309 173933 228427
rect 174051 228309 191773 228427
rect 191891 228309 191933 228427
rect 192051 228309 209773 228427
rect 209891 228309 209933 228427
rect 210051 228309 227773 228427
rect 227891 228309 227933 228427
rect 228051 228309 245773 228427
rect 245891 228309 245933 228427
rect 246051 228309 263773 228427
rect 263891 228309 263933 228427
rect 264051 228309 281773 228427
rect 281891 228309 281933 228427
rect 282051 228309 294111 228427
rect 294229 228309 294271 228427
rect 294389 228309 294405 228427
rect -2443 228293 294405 228309
rect -1483 226727 293445 226743
rect -1483 226609 -1467 226727
rect -1349 226609 -1307 226727
rect -1189 226609 9913 226727
rect 10031 226609 10073 226727
rect 10191 226609 27913 226727
rect 28031 226609 28073 226727
rect 28191 226609 45913 226727
rect 46031 226609 46073 226727
rect 46191 226609 63913 226727
rect 64031 226609 64073 226727
rect 64191 226609 81913 226727
rect 82031 226609 82073 226727
rect 82191 226609 99913 226727
rect 100031 226609 100073 226727
rect 100191 226609 117913 226727
rect 118031 226609 118073 226727
rect 118191 226609 135913 226727
rect 136031 226609 136073 226727
rect 136191 226609 153913 226727
rect 154031 226609 154073 226727
rect 154191 226609 171913 226727
rect 172031 226609 172073 226727
rect 172191 226609 189913 226727
rect 190031 226609 190073 226727
rect 190191 226609 207913 226727
rect 208031 226609 208073 226727
rect 208191 226609 225913 226727
rect 226031 226609 226073 226727
rect 226191 226609 243913 226727
rect 244031 226609 244073 226727
rect 244191 226609 261913 226727
rect 262031 226609 262073 226727
rect 262191 226609 279913 226727
rect 280031 226609 280073 226727
rect 280191 226609 293151 226727
rect 293269 226609 293311 226727
rect 293429 226609 293445 226727
rect -1483 226567 293445 226609
rect -1483 226449 -1467 226567
rect -1349 226449 -1307 226567
rect -1189 226449 9913 226567
rect 10031 226449 10073 226567
rect 10191 226449 27913 226567
rect 28031 226449 28073 226567
rect 28191 226449 45913 226567
rect 46031 226449 46073 226567
rect 46191 226449 63913 226567
rect 64031 226449 64073 226567
rect 64191 226449 81913 226567
rect 82031 226449 82073 226567
rect 82191 226449 99913 226567
rect 100031 226449 100073 226567
rect 100191 226449 117913 226567
rect 118031 226449 118073 226567
rect 118191 226449 135913 226567
rect 136031 226449 136073 226567
rect 136191 226449 153913 226567
rect 154031 226449 154073 226567
rect 154191 226449 171913 226567
rect 172031 226449 172073 226567
rect 172191 226449 189913 226567
rect 190031 226449 190073 226567
rect 190191 226449 207913 226567
rect 208031 226449 208073 226567
rect 208191 226449 225913 226567
rect 226031 226449 226073 226567
rect 226191 226449 243913 226567
rect 244031 226449 244073 226567
rect 244191 226449 261913 226567
rect 262031 226449 262073 226567
rect 262191 226449 279913 226567
rect 280031 226449 280073 226567
rect 280191 226449 293151 226567
rect 293269 226449 293311 226567
rect 293429 226449 293445 226567
rect -1483 226433 293445 226449
rect -4363 223307 296325 223323
rect -4363 223189 -3867 223307
rect -3749 223189 -3707 223307
rect -3589 223189 6493 223307
rect 6611 223189 6653 223307
rect 6771 223189 24493 223307
rect 24611 223189 24653 223307
rect 24771 223189 42493 223307
rect 42611 223189 42653 223307
rect 42771 223189 60493 223307
rect 60611 223189 60653 223307
rect 60771 223189 78493 223307
rect 78611 223189 78653 223307
rect 78771 223189 96493 223307
rect 96611 223189 96653 223307
rect 96771 223189 114493 223307
rect 114611 223189 114653 223307
rect 114771 223189 132493 223307
rect 132611 223189 132653 223307
rect 132771 223189 150493 223307
rect 150611 223189 150653 223307
rect 150771 223189 168493 223307
rect 168611 223189 168653 223307
rect 168771 223189 186493 223307
rect 186611 223189 186653 223307
rect 186771 223189 204493 223307
rect 204611 223189 204653 223307
rect 204771 223189 222493 223307
rect 222611 223189 222653 223307
rect 222771 223189 240493 223307
rect 240611 223189 240653 223307
rect 240771 223189 258493 223307
rect 258611 223189 258653 223307
rect 258771 223189 276493 223307
rect 276611 223189 276653 223307
rect 276771 223189 295551 223307
rect 295669 223189 295711 223307
rect 295829 223189 296325 223307
rect -4363 223147 296325 223189
rect -4363 223029 -3867 223147
rect -3749 223029 -3707 223147
rect -3589 223029 6493 223147
rect 6611 223029 6653 223147
rect 6771 223029 24493 223147
rect 24611 223029 24653 223147
rect 24771 223029 42493 223147
rect 42611 223029 42653 223147
rect 42771 223029 60493 223147
rect 60611 223029 60653 223147
rect 60771 223029 78493 223147
rect 78611 223029 78653 223147
rect 78771 223029 96493 223147
rect 96611 223029 96653 223147
rect 96771 223029 114493 223147
rect 114611 223029 114653 223147
rect 114771 223029 132493 223147
rect 132611 223029 132653 223147
rect 132771 223029 150493 223147
rect 150611 223029 150653 223147
rect 150771 223029 168493 223147
rect 168611 223029 168653 223147
rect 168771 223029 186493 223147
rect 186611 223029 186653 223147
rect 186771 223029 204493 223147
rect 204611 223029 204653 223147
rect 204771 223029 222493 223147
rect 222611 223029 222653 223147
rect 222771 223029 240493 223147
rect 240611 223029 240653 223147
rect 240771 223029 258493 223147
rect 258611 223029 258653 223147
rect 258771 223029 276493 223147
rect 276611 223029 276653 223147
rect 276771 223029 295551 223147
rect 295669 223029 295711 223147
rect 295829 223029 296325 223147
rect -4363 223013 296325 223029
rect -3403 221447 295365 221463
rect -3403 221329 -2907 221447
rect -2789 221329 -2747 221447
rect -2629 221329 4633 221447
rect 4751 221329 4793 221447
rect 4911 221329 22633 221447
rect 22751 221329 22793 221447
rect 22911 221329 40633 221447
rect 40751 221329 40793 221447
rect 40911 221329 58633 221447
rect 58751 221329 58793 221447
rect 58911 221329 76633 221447
rect 76751 221329 76793 221447
rect 76911 221329 94633 221447
rect 94751 221329 94793 221447
rect 94911 221329 112633 221447
rect 112751 221329 112793 221447
rect 112911 221329 130633 221447
rect 130751 221329 130793 221447
rect 130911 221329 148633 221447
rect 148751 221329 148793 221447
rect 148911 221329 166633 221447
rect 166751 221329 166793 221447
rect 166911 221329 184633 221447
rect 184751 221329 184793 221447
rect 184911 221329 202633 221447
rect 202751 221329 202793 221447
rect 202911 221329 220633 221447
rect 220751 221329 220793 221447
rect 220911 221329 238633 221447
rect 238751 221329 238793 221447
rect 238911 221329 256633 221447
rect 256751 221329 256793 221447
rect 256911 221329 274633 221447
rect 274751 221329 274793 221447
rect 274911 221329 294591 221447
rect 294709 221329 294751 221447
rect 294869 221329 295365 221447
rect -3403 221287 295365 221329
rect -3403 221169 -2907 221287
rect -2789 221169 -2747 221287
rect -2629 221169 4633 221287
rect 4751 221169 4793 221287
rect 4911 221169 22633 221287
rect 22751 221169 22793 221287
rect 22911 221169 40633 221287
rect 40751 221169 40793 221287
rect 40911 221169 58633 221287
rect 58751 221169 58793 221287
rect 58911 221169 76633 221287
rect 76751 221169 76793 221287
rect 76911 221169 94633 221287
rect 94751 221169 94793 221287
rect 94911 221169 112633 221287
rect 112751 221169 112793 221287
rect 112911 221169 130633 221287
rect 130751 221169 130793 221287
rect 130911 221169 148633 221287
rect 148751 221169 148793 221287
rect 148911 221169 166633 221287
rect 166751 221169 166793 221287
rect 166911 221169 184633 221287
rect 184751 221169 184793 221287
rect 184911 221169 202633 221287
rect 202751 221169 202793 221287
rect 202911 221169 220633 221287
rect 220751 221169 220793 221287
rect 220911 221169 238633 221287
rect 238751 221169 238793 221287
rect 238911 221169 256633 221287
rect 256751 221169 256793 221287
rect 256911 221169 274633 221287
rect 274751 221169 274793 221287
rect 274911 221169 294591 221287
rect 294709 221169 294751 221287
rect 294869 221169 295365 221287
rect -3403 221153 295365 221169
rect -2443 219587 294405 219603
rect -2443 219469 -1947 219587
rect -1829 219469 -1787 219587
rect -1669 219469 2773 219587
rect 2891 219469 2933 219587
rect 3051 219469 20773 219587
rect 20891 219469 20933 219587
rect 21051 219469 38773 219587
rect 38891 219469 38933 219587
rect 39051 219469 56773 219587
rect 56891 219469 56933 219587
rect 57051 219469 74773 219587
rect 74891 219469 74933 219587
rect 75051 219469 92773 219587
rect 92891 219469 92933 219587
rect 93051 219469 110773 219587
rect 110891 219469 110933 219587
rect 111051 219469 128773 219587
rect 128891 219469 128933 219587
rect 129051 219469 146773 219587
rect 146891 219469 146933 219587
rect 147051 219469 164773 219587
rect 164891 219469 164933 219587
rect 165051 219469 182773 219587
rect 182891 219469 182933 219587
rect 183051 219469 200773 219587
rect 200891 219469 200933 219587
rect 201051 219469 218773 219587
rect 218891 219469 218933 219587
rect 219051 219469 236773 219587
rect 236891 219469 236933 219587
rect 237051 219469 254773 219587
rect 254891 219469 254933 219587
rect 255051 219469 272773 219587
rect 272891 219469 272933 219587
rect 273051 219469 290773 219587
rect 290891 219469 290933 219587
rect 291051 219469 293631 219587
rect 293749 219469 293791 219587
rect 293909 219469 294405 219587
rect -2443 219427 294405 219469
rect -2443 219309 -1947 219427
rect -1829 219309 -1787 219427
rect -1669 219309 2773 219427
rect 2891 219309 2933 219427
rect 3051 219309 20773 219427
rect 20891 219309 20933 219427
rect 21051 219309 38773 219427
rect 38891 219309 38933 219427
rect 39051 219309 56773 219427
rect 56891 219309 56933 219427
rect 57051 219309 74773 219427
rect 74891 219309 74933 219427
rect 75051 219309 92773 219427
rect 92891 219309 92933 219427
rect 93051 219309 110773 219427
rect 110891 219309 110933 219427
rect 111051 219309 128773 219427
rect 128891 219309 128933 219427
rect 129051 219309 146773 219427
rect 146891 219309 146933 219427
rect 147051 219309 164773 219427
rect 164891 219309 164933 219427
rect 165051 219309 182773 219427
rect 182891 219309 182933 219427
rect 183051 219309 200773 219427
rect 200891 219309 200933 219427
rect 201051 219309 218773 219427
rect 218891 219309 218933 219427
rect 219051 219309 236773 219427
rect 236891 219309 236933 219427
rect 237051 219309 254773 219427
rect 254891 219309 254933 219427
rect 255051 219309 272773 219427
rect 272891 219309 272933 219427
rect 273051 219309 290773 219427
rect 290891 219309 290933 219427
rect 291051 219309 293631 219427
rect 293749 219309 293791 219427
rect 293909 219309 294405 219427
rect -2443 219293 294405 219309
rect -1483 217727 293445 217743
rect -1483 217609 -987 217727
rect -869 217609 -827 217727
rect -709 217609 913 217727
rect 1031 217609 1073 217727
rect 1191 217609 18913 217727
rect 19031 217609 19073 217727
rect 19191 217609 36913 217727
rect 37031 217609 37073 217727
rect 37191 217609 54913 217727
rect 55031 217609 55073 217727
rect 55191 217609 72913 217727
rect 73031 217609 73073 217727
rect 73191 217609 90913 217727
rect 91031 217609 91073 217727
rect 91191 217609 108913 217727
rect 109031 217609 109073 217727
rect 109191 217609 126913 217727
rect 127031 217609 127073 217727
rect 127191 217609 144913 217727
rect 145031 217609 145073 217727
rect 145191 217609 162913 217727
rect 163031 217609 163073 217727
rect 163191 217609 180913 217727
rect 181031 217609 181073 217727
rect 181191 217609 198913 217727
rect 199031 217609 199073 217727
rect 199191 217609 216913 217727
rect 217031 217609 217073 217727
rect 217191 217609 234913 217727
rect 235031 217609 235073 217727
rect 235191 217609 252913 217727
rect 253031 217609 253073 217727
rect 253191 217609 270913 217727
rect 271031 217609 271073 217727
rect 271191 217609 288913 217727
rect 289031 217609 289073 217727
rect 289191 217609 292671 217727
rect 292789 217609 292831 217727
rect 292949 217609 293445 217727
rect -1483 217567 293445 217609
rect -1483 217449 -987 217567
rect -869 217449 -827 217567
rect -709 217449 913 217567
rect 1031 217449 1073 217567
rect 1191 217449 18913 217567
rect 19031 217449 19073 217567
rect 19191 217449 36913 217567
rect 37031 217449 37073 217567
rect 37191 217449 54913 217567
rect 55031 217449 55073 217567
rect 55191 217449 72913 217567
rect 73031 217449 73073 217567
rect 73191 217449 90913 217567
rect 91031 217449 91073 217567
rect 91191 217449 108913 217567
rect 109031 217449 109073 217567
rect 109191 217449 126913 217567
rect 127031 217449 127073 217567
rect 127191 217449 144913 217567
rect 145031 217449 145073 217567
rect 145191 217449 162913 217567
rect 163031 217449 163073 217567
rect 163191 217449 180913 217567
rect 181031 217449 181073 217567
rect 181191 217449 198913 217567
rect 199031 217449 199073 217567
rect 199191 217449 216913 217567
rect 217031 217449 217073 217567
rect 217191 217449 234913 217567
rect 235031 217449 235073 217567
rect 235191 217449 252913 217567
rect 253031 217449 253073 217567
rect 253191 217449 270913 217567
rect 271031 217449 271073 217567
rect 271191 217449 288913 217567
rect 289031 217449 289073 217567
rect 289191 217449 292671 217567
rect 292789 217449 292831 217567
rect 292949 217449 293445 217567
rect -1483 217433 293445 217449
rect -4363 214307 296325 214323
rect -4363 214189 -4347 214307
rect -4229 214189 -4187 214307
rect -4069 214189 15493 214307
rect 15611 214189 15653 214307
rect 15771 214189 33493 214307
rect 33611 214189 33653 214307
rect 33771 214189 51493 214307
rect 51611 214189 51653 214307
rect 51771 214189 69493 214307
rect 69611 214189 69653 214307
rect 69771 214189 87493 214307
rect 87611 214189 87653 214307
rect 87771 214189 105493 214307
rect 105611 214189 105653 214307
rect 105771 214189 123493 214307
rect 123611 214189 123653 214307
rect 123771 214189 141493 214307
rect 141611 214189 141653 214307
rect 141771 214189 159493 214307
rect 159611 214189 159653 214307
rect 159771 214189 177493 214307
rect 177611 214189 177653 214307
rect 177771 214189 195493 214307
rect 195611 214189 195653 214307
rect 195771 214189 213493 214307
rect 213611 214189 213653 214307
rect 213771 214189 231493 214307
rect 231611 214189 231653 214307
rect 231771 214189 249493 214307
rect 249611 214189 249653 214307
rect 249771 214189 267493 214307
rect 267611 214189 267653 214307
rect 267771 214189 285493 214307
rect 285611 214189 285653 214307
rect 285771 214189 296031 214307
rect 296149 214189 296191 214307
rect 296309 214189 296325 214307
rect -4363 214147 296325 214189
rect -4363 214029 -4347 214147
rect -4229 214029 -4187 214147
rect -4069 214029 15493 214147
rect 15611 214029 15653 214147
rect 15771 214029 33493 214147
rect 33611 214029 33653 214147
rect 33771 214029 51493 214147
rect 51611 214029 51653 214147
rect 51771 214029 69493 214147
rect 69611 214029 69653 214147
rect 69771 214029 87493 214147
rect 87611 214029 87653 214147
rect 87771 214029 105493 214147
rect 105611 214029 105653 214147
rect 105771 214029 123493 214147
rect 123611 214029 123653 214147
rect 123771 214029 141493 214147
rect 141611 214029 141653 214147
rect 141771 214029 159493 214147
rect 159611 214029 159653 214147
rect 159771 214029 177493 214147
rect 177611 214029 177653 214147
rect 177771 214029 195493 214147
rect 195611 214029 195653 214147
rect 195771 214029 213493 214147
rect 213611 214029 213653 214147
rect 213771 214029 231493 214147
rect 231611 214029 231653 214147
rect 231771 214029 249493 214147
rect 249611 214029 249653 214147
rect 249771 214029 267493 214147
rect 267611 214029 267653 214147
rect 267771 214029 285493 214147
rect 285611 214029 285653 214147
rect 285771 214029 296031 214147
rect 296149 214029 296191 214147
rect 296309 214029 296325 214147
rect -4363 214013 296325 214029
rect -3403 212447 295365 212463
rect -3403 212329 -3387 212447
rect -3269 212329 -3227 212447
rect -3109 212329 13633 212447
rect 13751 212329 13793 212447
rect 13911 212329 31633 212447
rect 31751 212329 31793 212447
rect 31911 212329 49633 212447
rect 49751 212329 49793 212447
rect 49911 212329 67633 212447
rect 67751 212329 67793 212447
rect 67911 212329 85633 212447
rect 85751 212329 85793 212447
rect 85911 212329 103633 212447
rect 103751 212329 103793 212447
rect 103911 212329 121633 212447
rect 121751 212329 121793 212447
rect 121911 212329 139633 212447
rect 139751 212329 139793 212447
rect 139911 212329 157633 212447
rect 157751 212329 157793 212447
rect 157911 212329 175633 212447
rect 175751 212329 175793 212447
rect 175911 212329 193633 212447
rect 193751 212329 193793 212447
rect 193911 212329 211633 212447
rect 211751 212329 211793 212447
rect 211911 212329 229633 212447
rect 229751 212329 229793 212447
rect 229911 212329 247633 212447
rect 247751 212329 247793 212447
rect 247911 212329 265633 212447
rect 265751 212329 265793 212447
rect 265911 212329 283633 212447
rect 283751 212329 283793 212447
rect 283911 212329 295071 212447
rect 295189 212329 295231 212447
rect 295349 212329 295365 212447
rect -3403 212287 295365 212329
rect -3403 212169 -3387 212287
rect -3269 212169 -3227 212287
rect -3109 212169 13633 212287
rect 13751 212169 13793 212287
rect 13911 212169 31633 212287
rect 31751 212169 31793 212287
rect 31911 212169 49633 212287
rect 49751 212169 49793 212287
rect 49911 212169 67633 212287
rect 67751 212169 67793 212287
rect 67911 212169 85633 212287
rect 85751 212169 85793 212287
rect 85911 212169 103633 212287
rect 103751 212169 103793 212287
rect 103911 212169 121633 212287
rect 121751 212169 121793 212287
rect 121911 212169 139633 212287
rect 139751 212169 139793 212287
rect 139911 212169 157633 212287
rect 157751 212169 157793 212287
rect 157911 212169 175633 212287
rect 175751 212169 175793 212287
rect 175911 212169 193633 212287
rect 193751 212169 193793 212287
rect 193911 212169 211633 212287
rect 211751 212169 211793 212287
rect 211911 212169 229633 212287
rect 229751 212169 229793 212287
rect 229911 212169 247633 212287
rect 247751 212169 247793 212287
rect 247911 212169 265633 212287
rect 265751 212169 265793 212287
rect 265911 212169 283633 212287
rect 283751 212169 283793 212287
rect 283911 212169 295071 212287
rect 295189 212169 295231 212287
rect 295349 212169 295365 212287
rect -3403 212153 295365 212169
rect -2443 210587 294405 210603
rect -2443 210469 -2427 210587
rect -2309 210469 -2267 210587
rect -2149 210469 11773 210587
rect 11891 210469 11933 210587
rect 12051 210469 29773 210587
rect 29891 210469 29933 210587
rect 30051 210469 47773 210587
rect 47891 210469 47933 210587
rect 48051 210469 65773 210587
rect 65891 210469 65933 210587
rect 66051 210469 83773 210587
rect 83891 210469 83933 210587
rect 84051 210469 101773 210587
rect 101891 210469 101933 210587
rect 102051 210469 119773 210587
rect 119891 210469 119933 210587
rect 120051 210469 137773 210587
rect 137891 210469 137933 210587
rect 138051 210469 155773 210587
rect 155891 210469 155933 210587
rect 156051 210469 173773 210587
rect 173891 210469 173933 210587
rect 174051 210469 191773 210587
rect 191891 210469 191933 210587
rect 192051 210469 209773 210587
rect 209891 210469 209933 210587
rect 210051 210469 227773 210587
rect 227891 210469 227933 210587
rect 228051 210469 245773 210587
rect 245891 210469 245933 210587
rect 246051 210469 263773 210587
rect 263891 210469 263933 210587
rect 264051 210469 281773 210587
rect 281891 210469 281933 210587
rect 282051 210469 294111 210587
rect 294229 210469 294271 210587
rect 294389 210469 294405 210587
rect -2443 210427 294405 210469
rect -2443 210309 -2427 210427
rect -2309 210309 -2267 210427
rect -2149 210309 11773 210427
rect 11891 210309 11933 210427
rect 12051 210309 29773 210427
rect 29891 210309 29933 210427
rect 30051 210309 47773 210427
rect 47891 210309 47933 210427
rect 48051 210309 65773 210427
rect 65891 210309 65933 210427
rect 66051 210309 83773 210427
rect 83891 210309 83933 210427
rect 84051 210309 101773 210427
rect 101891 210309 101933 210427
rect 102051 210309 119773 210427
rect 119891 210309 119933 210427
rect 120051 210309 137773 210427
rect 137891 210309 137933 210427
rect 138051 210309 155773 210427
rect 155891 210309 155933 210427
rect 156051 210309 173773 210427
rect 173891 210309 173933 210427
rect 174051 210309 191773 210427
rect 191891 210309 191933 210427
rect 192051 210309 209773 210427
rect 209891 210309 209933 210427
rect 210051 210309 227773 210427
rect 227891 210309 227933 210427
rect 228051 210309 245773 210427
rect 245891 210309 245933 210427
rect 246051 210309 263773 210427
rect 263891 210309 263933 210427
rect 264051 210309 281773 210427
rect 281891 210309 281933 210427
rect 282051 210309 294111 210427
rect 294229 210309 294271 210427
rect 294389 210309 294405 210427
rect -2443 210293 294405 210309
rect -1483 208727 293445 208743
rect -1483 208609 -1467 208727
rect -1349 208609 -1307 208727
rect -1189 208609 9913 208727
rect 10031 208609 10073 208727
rect 10191 208609 27913 208727
rect 28031 208609 28073 208727
rect 28191 208609 45913 208727
rect 46031 208609 46073 208727
rect 46191 208609 63913 208727
rect 64031 208609 64073 208727
rect 64191 208609 81913 208727
rect 82031 208609 82073 208727
rect 82191 208609 99913 208727
rect 100031 208609 100073 208727
rect 100191 208609 117913 208727
rect 118031 208609 118073 208727
rect 118191 208609 135913 208727
rect 136031 208609 136073 208727
rect 136191 208609 153913 208727
rect 154031 208609 154073 208727
rect 154191 208609 171913 208727
rect 172031 208609 172073 208727
rect 172191 208609 189913 208727
rect 190031 208609 190073 208727
rect 190191 208609 207913 208727
rect 208031 208609 208073 208727
rect 208191 208609 225913 208727
rect 226031 208609 226073 208727
rect 226191 208609 243913 208727
rect 244031 208609 244073 208727
rect 244191 208609 261913 208727
rect 262031 208609 262073 208727
rect 262191 208609 279913 208727
rect 280031 208609 280073 208727
rect 280191 208609 293151 208727
rect 293269 208609 293311 208727
rect 293429 208609 293445 208727
rect -1483 208567 293445 208609
rect -1483 208449 -1467 208567
rect -1349 208449 -1307 208567
rect -1189 208449 9913 208567
rect 10031 208449 10073 208567
rect 10191 208449 27913 208567
rect 28031 208449 28073 208567
rect 28191 208449 45913 208567
rect 46031 208449 46073 208567
rect 46191 208449 63913 208567
rect 64031 208449 64073 208567
rect 64191 208449 81913 208567
rect 82031 208449 82073 208567
rect 82191 208449 99913 208567
rect 100031 208449 100073 208567
rect 100191 208449 117913 208567
rect 118031 208449 118073 208567
rect 118191 208449 135913 208567
rect 136031 208449 136073 208567
rect 136191 208449 153913 208567
rect 154031 208449 154073 208567
rect 154191 208449 171913 208567
rect 172031 208449 172073 208567
rect 172191 208449 189913 208567
rect 190031 208449 190073 208567
rect 190191 208449 207913 208567
rect 208031 208449 208073 208567
rect 208191 208449 225913 208567
rect 226031 208449 226073 208567
rect 226191 208449 243913 208567
rect 244031 208449 244073 208567
rect 244191 208449 261913 208567
rect 262031 208449 262073 208567
rect 262191 208449 279913 208567
rect 280031 208449 280073 208567
rect 280191 208449 293151 208567
rect 293269 208449 293311 208567
rect 293429 208449 293445 208567
rect -1483 208433 293445 208449
rect -4363 205307 296325 205323
rect -4363 205189 -3867 205307
rect -3749 205189 -3707 205307
rect -3589 205189 6493 205307
rect 6611 205189 6653 205307
rect 6771 205189 24493 205307
rect 24611 205189 24653 205307
rect 24771 205189 42493 205307
rect 42611 205189 42653 205307
rect 42771 205189 60493 205307
rect 60611 205189 60653 205307
rect 60771 205189 78493 205307
rect 78611 205189 78653 205307
rect 78771 205189 96493 205307
rect 96611 205189 96653 205307
rect 96771 205189 114493 205307
rect 114611 205189 114653 205307
rect 114771 205189 132493 205307
rect 132611 205189 132653 205307
rect 132771 205189 150493 205307
rect 150611 205189 150653 205307
rect 150771 205189 168493 205307
rect 168611 205189 168653 205307
rect 168771 205189 186493 205307
rect 186611 205189 186653 205307
rect 186771 205189 204493 205307
rect 204611 205189 204653 205307
rect 204771 205189 222493 205307
rect 222611 205189 222653 205307
rect 222771 205189 240493 205307
rect 240611 205189 240653 205307
rect 240771 205189 258493 205307
rect 258611 205189 258653 205307
rect 258771 205189 276493 205307
rect 276611 205189 276653 205307
rect 276771 205189 295551 205307
rect 295669 205189 295711 205307
rect 295829 205189 296325 205307
rect -4363 205147 296325 205189
rect -4363 205029 -3867 205147
rect -3749 205029 -3707 205147
rect -3589 205029 6493 205147
rect 6611 205029 6653 205147
rect 6771 205029 24493 205147
rect 24611 205029 24653 205147
rect 24771 205029 42493 205147
rect 42611 205029 42653 205147
rect 42771 205029 60493 205147
rect 60611 205029 60653 205147
rect 60771 205029 78493 205147
rect 78611 205029 78653 205147
rect 78771 205029 96493 205147
rect 96611 205029 96653 205147
rect 96771 205029 114493 205147
rect 114611 205029 114653 205147
rect 114771 205029 132493 205147
rect 132611 205029 132653 205147
rect 132771 205029 150493 205147
rect 150611 205029 150653 205147
rect 150771 205029 168493 205147
rect 168611 205029 168653 205147
rect 168771 205029 186493 205147
rect 186611 205029 186653 205147
rect 186771 205029 204493 205147
rect 204611 205029 204653 205147
rect 204771 205029 222493 205147
rect 222611 205029 222653 205147
rect 222771 205029 240493 205147
rect 240611 205029 240653 205147
rect 240771 205029 258493 205147
rect 258611 205029 258653 205147
rect 258771 205029 276493 205147
rect 276611 205029 276653 205147
rect 276771 205029 295551 205147
rect 295669 205029 295711 205147
rect 295829 205029 296325 205147
rect -4363 205013 296325 205029
rect -3403 203447 295365 203463
rect -3403 203329 -2907 203447
rect -2789 203329 -2747 203447
rect -2629 203329 4633 203447
rect 4751 203329 4793 203447
rect 4911 203329 22633 203447
rect 22751 203329 22793 203447
rect 22911 203329 40633 203447
rect 40751 203329 40793 203447
rect 40911 203329 58633 203447
rect 58751 203329 58793 203447
rect 58911 203329 76633 203447
rect 76751 203329 76793 203447
rect 76911 203329 94633 203447
rect 94751 203329 94793 203447
rect 94911 203329 112633 203447
rect 112751 203329 112793 203447
rect 112911 203329 130633 203447
rect 130751 203329 130793 203447
rect 130911 203329 148633 203447
rect 148751 203329 148793 203447
rect 148911 203329 166633 203447
rect 166751 203329 166793 203447
rect 166911 203329 184633 203447
rect 184751 203329 184793 203447
rect 184911 203329 202633 203447
rect 202751 203329 202793 203447
rect 202911 203329 220633 203447
rect 220751 203329 220793 203447
rect 220911 203329 238633 203447
rect 238751 203329 238793 203447
rect 238911 203329 256633 203447
rect 256751 203329 256793 203447
rect 256911 203329 274633 203447
rect 274751 203329 274793 203447
rect 274911 203329 294591 203447
rect 294709 203329 294751 203447
rect 294869 203329 295365 203447
rect -3403 203287 295365 203329
rect -3403 203169 -2907 203287
rect -2789 203169 -2747 203287
rect -2629 203169 4633 203287
rect 4751 203169 4793 203287
rect 4911 203169 22633 203287
rect 22751 203169 22793 203287
rect 22911 203169 40633 203287
rect 40751 203169 40793 203287
rect 40911 203169 58633 203287
rect 58751 203169 58793 203287
rect 58911 203169 76633 203287
rect 76751 203169 76793 203287
rect 76911 203169 94633 203287
rect 94751 203169 94793 203287
rect 94911 203169 112633 203287
rect 112751 203169 112793 203287
rect 112911 203169 130633 203287
rect 130751 203169 130793 203287
rect 130911 203169 148633 203287
rect 148751 203169 148793 203287
rect 148911 203169 166633 203287
rect 166751 203169 166793 203287
rect 166911 203169 184633 203287
rect 184751 203169 184793 203287
rect 184911 203169 202633 203287
rect 202751 203169 202793 203287
rect 202911 203169 220633 203287
rect 220751 203169 220793 203287
rect 220911 203169 238633 203287
rect 238751 203169 238793 203287
rect 238911 203169 256633 203287
rect 256751 203169 256793 203287
rect 256911 203169 274633 203287
rect 274751 203169 274793 203287
rect 274911 203169 294591 203287
rect 294709 203169 294751 203287
rect 294869 203169 295365 203287
rect -3403 203153 295365 203169
rect -2443 201587 294405 201603
rect -2443 201469 -1947 201587
rect -1829 201469 -1787 201587
rect -1669 201469 2773 201587
rect 2891 201469 2933 201587
rect 3051 201469 20773 201587
rect 20891 201469 20933 201587
rect 21051 201469 38773 201587
rect 38891 201469 38933 201587
rect 39051 201469 56773 201587
rect 56891 201469 56933 201587
rect 57051 201469 74773 201587
rect 74891 201469 74933 201587
rect 75051 201469 92773 201587
rect 92891 201469 92933 201587
rect 93051 201469 110773 201587
rect 110891 201469 110933 201587
rect 111051 201469 128773 201587
rect 128891 201469 128933 201587
rect 129051 201469 146773 201587
rect 146891 201469 146933 201587
rect 147051 201469 164773 201587
rect 164891 201469 164933 201587
rect 165051 201469 182773 201587
rect 182891 201469 182933 201587
rect 183051 201469 200773 201587
rect 200891 201469 200933 201587
rect 201051 201469 218773 201587
rect 218891 201469 218933 201587
rect 219051 201469 236773 201587
rect 236891 201469 236933 201587
rect 237051 201469 254773 201587
rect 254891 201469 254933 201587
rect 255051 201469 272773 201587
rect 272891 201469 272933 201587
rect 273051 201469 290773 201587
rect 290891 201469 290933 201587
rect 291051 201469 293631 201587
rect 293749 201469 293791 201587
rect 293909 201469 294405 201587
rect -2443 201427 294405 201469
rect -2443 201309 -1947 201427
rect -1829 201309 -1787 201427
rect -1669 201309 2773 201427
rect 2891 201309 2933 201427
rect 3051 201309 20773 201427
rect 20891 201309 20933 201427
rect 21051 201309 38773 201427
rect 38891 201309 38933 201427
rect 39051 201309 56773 201427
rect 56891 201309 56933 201427
rect 57051 201309 74773 201427
rect 74891 201309 74933 201427
rect 75051 201309 92773 201427
rect 92891 201309 92933 201427
rect 93051 201309 110773 201427
rect 110891 201309 110933 201427
rect 111051 201309 128773 201427
rect 128891 201309 128933 201427
rect 129051 201309 146773 201427
rect 146891 201309 146933 201427
rect 147051 201309 164773 201427
rect 164891 201309 164933 201427
rect 165051 201309 182773 201427
rect 182891 201309 182933 201427
rect 183051 201309 200773 201427
rect 200891 201309 200933 201427
rect 201051 201309 218773 201427
rect 218891 201309 218933 201427
rect 219051 201309 236773 201427
rect 236891 201309 236933 201427
rect 237051 201309 254773 201427
rect 254891 201309 254933 201427
rect 255051 201309 272773 201427
rect 272891 201309 272933 201427
rect 273051 201309 290773 201427
rect 290891 201309 290933 201427
rect 291051 201309 293631 201427
rect 293749 201309 293791 201427
rect 293909 201309 294405 201427
rect -2443 201293 294405 201309
rect -1483 199727 293445 199743
rect -1483 199609 -987 199727
rect -869 199609 -827 199727
rect -709 199609 913 199727
rect 1031 199609 1073 199727
rect 1191 199609 18913 199727
rect 19031 199609 19073 199727
rect 19191 199609 36913 199727
rect 37031 199609 37073 199727
rect 37191 199609 54913 199727
rect 55031 199609 55073 199727
rect 55191 199609 72913 199727
rect 73031 199609 73073 199727
rect 73191 199609 90913 199727
rect 91031 199609 91073 199727
rect 91191 199609 108913 199727
rect 109031 199609 109073 199727
rect 109191 199609 126913 199727
rect 127031 199609 127073 199727
rect 127191 199609 144913 199727
rect 145031 199609 145073 199727
rect 145191 199609 162913 199727
rect 163031 199609 163073 199727
rect 163191 199609 180913 199727
rect 181031 199609 181073 199727
rect 181191 199609 198913 199727
rect 199031 199609 199073 199727
rect 199191 199609 216913 199727
rect 217031 199609 217073 199727
rect 217191 199609 234913 199727
rect 235031 199609 235073 199727
rect 235191 199609 252913 199727
rect 253031 199609 253073 199727
rect 253191 199609 270913 199727
rect 271031 199609 271073 199727
rect 271191 199609 288913 199727
rect 289031 199609 289073 199727
rect 289191 199609 292671 199727
rect 292789 199609 292831 199727
rect 292949 199609 293445 199727
rect -1483 199567 293445 199609
rect -1483 199449 -987 199567
rect -869 199449 -827 199567
rect -709 199449 913 199567
rect 1031 199449 1073 199567
rect 1191 199449 18913 199567
rect 19031 199449 19073 199567
rect 19191 199449 36913 199567
rect 37031 199449 37073 199567
rect 37191 199449 54913 199567
rect 55031 199449 55073 199567
rect 55191 199449 72913 199567
rect 73031 199449 73073 199567
rect 73191 199449 90913 199567
rect 91031 199449 91073 199567
rect 91191 199449 108913 199567
rect 109031 199449 109073 199567
rect 109191 199449 126913 199567
rect 127031 199449 127073 199567
rect 127191 199449 144913 199567
rect 145031 199449 145073 199567
rect 145191 199449 162913 199567
rect 163031 199449 163073 199567
rect 163191 199449 180913 199567
rect 181031 199449 181073 199567
rect 181191 199449 198913 199567
rect 199031 199449 199073 199567
rect 199191 199449 216913 199567
rect 217031 199449 217073 199567
rect 217191 199449 234913 199567
rect 235031 199449 235073 199567
rect 235191 199449 252913 199567
rect 253031 199449 253073 199567
rect 253191 199449 270913 199567
rect 271031 199449 271073 199567
rect 271191 199449 288913 199567
rect 289031 199449 289073 199567
rect 289191 199449 292671 199567
rect 292789 199449 292831 199567
rect 292949 199449 293445 199567
rect -1483 199433 293445 199449
rect -4363 196307 296325 196323
rect -4363 196189 -4347 196307
rect -4229 196189 -4187 196307
rect -4069 196189 15493 196307
rect 15611 196189 15653 196307
rect 15771 196189 33493 196307
rect 33611 196189 33653 196307
rect 33771 196189 51493 196307
rect 51611 196189 51653 196307
rect 51771 196189 69493 196307
rect 69611 196189 69653 196307
rect 69771 196189 87493 196307
rect 87611 196189 87653 196307
rect 87771 196189 105493 196307
rect 105611 196189 105653 196307
rect 105771 196189 123493 196307
rect 123611 196189 123653 196307
rect 123771 196189 141493 196307
rect 141611 196189 141653 196307
rect 141771 196189 159493 196307
rect 159611 196189 159653 196307
rect 159771 196189 177493 196307
rect 177611 196189 177653 196307
rect 177771 196189 195493 196307
rect 195611 196189 195653 196307
rect 195771 196189 213493 196307
rect 213611 196189 213653 196307
rect 213771 196189 231493 196307
rect 231611 196189 231653 196307
rect 231771 196189 249493 196307
rect 249611 196189 249653 196307
rect 249771 196189 267493 196307
rect 267611 196189 267653 196307
rect 267771 196189 285493 196307
rect 285611 196189 285653 196307
rect 285771 196189 296031 196307
rect 296149 196189 296191 196307
rect 296309 196189 296325 196307
rect -4363 196147 296325 196189
rect -4363 196029 -4347 196147
rect -4229 196029 -4187 196147
rect -4069 196029 15493 196147
rect 15611 196029 15653 196147
rect 15771 196029 33493 196147
rect 33611 196029 33653 196147
rect 33771 196029 51493 196147
rect 51611 196029 51653 196147
rect 51771 196029 69493 196147
rect 69611 196029 69653 196147
rect 69771 196029 87493 196147
rect 87611 196029 87653 196147
rect 87771 196029 105493 196147
rect 105611 196029 105653 196147
rect 105771 196029 123493 196147
rect 123611 196029 123653 196147
rect 123771 196029 141493 196147
rect 141611 196029 141653 196147
rect 141771 196029 159493 196147
rect 159611 196029 159653 196147
rect 159771 196029 177493 196147
rect 177611 196029 177653 196147
rect 177771 196029 195493 196147
rect 195611 196029 195653 196147
rect 195771 196029 213493 196147
rect 213611 196029 213653 196147
rect 213771 196029 231493 196147
rect 231611 196029 231653 196147
rect 231771 196029 249493 196147
rect 249611 196029 249653 196147
rect 249771 196029 267493 196147
rect 267611 196029 267653 196147
rect 267771 196029 285493 196147
rect 285611 196029 285653 196147
rect 285771 196029 296031 196147
rect 296149 196029 296191 196147
rect 296309 196029 296325 196147
rect -4363 196013 296325 196029
rect -3403 194447 295365 194463
rect -3403 194329 -3387 194447
rect -3269 194329 -3227 194447
rect -3109 194329 13633 194447
rect 13751 194329 13793 194447
rect 13911 194329 31633 194447
rect 31751 194329 31793 194447
rect 31911 194329 49633 194447
rect 49751 194329 49793 194447
rect 49911 194329 67633 194447
rect 67751 194329 67793 194447
rect 67911 194329 85633 194447
rect 85751 194329 85793 194447
rect 85911 194329 103633 194447
rect 103751 194329 103793 194447
rect 103911 194329 121633 194447
rect 121751 194329 121793 194447
rect 121911 194329 139633 194447
rect 139751 194329 139793 194447
rect 139911 194329 157633 194447
rect 157751 194329 157793 194447
rect 157911 194329 175633 194447
rect 175751 194329 175793 194447
rect 175911 194329 193633 194447
rect 193751 194329 193793 194447
rect 193911 194329 211633 194447
rect 211751 194329 211793 194447
rect 211911 194329 229633 194447
rect 229751 194329 229793 194447
rect 229911 194329 247633 194447
rect 247751 194329 247793 194447
rect 247911 194329 265633 194447
rect 265751 194329 265793 194447
rect 265911 194329 283633 194447
rect 283751 194329 283793 194447
rect 283911 194329 295071 194447
rect 295189 194329 295231 194447
rect 295349 194329 295365 194447
rect -3403 194287 295365 194329
rect -3403 194169 -3387 194287
rect -3269 194169 -3227 194287
rect -3109 194169 13633 194287
rect 13751 194169 13793 194287
rect 13911 194169 31633 194287
rect 31751 194169 31793 194287
rect 31911 194169 49633 194287
rect 49751 194169 49793 194287
rect 49911 194169 67633 194287
rect 67751 194169 67793 194287
rect 67911 194169 85633 194287
rect 85751 194169 85793 194287
rect 85911 194169 103633 194287
rect 103751 194169 103793 194287
rect 103911 194169 121633 194287
rect 121751 194169 121793 194287
rect 121911 194169 139633 194287
rect 139751 194169 139793 194287
rect 139911 194169 157633 194287
rect 157751 194169 157793 194287
rect 157911 194169 175633 194287
rect 175751 194169 175793 194287
rect 175911 194169 193633 194287
rect 193751 194169 193793 194287
rect 193911 194169 211633 194287
rect 211751 194169 211793 194287
rect 211911 194169 229633 194287
rect 229751 194169 229793 194287
rect 229911 194169 247633 194287
rect 247751 194169 247793 194287
rect 247911 194169 265633 194287
rect 265751 194169 265793 194287
rect 265911 194169 283633 194287
rect 283751 194169 283793 194287
rect 283911 194169 295071 194287
rect 295189 194169 295231 194287
rect 295349 194169 295365 194287
rect -3403 194153 295365 194169
rect -2443 192587 294405 192603
rect -2443 192469 -2427 192587
rect -2309 192469 -2267 192587
rect -2149 192469 11773 192587
rect 11891 192469 11933 192587
rect 12051 192469 29773 192587
rect 29891 192469 29933 192587
rect 30051 192469 47773 192587
rect 47891 192469 47933 192587
rect 48051 192469 65773 192587
rect 65891 192469 65933 192587
rect 66051 192469 83773 192587
rect 83891 192469 83933 192587
rect 84051 192469 101773 192587
rect 101891 192469 101933 192587
rect 102051 192469 119773 192587
rect 119891 192469 119933 192587
rect 120051 192469 137773 192587
rect 137891 192469 137933 192587
rect 138051 192469 155773 192587
rect 155891 192469 155933 192587
rect 156051 192469 173773 192587
rect 173891 192469 173933 192587
rect 174051 192469 191773 192587
rect 191891 192469 191933 192587
rect 192051 192469 209773 192587
rect 209891 192469 209933 192587
rect 210051 192469 227773 192587
rect 227891 192469 227933 192587
rect 228051 192469 245773 192587
rect 245891 192469 245933 192587
rect 246051 192469 263773 192587
rect 263891 192469 263933 192587
rect 264051 192469 281773 192587
rect 281891 192469 281933 192587
rect 282051 192469 294111 192587
rect 294229 192469 294271 192587
rect 294389 192469 294405 192587
rect -2443 192427 294405 192469
rect -2443 192309 -2427 192427
rect -2309 192309 -2267 192427
rect -2149 192309 11773 192427
rect 11891 192309 11933 192427
rect 12051 192309 29773 192427
rect 29891 192309 29933 192427
rect 30051 192309 47773 192427
rect 47891 192309 47933 192427
rect 48051 192309 65773 192427
rect 65891 192309 65933 192427
rect 66051 192309 83773 192427
rect 83891 192309 83933 192427
rect 84051 192309 101773 192427
rect 101891 192309 101933 192427
rect 102051 192309 119773 192427
rect 119891 192309 119933 192427
rect 120051 192309 137773 192427
rect 137891 192309 137933 192427
rect 138051 192309 155773 192427
rect 155891 192309 155933 192427
rect 156051 192309 173773 192427
rect 173891 192309 173933 192427
rect 174051 192309 191773 192427
rect 191891 192309 191933 192427
rect 192051 192309 209773 192427
rect 209891 192309 209933 192427
rect 210051 192309 227773 192427
rect 227891 192309 227933 192427
rect 228051 192309 245773 192427
rect 245891 192309 245933 192427
rect 246051 192309 263773 192427
rect 263891 192309 263933 192427
rect 264051 192309 281773 192427
rect 281891 192309 281933 192427
rect 282051 192309 294111 192427
rect 294229 192309 294271 192427
rect 294389 192309 294405 192427
rect -2443 192293 294405 192309
rect -1483 190727 293445 190743
rect -1483 190609 -1467 190727
rect -1349 190609 -1307 190727
rect -1189 190609 9913 190727
rect 10031 190609 10073 190727
rect 10191 190609 27913 190727
rect 28031 190609 28073 190727
rect 28191 190609 45913 190727
rect 46031 190609 46073 190727
rect 46191 190609 63913 190727
rect 64031 190609 64073 190727
rect 64191 190609 81913 190727
rect 82031 190609 82073 190727
rect 82191 190609 99913 190727
rect 100031 190609 100073 190727
rect 100191 190609 117913 190727
rect 118031 190609 118073 190727
rect 118191 190609 135913 190727
rect 136031 190609 136073 190727
rect 136191 190609 153913 190727
rect 154031 190609 154073 190727
rect 154191 190609 171913 190727
rect 172031 190609 172073 190727
rect 172191 190609 189913 190727
rect 190031 190609 190073 190727
rect 190191 190609 207913 190727
rect 208031 190609 208073 190727
rect 208191 190609 225913 190727
rect 226031 190609 226073 190727
rect 226191 190609 243913 190727
rect 244031 190609 244073 190727
rect 244191 190609 261913 190727
rect 262031 190609 262073 190727
rect 262191 190609 279913 190727
rect 280031 190609 280073 190727
rect 280191 190609 293151 190727
rect 293269 190609 293311 190727
rect 293429 190609 293445 190727
rect -1483 190567 293445 190609
rect -1483 190449 -1467 190567
rect -1349 190449 -1307 190567
rect -1189 190449 9913 190567
rect 10031 190449 10073 190567
rect 10191 190449 27913 190567
rect 28031 190449 28073 190567
rect 28191 190449 45913 190567
rect 46031 190449 46073 190567
rect 46191 190449 63913 190567
rect 64031 190449 64073 190567
rect 64191 190449 81913 190567
rect 82031 190449 82073 190567
rect 82191 190449 99913 190567
rect 100031 190449 100073 190567
rect 100191 190449 117913 190567
rect 118031 190449 118073 190567
rect 118191 190449 135913 190567
rect 136031 190449 136073 190567
rect 136191 190449 153913 190567
rect 154031 190449 154073 190567
rect 154191 190449 171913 190567
rect 172031 190449 172073 190567
rect 172191 190449 189913 190567
rect 190031 190449 190073 190567
rect 190191 190449 207913 190567
rect 208031 190449 208073 190567
rect 208191 190449 225913 190567
rect 226031 190449 226073 190567
rect 226191 190449 243913 190567
rect 244031 190449 244073 190567
rect 244191 190449 261913 190567
rect 262031 190449 262073 190567
rect 262191 190449 279913 190567
rect 280031 190449 280073 190567
rect 280191 190449 293151 190567
rect 293269 190449 293311 190567
rect 293429 190449 293445 190567
rect -1483 190433 293445 190449
rect -4363 187307 296325 187323
rect -4363 187189 -3867 187307
rect -3749 187189 -3707 187307
rect -3589 187189 6493 187307
rect 6611 187189 6653 187307
rect 6771 187189 24493 187307
rect 24611 187189 24653 187307
rect 24771 187189 42493 187307
rect 42611 187189 42653 187307
rect 42771 187189 60493 187307
rect 60611 187189 60653 187307
rect 60771 187189 78493 187307
rect 78611 187189 78653 187307
rect 78771 187189 96493 187307
rect 96611 187189 96653 187307
rect 96771 187189 114493 187307
rect 114611 187189 114653 187307
rect 114771 187189 132493 187307
rect 132611 187189 132653 187307
rect 132771 187189 150493 187307
rect 150611 187189 150653 187307
rect 150771 187189 168493 187307
rect 168611 187189 168653 187307
rect 168771 187189 186493 187307
rect 186611 187189 186653 187307
rect 186771 187189 204493 187307
rect 204611 187189 204653 187307
rect 204771 187189 222493 187307
rect 222611 187189 222653 187307
rect 222771 187189 240493 187307
rect 240611 187189 240653 187307
rect 240771 187189 258493 187307
rect 258611 187189 258653 187307
rect 258771 187189 276493 187307
rect 276611 187189 276653 187307
rect 276771 187189 295551 187307
rect 295669 187189 295711 187307
rect 295829 187189 296325 187307
rect -4363 187147 296325 187189
rect -4363 187029 -3867 187147
rect -3749 187029 -3707 187147
rect -3589 187029 6493 187147
rect 6611 187029 6653 187147
rect 6771 187029 24493 187147
rect 24611 187029 24653 187147
rect 24771 187029 42493 187147
rect 42611 187029 42653 187147
rect 42771 187029 60493 187147
rect 60611 187029 60653 187147
rect 60771 187029 78493 187147
rect 78611 187029 78653 187147
rect 78771 187029 96493 187147
rect 96611 187029 96653 187147
rect 96771 187029 114493 187147
rect 114611 187029 114653 187147
rect 114771 187029 132493 187147
rect 132611 187029 132653 187147
rect 132771 187029 150493 187147
rect 150611 187029 150653 187147
rect 150771 187029 168493 187147
rect 168611 187029 168653 187147
rect 168771 187029 186493 187147
rect 186611 187029 186653 187147
rect 186771 187029 204493 187147
rect 204611 187029 204653 187147
rect 204771 187029 222493 187147
rect 222611 187029 222653 187147
rect 222771 187029 240493 187147
rect 240611 187029 240653 187147
rect 240771 187029 258493 187147
rect 258611 187029 258653 187147
rect 258771 187029 276493 187147
rect 276611 187029 276653 187147
rect 276771 187029 295551 187147
rect 295669 187029 295711 187147
rect 295829 187029 296325 187147
rect -4363 187013 296325 187029
rect -3403 185447 295365 185463
rect -3403 185329 -2907 185447
rect -2789 185329 -2747 185447
rect -2629 185329 4633 185447
rect 4751 185329 4793 185447
rect 4911 185329 22633 185447
rect 22751 185329 22793 185447
rect 22911 185329 40633 185447
rect 40751 185329 40793 185447
rect 40911 185329 58633 185447
rect 58751 185329 58793 185447
rect 58911 185329 76633 185447
rect 76751 185329 76793 185447
rect 76911 185329 94633 185447
rect 94751 185329 94793 185447
rect 94911 185329 112633 185447
rect 112751 185329 112793 185447
rect 112911 185329 130633 185447
rect 130751 185329 130793 185447
rect 130911 185329 148633 185447
rect 148751 185329 148793 185447
rect 148911 185329 166633 185447
rect 166751 185329 166793 185447
rect 166911 185329 184633 185447
rect 184751 185329 184793 185447
rect 184911 185329 202633 185447
rect 202751 185329 202793 185447
rect 202911 185329 220633 185447
rect 220751 185329 220793 185447
rect 220911 185329 238633 185447
rect 238751 185329 238793 185447
rect 238911 185329 256633 185447
rect 256751 185329 256793 185447
rect 256911 185329 274633 185447
rect 274751 185329 274793 185447
rect 274911 185329 294591 185447
rect 294709 185329 294751 185447
rect 294869 185329 295365 185447
rect -3403 185287 295365 185329
rect -3403 185169 -2907 185287
rect -2789 185169 -2747 185287
rect -2629 185169 4633 185287
rect 4751 185169 4793 185287
rect 4911 185169 22633 185287
rect 22751 185169 22793 185287
rect 22911 185169 40633 185287
rect 40751 185169 40793 185287
rect 40911 185169 58633 185287
rect 58751 185169 58793 185287
rect 58911 185169 76633 185287
rect 76751 185169 76793 185287
rect 76911 185169 94633 185287
rect 94751 185169 94793 185287
rect 94911 185169 112633 185287
rect 112751 185169 112793 185287
rect 112911 185169 130633 185287
rect 130751 185169 130793 185287
rect 130911 185169 148633 185287
rect 148751 185169 148793 185287
rect 148911 185169 166633 185287
rect 166751 185169 166793 185287
rect 166911 185169 184633 185287
rect 184751 185169 184793 185287
rect 184911 185169 202633 185287
rect 202751 185169 202793 185287
rect 202911 185169 220633 185287
rect 220751 185169 220793 185287
rect 220911 185169 238633 185287
rect 238751 185169 238793 185287
rect 238911 185169 256633 185287
rect 256751 185169 256793 185287
rect 256911 185169 274633 185287
rect 274751 185169 274793 185287
rect 274911 185169 294591 185287
rect 294709 185169 294751 185287
rect 294869 185169 295365 185287
rect -3403 185153 295365 185169
rect -2443 183587 294405 183603
rect -2443 183469 -1947 183587
rect -1829 183469 -1787 183587
rect -1669 183469 2773 183587
rect 2891 183469 2933 183587
rect 3051 183469 20773 183587
rect 20891 183469 20933 183587
rect 21051 183469 38773 183587
rect 38891 183469 38933 183587
rect 39051 183469 56773 183587
rect 56891 183469 56933 183587
rect 57051 183469 74773 183587
rect 74891 183469 74933 183587
rect 75051 183469 92773 183587
rect 92891 183469 92933 183587
rect 93051 183469 110773 183587
rect 110891 183469 110933 183587
rect 111051 183469 128773 183587
rect 128891 183469 128933 183587
rect 129051 183469 146773 183587
rect 146891 183469 146933 183587
rect 147051 183469 164773 183587
rect 164891 183469 164933 183587
rect 165051 183469 182773 183587
rect 182891 183469 182933 183587
rect 183051 183469 200773 183587
rect 200891 183469 200933 183587
rect 201051 183469 218773 183587
rect 218891 183469 218933 183587
rect 219051 183469 236773 183587
rect 236891 183469 236933 183587
rect 237051 183469 254773 183587
rect 254891 183469 254933 183587
rect 255051 183469 272773 183587
rect 272891 183469 272933 183587
rect 273051 183469 290773 183587
rect 290891 183469 290933 183587
rect 291051 183469 293631 183587
rect 293749 183469 293791 183587
rect 293909 183469 294405 183587
rect -2443 183427 294405 183469
rect -2443 183309 -1947 183427
rect -1829 183309 -1787 183427
rect -1669 183309 2773 183427
rect 2891 183309 2933 183427
rect 3051 183309 20773 183427
rect 20891 183309 20933 183427
rect 21051 183309 38773 183427
rect 38891 183309 38933 183427
rect 39051 183309 56773 183427
rect 56891 183309 56933 183427
rect 57051 183309 74773 183427
rect 74891 183309 74933 183427
rect 75051 183309 92773 183427
rect 92891 183309 92933 183427
rect 93051 183309 110773 183427
rect 110891 183309 110933 183427
rect 111051 183309 128773 183427
rect 128891 183309 128933 183427
rect 129051 183309 146773 183427
rect 146891 183309 146933 183427
rect 147051 183309 164773 183427
rect 164891 183309 164933 183427
rect 165051 183309 182773 183427
rect 182891 183309 182933 183427
rect 183051 183309 200773 183427
rect 200891 183309 200933 183427
rect 201051 183309 218773 183427
rect 218891 183309 218933 183427
rect 219051 183309 236773 183427
rect 236891 183309 236933 183427
rect 237051 183309 254773 183427
rect 254891 183309 254933 183427
rect 255051 183309 272773 183427
rect 272891 183309 272933 183427
rect 273051 183309 290773 183427
rect 290891 183309 290933 183427
rect 291051 183309 293631 183427
rect 293749 183309 293791 183427
rect 293909 183309 294405 183427
rect -2443 183293 294405 183309
rect -1483 181727 293445 181743
rect -1483 181609 -987 181727
rect -869 181609 -827 181727
rect -709 181609 913 181727
rect 1031 181609 1073 181727
rect 1191 181609 18913 181727
rect 19031 181609 19073 181727
rect 19191 181609 36913 181727
rect 37031 181609 37073 181727
rect 37191 181609 54913 181727
rect 55031 181609 55073 181727
rect 55191 181609 72913 181727
rect 73031 181609 73073 181727
rect 73191 181609 90913 181727
rect 91031 181609 91073 181727
rect 91191 181609 108913 181727
rect 109031 181609 109073 181727
rect 109191 181609 126913 181727
rect 127031 181609 127073 181727
rect 127191 181609 144913 181727
rect 145031 181609 145073 181727
rect 145191 181609 162913 181727
rect 163031 181609 163073 181727
rect 163191 181609 180913 181727
rect 181031 181609 181073 181727
rect 181191 181609 198913 181727
rect 199031 181609 199073 181727
rect 199191 181609 216913 181727
rect 217031 181609 217073 181727
rect 217191 181609 234913 181727
rect 235031 181609 235073 181727
rect 235191 181609 252913 181727
rect 253031 181609 253073 181727
rect 253191 181609 270913 181727
rect 271031 181609 271073 181727
rect 271191 181609 288913 181727
rect 289031 181609 289073 181727
rect 289191 181609 292671 181727
rect 292789 181609 292831 181727
rect 292949 181609 293445 181727
rect -1483 181567 293445 181609
rect -1483 181449 -987 181567
rect -869 181449 -827 181567
rect -709 181449 913 181567
rect 1031 181449 1073 181567
rect 1191 181449 18913 181567
rect 19031 181449 19073 181567
rect 19191 181449 36913 181567
rect 37031 181449 37073 181567
rect 37191 181449 54913 181567
rect 55031 181449 55073 181567
rect 55191 181449 72913 181567
rect 73031 181449 73073 181567
rect 73191 181449 90913 181567
rect 91031 181449 91073 181567
rect 91191 181449 108913 181567
rect 109031 181449 109073 181567
rect 109191 181449 126913 181567
rect 127031 181449 127073 181567
rect 127191 181449 144913 181567
rect 145031 181449 145073 181567
rect 145191 181449 162913 181567
rect 163031 181449 163073 181567
rect 163191 181449 180913 181567
rect 181031 181449 181073 181567
rect 181191 181449 198913 181567
rect 199031 181449 199073 181567
rect 199191 181449 216913 181567
rect 217031 181449 217073 181567
rect 217191 181449 234913 181567
rect 235031 181449 235073 181567
rect 235191 181449 252913 181567
rect 253031 181449 253073 181567
rect 253191 181449 270913 181567
rect 271031 181449 271073 181567
rect 271191 181449 288913 181567
rect 289031 181449 289073 181567
rect 289191 181449 292671 181567
rect 292789 181449 292831 181567
rect 292949 181449 293445 181567
rect -1483 181433 293445 181449
rect -4363 178307 296325 178323
rect -4363 178189 -4347 178307
rect -4229 178189 -4187 178307
rect -4069 178189 15493 178307
rect 15611 178189 15653 178307
rect 15771 178189 33493 178307
rect 33611 178189 33653 178307
rect 33771 178189 51493 178307
rect 51611 178189 51653 178307
rect 51771 178189 69493 178307
rect 69611 178189 69653 178307
rect 69771 178189 87493 178307
rect 87611 178189 87653 178307
rect 87771 178189 105493 178307
rect 105611 178189 105653 178307
rect 105771 178189 123493 178307
rect 123611 178189 123653 178307
rect 123771 178189 141493 178307
rect 141611 178189 141653 178307
rect 141771 178189 159493 178307
rect 159611 178189 159653 178307
rect 159771 178189 177493 178307
rect 177611 178189 177653 178307
rect 177771 178189 195493 178307
rect 195611 178189 195653 178307
rect 195771 178189 213493 178307
rect 213611 178189 213653 178307
rect 213771 178189 231493 178307
rect 231611 178189 231653 178307
rect 231771 178189 249493 178307
rect 249611 178189 249653 178307
rect 249771 178189 267493 178307
rect 267611 178189 267653 178307
rect 267771 178189 285493 178307
rect 285611 178189 285653 178307
rect 285771 178189 296031 178307
rect 296149 178189 296191 178307
rect 296309 178189 296325 178307
rect -4363 178147 296325 178189
rect -4363 178029 -4347 178147
rect -4229 178029 -4187 178147
rect -4069 178029 15493 178147
rect 15611 178029 15653 178147
rect 15771 178029 33493 178147
rect 33611 178029 33653 178147
rect 33771 178029 51493 178147
rect 51611 178029 51653 178147
rect 51771 178029 69493 178147
rect 69611 178029 69653 178147
rect 69771 178029 87493 178147
rect 87611 178029 87653 178147
rect 87771 178029 105493 178147
rect 105611 178029 105653 178147
rect 105771 178029 123493 178147
rect 123611 178029 123653 178147
rect 123771 178029 141493 178147
rect 141611 178029 141653 178147
rect 141771 178029 159493 178147
rect 159611 178029 159653 178147
rect 159771 178029 177493 178147
rect 177611 178029 177653 178147
rect 177771 178029 195493 178147
rect 195611 178029 195653 178147
rect 195771 178029 213493 178147
rect 213611 178029 213653 178147
rect 213771 178029 231493 178147
rect 231611 178029 231653 178147
rect 231771 178029 249493 178147
rect 249611 178029 249653 178147
rect 249771 178029 267493 178147
rect 267611 178029 267653 178147
rect 267771 178029 285493 178147
rect 285611 178029 285653 178147
rect 285771 178029 296031 178147
rect 296149 178029 296191 178147
rect 296309 178029 296325 178147
rect -4363 178013 296325 178029
rect -3403 176447 295365 176463
rect -3403 176329 -3387 176447
rect -3269 176329 -3227 176447
rect -3109 176329 13633 176447
rect 13751 176329 13793 176447
rect 13911 176329 31633 176447
rect 31751 176329 31793 176447
rect 31911 176329 49633 176447
rect 49751 176329 49793 176447
rect 49911 176329 67633 176447
rect 67751 176329 67793 176447
rect 67911 176329 85633 176447
rect 85751 176329 85793 176447
rect 85911 176329 103633 176447
rect 103751 176329 103793 176447
rect 103911 176329 121633 176447
rect 121751 176329 121793 176447
rect 121911 176329 139633 176447
rect 139751 176329 139793 176447
rect 139911 176329 157633 176447
rect 157751 176329 157793 176447
rect 157911 176329 175633 176447
rect 175751 176329 175793 176447
rect 175911 176329 193633 176447
rect 193751 176329 193793 176447
rect 193911 176329 211633 176447
rect 211751 176329 211793 176447
rect 211911 176329 229633 176447
rect 229751 176329 229793 176447
rect 229911 176329 247633 176447
rect 247751 176329 247793 176447
rect 247911 176329 265633 176447
rect 265751 176329 265793 176447
rect 265911 176329 283633 176447
rect 283751 176329 283793 176447
rect 283911 176329 295071 176447
rect 295189 176329 295231 176447
rect 295349 176329 295365 176447
rect -3403 176287 295365 176329
rect -3403 176169 -3387 176287
rect -3269 176169 -3227 176287
rect -3109 176169 13633 176287
rect 13751 176169 13793 176287
rect 13911 176169 31633 176287
rect 31751 176169 31793 176287
rect 31911 176169 49633 176287
rect 49751 176169 49793 176287
rect 49911 176169 67633 176287
rect 67751 176169 67793 176287
rect 67911 176169 85633 176287
rect 85751 176169 85793 176287
rect 85911 176169 103633 176287
rect 103751 176169 103793 176287
rect 103911 176169 121633 176287
rect 121751 176169 121793 176287
rect 121911 176169 139633 176287
rect 139751 176169 139793 176287
rect 139911 176169 157633 176287
rect 157751 176169 157793 176287
rect 157911 176169 175633 176287
rect 175751 176169 175793 176287
rect 175911 176169 193633 176287
rect 193751 176169 193793 176287
rect 193911 176169 211633 176287
rect 211751 176169 211793 176287
rect 211911 176169 229633 176287
rect 229751 176169 229793 176287
rect 229911 176169 247633 176287
rect 247751 176169 247793 176287
rect 247911 176169 265633 176287
rect 265751 176169 265793 176287
rect 265911 176169 283633 176287
rect 283751 176169 283793 176287
rect 283911 176169 295071 176287
rect 295189 176169 295231 176287
rect 295349 176169 295365 176287
rect -3403 176153 295365 176169
rect -2443 174587 294405 174603
rect -2443 174469 -2427 174587
rect -2309 174469 -2267 174587
rect -2149 174469 11773 174587
rect 11891 174469 11933 174587
rect 12051 174469 29773 174587
rect 29891 174469 29933 174587
rect 30051 174469 47773 174587
rect 47891 174469 47933 174587
rect 48051 174469 65773 174587
rect 65891 174469 65933 174587
rect 66051 174469 83773 174587
rect 83891 174469 83933 174587
rect 84051 174469 101773 174587
rect 101891 174469 101933 174587
rect 102051 174469 119773 174587
rect 119891 174469 119933 174587
rect 120051 174469 137773 174587
rect 137891 174469 137933 174587
rect 138051 174469 155773 174587
rect 155891 174469 155933 174587
rect 156051 174469 173773 174587
rect 173891 174469 173933 174587
rect 174051 174469 191773 174587
rect 191891 174469 191933 174587
rect 192051 174469 209773 174587
rect 209891 174469 209933 174587
rect 210051 174469 227773 174587
rect 227891 174469 227933 174587
rect 228051 174469 245773 174587
rect 245891 174469 245933 174587
rect 246051 174469 263773 174587
rect 263891 174469 263933 174587
rect 264051 174469 281773 174587
rect 281891 174469 281933 174587
rect 282051 174469 294111 174587
rect 294229 174469 294271 174587
rect 294389 174469 294405 174587
rect -2443 174427 294405 174469
rect -2443 174309 -2427 174427
rect -2309 174309 -2267 174427
rect -2149 174309 11773 174427
rect 11891 174309 11933 174427
rect 12051 174309 29773 174427
rect 29891 174309 29933 174427
rect 30051 174309 47773 174427
rect 47891 174309 47933 174427
rect 48051 174309 65773 174427
rect 65891 174309 65933 174427
rect 66051 174309 83773 174427
rect 83891 174309 83933 174427
rect 84051 174309 101773 174427
rect 101891 174309 101933 174427
rect 102051 174309 119773 174427
rect 119891 174309 119933 174427
rect 120051 174309 137773 174427
rect 137891 174309 137933 174427
rect 138051 174309 155773 174427
rect 155891 174309 155933 174427
rect 156051 174309 173773 174427
rect 173891 174309 173933 174427
rect 174051 174309 191773 174427
rect 191891 174309 191933 174427
rect 192051 174309 209773 174427
rect 209891 174309 209933 174427
rect 210051 174309 227773 174427
rect 227891 174309 227933 174427
rect 228051 174309 245773 174427
rect 245891 174309 245933 174427
rect 246051 174309 263773 174427
rect 263891 174309 263933 174427
rect 264051 174309 281773 174427
rect 281891 174309 281933 174427
rect 282051 174309 294111 174427
rect 294229 174309 294271 174427
rect 294389 174309 294405 174427
rect -2443 174293 294405 174309
rect -1483 172727 293445 172743
rect -1483 172609 -1467 172727
rect -1349 172609 -1307 172727
rect -1189 172609 9913 172727
rect 10031 172609 10073 172727
rect 10191 172609 27913 172727
rect 28031 172609 28073 172727
rect 28191 172609 45913 172727
rect 46031 172609 46073 172727
rect 46191 172609 63913 172727
rect 64031 172609 64073 172727
rect 64191 172609 81913 172727
rect 82031 172609 82073 172727
rect 82191 172609 99913 172727
rect 100031 172609 100073 172727
rect 100191 172609 117913 172727
rect 118031 172609 118073 172727
rect 118191 172609 135913 172727
rect 136031 172609 136073 172727
rect 136191 172609 153913 172727
rect 154031 172609 154073 172727
rect 154191 172609 171913 172727
rect 172031 172609 172073 172727
rect 172191 172609 189913 172727
rect 190031 172609 190073 172727
rect 190191 172609 207913 172727
rect 208031 172609 208073 172727
rect 208191 172609 225913 172727
rect 226031 172609 226073 172727
rect 226191 172609 243913 172727
rect 244031 172609 244073 172727
rect 244191 172609 261913 172727
rect 262031 172609 262073 172727
rect 262191 172609 279913 172727
rect 280031 172609 280073 172727
rect 280191 172609 293151 172727
rect 293269 172609 293311 172727
rect 293429 172609 293445 172727
rect -1483 172567 293445 172609
rect -1483 172449 -1467 172567
rect -1349 172449 -1307 172567
rect -1189 172449 9913 172567
rect 10031 172449 10073 172567
rect 10191 172449 27913 172567
rect 28031 172449 28073 172567
rect 28191 172449 45913 172567
rect 46031 172449 46073 172567
rect 46191 172449 63913 172567
rect 64031 172449 64073 172567
rect 64191 172449 81913 172567
rect 82031 172449 82073 172567
rect 82191 172449 99913 172567
rect 100031 172449 100073 172567
rect 100191 172449 117913 172567
rect 118031 172449 118073 172567
rect 118191 172449 135913 172567
rect 136031 172449 136073 172567
rect 136191 172449 153913 172567
rect 154031 172449 154073 172567
rect 154191 172449 171913 172567
rect 172031 172449 172073 172567
rect 172191 172449 189913 172567
rect 190031 172449 190073 172567
rect 190191 172449 207913 172567
rect 208031 172449 208073 172567
rect 208191 172449 225913 172567
rect 226031 172449 226073 172567
rect 226191 172449 243913 172567
rect 244031 172449 244073 172567
rect 244191 172449 261913 172567
rect 262031 172449 262073 172567
rect 262191 172449 279913 172567
rect 280031 172449 280073 172567
rect 280191 172449 293151 172567
rect 293269 172449 293311 172567
rect 293429 172449 293445 172567
rect -1483 172433 293445 172449
rect -4363 169307 296325 169323
rect -4363 169189 -3867 169307
rect -3749 169189 -3707 169307
rect -3589 169189 6493 169307
rect 6611 169189 6653 169307
rect 6771 169189 24493 169307
rect 24611 169189 24653 169307
rect 24771 169189 42493 169307
rect 42611 169189 42653 169307
rect 42771 169189 60493 169307
rect 60611 169189 60653 169307
rect 60771 169189 78493 169307
rect 78611 169189 78653 169307
rect 78771 169189 96493 169307
rect 96611 169189 96653 169307
rect 96771 169189 114493 169307
rect 114611 169189 114653 169307
rect 114771 169189 132493 169307
rect 132611 169189 132653 169307
rect 132771 169189 150493 169307
rect 150611 169189 150653 169307
rect 150771 169189 168493 169307
rect 168611 169189 168653 169307
rect 168771 169189 186493 169307
rect 186611 169189 186653 169307
rect 186771 169189 204493 169307
rect 204611 169189 204653 169307
rect 204771 169189 222493 169307
rect 222611 169189 222653 169307
rect 222771 169189 240493 169307
rect 240611 169189 240653 169307
rect 240771 169189 258493 169307
rect 258611 169189 258653 169307
rect 258771 169189 276493 169307
rect 276611 169189 276653 169307
rect 276771 169189 295551 169307
rect 295669 169189 295711 169307
rect 295829 169189 296325 169307
rect -4363 169147 296325 169189
rect -4363 169029 -3867 169147
rect -3749 169029 -3707 169147
rect -3589 169029 6493 169147
rect 6611 169029 6653 169147
rect 6771 169029 24493 169147
rect 24611 169029 24653 169147
rect 24771 169029 42493 169147
rect 42611 169029 42653 169147
rect 42771 169029 60493 169147
rect 60611 169029 60653 169147
rect 60771 169029 78493 169147
rect 78611 169029 78653 169147
rect 78771 169029 96493 169147
rect 96611 169029 96653 169147
rect 96771 169029 114493 169147
rect 114611 169029 114653 169147
rect 114771 169029 132493 169147
rect 132611 169029 132653 169147
rect 132771 169029 150493 169147
rect 150611 169029 150653 169147
rect 150771 169029 168493 169147
rect 168611 169029 168653 169147
rect 168771 169029 186493 169147
rect 186611 169029 186653 169147
rect 186771 169029 204493 169147
rect 204611 169029 204653 169147
rect 204771 169029 222493 169147
rect 222611 169029 222653 169147
rect 222771 169029 240493 169147
rect 240611 169029 240653 169147
rect 240771 169029 258493 169147
rect 258611 169029 258653 169147
rect 258771 169029 276493 169147
rect 276611 169029 276653 169147
rect 276771 169029 295551 169147
rect 295669 169029 295711 169147
rect 295829 169029 296325 169147
rect -4363 169013 296325 169029
rect -3403 167447 295365 167463
rect -3403 167329 -2907 167447
rect -2789 167329 -2747 167447
rect -2629 167329 4633 167447
rect 4751 167329 4793 167447
rect 4911 167329 22633 167447
rect 22751 167329 22793 167447
rect 22911 167329 40633 167447
rect 40751 167329 40793 167447
rect 40911 167329 58633 167447
rect 58751 167329 58793 167447
rect 58911 167329 76633 167447
rect 76751 167329 76793 167447
rect 76911 167329 94633 167447
rect 94751 167329 94793 167447
rect 94911 167329 112633 167447
rect 112751 167329 112793 167447
rect 112911 167329 130633 167447
rect 130751 167329 130793 167447
rect 130911 167329 148633 167447
rect 148751 167329 148793 167447
rect 148911 167329 166633 167447
rect 166751 167329 166793 167447
rect 166911 167329 184633 167447
rect 184751 167329 184793 167447
rect 184911 167329 202633 167447
rect 202751 167329 202793 167447
rect 202911 167329 220633 167447
rect 220751 167329 220793 167447
rect 220911 167329 238633 167447
rect 238751 167329 238793 167447
rect 238911 167329 256633 167447
rect 256751 167329 256793 167447
rect 256911 167329 274633 167447
rect 274751 167329 274793 167447
rect 274911 167329 294591 167447
rect 294709 167329 294751 167447
rect 294869 167329 295365 167447
rect -3403 167287 295365 167329
rect -3403 167169 -2907 167287
rect -2789 167169 -2747 167287
rect -2629 167169 4633 167287
rect 4751 167169 4793 167287
rect 4911 167169 22633 167287
rect 22751 167169 22793 167287
rect 22911 167169 40633 167287
rect 40751 167169 40793 167287
rect 40911 167169 58633 167287
rect 58751 167169 58793 167287
rect 58911 167169 76633 167287
rect 76751 167169 76793 167287
rect 76911 167169 94633 167287
rect 94751 167169 94793 167287
rect 94911 167169 112633 167287
rect 112751 167169 112793 167287
rect 112911 167169 130633 167287
rect 130751 167169 130793 167287
rect 130911 167169 148633 167287
rect 148751 167169 148793 167287
rect 148911 167169 166633 167287
rect 166751 167169 166793 167287
rect 166911 167169 184633 167287
rect 184751 167169 184793 167287
rect 184911 167169 202633 167287
rect 202751 167169 202793 167287
rect 202911 167169 220633 167287
rect 220751 167169 220793 167287
rect 220911 167169 238633 167287
rect 238751 167169 238793 167287
rect 238911 167169 256633 167287
rect 256751 167169 256793 167287
rect 256911 167169 274633 167287
rect 274751 167169 274793 167287
rect 274911 167169 294591 167287
rect 294709 167169 294751 167287
rect 294869 167169 295365 167287
rect -3403 167153 295365 167169
rect -2443 165587 294405 165603
rect -2443 165469 -1947 165587
rect -1829 165469 -1787 165587
rect -1669 165469 2773 165587
rect 2891 165469 2933 165587
rect 3051 165469 20773 165587
rect 20891 165469 20933 165587
rect 21051 165469 38773 165587
rect 38891 165469 38933 165587
rect 39051 165469 56773 165587
rect 56891 165469 56933 165587
rect 57051 165469 74773 165587
rect 74891 165469 74933 165587
rect 75051 165469 92773 165587
rect 92891 165469 92933 165587
rect 93051 165469 110773 165587
rect 110891 165469 110933 165587
rect 111051 165469 128773 165587
rect 128891 165469 128933 165587
rect 129051 165469 146773 165587
rect 146891 165469 146933 165587
rect 147051 165469 164773 165587
rect 164891 165469 164933 165587
rect 165051 165469 182773 165587
rect 182891 165469 182933 165587
rect 183051 165469 200773 165587
rect 200891 165469 200933 165587
rect 201051 165469 218773 165587
rect 218891 165469 218933 165587
rect 219051 165469 236773 165587
rect 236891 165469 236933 165587
rect 237051 165469 254773 165587
rect 254891 165469 254933 165587
rect 255051 165469 272773 165587
rect 272891 165469 272933 165587
rect 273051 165469 290773 165587
rect 290891 165469 290933 165587
rect 291051 165469 293631 165587
rect 293749 165469 293791 165587
rect 293909 165469 294405 165587
rect -2443 165427 294405 165469
rect -2443 165309 -1947 165427
rect -1829 165309 -1787 165427
rect -1669 165309 2773 165427
rect 2891 165309 2933 165427
rect 3051 165309 20773 165427
rect 20891 165309 20933 165427
rect 21051 165309 38773 165427
rect 38891 165309 38933 165427
rect 39051 165309 56773 165427
rect 56891 165309 56933 165427
rect 57051 165309 74773 165427
rect 74891 165309 74933 165427
rect 75051 165309 92773 165427
rect 92891 165309 92933 165427
rect 93051 165309 110773 165427
rect 110891 165309 110933 165427
rect 111051 165309 128773 165427
rect 128891 165309 128933 165427
rect 129051 165309 146773 165427
rect 146891 165309 146933 165427
rect 147051 165309 164773 165427
rect 164891 165309 164933 165427
rect 165051 165309 182773 165427
rect 182891 165309 182933 165427
rect 183051 165309 200773 165427
rect 200891 165309 200933 165427
rect 201051 165309 218773 165427
rect 218891 165309 218933 165427
rect 219051 165309 236773 165427
rect 236891 165309 236933 165427
rect 237051 165309 254773 165427
rect 254891 165309 254933 165427
rect 255051 165309 272773 165427
rect 272891 165309 272933 165427
rect 273051 165309 290773 165427
rect 290891 165309 290933 165427
rect 291051 165309 293631 165427
rect 293749 165309 293791 165427
rect 293909 165309 294405 165427
rect -2443 165293 294405 165309
rect -1483 163727 293445 163743
rect -1483 163609 -987 163727
rect -869 163609 -827 163727
rect -709 163609 913 163727
rect 1031 163609 1073 163727
rect 1191 163609 18913 163727
rect 19031 163609 19073 163727
rect 19191 163609 36913 163727
rect 37031 163609 37073 163727
rect 37191 163609 54913 163727
rect 55031 163609 55073 163727
rect 55191 163609 72913 163727
rect 73031 163609 73073 163727
rect 73191 163609 90913 163727
rect 91031 163609 91073 163727
rect 91191 163609 108913 163727
rect 109031 163609 109073 163727
rect 109191 163609 126913 163727
rect 127031 163609 127073 163727
rect 127191 163609 144913 163727
rect 145031 163609 145073 163727
rect 145191 163609 162913 163727
rect 163031 163609 163073 163727
rect 163191 163609 180913 163727
rect 181031 163609 181073 163727
rect 181191 163609 198913 163727
rect 199031 163609 199073 163727
rect 199191 163609 216913 163727
rect 217031 163609 217073 163727
rect 217191 163609 234913 163727
rect 235031 163609 235073 163727
rect 235191 163609 252913 163727
rect 253031 163609 253073 163727
rect 253191 163609 270913 163727
rect 271031 163609 271073 163727
rect 271191 163609 288913 163727
rect 289031 163609 289073 163727
rect 289191 163609 292671 163727
rect 292789 163609 292831 163727
rect 292949 163609 293445 163727
rect -1483 163567 293445 163609
rect -1483 163449 -987 163567
rect -869 163449 -827 163567
rect -709 163449 913 163567
rect 1031 163449 1073 163567
rect 1191 163449 18913 163567
rect 19031 163449 19073 163567
rect 19191 163449 36913 163567
rect 37031 163449 37073 163567
rect 37191 163449 54913 163567
rect 55031 163449 55073 163567
rect 55191 163449 72913 163567
rect 73031 163449 73073 163567
rect 73191 163449 90913 163567
rect 91031 163449 91073 163567
rect 91191 163449 108913 163567
rect 109031 163449 109073 163567
rect 109191 163449 126913 163567
rect 127031 163449 127073 163567
rect 127191 163449 144913 163567
rect 145031 163449 145073 163567
rect 145191 163449 162913 163567
rect 163031 163449 163073 163567
rect 163191 163449 180913 163567
rect 181031 163449 181073 163567
rect 181191 163449 198913 163567
rect 199031 163449 199073 163567
rect 199191 163449 216913 163567
rect 217031 163449 217073 163567
rect 217191 163449 234913 163567
rect 235031 163449 235073 163567
rect 235191 163449 252913 163567
rect 253031 163449 253073 163567
rect 253191 163449 270913 163567
rect 271031 163449 271073 163567
rect 271191 163449 288913 163567
rect 289031 163449 289073 163567
rect 289191 163449 292671 163567
rect 292789 163449 292831 163567
rect 292949 163449 293445 163567
rect -1483 163433 293445 163449
rect -4363 160307 296325 160323
rect -4363 160189 -4347 160307
rect -4229 160189 -4187 160307
rect -4069 160189 15493 160307
rect 15611 160189 15653 160307
rect 15771 160189 33493 160307
rect 33611 160189 33653 160307
rect 33771 160189 51493 160307
rect 51611 160189 51653 160307
rect 51771 160189 69493 160307
rect 69611 160189 69653 160307
rect 69771 160189 87493 160307
rect 87611 160189 87653 160307
rect 87771 160189 105493 160307
rect 105611 160189 105653 160307
rect 105771 160189 123493 160307
rect 123611 160189 123653 160307
rect 123771 160189 141493 160307
rect 141611 160189 141653 160307
rect 141771 160189 159493 160307
rect 159611 160189 159653 160307
rect 159771 160189 177493 160307
rect 177611 160189 177653 160307
rect 177771 160189 195493 160307
rect 195611 160189 195653 160307
rect 195771 160189 213493 160307
rect 213611 160189 213653 160307
rect 213771 160189 231493 160307
rect 231611 160189 231653 160307
rect 231771 160189 249493 160307
rect 249611 160189 249653 160307
rect 249771 160189 267493 160307
rect 267611 160189 267653 160307
rect 267771 160189 285493 160307
rect 285611 160189 285653 160307
rect 285771 160189 296031 160307
rect 296149 160189 296191 160307
rect 296309 160189 296325 160307
rect -4363 160147 296325 160189
rect -4363 160029 -4347 160147
rect -4229 160029 -4187 160147
rect -4069 160029 15493 160147
rect 15611 160029 15653 160147
rect 15771 160029 33493 160147
rect 33611 160029 33653 160147
rect 33771 160029 51493 160147
rect 51611 160029 51653 160147
rect 51771 160029 69493 160147
rect 69611 160029 69653 160147
rect 69771 160029 87493 160147
rect 87611 160029 87653 160147
rect 87771 160029 105493 160147
rect 105611 160029 105653 160147
rect 105771 160029 123493 160147
rect 123611 160029 123653 160147
rect 123771 160029 141493 160147
rect 141611 160029 141653 160147
rect 141771 160029 159493 160147
rect 159611 160029 159653 160147
rect 159771 160029 177493 160147
rect 177611 160029 177653 160147
rect 177771 160029 195493 160147
rect 195611 160029 195653 160147
rect 195771 160029 213493 160147
rect 213611 160029 213653 160147
rect 213771 160029 231493 160147
rect 231611 160029 231653 160147
rect 231771 160029 249493 160147
rect 249611 160029 249653 160147
rect 249771 160029 267493 160147
rect 267611 160029 267653 160147
rect 267771 160029 285493 160147
rect 285611 160029 285653 160147
rect 285771 160029 296031 160147
rect 296149 160029 296191 160147
rect 296309 160029 296325 160147
rect -4363 160013 296325 160029
rect -3403 158447 295365 158463
rect -3403 158329 -3387 158447
rect -3269 158329 -3227 158447
rect -3109 158329 13633 158447
rect 13751 158329 13793 158447
rect 13911 158329 31633 158447
rect 31751 158329 31793 158447
rect 31911 158329 49633 158447
rect 49751 158329 49793 158447
rect 49911 158329 67633 158447
rect 67751 158329 67793 158447
rect 67911 158329 85633 158447
rect 85751 158329 85793 158447
rect 85911 158329 103633 158447
rect 103751 158329 103793 158447
rect 103911 158329 121633 158447
rect 121751 158329 121793 158447
rect 121911 158329 139633 158447
rect 139751 158329 139793 158447
rect 139911 158329 157633 158447
rect 157751 158329 157793 158447
rect 157911 158329 175633 158447
rect 175751 158329 175793 158447
rect 175911 158329 193633 158447
rect 193751 158329 193793 158447
rect 193911 158329 211633 158447
rect 211751 158329 211793 158447
rect 211911 158329 229633 158447
rect 229751 158329 229793 158447
rect 229911 158329 247633 158447
rect 247751 158329 247793 158447
rect 247911 158329 265633 158447
rect 265751 158329 265793 158447
rect 265911 158329 283633 158447
rect 283751 158329 283793 158447
rect 283911 158329 295071 158447
rect 295189 158329 295231 158447
rect 295349 158329 295365 158447
rect -3403 158287 295365 158329
rect -3403 158169 -3387 158287
rect -3269 158169 -3227 158287
rect -3109 158169 13633 158287
rect 13751 158169 13793 158287
rect 13911 158169 31633 158287
rect 31751 158169 31793 158287
rect 31911 158169 49633 158287
rect 49751 158169 49793 158287
rect 49911 158169 67633 158287
rect 67751 158169 67793 158287
rect 67911 158169 85633 158287
rect 85751 158169 85793 158287
rect 85911 158169 103633 158287
rect 103751 158169 103793 158287
rect 103911 158169 121633 158287
rect 121751 158169 121793 158287
rect 121911 158169 139633 158287
rect 139751 158169 139793 158287
rect 139911 158169 157633 158287
rect 157751 158169 157793 158287
rect 157911 158169 175633 158287
rect 175751 158169 175793 158287
rect 175911 158169 193633 158287
rect 193751 158169 193793 158287
rect 193911 158169 211633 158287
rect 211751 158169 211793 158287
rect 211911 158169 229633 158287
rect 229751 158169 229793 158287
rect 229911 158169 247633 158287
rect 247751 158169 247793 158287
rect 247911 158169 265633 158287
rect 265751 158169 265793 158287
rect 265911 158169 283633 158287
rect 283751 158169 283793 158287
rect 283911 158169 295071 158287
rect 295189 158169 295231 158287
rect 295349 158169 295365 158287
rect -3403 158153 295365 158169
rect -2443 156587 294405 156603
rect -2443 156469 -2427 156587
rect -2309 156469 -2267 156587
rect -2149 156469 11773 156587
rect 11891 156469 11933 156587
rect 12051 156469 29773 156587
rect 29891 156469 29933 156587
rect 30051 156469 47773 156587
rect 47891 156469 47933 156587
rect 48051 156469 65773 156587
rect 65891 156469 65933 156587
rect 66051 156469 83773 156587
rect 83891 156469 83933 156587
rect 84051 156469 101773 156587
rect 101891 156469 101933 156587
rect 102051 156469 119773 156587
rect 119891 156469 119933 156587
rect 120051 156469 137773 156587
rect 137891 156469 137933 156587
rect 138051 156469 155773 156587
rect 155891 156469 155933 156587
rect 156051 156469 173773 156587
rect 173891 156469 173933 156587
rect 174051 156469 191773 156587
rect 191891 156469 191933 156587
rect 192051 156469 209773 156587
rect 209891 156469 209933 156587
rect 210051 156469 227773 156587
rect 227891 156469 227933 156587
rect 228051 156469 245773 156587
rect 245891 156469 245933 156587
rect 246051 156469 263773 156587
rect 263891 156469 263933 156587
rect 264051 156469 281773 156587
rect 281891 156469 281933 156587
rect 282051 156469 294111 156587
rect 294229 156469 294271 156587
rect 294389 156469 294405 156587
rect -2443 156427 294405 156469
rect -2443 156309 -2427 156427
rect -2309 156309 -2267 156427
rect -2149 156309 11773 156427
rect 11891 156309 11933 156427
rect 12051 156309 29773 156427
rect 29891 156309 29933 156427
rect 30051 156309 47773 156427
rect 47891 156309 47933 156427
rect 48051 156309 65773 156427
rect 65891 156309 65933 156427
rect 66051 156309 83773 156427
rect 83891 156309 83933 156427
rect 84051 156309 101773 156427
rect 101891 156309 101933 156427
rect 102051 156309 119773 156427
rect 119891 156309 119933 156427
rect 120051 156309 137773 156427
rect 137891 156309 137933 156427
rect 138051 156309 155773 156427
rect 155891 156309 155933 156427
rect 156051 156309 173773 156427
rect 173891 156309 173933 156427
rect 174051 156309 191773 156427
rect 191891 156309 191933 156427
rect 192051 156309 209773 156427
rect 209891 156309 209933 156427
rect 210051 156309 227773 156427
rect 227891 156309 227933 156427
rect 228051 156309 245773 156427
rect 245891 156309 245933 156427
rect 246051 156309 263773 156427
rect 263891 156309 263933 156427
rect 264051 156309 281773 156427
rect 281891 156309 281933 156427
rect 282051 156309 294111 156427
rect 294229 156309 294271 156427
rect 294389 156309 294405 156427
rect -2443 156293 294405 156309
rect -1483 154727 293445 154743
rect -1483 154609 -1467 154727
rect -1349 154609 -1307 154727
rect -1189 154609 9913 154727
rect 10031 154609 10073 154727
rect 10191 154609 27913 154727
rect 28031 154609 28073 154727
rect 28191 154609 45913 154727
rect 46031 154609 46073 154727
rect 46191 154609 63913 154727
rect 64031 154609 64073 154727
rect 64191 154609 81913 154727
rect 82031 154609 82073 154727
rect 82191 154609 99913 154727
rect 100031 154609 100073 154727
rect 100191 154609 117913 154727
rect 118031 154609 118073 154727
rect 118191 154609 135913 154727
rect 136031 154609 136073 154727
rect 136191 154609 153913 154727
rect 154031 154609 154073 154727
rect 154191 154609 171913 154727
rect 172031 154609 172073 154727
rect 172191 154609 189913 154727
rect 190031 154609 190073 154727
rect 190191 154609 207913 154727
rect 208031 154609 208073 154727
rect 208191 154609 225913 154727
rect 226031 154609 226073 154727
rect 226191 154609 243913 154727
rect 244031 154609 244073 154727
rect 244191 154609 261913 154727
rect 262031 154609 262073 154727
rect 262191 154609 279913 154727
rect 280031 154609 280073 154727
rect 280191 154609 293151 154727
rect 293269 154609 293311 154727
rect 293429 154609 293445 154727
rect -1483 154567 293445 154609
rect -1483 154449 -1467 154567
rect -1349 154449 -1307 154567
rect -1189 154449 9913 154567
rect 10031 154449 10073 154567
rect 10191 154449 27913 154567
rect 28031 154449 28073 154567
rect 28191 154449 45913 154567
rect 46031 154449 46073 154567
rect 46191 154449 63913 154567
rect 64031 154449 64073 154567
rect 64191 154449 81913 154567
rect 82031 154449 82073 154567
rect 82191 154449 99913 154567
rect 100031 154449 100073 154567
rect 100191 154449 117913 154567
rect 118031 154449 118073 154567
rect 118191 154449 135913 154567
rect 136031 154449 136073 154567
rect 136191 154449 153913 154567
rect 154031 154449 154073 154567
rect 154191 154449 171913 154567
rect 172031 154449 172073 154567
rect 172191 154449 189913 154567
rect 190031 154449 190073 154567
rect 190191 154449 207913 154567
rect 208031 154449 208073 154567
rect 208191 154449 225913 154567
rect 226031 154449 226073 154567
rect 226191 154449 243913 154567
rect 244031 154449 244073 154567
rect 244191 154449 261913 154567
rect 262031 154449 262073 154567
rect 262191 154449 279913 154567
rect 280031 154449 280073 154567
rect 280191 154449 293151 154567
rect 293269 154449 293311 154567
rect 293429 154449 293445 154567
rect -1483 154433 293445 154449
rect -4363 151307 296325 151323
rect -4363 151189 -3867 151307
rect -3749 151189 -3707 151307
rect -3589 151189 6493 151307
rect 6611 151189 6653 151307
rect 6771 151189 24493 151307
rect 24611 151189 24653 151307
rect 24771 151189 42493 151307
rect 42611 151189 42653 151307
rect 42771 151189 60493 151307
rect 60611 151189 60653 151307
rect 60771 151189 78493 151307
rect 78611 151189 78653 151307
rect 78771 151189 96493 151307
rect 96611 151189 96653 151307
rect 96771 151189 114493 151307
rect 114611 151189 114653 151307
rect 114771 151189 132493 151307
rect 132611 151189 132653 151307
rect 132771 151189 150493 151307
rect 150611 151189 150653 151307
rect 150771 151189 168493 151307
rect 168611 151189 168653 151307
rect 168771 151189 186493 151307
rect 186611 151189 186653 151307
rect 186771 151189 204493 151307
rect 204611 151189 204653 151307
rect 204771 151189 222493 151307
rect 222611 151189 222653 151307
rect 222771 151189 240493 151307
rect 240611 151189 240653 151307
rect 240771 151189 258493 151307
rect 258611 151189 258653 151307
rect 258771 151189 276493 151307
rect 276611 151189 276653 151307
rect 276771 151189 295551 151307
rect 295669 151189 295711 151307
rect 295829 151189 296325 151307
rect -4363 151147 296325 151189
rect -4363 151029 -3867 151147
rect -3749 151029 -3707 151147
rect -3589 151029 6493 151147
rect 6611 151029 6653 151147
rect 6771 151029 24493 151147
rect 24611 151029 24653 151147
rect 24771 151029 42493 151147
rect 42611 151029 42653 151147
rect 42771 151029 60493 151147
rect 60611 151029 60653 151147
rect 60771 151029 78493 151147
rect 78611 151029 78653 151147
rect 78771 151029 96493 151147
rect 96611 151029 96653 151147
rect 96771 151029 114493 151147
rect 114611 151029 114653 151147
rect 114771 151029 132493 151147
rect 132611 151029 132653 151147
rect 132771 151029 150493 151147
rect 150611 151029 150653 151147
rect 150771 151029 168493 151147
rect 168611 151029 168653 151147
rect 168771 151029 186493 151147
rect 186611 151029 186653 151147
rect 186771 151029 204493 151147
rect 204611 151029 204653 151147
rect 204771 151029 222493 151147
rect 222611 151029 222653 151147
rect 222771 151029 240493 151147
rect 240611 151029 240653 151147
rect 240771 151029 258493 151147
rect 258611 151029 258653 151147
rect 258771 151029 276493 151147
rect 276611 151029 276653 151147
rect 276771 151029 295551 151147
rect 295669 151029 295711 151147
rect 295829 151029 296325 151147
rect -4363 151013 296325 151029
rect -3403 149447 295365 149463
rect -3403 149329 -2907 149447
rect -2789 149329 -2747 149447
rect -2629 149329 4633 149447
rect 4751 149329 4793 149447
rect 4911 149329 22633 149447
rect 22751 149329 22793 149447
rect 22911 149329 40633 149447
rect 40751 149329 40793 149447
rect 40911 149329 58633 149447
rect 58751 149329 58793 149447
rect 58911 149329 76633 149447
rect 76751 149329 76793 149447
rect 76911 149329 94633 149447
rect 94751 149329 94793 149447
rect 94911 149329 112633 149447
rect 112751 149329 112793 149447
rect 112911 149329 130633 149447
rect 130751 149329 130793 149447
rect 130911 149329 148633 149447
rect 148751 149329 148793 149447
rect 148911 149329 166633 149447
rect 166751 149329 166793 149447
rect 166911 149329 184633 149447
rect 184751 149329 184793 149447
rect 184911 149329 202633 149447
rect 202751 149329 202793 149447
rect 202911 149329 220633 149447
rect 220751 149329 220793 149447
rect 220911 149329 238633 149447
rect 238751 149329 238793 149447
rect 238911 149329 256633 149447
rect 256751 149329 256793 149447
rect 256911 149329 274633 149447
rect 274751 149329 274793 149447
rect 274911 149329 294591 149447
rect 294709 149329 294751 149447
rect 294869 149329 295365 149447
rect -3403 149287 295365 149329
rect -3403 149169 -2907 149287
rect -2789 149169 -2747 149287
rect -2629 149169 4633 149287
rect 4751 149169 4793 149287
rect 4911 149169 22633 149287
rect 22751 149169 22793 149287
rect 22911 149169 40633 149287
rect 40751 149169 40793 149287
rect 40911 149169 58633 149287
rect 58751 149169 58793 149287
rect 58911 149169 76633 149287
rect 76751 149169 76793 149287
rect 76911 149169 94633 149287
rect 94751 149169 94793 149287
rect 94911 149169 112633 149287
rect 112751 149169 112793 149287
rect 112911 149169 130633 149287
rect 130751 149169 130793 149287
rect 130911 149169 148633 149287
rect 148751 149169 148793 149287
rect 148911 149169 166633 149287
rect 166751 149169 166793 149287
rect 166911 149169 184633 149287
rect 184751 149169 184793 149287
rect 184911 149169 202633 149287
rect 202751 149169 202793 149287
rect 202911 149169 220633 149287
rect 220751 149169 220793 149287
rect 220911 149169 238633 149287
rect 238751 149169 238793 149287
rect 238911 149169 256633 149287
rect 256751 149169 256793 149287
rect 256911 149169 274633 149287
rect 274751 149169 274793 149287
rect 274911 149169 294591 149287
rect 294709 149169 294751 149287
rect 294869 149169 295365 149287
rect -3403 149153 295365 149169
rect -2443 147587 294405 147603
rect -2443 147469 -1947 147587
rect -1829 147469 -1787 147587
rect -1669 147469 2773 147587
rect 2891 147469 2933 147587
rect 3051 147469 20773 147587
rect 20891 147469 20933 147587
rect 21051 147469 38773 147587
rect 38891 147469 38933 147587
rect 39051 147469 56773 147587
rect 56891 147469 56933 147587
rect 57051 147469 74773 147587
rect 74891 147469 74933 147587
rect 75051 147469 92773 147587
rect 92891 147469 92933 147587
rect 93051 147469 110773 147587
rect 110891 147469 110933 147587
rect 111051 147469 128773 147587
rect 128891 147469 128933 147587
rect 129051 147469 146773 147587
rect 146891 147469 146933 147587
rect 147051 147469 164773 147587
rect 164891 147469 164933 147587
rect 165051 147469 182773 147587
rect 182891 147469 182933 147587
rect 183051 147469 200773 147587
rect 200891 147469 200933 147587
rect 201051 147469 218773 147587
rect 218891 147469 218933 147587
rect 219051 147469 236773 147587
rect 236891 147469 236933 147587
rect 237051 147469 254773 147587
rect 254891 147469 254933 147587
rect 255051 147469 272773 147587
rect 272891 147469 272933 147587
rect 273051 147469 290773 147587
rect 290891 147469 290933 147587
rect 291051 147469 293631 147587
rect 293749 147469 293791 147587
rect 293909 147469 294405 147587
rect -2443 147427 294405 147469
rect -2443 147309 -1947 147427
rect -1829 147309 -1787 147427
rect -1669 147309 2773 147427
rect 2891 147309 2933 147427
rect 3051 147309 20773 147427
rect 20891 147309 20933 147427
rect 21051 147309 38773 147427
rect 38891 147309 38933 147427
rect 39051 147309 56773 147427
rect 56891 147309 56933 147427
rect 57051 147309 74773 147427
rect 74891 147309 74933 147427
rect 75051 147309 92773 147427
rect 92891 147309 92933 147427
rect 93051 147309 110773 147427
rect 110891 147309 110933 147427
rect 111051 147309 128773 147427
rect 128891 147309 128933 147427
rect 129051 147309 146773 147427
rect 146891 147309 146933 147427
rect 147051 147309 164773 147427
rect 164891 147309 164933 147427
rect 165051 147309 182773 147427
rect 182891 147309 182933 147427
rect 183051 147309 200773 147427
rect 200891 147309 200933 147427
rect 201051 147309 218773 147427
rect 218891 147309 218933 147427
rect 219051 147309 236773 147427
rect 236891 147309 236933 147427
rect 237051 147309 254773 147427
rect 254891 147309 254933 147427
rect 255051 147309 272773 147427
rect 272891 147309 272933 147427
rect 273051 147309 290773 147427
rect 290891 147309 290933 147427
rect 291051 147309 293631 147427
rect 293749 147309 293791 147427
rect 293909 147309 294405 147427
rect -2443 147293 294405 147309
rect -1483 145727 293445 145743
rect -1483 145609 -987 145727
rect -869 145609 -827 145727
rect -709 145609 913 145727
rect 1031 145609 1073 145727
rect 1191 145609 18913 145727
rect 19031 145609 19073 145727
rect 19191 145609 36913 145727
rect 37031 145609 37073 145727
rect 37191 145609 54913 145727
rect 55031 145609 55073 145727
rect 55191 145609 72913 145727
rect 73031 145609 73073 145727
rect 73191 145609 90913 145727
rect 91031 145609 91073 145727
rect 91191 145609 108913 145727
rect 109031 145609 109073 145727
rect 109191 145609 126913 145727
rect 127031 145609 127073 145727
rect 127191 145609 144913 145727
rect 145031 145609 145073 145727
rect 145191 145609 162913 145727
rect 163031 145609 163073 145727
rect 163191 145609 180913 145727
rect 181031 145609 181073 145727
rect 181191 145609 198913 145727
rect 199031 145609 199073 145727
rect 199191 145609 216913 145727
rect 217031 145609 217073 145727
rect 217191 145609 234913 145727
rect 235031 145609 235073 145727
rect 235191 145609 252913 145727
rect 253031 145609 253073 145727
rect 253191 145609 270913 145727
rect 271031 145609 271073 145727
rect 271191 145609 288913 145727
rect 289031 145609 289073 145727
rect 289191 145609 292671 145727
rect 292789 145609 292831 145727
rect 292949 145609 293445 145727
rect -1483 145567 293445 145609
rect -1483 145449 -987 145567
rect -869 145449 -827 145567
rect -709 145449 913 145567
rect 1031 145449 1073 145567
rect 1191 145449 18913 145567
rect 19031 145449 19073 145567
rect 19191 145449 36913 145567
rect 37031 145449 37073 145567
rect 37191 145449 54913 145567
rect 55031 145449 55073 145567
rect 55191 145449 72913 145567
rect 73031 145449 73073 145567
rect 73191 145449 90913 145567
rect 91031 145449 91073 145567
rect 91191 145449 108913 145567
rect 109031 145449 109073 145567
rect 109191 145449 126913 145567
rect 127031 145449 127073 145567
rect 127191 145449 144913 145567
rect 145031 145449 145073 145567
rect 145191 145449 162913 145567
rect 163031 145449 163073 145567
rect 163191 145449 180913 145567
rect 181031 145449 181073 145567
rect 181191 145449 198913 145567
rect 199031 145449 199073 145567
rect 199191 145449 216913 145567
rect 217031 145449 217073 145567
rect 217191 145449 234913 145567
rect 235031 145449 235073 145567
rect 235191 145449 252913 145567
rect 253031 145449 253073 145567
rect 253191 145449 270913 145567
rect 271031 145449 271073 145567
rect 271191 145449 288913 145567
rect 289031 145449 289073 145567
rect 289191 145449 292671 145567
rect 292789 145449 292831 145567
rect 292949 145449 293445 145567
rect -1483 145433 293445 145449
rect -4363 142307 296325 142323
rect -4363 142189 -4347 142307
rect -4229 142189 -4187 142307
rect -4069 142189 15493 142307
rect 15611 142189 15653 142307
rect 15771 142189 33493 142307
rect 33611 142189 33653 142307
rect 33771 142189 51493 142307
rect 51611 142189 51653 142307
rect 51771 142189 69493 142307
rect 69611 142189 69653 142307
rect 69771 142189 87493 142307
rect 87611 142189 87653 142307
rect 87771 142189 105493 142307
rect 105611 142189 105653 142307
rect 105771 142189 123493 142307
rect 123611 142189 123653 142307
rect 123771 142189 141493 142307
rect 141611 142189 141653 142307
rect 141771 142189 159493 142307
rect 159611 142189 159653 142307
rect 159771 142189 177493 142307
rect 177611 142189 177653 142307
rect 177771 142189 195493 142307
rect 195611 142189 195653 142307
rect 195771 142189 213493 142307
rect 213611 142189 213653 142307
rect 213771 142189 231493 142307
rect 231611 142189 231653 142307
rect 231771 142189 249493 142307
rect 249611 142189 249653 142307
rect 249771 142189 267493 142307
rect 267611 142189 267653 142307
rect 267771 142189 285493 142307
rect 285611 142189 285653 142307
rect 285771 142189 296031 142307
rect 296149 142189 296191 142307
rect 296309 142189 296325 142307
rect -4363 142147 296325 142189
rect -4363 142029 -4347 142147
rect -4229 142029 -4187 142147
rect -4069 142029 15493 142147
rect 15611 142029 15653 142147
rect 15771 142029 33493 142147
rect 33611 142029 33653 142147
rect 33771 142029 51493 142147
rect 51611 142029 51653 142147
rect 51771 142029 69493 142147
rect 69611 142029 69653 142147
rect 69771 142029 87493 142147
rect 87611 142029 87653 142147
rect 87771 142029 105493 142147
rect 105611 142029 105653 142147
rect 105771 142029 123493 142147
rect 123611 142029 123653 142147
rect 123771 142029 141493 142147
rect 141611 142029 141653 142147
rect 141771 142029 159493 142147
rect 159611 142029 159653 142147
rect 159771 142029 177493 142147
rect 177611 142029 177653 142147
rect 177771 142029 195493 142147
rect 195611 142029 195653 142147
rect 195771 142029 213493 142147
rect 213611 142029 213653 142147
rect 213771 142029 231493 142147
rect 231611 142029 231653 142147
rect 231771 142029 249493 142147
rect 249611 142029 249653 142147
rect 249771 142029 267493 142147
rect 267611 142029 267653 142147
rect 267771 142029 285493 142147
rect 285611 142029 285653 142147
rect 285771 142029 296031 142147
rect 296149 142029 296191 142147
rect 296309 142029 296325 142147
rect -4363 142013 296325 142029
rect -3403 140447 295365 140463
rect -3403 140329 -3387 140447
rect -3269 140329 -3227 140447
rect -3109 140329 13633 140447
rect 13751 140329 13793 140447
rect 13911 140329 31633 140447
rect 31751 140329 31793 140447
rect 31911 140329 49633 140447
rect 49751 140329 49793 140447
rect 49911 140329 67633 140447
rect 67751 140329 67793 140447
rect 67911 140329 85633 140447
rect 85751 140329 85793 140447
rect 85911 140329 103633 140447
rect 103751 140329 103793 140447
rect 103911 140329 121633 140447
rect 121751 140329 121793 140447
rect 121911 140329 139633 140447
rect 139751 140329 139793 140447
rect 139911 140329 157633 140447
rect 157751 140329 157793 140447
rect 157911 140329 175633 140447
rect 175751 140329 175793 140447
rect 175911 140329 193633 140447
rect 193751 140329 193793 140447
rect 193911 140329 211633 140447
rect 211751 140329 211793 140447
rect 211911 140329 229633 140447
rect 229751 140329 229793 140447
rect 229911 140329 247633 140447
rect 247751 140329 247793 140447
rect 247911 140329 265633 140447
rect 265751 140329 265793 140447
rect 265911 140329 283633 140447
rect 283751 140329 283793 140447
rect 283911 140329 295071 140447
rect 295189 140329 295231 140447
rect 295349 140329 295365 140447
rect -3403 140287 295365 140329
rect -3403 140169 -3387 140287
rect -3269 140169 -3227 140287
rect -3109 140169 13633 140287
rect 13751 140169 13793 140287
rect 13911 140169 31633 140287
rect 31751 140169 31793 140287
rect 31911 140169 49633 140287
rect 49751 140169 49793 140287
rect 49911 140169 67633 140287
rect 67751 140169 67793 140287
rect 67911 140169 85633 140287
rect 85751 140169 85793 140287
rect 85911 140169 103633 140287
rect 103751 140169 103793 140287
rect 103911 140169 121633 140287
rect 121751 140169 121793 140287
rect 121911 140169 139633 140287
rect 139751 140169 139793 140287
rect 139911 140169 157633 140287
rect 157751 140169 157793 140287
rect 157911 140169 175633 140287
rect 175751 140169 175793 140287
rect 175911 140169 193633 140287
rect 193751 140169 193793 140287
rect 193911 140169 211633 140287
rect 211751 140169 211793 140287
rect 211911 140169 229633 140287
rect 229751 140169 229793 140287
rect 229911 140169 247633 140287
rect 247751 140169 247793 140287
rect 247911 140169 265633 140287
rect 265751 140169 265793 140287
rect 265911 140169 283633 140287
rect 283751 140169 283793 140287
rect 283911 140169 295071 140287
rect 295189 140169 295231 140287
rect 295349 140169 295365 140287
rect -3403 140153 295365 140169
rect -2443 138587 294405 138603
rect -2443 138469 -2427 138587
rect -2309 138469 -2267 138587
rect -2149 138469 11773 138587
rect 11891 138469 11933 138587
rect 12051 138469 29773 138587
rect 29891 138469 29933 138587
rect 30051 138469 47773 138587
rect 47891 138469 47933 138587
rect 48051 138469 65773 138587
rect 65891 138469 65933 138587
rect 66051 138469 83773 138587
rect 83891 138469 83933 138587
rect 84051 138469 101773 138587
rect 101891 138469 101933 138587
rect 102051 138469 119773 138587
rect 119891 138469 119933 138587
rect 120051 138469 137773 138587
rect 137891 138469 137933 138587
rect 138051 138469 155773 138587
rect 155891 138469 155933 138587
rect 156051 138469 173773 138587
rect 173891 138469 173933 138587
rect 174051 138469 191773 138587
rect 191891 138469 191933 138587
rect 192051 138469 209773 138587
rect 209891 138469 209933 138587
rect 210051 138469 227773 138587
rect 227891 138469 227933 138587
rect 228051 138469 245773 138587
rect 245891 138469 245933 138587
rect 246051 138469 263773 138587
rect 263891 138469 263933 138587
rect 264051 138469 281773 138587
rect 281891 138469 281933 138587
rect 282051 138469 294111 138587
rect 294229 138469 294271 138587
rect 294389 138469 294405 138587
rect -2443 138427 294405 138469
rect -2443 138309 -2427 138427
rect -2309 138309 -2267 138427
rect -2149 138309 11773 138427
rect 11891 138309 11933 138427
rect 12051 138309 29773 138427
rect 29891 138309 29933 138427
rect 30051 138309 47773 138427
rect 47891 138309 47933 138427
rect 48051 138309 65773 138427
rect 65891 138309 65933 138427
rect 66051 138309 83773 138427
rect 83891 138309 83933 138427
rect 84051 138309 101773 138427
rect 101891 138309 101933 138427
rect 102051 138309 119773 138427
rect 119891 138309 119933 138427
rect 120051 138309 137773 138427
rect 137891 138309 137933 138427
rect 138051 138309 155773 138427
rect 155891 138309 155933 138427
rect 156051 138309 173773 138427
rect 173891 138309 173933 138427
rect 174051 138309 191773 138427
rect 191891 138309 191933 138427
rect 192051 138309 209773 138427
rect 209891 138309 209933 138427
rect 210051 138309 227773 138427
rect 227891 138309 227933 138427
rect 228051 138309 245773 138427
rect 245891 138309 245933 138427
rect 246051 138309 263773 138427
rect 263891 138309 263933 138427
rect 264051 138309 281773 138427
rect 281891 138309 281933 138427
rect 282051 138309 294111 138427
rect 294229 138309 294271 138427
rect 294389 138309 294405 138427
rect -2443 138293 294405 138309
rect -1483 136727 293445 136743
rect -1483 136609 -1467 136727
rect -1349 136609 -1307 136727
rect -1189 136609 9913 136727
rect 10031 136609 10073 136727
rect 10191 136609 27913 136727
rect 28031 136609 28073 136727
rect 28191 136609 45913 136727
rect 46031 136609 46073 136727
rect 46191 136609 63913 136727
rect 64031 136609 64073 136727
rect 64191 136609 81913 136727
rect 82031 136609 82073 136727
rect 82191 136609 99913 136727
rect 100031 136609 100073 136727
rect 100191 136609 117913 136727
rect 118031 136609 118073 136727
rect 118191 136609 135913 136727
rect 136031 136609 136073 136727
rect 136191 136609 153913 136727
rect 154031 136609 154073 136727
rect 154191 136609 171913 136727
rect 172031 136609 172073 136727
rect 172191 136609 189913 136727
rect 190031 136609 190073 136727
rect 190191 136609 207913 136727
rect 208031 136609 208073 136727
rect 208191 136609 225913 136727
rect 226031 136609 226073 136727
rect 226191 136609 243913 136727
rect 244031 136609 244073 136727
rect 244191 136609 261913 136727
rect 262031 136609 262073 136727
rect 262191 136609 279913 136727
rect 280031 136609 280073 136727
rect 280191 136609 293151 136727
rect 293269 136609 293311 136727
rect 293429 136609 293445 136727
rect -1483 136567 293445 136609
rect -1483 136449 -1467 136567
rect -1349 136449 -1307 136567
rect -1189 136449 9913 136567
rect 10031 136449 10073 136567
rect 10191 136449 27913 136567
rect 28031 136449 28073 136567
rect 28191 136449 45913 136567
rect 46031 136449 46073 136567
rect 46191 136449 63913 136567
rect 64031 136449 64073 136567
rect 64191 136449 81913 136567
rect 82031 136449 82073 136567
rect 82191 136449 99913 136567
rect 100031 136449 100073 136567
rect 100191 136449 117913 136567
rect 118031 136449 118073 136567
rect 118191 136449 135913 136567
rect 136031 136449 136073 136567
rect 136191 136449 153913 136567
rect 154031 136449 154073 136567
rect 154191 136449 171913 136567
rect 172031 136449 172073 136567
rect 172191 136449 189913 136567
rect 190031 136449 190073 136567
rect 190191 136449 207913 136567
rect 208031 136449 208073 136567
rect 208191 136449 225913 136567
rect 226031 136449 226073 136567
rect 226191 136449 243913 136567
rect 244031 136449 244073 136567
rect 244191 136449 261913 136567
rect 262031 136449 262073 136567
rect 262191 136449 279913 136567
rect 280031 136449 280073 136567
rect 280191 136449 293151 136567
rect 293269 136449 293311 136567
rect 293429 136449 293445 136567
rect -1483 136433 293445 136449
rect -4363 133307 296325 133323
rect -4363 133189 -3867 133307
rect -3749 133189 -3707 133307
rect -3589 133189 6493 133307
rect 6611 133189 6653 133307
rect 6771 133189 24493 133307
rect 24611 133189 24653 133307
rect 24771 133189 42493 133307
rect 42611 133189 42653 133307
rect 42771 133189 60493 133307
rect 60611 133189 60653 133307
rect 60771 133189 78493 133307
rect 78611 133189 78653 133307
rect 78771 133189 96493 133307
rect 96611 133189 96653 133307
rect 96771 133189 114493 133307
rect 114611 133189 114653 133307
rect 114771 133189 132493 133307
rect 132611 133189 132653 133307
rect 132771 133189 150493 133307
rect 150611 133189 150653 133307
rect 150771 133189 168493 133307
rect 168611 133189 168653 133307
rect 168771 133189 186493 133307
rect 186611 133189 186653 133307
rect 186771 133189 204493 133307
rect 204611 133189 204653 133307
rect 204771 133189 222493 133307
rect 222611 133189 222653 133307
rect 222771 133189 240493 133307
rect 240611 133189 240653 133307
rect 240771 133189 258493 133307
rect 258611 133189 258653 133307
rect 258771 133189 276493 133307
rect 276611 133189 276653 133307
rect 276771 133189 295551 133307
rect 295669 133189 295711 133307
rect 295829 133189 296325 133307
rect -4363 133147 296325 133189
rect -4363 133029 -3867 133147
rect -3749 133029 -3707 133147
rect -3589 133029 6493 133147
rect 6611 133029 6653 133147
rect 6771 133029 24493 133147
rect 24611 133029 24653 133147
rect 24771 133029 42493 133147
rect 42611 133029 42653 133147
rect 42771 133029 60493 133147
rect 60611 133029 60653 133147
rect 60771 133029 78493 133147
rect 78611 133029 78653 133147
rect 78771 133029 96493 133147
rect 96611 133029 96653 133147
rect 96771 133029 114493 133147
rect 114611 133029 114653 133147
rect 114771 133029 132493 133147
rect 132611 133029 132653 133147
rect 132771 133029 150493 133147
rect 150611 133029 150653 133147
rect 150771 133029 168493 133147
rect 168611 133029 168653 133147
rect 168771 133029 186493 133147
rect 186611 133029 186653 133147
rect 186771 133029 204493 133147
rect 204611 133029 204653 133147
rect 204771 133029 222493 133147
rect 222611 133029 222653 133147
rect 222771 133029 240493 133147
rect 240611 133029 240653 133147
rect 240771 133029 258493 133147
rect 258611 133029 258653 133147
rect 258771 133029 276493 133147
rect 276611 133029 276653 133147
rect 276771 133029 295551 133147
rect 295669 133029 295711 133147
rect 295829 133029 296325 133147
rect -4363 133013 296325 133029
rect -3403 131447 295365 131463
rect -3403 131329 -2907 131447
rect -2789 131329 -2747 131447
rect -2629 131329 4633 131447
rect 4751 131329 4793 131447
rect 4911 131329 22633 131447
rect 22751 131329 22793 131447
rect 22911 131329 40633 131447
rect 40751 131329 40793 131447
rect 40911 131329 58633 131447
rect 58751 131329 58793 131447
rect 58911 131329 76633 131447
rect 76751 131329 76793 131447
rect 76911 131329 94633 131447
rect 94751 131329 94793 131447
rect 94911 131329 112633 131447
rect 112751 131329 112793 131447
rect 112911 131329 130633 131447
rect 130751 131329 130793 131447
rect 130911 131329 148633 131447
rect 148751 131329 148793 131447
rect 148911 131329 166633 131447
rect 166751 131329 166793 131447
rect 166911 131329 184633 131447
rect 184751 131329 184793 131447
rect 184911 131329 202633 131447
rect 202751 131329 202793 131447
rect 202911 131329 220633 131447
rect 220751 131329 220793 131447
rect 220911 131329 238633 131447
rect 238751 131329 238793 131447
rect 238911 131329 256633 131447
rect 256751 131329 256793 131447
rect 256911 131329 274633 131447
rect 274751 131329 274793 131447
rect 274911 131329 294591 131447
rect 294709 131329 294751 131447
rect 294869 131329 295365 131447
rect -3403 131287 295365 131329
rect -3403 131169 -2907 131287
rect -2789 131169 -2747 131287
rect -2629 131169 4633 131287
rect 4751 131169 4793 131287
rect 4911 131169 22633 131287
rect 22751 131169 22793 131287
rect 22911 131169 40633 131287
rect 40751 131169 40793 131287
rect 40911 131169 58633 131287
rect 58751 131169 58793 131287
rect 58911 131169 76633 131287
rect 76751 131169 76793 131287
rect 76911 131169 94633 131287
rect 94751 131169 94793 131287
rect 94911 131169 112633 131287
rect 112751 131169 112793 131287
rect 112911 131169 130633 131287
rect 130751 131169 130793 131287
rect 130911 131169 148633 131287
rect 148751 131169 148793 131287
rect 148911 131169 166633 131287
rect 166751 131169 166793 131287
rect 166911 131169 184633 131287
rect 184751 131169 184793 131287
rect 184911 131169 202633 131287
rect 202751 131169 202793 131287
rect 202911 131169 220633 131287
rect 220751 131169 220793 131287
rect 220911 131169 238633 131287
rect 238751 131169 238793 131287
rect 238911 131169 256633 131287
rect 256751 131169 256793 131287
rect 256911 131169 274633 131287
rect 274751 131169 274793 131287
rect 274911 131169 294591 131287
rect 294709 131169 294751 131287
rect 294869 131169 295365 131287
rect -3403 131153 295365 131169
rect -2443 129587 294405 129603
rect -2443 129469 -1947 129587
rect -1829 129469 -1787 129587
rect -1669 129469 2773 129587
rect 2891 129469 2933 129587
rect 3051 129469 20773 129587
rect 20891 129469 20933 129587
rect 21051 129469 38773 129587
rect 38891 129469 38933 129587
rect 39051 129469 56773 129587
rect 56891 129469 56933 129587
rect 57051 129469 74773 129587
rect 74891 129469 74933 129587
rect 75051 129469 92773 129587
rect 92891 129469 92933 129587
rect 93051 129469 110773 129587
rect 110891 129469 110933 129587
rect 111051 129469 128773 129587
rect 128891 129469 128933 129587
rect 129051 129469 146773 129587
rect 146891 129469 146933 129587
rect 147051 129469 164773 129587
rect 164891 129469 164933 129587
rect 165051 129469 182773 129587
rect 182891 129469 182933 129587
rect 183051 129469 200773 129587
rect 200891 129469 200933 129587
rect 201051 129469 218773 129587
rect 218891 129469 218933 129587
rect 219051 129469 236773 129587
rect 236891 129469 236933 129587
rect 237051 129469 254773 129587
rect 254891 129469 254933 129587
rect 255051 129469 272773 129587
rect 272891 129469 272933 129587
rect 273051 129469 290773 129587
rect 290891 129469 290933 129587
rect 291051 129469 293631 129587
rect 293749 129469 293791 129587
rect 293909 129469 294405 129587
rect -2443 129427 294405 129469
rect -2443 129309 -1947 129427
rect -1829 129309 -1787 129427
rect -1669 129309 2773 129427
rect 2891 129309 2933 129427
rect 3051 129309 20773 129427
rect 20891 129309 20933 129427
rect 21051 129309 38773 129427
rect 38891 129309 38933 129427
rect 39051 129309 56773 129427
rect 56891 129309 56933 129427
rect 57051 129309 74773 129427
rect 74891 129309 74933 129427
rect 75051 129309 92773 129427
rect 92891 129309 92933 129427
rect 93051 129309 110773 129427
rect 110891 129309 110933 129427
rect 111051 129309 128773 129427
rect 128891 129309 128933 129427
rect 129051 129309 146773 129427
rect 146891 129309 146933 129427
rect 147051 129309 164773 129427
rect 164891 129309 164933 129427
rect 165051 129309 182773 129427
rect 182891 129309 182933 129427
rect 183051 129309 200773 129427
rect 200891 129309 200933 129427
rect 201051 129309 218773 129427
rect 218891 129309 218933 129427
rect 219051 129309 236773 129427
rect 236891 129309 236933 129427
rect 237051 129309 254773 129427
rect 254891 129309 254933 129427
rect 255051 129309 272773 129427
rect 272891 129309 272933 129427
rect 273051 129309 290773 129427
rect 290891 129309 290933 129427
rect 291051 129309 293631 129427
rect 293749 129309 293791 129427
rect 293909 129309 294405 129427
rect -2443 129293 294405 129309
rect -1483 127727 293445 127743
rect -1483 127609 -987 127727
rect -869 127609 -827 127727
rect -709 127609 913 127727
rect 1031 127609 1073 127727
rect 1191 127609 18913 127727
rect 19031 127609 19073 127727
rect 19191 127609 36913 127727
rect 37031 127609 37073 127727
rect 37191 127609 54913 127727
rect 55031 127609 55073 127727
rect 55191 127609 72913 127727
rect 73031 127609 73073 127727
rect 73191 127609 90913 127727
rect 91031 127609 91073 127727
rect 91191 127609 108913 127727
rect 109031 127609 109073 127727
rect 109191 127609 126913 127727
rect 127031 127609 127073 127727
rect 127191 127609 144913 127727
rect 145031 127609 145073 127727
rect 145191 127609 162913 127727
rect 163031 127609 163073 127727
rect 163191 127609 180913 127727
rect 181031 127609 181073 127727
rect 181191 127609 198913 127727
rect 199031 127609 199073 127727
rect 199191 127609 216913 127727
rect 217031 127609 217073 127727
rect 217191 127609 234913 127727
rect 235031 127609 235073 127727
rect 235191 127609 252913 127727
rect 253031 127609 253073 127727
rect 253191 127609 270913 127727
rect 271031 127609 271073 127727
rect 271191 127609 288913 127727
rect 289031 127609 289073 127727
rect 289191 127609 292671 127727
rect 292789 127609 292831 127727
rect 292949 127609 293445 127727
rect -1483 127567 293445 127609
rect -1483 127449 -987 127567
rect -869 127449 -827 127567
rect -709 127449 913 127567
rect 1031 127449 1073 127567
rect 1191 127449 18913 127567
rect 19031 127449 19073 127567
rect 19191 127449 36913 127567
rect 37031 127449 37073 127567
rect 37191 127449 54913 127567
rect 55031 127449 55073 127567
rect 55191 127449 72913 127567
rect 73031 127449 73073 127567
rect 73191 127449 90913 127567
rect 91031 127449 91073 127567
rect 91191 127449 108913 127567
rect 109031 127449 109073 127567
rect 109191 127449 126913 127567
rect 127031 127449 127073 127567
rect 127191 127449 144913 127567
rect 145031 127449 145073 127567
rect 145191 127449 162913 127567
rect 163031 127449 163073 127567
rect 163191 127449 180913 127567
rect 181031 127449 181073 127567
rect 181191 127449 198913 127567
rect 199031 127449 199073 127567
rect 199191 127449 216913 127567
rect 217031 127449 217073 127567
rect 217191 127449 234913 127567
rect 235031 127449 235073 127567
rect 235191 127449 252913 127567
rect 253031 127449 253073 127567
rect 253191 127449 270913 127567
rect 271031 127449 271073 127567
rect 271191 127449 288913 127567
rect 289031 127449 289073 127567
rect 289191 127449 292671 127567
rect 292789 127449 292831 127567
rect 292949 127449 293445 127567
rect -1483 127433 293445 127449
rect -4363 124307 296325 124323
rect -4363 124189 -4347 124307
rect -4229 124189 -4187 124307
rect -4069 124189 15493 124307
rect 15611 124189 15653 124307
rect 15771 124189 33493 124307
rect 33611 124189 33653 124307
rect 33771 124189 51493 124307
rect 51611 124189 51653 124307
rect 51771 124189 69493 124307
rect 69611 124189 69653 124307
rect 69771 124189 87493 124307
rect 87611 124189 87653 124307
rect 87771 124189 105493 124307
rect 105611 124189 105653 124307
rect 105771 124189 123493 124307
rect 123611 124189 123653 124307
rect 123771 124189 141493 124307
rect 141611 124189 141653 124307
rect 141771 124189 159493 124307
rect 159611 124189 159653 124307
rect 159771 124189 177493 124307
rect 177611 124189 177653 124307
rect 177771 124189 195493 124307
rect 195611 124189 195653 124307
rect 195771 124189 213493 124307
rect 213611 124189 213653 124307
rect 213771 124189 231493 124307
rect 231611 124189 231653 124307
rect 231771 124189 249493 124307
rect 249611 124189 249653 124307
rect 249771 124189 267493 124307
rect 267611 124189 267653 124307
rect 267771 124189 285493 124307
rect 285611 124189 285653 124307
rect 285771 124189 296031 124307
rect 296149 124189 296191 124307
rect 296309 124189 296325 124307
rect -4363 124147 296325 124189
rect -4363 124029 -4347 124147
rect -4229 124029 -4187 124147
rect -4069 124029 15493 124147
rect 15611 124029 15653 124147
rect 15771 124029 33493 124147
rect 33611 124029 33653 124147
rect 33771 124029 51493 124147
rect 51611 124029 51653 124147
rect 51771 124029 69493 124147
rect 69611 124029 69653 124147
rect 69771 124029 87493 124147
rect 87611 124029 87653 124147
rect 87771 124029 105493 124147
rect 105611 124029 105653 124147
rect 105771 124029 123493 124147
rect 123611 124029 123653 124147
rect 123771 124029 141493 124147
rect 141611 124029 141653 124147
rect 141771 124029 159493 124147
rect 159611 124029 159653 124147
rect 159771 124029 177493 124147
rect 177611 124029 177653 124147
rect 177771 124029 195493 124147
rect 195611 124029 195653 124147
rect 195771 124029 213493 124147
rect 213611 124029 213653 124147
rect 213771 124029 231493 124147
rect 231611 124029 231653 124147
rect 231771 124029 249493 124147
rect 249611 124029 249653 124147
rect 249771 124029 267493 124147
rect 267611 124029 267653 124147
rect 267771 124029 285493 124147
rect 285611 124029 285653 124147
rect 285771 124029 296031 124147
rect 296149 124029 296191 124147
rect 296309 124029 296325 124147
rect -4363 124013 296325 124029
rect -3403 122447 295365 122463
rect -3403 122329 -3387 122447
rect -3269 122329 -3227 122447
rect -3109 122329 13633 122447
rect 13751 122329 13793 122447
rect 13911 122329 31633 122447
rect 31751 122329 31793 122447
rect 31911 122329 49633 122447
rect 49751 122329 49793 122447
rect 49911 122329 67633 122447
rect 67751 122329 67793 122447
rect 67911 122329 85633 122447
rect 85751 122329 85793 122447
rect 85911 122329 103633 122447
rect 103751 122329 103793 122447
rect 103911 122329 121633 122447
rect 121751 122329 121793 122447
rect 121911 122329 139633 122447
rect 139751 122329 139793 122447
rect 139911 122329 157633 122447
rect 157751 122329 157793 122447
rect 157911 122329 175633 122447
rect 175751 122329 175793 122447
rect 175911 122329 193633 122447
rect 193751 122329 193793 122447
rect 193911 122329 211633 122447
rect 211751 122329 211793 122447
rect 211911 122329 229633 122447
rect 229751 122329 229793 122447
rect 229911 122329 247633 122447
rect 247751 122329 247793 122447
rect 247911 122329 265633 122447
rect 265751 122329 265793 122447
rect 265911 122329 283633 122447
rect 283751 122329 283793 122447
rect 283911 122329 295071 122447
rect 295189 122329 295231 122447
rect 295349 122329 295365 122447
rect -3403 122287 295365 122329
rect -3403 122169 -3387 122287
rect -3269 122169 -3227 122287
rect -3109 122169 13633 122287
rect 13751 122169 13793 122287
rect 13911 122169 31633 122287
rect 31751 122169 31793 122287
rect 31911 122169 49633 122287
rect 49751 122169 49793 122287
rect 49911 122169 67633 122287
rect 67751 122169 67793 122287
rect 67911 122169 85633 122287
rect 85751 122169 85793 122287
rect 85911 122169 103633 122287
rect 103751 122169 103793 122287
rect 103911 122169 121633 122287
rect 121751 122169 121793 122287
rect 121911 122169 139633 122287
rect 139751 122169 139793 122287
rect 139911 122169 157633 122287
rect 157751 122169 157793 122287
rect 157911 122169 175633 122287
rect 175751 122169 175793 122287
rect 175911 122169 193633 122287
rect 193751 122169 193793 122287
rect 193911 122169 211633 122287
rect 211751 122169 211793 122287
rect 211911 122169 229633 122287
rect 229751 122169 229793 122287
rect 229911 122169 247633 122287
rect 247751 122169 247793 122287
rect 247911 122169 265633 122287
rect 265751 122169 265793 122287
rect 265911 122169 283633 122287
rect 283751 122169 283793 122287
rect 283911 122169 295071 122287
rect 295189 122169 295231 122287
rect 295349 122169 295365 122287
rect -3403 122153 295365 122169
rect -2443 120587 294405 120603
rect -2443 120469 -2427 120587
rect -2309 120469 -2267 120587
rect -2149 120469 11773 120587
rect 11891 120469 11933 120587
rect 12051 120469 29773 120587
rect 29891 120469 29933 120587
rect 30051 120469 47773 120587
rect 47891 120469 47933 120587
rect 48051 120469 65773 120587
rect 65891 120469 65933 120587
rect 66051 120469 83773 120587
rect 83891 120469 83933 120587
rect 84051 120469 101773 120587
rect 101891 120469 101933 120587
rect 102051 120469 119773 120587
rect 119891 120469 119933 120587
rect 120051 120469 137773 120587
rect 137891 120469 137933 120587
rect 138051 120469 155773 120587
rect 155891 120469 155933 120587
rect 156051 120469 173773 120587
rect 173891 120469 173933 120587
rect 174051 120469 191773 120587
rect 191891 120469 191933 120587
rect 192051 120469 209773 120587
rect 209891 120469 209933 120587
rect 210051 120469 227773 120587
rect 227891 120469 227933 120587
rect 228051 120469 245773 120587
rect 245891 120469 245933 120587
rect 246051 120469 263773 120587
rect 263891 120469 263933 120587
rect 264051 120469 281773 120587
rect 281891 120469 281933 120587
rect 282051 120469 294111 120587
rect 294229 120469 294271 120587
rect 294389 120469 294405 120587
rect -2443 120427 294405 120469
rect -2443 120309 -2427 120427
rect -2309 120309 -2267 120427
rect -2149 120309 11773 120427
rect 11891 120309 11933 120427
rect 12051 120309 29773 120427
rect 29891 120309 29933 120427
rect 30051 120309 47773 120427
rect 47891 120309 47933 120427
rect 48051 120309 65773 120427
rect 65891 120309 65933 120427
rect 66051 120309 83773 120427
rect 83891 120309 83933 120427
rect 84051 120309 101773 120427
rect 101891 120309 101933 120427
rect 102051 120309 119773 120427
rect 119891 120309 119933 120427
rect 120051 120309 137773 120427
rect 137891 120309 137933 120427
rect 138051 120309 155773 120427
rect 155891 120309 155933 120427
rect 156051 120309 173773 120427
rect 173891 120309 173933 120427
rect 174051 120309 191773 120427
rect 191891 120309 191933 120427
rect 192051 120309 209773 120427
rect 209891 120309 209933 120427
rect 210051 120309 227773 120427
rect 227891 120309 227933 120427
rect 228051 120309 245773 120427
rect 245891 120309 245933 120427
rect 246051 120309 263773 120427
rect 263891 120309 263933 120427
rect 264051 120309 281773 120427
rect 281891 120309 281933 120427
rect 282051 120309 294111 120427
rect 294229 120309 294271 120427
rect 294389 120309 294405 120427
rect -2443 120293 294405 120309
rect -1483 118727 293445 118743
rect -1483 118609 -1467 118727
rect -1349 118609 -1307 118727
rect -1189 118609 9913 118727
rect 10031 118609 10073 118727
rect 10191 118609 27913 118727
rect 28031 118609 28073 118727
rect 28191 118609 45913 118727
rect 46031 118609 46073 118727
rect 46191 118609 63913 118727
rect 64031 118609 64073 118727
rect 64191 118609 81913 118727
rect 82031 118609 82073 118727
rect 82191 118609 99913 118727
rect 100031 118609 100073 118727
rect 100191 118609 117913 118727
rect 118031 118609 118073 118727
rect 118191 118609 135913 118727
rect 136031 118609 136073 118727
rect 136191 118609 153913 118727
rect 154031 118609 154073 118727
rect 154191 118609 171913 118727
rect 172031 118609 172073 118727
rect 172191 118609 189913 118727
rect 190031 118609 190073 118727
rect 190191 118609 207913 118727
rect 208031 118609 208073 118727
rect 208191 118609 225913 118727
rect 226031 118609 226073 118727
rect 226191 118609 243913 118727
rect 244031 118609 244073 118727
rect 244191 118609 261913 118727
rect 262031 118609 262073 118727
rect 262191 118609 279913 118727
rect 280031 118609 280073 118727
rect 280191 118609 293151 118727
rect 293269 118609 293311 118727
rect 293429 118609 293445 118727
rect -1483 118567 293445 118609
rect -1483 118449 -1467 118567
rect -1349 118449 -1307 118567
rect -1189 118449 9913 118567
rect 10031 118449 10073 118567
rect 10191 118449 27913 118567
rect 28031 118449 28073 118567
rect 28191 118449 45913 118567
rect 46031 118449 46073 118567
rect 46191 118449 63913 118567
rect 64031 118449 64073 118567
rect 64191 118449 81913 118567
rect 82031 118449 82073 118567
rect 82191 118449 99913 118567
rect 100031 118449 100073 118567
rect 100191 118449 117913 118567
rect 118031 118449 118073 118567
rect 118191 118449 135913 118567
rect 136031 118449 136073 118567
rect 136191 118449 153913 118567
rect 154031 118449 154073 118567
rect 154191 118449 171913 118567
rect 172031 118449 172073 118567
rect 172191 118449 189913 118567
rect 190031 118449 190073 118567
rect 190191 118449 207913 118567
rect 208031 118449 208073 118567
rect 208191 118449 225913 118567
rect 226031 118449 226073 118567
rect 226191 118449 243913 118567
rect 244031 118449 244073 118567
rect 244191 118449 261913 118567
rect 262031 118449 262073 118567
rect 262191 118449 279913 118567
rect 280031 118449 280073 118567
rect 280191 118449 293151 118567
rect 293269 118449 293311 118567
rect 293429 118449 293445 118567
rect -1483 118433 293445 118449
rect -4363 115307 296325 115323
rect -4363 115189 -3867 115307
rect -3749 115189 -3707 115307
rect -3589 115189 6493 115307
rect 6611 115189 6653 115307
rect 6771 115189 24493 115307
rect 24611 115189 24653 115307
rect 24771 115189 42493 115307
rect 42611 115189 42653 115307
rect 42771 115189 60493 115307
rect 60611 115189 60653 115307
rect 60771 115189 78493 115307
rect 78611 115189 78653 115307
rect 78771 115189 96493 115307
rect 96611 115189 96653 115307
rect 96771 115189 114493 115307
rect 114611 115189 114653 115307
rect 114771 115189 132493 115307
rect 132611 115189 132653 115307
rect 132771 115189 150493 115307
rect 150611 115189 150653 115307
rect 150771 115189 168493 115307
rect 168611 115189 168653 115307
rect 168771 115189 186493 115307
rect 186611 115189 186653 115307
rect 186771 115189 204493 115307
rect 204611 115189 204653 115307
rect 204771 115189 222493 115307
rect 222611 115189 222653 115307
rect 222771 115189 240493 115307
rect 240611 115189 240653 115307
rect 240771 115189 258493 115307
rect 258611 115189 258653 115307
rect 258771 115189 276493 115307
rect 276611 115189 276653 115307
rect 276771 115189 295551 115307
rect 295669 115189 295711 115307
rect 295829 115189 296325 115307
rect -4363 115147 296325 115189
rect -4363 115029 -3867 115147
rect -3749 115029 -3707 115147
rect -3589 115029 6493 115147
rect 6611 115029 6653 115147
rect 6771 115029 24493 115147
rect 24611 115029 24653 115147
rect 24771 115029 42493 115147
rect 42611 115029 42653 115147
rect 42771 115029 60493 115147
rect 60611 115029 60653 115147
rect 60771 115029 78493 115147
rect 78611 115029 78653 115147
rect 78771 115029 96493 115147
rect 96611 115029 96653 115147
rect 96771 115029 114493 115147
rect 114611 115029 114653 115147
rect 114771 115029 132493 115147
rect 132611 115029 132653 115147
rect 132771 115029 150493 115147
rect 150611 115029 150653 115147
rect 150771 115029 168493 115147
rect 168611 115029 168653 115147
rect 168771 115029 186493 115147
rect 186611 115029 186653 115147
rect 186771 115029 204493 115147
rect 204611 115029 204653 115147
rect 204771 115029 222493 115147
rect 222611 115029 222653 115147
rect 222771 115029 240493 115147
rect 240611 115029 240653 115147
rect 240771 115029 258493 115147
rect 258611 115029 258653 115147
rect 258771 115029 276493 115147
rect 276611 115029 276653 115147
rect 276771 115029 295551 115147
rect 295669 115029 295711 115147
rect 295829 115029 296325 115147
rect -4363 115013 296325 115029
rect -3403 113447 295365 113463
rect -3403 113329 -2907 113447
rect -2789 113329 -2747 113447
rect -2629 113329 4633 113447
rect 4751 113329 4793 113447
rect 4911 113329 22633 113447
rect 22751 113329 22793 113447
rect 22911 113329 40633 113447
rect 40751 113329 40793 113447
rect 40911 113329 58633 113447
rect 58751 113329 58793 113447
rect 58911 113329 76633 113447
rect 76751 113329 76793 113447
rect 76911 113329 94633 113447
rect 94751 113329 94793 113447
rect 94911 113329 112633 113447
rect 112751 113329 112793 113447
rect 112911 113329 130633 113447
rect 130751 113329 130793 113447
rect 130911 113329 148633 113447
rect 148751 113329 148793 113447
rect 148911 113329 166633 113447
rect 166751 113329 166793 113447
rect 166911 113329 184633 113447
rect 184751 113329 184793 113447
rect 184911 113329 202633 113447
rect 202751 113329 202793 113447
rect 202911 113329 220633 113447
rect 220751 113329 220793 113447
rect 220911 113329 238633 113447
rect 238751 113329 238793 113447
rect 238911 113329 256633 113447
rect 256751 113329 256793 113447
rect 256911 113329 274633 113447
rect 274751 113329 274793 113447
rect 274911 113329 294591 113447
rect 294709 113329 294751 113447
rect 294869 113329 295365 113447
rect -3403 113287 295365 113329
rect -3403 113169 -2907 113287
rect -2789 113169 -2747 113287
rect -2629 113169 4633 113287
rect 4751 113169 4793 113287
rect 4911 113169 22633 113287
rect 22751 113169 22793 113287
rect 22911 113169 40633 113287
rect 40751 113169 40793 113287
rect 40911 113169 58633 113287
rect 58751 113169 58793 113287
rect 58911 113169 76633 113287
rect 76751 113169 76793 113287
rect 76911 113169 94633 113287
rect 94751 113169 94793 113287
rect 94911 113169 112633 113287
rect 112751 113169 112793 113287
rect 112911 113169 130633 113287
rect 130751 113169 130793 113287
rect 130911 113169 148633 113287
rect 148751 113169 148793 113287
rect 148911 113169 166633 113287
rect 166751 113169 166793 113287
rect 166911 113169 184633 113287
rect 184751 113169 184793 113287
rect 184911 113169 202633 113287
rect 202751 113169 202793 113287
rect 202911 113169 220633 113287
rect 220751 113169 220793 113287
rect 220911 113169 238633 113287
rect 238751 113169 238793 113287
rect 238911 113169 256633 113287
rect 256751 113169 256793 113287
rect 256911 113169 274633 113287
rect 274751 113169 274793 113287
rect 274911 113169 294591 113287
rect 294709 113169 294751 113287
rect 294869 113169 295365 113287
rect -3403 113153 295365 113169
rect -2443 111587 294405 111603
rect -2443 111469 -1947 111587
rect -1829 111469 -1787 111587
rect -1669 111469 2773 111587
rect 2891 111469 2933 111587
rect 3051 111469 20773 111587
rect 20891 111469 20933 111587
rect 21051 111469 38773 111587
rect 38891 111469 38933 111587
rect 39051 111469 56773 111587
rect 56891 111469 56933 111587
rect 57051 111469 74773 111587
rect 74891 111469 74933 111587
rect 75051 111469 92773 111587
rect 92891 111469 92933 111587
rect 93051 111469 110773 111587
rect 110891 111469 110933 111587
rect 111051 111469 128773 111587
rect 128891 111469 128933 111587
rect 129051 111469 146773 111587
rect 146891 111469 146933 111587
rect 147051 111469 164773 111587
rect 164891 111469 164933 111587
rect 165051 111469 182773 111587
rect 182891 111469 182933 111587
rect 183051 111469 200773 111587
rect 200891 111469 200933 111587
rect 201051 111469 218773 111587
rect 218891 111469 218933 111587
rect 219051 111469 236773 111587
rect 236891 111469 236933 111587
rect 237051 111469 254773 111587
rect 254891 111469 254933 111587
rect 255051 111469 272773 111587
rect 272891 111469 272933 111587
rect 273051 111469 290773 111587
rect 290891 111469 290933 111587
rect 291051 111469 293631 111587
rect 293749 111469 293791 111587
rect 293909 111469 294405 111587
rect -2443 111427 294405 111469
rect -2443 111309 -1947 111427
rect -1829 111309 -1787 111427
rect -1669 111309 2773 111427
rect 2891 111309 2933 111427
rect 3051 111309 20773 111427
rect 20891 111309 20933 111427
rect 21051 111309 38773 111427
rect 38891 111309 38933 111427
rect 39051 111309 56773 111427
rect 56891 111309 56933 111427
rect 57051 111309 74773 111427
rect 74891 111309 74933 111427
rect 75051 111309 92773 111427
rect 92891 111309 92933 111427
rect 93051 111309 110773 111427
rect 110891 111309 110933 111427
rect 111051 111309 128773 111427
rect 128891 111309 128933 111427
rect 129051 111309 146773 111427
rect 146891 111309 146933 111427
rect 147051 111309 164773 111427
rect 164891 111309 164933 111427
rect 165051 111309 182773 111427
rect 182891 111309 182933 111427
rect 183051 111309 200773 111427
rect 200891 111309 200933 111427
rect 201051 111309 218773 111427
rect 218891 111309 218933 111427
rect 219051 111309 236773 111427
rect 236891 111309 236933 111427
rect 237051 111309 254773 111427
rect 254891 111309 254933 111427
rect 255051 111309 272773 111427
rect 272891 111309 272933 111427
rect 273051 111309 290773 111427
rect 290891 111309 290933 111427
rect 291051 111309 293631 111427
rect 293749 111309 293791 111427
rect 293909 111309 294405 111427
rect -2443 111293 294405 111309
rect -1483 109727 293445 109743
rect -1483 109609 -987 109727
rect -869 109609 -827 109727
rect -709 109609 913 109727
rect 1031 109609 1073 109727
rect 1191 109609 18913 109727
rect 19031 109609 19073 109727
rect 19191 109609 36913 109727
rect 37031 109609 37073 109727
rect 37191 109609 54913 109727
rect 55031 109609 55073 109727
rect 55191 109609 72913 109727
rect 73031 109609 73073 109727
rect 73191 109609 90913 109727
rect 91031 109609 91073 109727
rect 91191 109609 108913 109727
rect 109031 109609 109073 109727
rect 109191 109609 126913 109727
rect 127031 109609 127073 109727
rect 127191 109609 144913 109727
rect 145031 109609 145073 109727
rect 145191 109609 162913 109727
rect 163031 109609 163073 109727
rect 163191 109609 180913 109727
rect 181031 109609 181073 109727
rect 181191 109609 198913 109727
rect 199031 109609 199073 109727
rect 199191 109609 216913 109727
rect 217031 109609 217073 109727
rect 217191 109609 234913 109727
rect 235031 109609 235073 109727
rect 235191 109609 252913 109727
rect 253031 109609 253073 109727
rect 253191 109609 270913 109727
rect 271031 109609 271073 109727
rect 271191 109609 288913 109727
rect 289031 109609 289073 109727
rect 289191 109609 292671 109727
rect 292789 109609 292831 109727
rect 292949 109609 293445 109727
rect -1483 109567 293445 109609
rect -1483 109449 -987 109567
rect -869 109449 -827 109567
rect -709 109449 913 109567
rect 1031 109449 1073 109567
rect 1191 109449 18913 109567
rect 19031 109449 19073 109567
rect 19191 109449 36913 109567
rect 37031 109449 37073 109567
rect 37191 109449 54913 109567
rect 55031 109449 55073 109567
rect 55191 109449 72913 109567
rect 73031 109449 73073 109567
rect 73191 109449 90913 109567
rect 91031 109449 91073 109567
rect 91191 109449 108913 109567
rect 109031 109449 109073 109567
rect 109191 109449 126913 109567
rect 127031 109449 127073 109567
rect 127191 109449 144913 109567
rect 145031 109449 145073 109567
rect 145191 109449 162913 109567
rect 163031 109449 163073 109567
rect 163191 109449 180913 109567
rect 181031 109449 181073 109567
rect 181191 109449 198913 109567
rect 199031 109449 199073 109567
rect 199191 109449 216913 109567
rect 217031 109449 217073 109567
rect 217191 109449 234913 109567
rect 235031 109449 235073 109567
rect 235191 109449 252913 109567
rect 253031 109449 253073 109567
rect 253191 109449 270913 109567
rect 271031 109449 271073 109567
rect 271191 109449 288913 109567
rect 289031 109449 289073 109567
rect 289191 109449 292671 109567
rect 292789 109449 292831 109567
rect 292949 109449 293445 109567
rect -1483 109433 293445 109449
rect -4363 106307 296325 106323
rect -4363 106189 -4347 106307
rect -4229 106189 -4187 106307
rect -4069 106189 15493 106307
rect 15611 106189 15653 106307
rect 15771 106189 33493 106307
rect 33611 106189 33653 106307
rect 33771 106189 51493 106307
rect 51611 106189 51653 106307
rect 51771 106189 69493 106307
rect 69611 106189 69653 106307
rect 69771 106189 87493 106307
rect 87611 106189 87653 106307
rect 87771 106189 105493 106307
rect 105611 106189 105653 106307
rect 105771 106189 123493 106307
rect 123611 106189 123653 106307
rect 123771 106189 141493 106307
rect 141611 106189 141653 106307
rect 141771 106189 159493 106307
rect 159611 106189 159653 106307
rect 159771 106189 177493 106307
rect 177611 106189 177653 106307
rect 177771 106189 195493 106307
rect 195611 106189 195653 106307
rect 195771 106189 213493 106307
rect 213611 106189 213653 106307
rect 213771 106189 231493 106307
rect 231611 106189 231653 106307
rect 231771 106189 249493 106307
rect 249611 106189 249653 106307
rect 249771 106189 267493 106307
rect 267611 106189 267653 106307
rect 267771 106189 285493 106307
rect 285611 106189 285653 106307
rect 285771 106189 296031 106307
rect 296149 106189 296191 106307
rect 296309 106189 296325 106307
rect -4363 106147 296325 106189
rect -4363 106029 -4347 106147
rect -4229 106029 -4187 106147
rect -4069 106029 15493 106147
rect 15611 106029 15653 106147
rect 15771 106029 33493 106147
rect 33611 106029 33653 106147
rect 33771 106029 51493 106147
rect 51611 106029 51653 106147
rect 51771 106029 69493 106147
rect 69611 106029 69653 106147
rect 69771 106029 87493 106147
rect 87611 106029 87653 106147
rect 87771 106029 105493 106147
rect 105611 106029 105653 106147
rect 105771 106029 123493 106147
rect 123611 106029 123653 106147
rect 123771 106029 141493 106147
rect 141611 106029 141653 106147
rect 141771 106029 159493 106147
rect 159611 106029 159653 106147
rect 159771 106029 177493 106147
rect 177611 106029 177653 106147
rect 177771 106029 195493 106147
rect 195611 106029 195653 106147
rect 195771 106029 213493 106147
rect 213611 106029 213653 106147
rect 213771 106029 231493 106147
rect 231611 106029 231653 106147
rect 231771 106029 249493 106147
rect 249611 106029 249653 106147
rect 249771 106029 267493 106147
rect 267611 106029 267653 106147
rect 267771 106029 285493 106147
rect 285611 106029 285653 106147
rect 285771 106029 296031 106147
rect 296149 106029 296191 106147
rect 296309 106029 296325 106147
rect -4363 106013 296325 106029
rect -3403 104447 295365 104463
rect -3403 104329 -3387 104447
rect -3269 104329 -3227 104447
rect -3109 104329 13633 104447
rect 13751 104329 13793 104447
rect 13911 104329 31633 104447
rect 31751 104329 31793 104447
rect 31911 104329 49633 104447
rect 49751 104329 49793 104447
rect 49911 104329 67633 104447
rect 67751 104329 67793 104447
rect 67911 104329 85633 104447
rect 85751 104329 85793 104447
rect 85911 104329 103633 104447
rect 103751 104329 103793 104447
rect 103911 104329 121633 104447
rect 121751 104329 121793 104447
rect 121911 104329 139633 104447
rect 139751 104329 139793 104447
rect 139911 104329 157633 104447
rect 157751 104329 157793 104447
rect 157911 104329 175633 104447
rect 175751 104329 175793 104447
rect 175911 104329 193633 104447
rect 193751 104329 193793 104447
rect 193911 104329 211633 104447
rect 211751 104329 211793 104447
rect 211911 104329 229633 104447
rect 229751 104329 229793 104447
rect 229911 104329 247633 104447
rect 247751 104329 247793 104447
rect 247911 104329 265633 104447
rect 265751 104329 265793 104447
rect 265911 104329 283633 104447
rect 283751 104329 283793 104447
rect 283911 104329 295071 104447
rect 295189 104329 295231 104447
rect 295349 104329 295365 104447
rect -3403 104287 295365 104329
rect -3403 104169 -3387 104287
rect -3269 104169 -3227 104287
rect -3109 104169 13633 104287
rect 13751 104169 13793 104287
rect 13911 104169 31633 104287
rect 31751 104169 31793 104287
rect 31911 104169 49633 104287
rect 49751 104169 49793 104287
rect 49911 104169 67633 104287
rect 67751 104169 67793 104287
rect 67911 104169 85633 104287
rect 85751 104169 85793 104287
rect 85911 104169 103633 104287
rect 103751 104169 103793 104287
rect 103911 104169 121633 104287
rect 121751 104169 121793 104287
rect 121911 104169 139633 104287
rect 139751 104169 139793 104287
rect 139911 104169 157633 104287
rect 157751 104169 157793 104287
rect 157911 104169 175633 104287
rect 175751 104169 175793 104287
rect 175911 104169 193633 104287
rect 193751 104169 193793 104287
rect 193911 104169 211633 104287
rect 211751 104169 211793 104287
rect 211911 104169 229633 104287
rect 229751 104169 229793 104287
rect 229911 104169 247633 104287
rect 247751 104169 247793 104287
rect 247911 104169 265633 104287
rect 265751 104169 265793 104287
rect 265911 104169 283633 104287
rect 283751 104169 283793 104287
rect 283911 104169 295071 104287
rect 295189 104169 295231 104287
rect 295349 104169 295365 104287
rect -3403 104153 295365 104169
rect -2443 102587 294405 102603
rect -2443 102469 -2427 102587
rect -2309 102469 -2267 102587
rect -2149 102469 11773 102587
rect 11891 102469 11933 102587
rect 12051 102469 29773 102587
rect 29891 102469 29933 102587
rect 30051 102469 47773 102587
rect 47891 102469 47933 102587
rect 48051 102469 65773 102587
rect 65891 102469 65933 102587
rect 66051 102469 83773 102587
rect 83891 102469 83933 102587
rect 84051 102469 101773 102587
rect 101891 102469 101933 102587
rect 102051 102469 119773 102587
rect 119891 102469 119933 102587
rect 120051 102469 137773 102587
rect 137891 102469 137933 102587
rect 138051 102469 155773 102587
rect 155891 102469 155933 102587
rect 156051 102469 173773 102587
rect 173891 102469 173933 102587
rect 174051 102469 191773 102587
rect 191891 102469 191933 102587
rect 192051 102469 209773 102587
rect 209891 102469 209933 102587
rect 210051 102469 227773 102587
rect 227891 102469 227933 102587
rect 228051 102469 245773 102587
rect 245891 102469 245933 102587
rect 246051 102469 263773 102587
rect 263891 102469 263933 102587
rect 264051 102469 281773 102587
rect 281891 102469 281933 102587
rect 282051 102469 294111 102587
rect 294229 102469 294271 102587
rect 294389 102469 294405 102587
rect -2443 102427 294405 102469
rect -2443 102309 -2427 102427
rect -2309 102309 -2267 102427
rect -2149 102309 11773 102427
rect 11891 102309 11933 102427
rect 12051 102309 29773 102427
rect 29891 102309 29933 102427
rect 30051 102309 47773 102427
rect 47891 102309 47933 102427
rect 48051 102309 65773 102427
rect 65891 102309 65933 102427
rect 66051 102309 83773 102427
rect 83891 102309 83933 102427
rect 84051 102309 101773 102427
rect 101891 102309 101933 102427
rect 102051 102309 119773 102427
rect 119891 102309 119933 102427
rect 120051 102309 137773 102427
rect 137891 102309 137933 102427
rect 138051 102309 155773 102427
rect 155891 102309 155933 102427
rect 156051 102309 173773 102427
rect 173891 102309 173933 102427
rect 174051 102309 191773 102427
rect 191891 102309 191933 102427
rect 192051 102309 209773 102427
rect 209891 102309 209933 102427
rect 210051 102309 227773 102427
rect 227891 102309 227933 102427
rect 228051 102309 245773 102427
rect 245891 102309 245933 102427
rect 246051 102309 263773 102427
rect 263891 102309 263933 102427
rect 264051 102309 281773 102427
rect 281891 102309 281933 102427
rect 282051 102309 294111 102427
rect 294229 102309 294271 102427
rect 294389 102309 294405 102427
rect -2443 102293 294405 102309
rect -1483 100727 293445 100743
rect -1483 100609 -1467 100727
rect -1349 100609 -1307 100727
rect -1189 100609 9913 100727
rect 10031 100609 10073 100727
rect 10191 100609 27913 100727
rect 28031 100609 28073 100727
rect 28191 100609 45913 100727
rect 46031 100609 46073 100727
rect 46191 100609 63913 100727
rect 64031 100609 64073 100727
rect 64191 100609 81913 100727
rect 82031 100609 82073 100727
rect 82191 100609 99913 100727
rect 100031 100609 100073 100727
rect 100191 100609 117913 100727
rect 118031 100609 118073 100727
rect 118191 100609 135913 100727
rect 136031 100609 136073 100727
rect 136191 100609 153913 100727
rect 154031 100609 154073 100727
rect 154191 100609 171913 100727
rect 172031 100609 172073 100727
rect 172191 100609 189913 100727
rect 190031 100609 190073 100727
rect 190191 100609 207913 100727
rect 208031 100609 208073 100727
rect 208191 100609 225913 100727
rect 226031 100609 226073 100727
rect 226191 100609 243913 100727
rect 244031 100609 244073 100727
rect 244191 100609 261913 100727
rect 262031 100609 262073 100727
rect 262191 100609 279913 100727
rect 280031 100609 280073 100727
rect 280191 100609 293151 100727
rect 293269 100609 293311 100727
rect 293429 100609 293445 100727
rect -1483 100567 293445 100609
rect -1483 100449 -1467 100567
rect -1349 100449 -1307 100567
rect -1189 100449 9913 100567
rect 10031 100449 10073 100567
rect 10191 100449 27913 100567
rect 28031 100449 28073 100567
rect 28191 100449 45913 100567
rect 46031 100449 46073 100567
rect 46191 100449 63913 100567
rect 64031 100449 64073 100567
rect 64191 100449 81913 100567
rect 82031 100449 82073 100567
rect 82191 100449 99913 100567
rect 100031 100449 100073 100567
rect 100191 100449 117913 100567
rect 118031 100449 118073 100567
rect 118191 100449 135913 100567
rect 136031 100449 136073 100567
rect 136191 100449 153913 100567
rect 154031 100449 154073 100567
rect 154191 100449 171913 100567
rect 172031 100449 172073 100567
rect 172191 100449 189913 100567
rect 190031 100449 190073 100567
rect 190191 100449 207913 100567
rect 208031 100449 208073 100567
rect 208191 100449 225913 100567
rect 226031 100449 226073 100567
rect 226191 100449 243913 100567
rect 244031 100449 244073 100567
rect 244191 100449 261913 100567
rect 262031 100449 262073 100567
rect 262191 100449 279913 100567
rect 280031 100449 280073 100567
rect 280191 100449 293151 100567
rect 293269 100449 293311 100567
rect 293429 100449 293445 100567
rect -1483 100433 293445 100449
rect -4363 97307 296325 97323
rect -4363 97189 -3867 97307
rect -3749 97189 -3707 97307
rect -3589 97189 6493 97307
rect 6611 97189 6653 97307
rect 6771 97189 24493 97307
rect 24611 97189 24653 97307
rect 24771 97189 42493 97307
rect 42611 97189 42653 97307
rect 42771 97189 60493 97307
rect 60611 97189 60653 97307
rect 60771 97189 78493 97307
rect 78611 97189 78653 97307
rect 78771 97189 96493 97307
rect 96611 97189 96653 97307
rect 96771 97189 114493 97307
rect 114611 97189 114653 97307
rect 114771 97189 132493 97307
rect 132611 97189 132653 97307
rect 132771 97189 150493 97307
rect 150611 97189 150653 97307
rect 150771 97189 168493 97307
rect 168611 97189 168653 97307
rect 168771 97189 186493 97307
rect 186611 97189 186653 97307
rect 186771 97189 204493 97307
rect 204611 97189 204653 97307
rect 204771 97189 222493 97307
rect 222611 97189 222653 97307
rect 222771 97189 240493 97307
rect 240611 97189 240653 97307
rect 240771 97189 258493 97307
rect 258611 97189 258653 97307
rect 258771 97189 276493 97307
rect 276611 97189 276653 97307
rect 276771 97189 295551 97307
rect 295669 97189 295711 97307
rect 295829 97189 296325 97307
rect -4363 97147 296325 97189
rect -4363 97029 -3867 97147
rect -3749 97029 -3707 97147
rect -3589 97029 6493 97147
rect 6611 97029 6653 97147
rect 6771 97029 24493 97147
rect 24611 97029 24653 97147
rect 24771 97029 42493 97147
rect 42611 97029 42653 97147
rect 42771 97029 60493 97147
rect 60611 97029 60653 97147
rect 60771 97029 78493 97147
rect 78611 97029 78653 97147
rect 78771 97029 96493 97147
rect 96611 97029 96653 97147
rect 96771 97029 114493 97147
rect 114611 97029 114653 97147
rect 114771 97029 132493 97147
rect 132611 97029 132653 97147
rect 132771 97029 150493 97147
rect 150611 97029 150653 97147
rect 150771 97029 168493 97147
rect 168611 97029 168653 97147
rect 168771 97029 186493 97147
rect 186611 97029 186653 97147
rect 186771 97029 204493 97147
rect 204611 97029 204653 97147
rect 204771 97029 222493 97147
rect 222611 97029 222653 97147
rect 222771 97029 240493 97147
rect 240611 97029 240653 97147
rect 240771 97029 258493 97147
rect 258611 97029 258653 97147
rect 258771 97029 276493 97147
rect 276611 97029 276653 97147
rect 276771 97029 295551 97147
rect 295669 97029 295711 97147
rect 295829 97029 296325 97147
rect -4363 97013 296325 97029
rect -3403 95447 295365 95463
rect -3403 95329 -2907 95447
rect -2789 95329 -2747 95447
rect -2629 95329 4633 95447
rect 4751 95329 4793 95447
rect 4911 95329 22633 95447
rect 22751 95329 22793 95447
rect 22911 95329 40633 95447
rect 40751 95329 40793 95447
rect 40911 95329 58633 95447
rect 58751 95329 58793 95447
rect 58911 95329 76633 95447
rect 76751 95329 76793 95447
rect 76911 95329 94633 95447
rect 94751 95329 94793 95447
rect 94911 95329 112633 95447
rect 112751 95329 112793 95447
rect 112911 95329 130633 95447
rect 130751 95329 130793 95447
rect 130911 95329 148633 95447
rect 148751 95329 148793 95447
rect 148911 95329 166633 95447
rect 166751 95329 166793 95447
rect 166911 95329 184633 95447
rect 184751 95329 184793 95447
rect 184911 95329 202633 95447
rect 202751 95329 202793 95447
rect 202911 95329 220633 95447
rect 220751 95329 220793 95447
rect 220911 95329 238633 95447
rect 238751 95329 238793 95447
rect 238911 95329 256633 95447
rect 256751 95329 256793 95447
rect 256911 95329 274633 95447
rect 274751 95329 274793 95447
rect 274911 95329 294591 95447
rect 294709 95329 294751 95447
rect 294869 95329 295365 95447
rect -3403 95287 295365 95329
rect -3403 95169 -2907 95287
rect -2789 95169 -2747 95287
rect -2629 95169 4633 95287
rect 4751 95169 4793 95287
rect 4911 95169 22633 95287
rect 22751 95169 22793 95287
rect 22911 95169 40633 95287
rect 40751 95169 40793 95287
rect 40911 95169 58633 95287
rect 58751 95169 58793 95287
rect 58911 95169 76633 95287
rect 76751 95169 76793 95287
rect 76911 95169 94633 95287
rect 94751 95169 94793 95287
rect 94911 95169 112633 95287
rect 112751 95169 112793 95287
rect 112911 95169 130633 95287
rect 130751 95169 130793 95287
rect 130911 95169 148633 95287
rect 148751 95169 148793 95287
rect 148911 95169 166633 95287
rect 166751 95169 166793 95287
rect 166911 95169 184633 95287
rect 184751 95169 184793 95287
rect 184911 95169 202633 95287
rect 202751 95169 202793 95287
rect 202911 95169 220633 95287
rect 220751 95169 220793 95287
rect 220911 95169 238633 95287
rect 238751 95169 238793 95287
rect 238911 95169 256633 95287
rect 256751 95169 256793 95287
rect 256911 95169 274633 95287
rect 274751 95169 274793 95287
rect 274911 95169 294591 95287
rect 294709 95169 294751 95287
rect 294869 95169 295365 95287
rect -3403 95153 295365 95169
rect -2443 93587 294405 93603
rect -2443 93469 -1947 93587
rect -1829 93469 -1787 93587
rect -1669 93469 2773 93587
rect 2891 93469 2933 93587
rect 3051 93469 20773 93587
rect 20891 93469 20933 93587
rect 21051 93469 38773 93587
rect 38891 93469 38933 93587
rect 39051 93469 56773 93587
rect 56891 93469 56933 93587
rect 57051 93469 74773 93587
rect 74891 93469 74933 93587
rect 75051 93469 92773 93587
rect 92891 93469 92933 93587
rect 93051 93469 110773 93587
rect 110891 93469 110933 93587
rect 111051 93469 128773 93587
rect 128891 93469 128933 93587
rect 129051 93469 146773 93587
rect 146891 93469 146933 93587
rect 147051 93469 164773 93587
rect 164891 93469 164933 93587
rect 165051 93469 182773 93587
rect 182891 93469 182933 93587
rect 183051 93469 200773 93587
rect 200891 93469 200933 93587
rect 201051 93469 218773 93587
rect 218891 93469 218933 93587
rect 219051 93469 236773 93587
rect 236891 93469 236933 93587
rect 237051 93469 254773 93587
rect 254891 93469 254933 93587
rect 255051 93469 272773 93587
rect 272891 93469 272933 93587
rect 273051 93469 290773 93587
rect 290891 93469 290933 93587
rect 291051 93469 293631 93587
rect 293749 93469 293791 93587
rect 293909 93469 294405 93587
rect -2443 93427 294405 93469
rect -2443 93309 -1947 93427
rect -1829 93309 -1787 93427
rect -1669 93309 2773 93427
rect 2891 93309 2933 93427
rect 3051 93309 20773 93427
rect 20891 93309 20933 93427
rect 21051 93309 38773 93427
rect 38891 93309 38933 93427
rect 39051 93309 56773 93427
rect 56891 93309 56933 93427
rect 57051 93309 74773 93427
rect 74891 93309 74933 93427
rect 75051 93309 92773 93427
rect 92891 93309 92933 93427
rect 93051 93309 110773 93427
rect 110891 93309 110933 93427
rect 111051 93309 128773 93427
rect 128891 93309 128933 93427
rect 129051 93309 146773 93427
rect 146891 93309 146933 93427
rect 147051 93309 164773 93427
rect 164891 93309 164933 93427
rect 165051 93309 182773 93427
rect 182891 93309 182933 93427
rect 183051 93309 200773 93427
rect 200891 93309 200933 93427
rect 201051 93309 218773 93427
rect 218891 93309 218933 93427
rect 219051 93309 236773 93427
rect 236891 93309 236933 93427
rect 237051 93309 254773 93427
rect 254891 93309 254933 93427
rect 255051 93309 272773 93427
rect 272891 93309 272933 93427
rect 273051 93309 290773 93427
rect 290891 93309 290933 93427
rect 291051 93309 293631 93427
rect 293749 93309 293791 93427
rect 293909 93309 294405 93427
rect -2443 93293 294405 93309
rect -1483 91727 293445 91743
rect -1483 91609 -987 91727
rect -869 91609 -827 91727
rect -709 91609 913 91727
rect 1031 91609 1073 91727
rect 1191 91609 18913 91727
rect 19031 91609 19073 91727
rect 19191 91609 36913 91727
rect 37031 91609 37073 91727
rect 37191 91609 54913 91727
rect 55031 91609 55073 91727
rect 55191 91609 72913 91727
rect 73031 91609 73073 91727
rect 73191 91609 90913 91727
rect 91031 91609 91073 91727
rect 91191 91609 108913 91727
rect 109031 91609 109073 91727
rect 109191 91609 126913 91727
rect 127031 91609 127073 91727
rect 127191 91609 144913 91727
rect 145031 91609 145073 91727
rect 145191 91609 162913 91727
rect 163031 91609 163073 91727
rect 163191 91609 180913 91727
rect 181031 91609 181073 91727
rect 181191 91609 198913 91727
rect 199031 91609 199073 91727
rect 199191 91609 216913 91727
rect 217031 91609 217073 91727
rect 217191 91609 234913 91727
rect 235031 91609 235073 91727
rect 235191 91609 252913 91727
rect 253031 91609 253073 91727
rect 253191 91609 270913 91727
rect 271031 91609 271073 91727
rect 271191 91609 288913 91727
rect 289031 91609 289073 91727
rect 289191 91609 292671 91727
rect 292789 91609 292831 91727
rect 292949 91609 293445 91727
rect -1483 91567 293445 91609
rect -1483 91449 -987 91567
rect -869 91449 -827 91567
rect -709 91449 913 91567
rect 1031 91449 1073 91567
rect 1191 91449 18913 91567
rect 19031 91449 19073 91567
rect 19191 91449 36913 91567
rect 37031 91449 37073 91567
rect 37191 91449 54913 91567
rect 55031 91449 55073 91567
rect 55191 91449 72913 91567
rect 73031 91449 73073 91567
rect 73191 91449 90913 91567
rect 91031 91449 91073 91567
rect 91191 91449 108913 91567
rect 109031 91449 109073 91567
rect 109191 91449 126913 91567
rect 127031 91449 127073 91567
rect 127191 91449 144913 91567
rect 145031 91449 145073 91567
rect 145191 91449 162913 91567
rect 163031 91449 163073 91567
rect 163191 91449 180913 91567
rect 181031 91449 181073 91567
rect 181191 91449 198913 91567
rect 199031 91449 199073 91567
rect 199191 91449 216913 91567
rect 217031 91449 217073 91567
rect 217191 91449 234913 91567
rect 235031 91449 235073 91567
rect 235191 91449 252913 91567
rect 253031 91449 253073 91567
rect 253191 91449 270913 91567
rect 271031 91449 271073 91567
rect 271191 91449 288913 91567
rect 289031 91449 289073 91567
rect 289191 91449 292671 91567
rect 292789 91449 292831 91567
rect 292949 91449 293445 91567
rect -1483 91433 293445 91449
rect -4363 88307 296325 88323
rect -4363 88189 -4347 88307
rect -4229 88189 -4187 88307
rect -4069 88189 15493 88307
rect 15611 88189 15653 88307
rect 15771 88189 33493 88307
rect 33611 88189 33653 88307
rect 33771 88189 51493 88307
rect 51611 88189 51653 88307
rect 51771 88189 69493 88307
rect 69611 88189 69653 88307
rect 69771 88189 87493 88307
rect 87611 88189 87653 88307
rect 87771 88189 105493 88307
rect 105611 88189 105653 88307
rect 105771 88189 123493 88307
rect 123611 88189 123653 88307
rect 123771 88189 141493 88307
rect 141611 88189 141653 88307
rect 141771 88189 159493 88307
rect 159611 88189 159653 88307
rect 159771 88189 177493 88307
rect 177611 88189 177653 88307
rect 177771 88189 195493 88307
rect 195611 88189 195653 88307
rect 195771 88189 213493 88307
rect 213611 88189 213653 88307
rect 213771 88189 231493 88307
rect 231611 88189 231653 88307
rect 231771 88189 249493 88307
rect 249611 88189 249653 88307
rect 249771 88189 267493 88307
rect 267611 88189 267653 88307
rect 267771 88189 285493 88307
rect 285611 88189 285653 88307
rect 285771 88189 296031 88307
rect 296149 88189 296191 88307
rect 296309 88189 296325 88307
rect -4363 88147 296325 88189
rect -4363 88029 -4347 88147
rect -4229 88029 -4187 88147
rect -4069 88029 15493 88147
rect 15611 88029 15653 88147
rect 15771 88029 33493 88147
rect 33611 88029 33653 88147
rect 33771 88029 51493 88147
rect 51611 88029 51653 88147
rect 51771 88029 69493 88147
rect 69611 88029 69653 88147
rect 69771 88029 87493 88147
rect 87611 88029 87653 88147
rect 87771 88029 105493 88147
rect 105611 88029 105653 88147
rect 105771 88029 123493 88147
rect 123611 88029 123653 88147
rect 123771 88029 141493 88147
rect 141611 88029 141653 88147
rect 141771 88029 159493 88147
rect 159611 88029 159653 88147
rect 159771 88029 177493 88147
rect 177611 88029 177653 88147
rect 177771 88029 195493 88147
rect 195611 88029 195653 88147
rect 195771 88029 213493 88147
rect 213611 88029 213653 88147
rect 213771 88029 231493 88147
rect 231611 88029 231653 88147
rect 231771 88029 249493 88147
rect 249611 88029 249653 88147
rect 249771 88029 267493 88147
rect 267611 88029 267653 88147
rect 267771 88029 285493 88147
rect 285611 88029 285653 88147
rect 285771 88029 296031 88147
rect 296149 88029 296191 88147
rect 296309 88029 296325 88147
rect -4363 88013 296325 88029
rect -3403 86447 295365 86463
rect -3403 86329 -3387 86447
rect -3269 86329 -3227 86447
rect -3109 86329 13633 86447
rect 13751 86329 13793 86447
rect 13911 86329 31633 86447
rect 31751 86329 31793 86447
rect 31911 86329 49633 86447
rect 49751 86329 49793 86447
rect 49911 86329 67633 86447
rect 67751 86329 67793 86447
rect 67911 86329 85633 86447
rect 85751 86329 85793 86447
rect 85911 86329 103633 86447
rect 103751 86329 103793 86447
rect 103911 86329 121633 86447
rect 121751 86329 121793 86447
rect 121911 86329 139633 86447
rect 139751 86329 139793 86447
rect 139911 86329 157633 86447
rect 157751 86329 157793 86447
rect 157911 86329 175633 86447
rect 175751 86329 175793 86447
rect 175911 86329 193633 86447
rect 193751 86329 193793 86447
rect 193911 86329 211633 86447
rect 211751 86329 211793 86447
rect 211911 86329 229633 86447
rect 229751 86329 229793 86447
rect 229911 86329 247633 86447
rect 247751 86329 247793 86447
rect 247911 86329 265633 86447
rect 265751 86329 265793 86447
rect 265911 86329 283633 86447
rect 283751 86329 283793 86447
rect 283911 86329 295071 86447
rect 295189 86329 295231 86447
rect 295349 86329 295365 86447
rect -3403 86287 295365 86329
rect -3403 86169 -3387 86287
rect -3269 86169 -3227 86287
rect -3109 86169 13633 86287
rect 13751 86169 13793 86287
rect 13911 86169 31633 86287
rect 31751 86169 31793 86287
rect 31911 86169 49633 86287
rect 49751 86169 49793 86287
rect 49911 86169 67633 86287
rect 67751 86169 67793 86287
rect 67911 86169 85633 86287
rect 85751 86169 85793 86287
rect 85911 86169 103633 86287
rect 103751 86169 103793 86287
rect 103911 86169 121633 86287
rect 121751 86169 121793 86287
rect 121911 86169 139633 86287
rect 139751 86169 139793 86287
rect 139911 86169 157633 86287
rect 157751 86169 157793 86287
rect 157911 86169 175633 86287
rect 175751 86169 175793 86287
rect 175911 86169 193633 86287
rect 193751 86169 193793 86287
rect 193911 86169 211633 86287
rect 211751 86169 211793 86287
rect 211911 86169 229633 86287
rect 229751 86169 229793 86287
rect 229911 86169 247633 86287
rect 247751 86169 247793 86287
rect 247911 86169 265633 86287
rect 265751 86169 265793 86287
rect 265911 86169 283633 86287
rect 283751 86169 283793 86287
rect 283911 86169 295071 86287
rect 295189 86169 295231 86287
rect 295349 86169 295365 86287
rect -3403 86153 295365 86169
rect -2443 84587 294405 84603
rect -2443 84469 -2427 84587
rect -2309 84469 -2267 84587
rect -2149 84469 11773 84587
rect 11891 84469 11933 84587
rect 12051 84469 29773 84587
rect 29891 84469 29933 84587
rect 30051 84469 47773 84587
rect 47891 84469 47933 84587
rect 48051 84469 65773 84587
rect 65891 84469 65933 84587
rect 66051 84469 83773 84587
rect 83891 84469 83933 84587
rect 84051 84469 101773 84587
rect 101891 84469 101933 84587
rect 102051 84469 119773 84587
rect 119891 84469 119933 84587
rect 120051 84469 137773 84587
rect 137891 84469 137933 84587
rect 138051 84469 155773 84587
rect 155891 84469 155933 84587
rect 156051 84469 173773 84587
rect 173891 84469 173933 84587
rect 174051 84469 191773 84587
rect 191891 84469 191933 84587
rect 192051 84469 209773 84587
rect 209891 84469 209933 84587
rect 210051 84469 227773 84587
rect 227891 84469 227933 84587
rect 228051 84469 245773 84587
rect 245891 84469 245933 84587
rect 246051 84469 263773 84587
rect 263891 84469 263933 84587
rect 264051 84469 281773 84587
rect 281891 84469 281933 84587
rect 282051 84469 294111 84587
rect 294229 84469 294271 84587
rect 294389 84469 294405 84587
rect -2443 84427 294405 84469
rect -2443 84309 -2427 84427
rect -2309 84309 -2267 84427
rect -2149 84309 11773 84427
rect 11891 84309 11933 84427
rect 12051 84309 29773 84427
rect 29891 84309 29933 84427
rect 30051 84309 47773 84427
rect 47891 84309 47933 84427
rect 48051 84309 65773 84427
rect 65891 84309 65933 84427
rect 66051 84309 83773 84427
rect 83891 84309 83933 84427
rect 84051 84309 101773 84427
rect 101891 84309 101933 84427
rect 102051 84309 119773 84427
rect 119891 84309 119933 84427
rect 120051 84309 137773 84427
rect 137891 84309 137933 84427
rect 138051 84309 155773 84427
rect 155891 84309 155933 84427
rect 156051 84309 173773 84427
rect 173891 84309 173933 84427
rect 174051 84309 191773 84427
rect 191891 84309 191933 84427
rect 192051 84309 209773 84427
rect 209891 84309 209933 84427
rect 210051 84309 227773 84427
rect 227891 84309 227933 84427
rect 228051 84309 245773 84427
rect 245891 84309 245933 84427
rect 246051 84309 263773 84427
rect 263891 84309 263933 84427
rect 264051 84309 281773 84427
rect 281891 84309 281933 84427
rect 282051 84309 294111 84427
rect 294229 84309 294271 84427
rect 294389 84309 294405 84427
rect -2443 84293 294405 84309
rect -1483 82727 293445 82743
rect -1483 82609 -1467 82727
rect -1349 82609 -1307 82727
rect -1189 82609 9913 82727
rect 10031 82609 10073 82727
rect 10191 82609 27913 82727
rect 28031 82609 28073 82727
rect 28191 82609 45913 82727
rect 46031 82609 46073 82727
rect 46191 82609 63913 82727
rect 64031 82609 64073 82727
rect 64191 82609 81913 82727
rect 82031 82609 82073 82727
rect 82191 82609 99913 82727
rect 100031 82609 100073 82727
rect 100191 82609 117913 82727
rect 118031 82609 118073 82727
rect 118191 82609 135913 82727
rect 136031 82609 136073 82727
rect 136191 82609 153913 82727
rect 154031 82609 154073 82727
rect 154191 82609 171913 82727
rect 172031 82609 172073 82727
rect 172191 82609 189913 82727
rect 190031 82609 190073 82727
rect 190191 82609 207913 82727
rect 208031 82609 208073 82727
rect 208191 82609 225913 82727
rect 226031 82609 226073 82727
rect 226191 82609 243913 82727
rect 244031 82609 244073 82727
rect 244191 82609 261913 82727
rect 262031 82609 262073 82727
rect 262191 82609 279913 82727
rect 280031 82609 280073 82727
rect 280191 82609 293151 82727
rect 293269 82609 293311 82727
rect 293429 82609 293445 82727
rect -1483 82567 293445 82609
rect -1483 82449 -1467 82567
rect -1349 82449 -1307 82567
rect -1189 82449 9913 82567
rect 10031 82449 10073 82567
rect 10191 82449 27913 82567
rect 28031 82449 28073 82567
rect 28191 82449 45913 82567
rect 46031 82449 46073 82567
rect 46191 82449 63913 82567
rect 64031 82449 64073 82567
rect 64191 82449 81913 82567
rect 82031 82449 82073 82567
rect 82191 82449 99913 82567
rect 100031 82449 100073 82567
rect 100191 82449 117913 82567
rect 118031 82449 118073 82567
rect 118191 82449 135913 82567
rect 136031 82449 136073 82567
rect 136191 82449 153913 82567
rect 154031 82449 154073 82567
rect 154191 82449 171913 82567
rect 172031 82449 172073 82567
rect 172191 82449 189913 82567
rect 190031 82449 190073 82567
rect 190191 82449 207913 82567
rect 208031 82449 208073 82567
rect 208191 82449 225913 82567
rect 226031 82449 226073 82567
rect 226191 82449 243913 82567
rect 244031 82449 244073 82567
rect 244191 82449 261913 82567
rect 262031 82449 262073 82567
rect 262191 82449 279913 82567
rect 280031 82449 280073 82567
rect 280191 82449 293151 82567
rect 293269 82449 293311 82567
rect 293429 82449 293445 82567
rect -1483 82433 293445 82449
rect -4363 79307 296325 79323
rect -4363 79189 -3867 79307
rect -3749 79189 -3707 79307
rect -3589 79189 6493 79307
rect 6611 79189 6653 79307
rect 6771 79189 24493 79307
rect 24611 79189 24653 79307
rect 24771 79189 42493 79307
rect 42611 79189 42653 79307
rect 42771 79189 60493 79307
rect 60611 79189 60653 79307
rect 60771 79189 78493 79307
rect 78611 79189 78653 79307
rect 78771 79189 96493 79307
rect 96611 79189 96653 79307
rect 96771 79189 114493 79307
rect 114611 79189 114653 79307
rect 114771 79189 132493 79307
rect 132611 79189 132653 79307
rect 132771 79189 150493 79307
rect 150611 79189 150653 79307
rect 150771 79189 168493 79307
rect 168611 79189 168653 79307
rect 168771 79189 186493 79307
rect 186611 79189 186653 79307
rect 186771 79189 204493 79307
rect 204611 79189 204653 79307
rect 204771 79189 222493 79307
rect 222611 79189 222653 79307
rect 222771 79189 240493 79307
rect 240611 79189 240653 79307
rect 240771 79189 258493 79307
rect 258611 79189 258653 79307
rect 258771 79189 276493 79307
rect 276611 79189 276653 79307
rect 276771 79189 295551 79307
rect 295669 79189 295711 79307
rect 295829 79189 296325 79307
rect -4363 79147 296325 79189
rect -4363 79029 -3867 79147
rect -3749 79029 -3707 79147
rect -3589 79029 6493 79147
rect 6611 79029 6653 79147
rect 6771 79029 24493 79147
rect 24611 79029 24653 79147
rect 24771 79029 42493 79147
rect 42611 79029 42653 79147
rect 42771 79029 60493 79147
rect 60611 79029 60653 79147
rect 60771 79029 78493 79147
rect 78611 79029 78653 79147
rect 78771 79029 96493 79147
rect 96611 79029 96653 79147
rect 96771 79029 114493 79147
rect 114611 79029 114653 79147
rect 114771 79029 132493 79147
rect 132611 79029 132653 79147
rect 132771 79029 150493 79147
rect 150611 79029 150653 79147
rect 150771 79029 168493 79147
rect 168611 79029 168653 79147
rect 168771 79029 186493 79147
rect 186611 79029 186653 79147
rect 186771 79029 204493 79147
rect 204611 79029 204653 79147
rect 204771 79029 222493 79147
rect 222611 79029 222653 79147
rect 222771 79029 240493 79147
rect 240611 79029 240653 79147
rect 240771 79029 258493 79147
rect 258611 79029 258653 79147
rect 258771 79029 276493 79147
rect 276611 79029 276653 79147
rect 276771 79029 295551 79147
rect 295669 79029 295711 79147
rect 295829 79029 296325 79147
rect -4363 79013 296325 79029
rect -3403 77447 295365 77463
rect -3403 77329 -2907 77447
rect -2789 77329 -2747 77447
rect -2629 77329 4633 77447
rect 4751 77329 4793 77447
rect 4911 77329 22633 77447
rect 22751 77329 22793 77447
rect 22911 77329 40633 77447
rect 40751 77329 40793 77447
rect 40911 77329 58633 77447
rect 58751 77329 58793 77447
rect 58911 77329 76633 77447
rect 76751 77329 76793 77447
rect 76911 77329 94633 77447
rect 94751 77329 94793 77447
rect 94911 77329 112633 77447
rect 112751 77329 112793 77447
rect 112911 77329 130633 77447
rect 130751 77329 130793 77447
rect 130911 77329 148633 77447
rect 148751 77329 148793 77447
rect 148911 77329 166633 77447
rect 166751 77329 166793 77447
rect 166911 77329 184633 77447
rect 184751 77329 184793 77447
rect 184911 77329 202633 77447
rect 202751 77329 202793 77447
rect 202911 77329 220633 77447
rect 220751 77329 220793 77447
rect 220911 77329 238633 77447
rect 238751 77329 238793 77447
rect 238911 77329 256633 77447
rect 256751 77329 256793 77447
rect 256911 77329 274633 77447
rect 274751 77329 274793 77447
rect 274911 77329 294591 77447
rect 294709 77329 294751 77447
rect 294869 77329 295365 77447
rect -3403 77287 295365 77329
rect -3403 77169 -2907 77287
rect -2789 77169 -2747 77287
rect -2629 77169 4633 77287
rect 4751 77169 4793 77287
rect 4911 77169 22633 77287
rect 22751 77169 22793 77287
rect 22911 77169 40633 77287
rect 40751 77169 40793 77287
rect 40911 77169 58633 77287
rect 58751 77169 58793 77287
rect 58911 77169 76633 77287
rect 76751 77169 76793 77287
rect 76911 77169 94633 77287
rect 94751 77169 94793 77287
rect 94911 77169 112633 77287
rect 112751 77169 112793 77287
rect 112911 77169 130633 77287
rect 130751 77169 130793 77287
rect 130911 77169 148633 77287
rect 148751 77169 148793 77287
rect 148911 77169 166633 77287
rect 166751 77169 166793 77287
rect 166911 77169 184633 77287
rect 184751 77169 184793 77287
rect 184911 77169 202633 77287
rect 202751 77169 202793 77287
rect 202911 77169 220633 77287
rect 220751 77169 220793 77287
rect 220911 77169 238633 77287
rect 238751 77169 238793 77287
rect 238911 77169 256633 77287
rect 256751 77169 256793 77287
rect 256911 77169 274633 77287
rect 274751 77169 274793 77287
rect 274911 77169 294591 77287
rect 294709 77169 294751 77287
rect 294869 77169 295365 77287
rect -3403 77153 295365 77169
rect -2443 75587 294405 75603
rect -2443 75469 -1947 75587
rect -1829 75469 -1787 75587
rect -1669 75469 2773 75587
rect 2891 75469 2933 75587
rect 3051 75469 20773 75587
rect 20891 75469 20933 75587
rect 21051 75469 38773 75587
rect 38891 75469 38933 75587
rect 39051 75469 56773 75587
rect 56891 75469 56933 75587
rect 57051 75469 74773 75587
rect 74891 75469 74933 75587
rect 75051 75469 92773 75587
rect 92891 75469 92933 75587
rect 93051 75469 110773 75587
rect 110891 75469 110933 75587
rect 111051 75469 128773 75587
rect 128891 75469 128933 75587
rect 129051 75469 146773 75587
rect 146891 75469 146933 75587
rect 147051 75469 164773 75587
rect 164891 75469 164933 75587
rect 165051 75469 182773 75587
rect 182891 75469 182933 75587
rect 183051 75469 200773 75587
rect 200891 75469 200933 75587
rect 201051 75469 218773 75587
rect 218891 75469 218933 75587
rect 219051 75469 236773 75587
rect 236891 75469 236933 75587
rect 237051 75469 254773 75587
rect 254891 75469 254933 75587
rect 255051 75469 272773 75587
rect 272891 75469 272933 75587
rect 273051 75469 290773 75587
rect 290891 75469 290933 75587
rect 291051 75469 293631 75587
rect 293749 75469 293791 75587
rect 293909 75469 294405 75587
rect -2443 75427 294405 75469
rect -2443 75309 -1947 75427
rect -1829 75309 -1787 75427
rect -1669 75309 2773 75427
rect 2891 75309 2933 75427
rect 3051 75309 20773 75427
rect 20891 75309 20933 75427
rect 21051 75309 38773 75427
rect 38891 75309 38933 75427
rect 39051 75309 56773 75427
rect 56891 75309 56933 75427
rect 57051 75309 74773 75427
rect 74891 75309 74933 75427
rect 75051 75309 92773 75427
rect 92891 75309 92933 75427
rect 93051 75309 110773 75427
rect 110891 75309 110933 75427
rect 111051 75309 128773 75427
rect 128891 75309 128933 75427
rect 129051 75309 146773 75427
rect 146891 75309 146933 75427
rect 147051 75309 164773 75427
rect 164891 75309 164933 75427
rect 165051 75309 182773 75427
rect 182891 75309 182933 75427
rect 183051 75309 200773 75427
rect 200891 75309 200933 75427
rect 201051 75309 218773 75427
rect 218891 75309 218933 75427
rect 219051 75309 236773 75427
rect 236891 75309 236933 75427
rect 237051 75309 254773 75427
rect 254891 75309 254933 75427
rect 255051 75309 272773 75427
rect 272891 75309 272933 75427
rect 273051 75309 290773 75427
rect 290891 75309 290933 75427
rect 291051 75309 293631 75427
rect 293749 75309 293791 75427
rect 293909 75309 294405 75427
rect -2443 75293 294405 75309
rect -1483 73727 293445 73743
rect -1483 73609 -987 73727
rect -869 73609 -827 73727
rect -709 73609 913 73727
rect 1031 73609 1073 73727
rect 1191 73609 18913 73727
rect 19031 73609 19073 73727
rect 19191 73609 36913 73727
rect 37031 73609 37073 73727
rect 37191 73609 54913 73727
rect 55031 73609 55073 73727
rect 55191 73609 72913 73727
rect 73031 73609 73073 73727
rect 73191 73609 90913 73727
rect 91031 73609 91073 73727
rect 91191 73609 108913 73727
rect 109031 73609 109073 73727
rect 109191 73609 126913 73727
rect 127031 73609 127073 73727
rect 127191 73609 144913 73727
rect 145031 73609 145073 73727
rect 145191 73609 162913 73727
rect 163031 73609 163073 73727
rect 163191 73609 180913 73727
rect 181031 73609 181073 73727
rect 181191 73609 198913 73727
rect 199031 73609 199073 73727
rect 199191 73609 216913 73727
rect 217031 73609 217073 73727
rect 217191 73609 234913 73727
rect 235031 73609 235073 73727
rect 235191 73609 252913 73727
rect 253031 73609 253073 73727
rect 253191 73609 270913 73727
rect 271031 73609 271073 73727
rect 271191 73609 288913 73727
rect 289031 73609 289073 73727
rect 289191 73609 292671 73727
rect 292789 73609 292831 73727
rect 292949 73609 293445 73727
rect -1483 73567 293445 73609
rect -1483 73449 -987 73567
rect -869 73449 -827 73567
rect -709 73449 913 73567
rect 1031 73449 1073 73567
rect 1191 73449 18913 73567
rect 19031 73449 19073 73567
rect 19191 73449 36913 73567
rect 37031 73449 37073 73567
rect 37191 73449 54913 73567
rect 55031 73449 55073 73567
rect 55191 73449 72913 73567
rect 73031 73449 73073 73567
rect 73191 73449 90913 73567
rect 91031 73449 91073 73567
rect 91191 73449 108913 73567
rect 109031 73449 109073 73567
rect 109191 73449 126913 73567
rect 127031 73449 127073 73567
rect 127191 73449 144913 73567
rect 145031 73449 145073 73567
rect 145191 73449 162913 73567
rect 163031 73449 163073 73567
rect 163191 73449 180913 73567
rect 181031 73449 181073 73567
rect 181191 73449 198913 73567
rect 199031 73449 199073 73567
rect 199191 73449 216913 73567
rect 217031 73449 217073 73567
rect 217191 73449 234913 73567
rect 235031 73449 235073 73567
rect 235191 73449 252913 73567
rect 253031 73449 253073 73567
rect 253191 73449 270913 73567
rect 271031 73449 271073 73567
rect 271191 73449 288913 73567
rect 289031 73449 289073 73567
rect 289191 73449 292671 73567
rect 292789 73449 292831 73567
rect 292949 73449 293445 73567
rect -1483 73433 293445 73449
rect -4363 70307 296325 70323
rect -4363 70189 -4347 70307
rect -4229 70189 -4187 70307
rect -4069 70189 15493 70307
rect 15611 70189 15653 70307
rect 15771 70189 33493 70307
rect 33611 70189 33653 70307
rect 33771 70189 51493 70307
rect 51611 70189 51653 70307
rect 51771 70189 69493 70307
rect 69611 70189 69653 70307
rect 69771 70189 87493 70307
rect 87611 70189 87653 70307
rect 87771 70189 105493 70307
rect 105611 70189 105653 70307
rect 105771 70189 123493 70307
rect 123611 70189 123653 70307
rect 123771 70189 141493 70307
rect 141611 70189 141653 70307
rect 141771 70189 159493 70307
rect 159611 70189 159653 70307
rect 159771 70189 177493 70307
rect 177611 70189 177653 70307
rect 177771 70189 195493 70307
rect 195611 70189 195653 70307
rect 195771 70189 213493 70307
rect 213611 70189 213653 70307
rect 213771 70189 231493 70307
rect 231611 70189 231653 70307
rect 231771 70189 249493 70307
rect 249611 70189 249653 70307
rect 249771 70189 267493 70307
rect 267611 70189 267653 70307
rect 267771 70189 285493 70307
rect 285611 70189 285653 70307
rect 285771 70189 296031 70307
rect 296149 70189 296191 70307
rect 296309 70189 296325 70307
rect -4363 70147 296325 70189
rect -4363 70029 -4347 70147
rect -4229 70029 -4187 70147
rect -4069 70029 15493 70147
rect 15611 70029 15653 70147
rect 15771 70029 33493 70147
rect 33611 70029 33653 70147
rect 33771 70029 51493 70147
rect 51611 70029 51653 70147
rect 51771 70029 69493 70147
rect 69611 70029 69653 70147
rect 69771 70029 87493 70147
rect 87611 70029 87653 70147
rect 87771 70029 105493 70147
rect 105611 70029 105653 70147
rect 105771 70029 123493 70147
rect 123611 70029 123653 70147
rect 123771 70029 141493 70147
rect 141611 70029 141653 70147
rect 141771 70029 159493 70147
rect 159611 70029 159653 70147
rect 159771 70029 177493 70147
rect 177611 70029 177653 70147
rect 177771 70029 195493 70147
rect 195611 70029 195653 70147
rect 195771 70029 213493 70147
rect 213611 70029 213653 70147
rect 213771 70029 231493 70147
rect 231611 70029 231653 70147
rect 231771 70029 249493 70147
rect 249611 70029 249653 70147
rect 249771 70029 267493 70147
rect 267611 70029 267653 70147
rect 267771 70029 285493 70147
rect 285611 70029 285653 70147
rect 285771 70029 296031 70147
rect 296149 70029 296191 70147
rect 296309 70029 296325 70147
rect -4363 70013 296325 70029
rect -3403 68447 295365 68463
rect -3403 68329 -3387 68447
rect -3269 68329 -3227 68447
rect -3109 68329 13633 68447
rect 13751 68329 13793 68447
rect 13911 68329 31633 68447
rect 31751 68329 31793 68447
rect 31911 68329 49633 68447
rect 49751 68329 49793 68447
rect 49911 68329 67633 68447
rect 67751 68329 67793 68447
rect 67911 68329 85633 68447
rect 85751 68329 85793 68447
rect 85911 68329 103633 68447
rect 103751 68329 103793 68447
rect 103911 68329 121633 68447
rect 121751 68329 121793 68447
rect 121911 68329 139633 68447
rect 139751 68329 139793 68447
rect 139911 68329 157633 68447
rect 157751 68329 157793 68447
rect 157911 68329 175633 68447
rect 175751 68329 175793 68447
rect 175911 68329 193633 68447
rect 193751 68329 193793 68447
rect 193911 68329 211633 68447
rect 211751 68329 211793 68447
rect 211911 68329 229633 68447
rect 229751 68329 229793 68447
rect 229911 68329 247633 68447
rect 247751 68329 247793 68447
rect 247911 68329 265633 68447
rect 265751 68329 265793 68447
rect 265911 68329 283633 68447
rect 283751 68329 283793 68447
rect 283911 68329 295071 68447
rect 295189 68329 295231 68447
rect 295349 68329 295365 68447
rect -3403 68287 295365 68329
rect -3403 68169 -3387 68287
rect -3269 68169 -3227 68287
rect -3109 68169 13633 68287
rect 13751 68169 13793 68287
rect 13911 68169 31633 68287
rect 31751 68169 31793 68287
rect 31911 68169 49633 68287
rect 49751 68169 49793 68287
rect 49911 68169 67633 68287
rect 67751 68169 67793 68287
rect 67911 68169 85633 68287
rect 85751 68169 85793 68287
rect 85911 68169 103633 68287
rect 103751 68169 103793 68287
rect 103911 68169 121633 68287
rect 121751 68169 121793 68287
rect 121911 68169 139633 68287
rect 139751 68169 139793 68287
rect 139911 68169 157633 68287
rect 157751 68169 157793 68287
rect 157911 68169 175633 68287
rect 175751 68169 175793 68287
rect 175911 68169 193633 68287
rect 193751 68169 193793 68287
rect 193911 68169 211633 68287
rect 211751 68169 211793 68287
rect 211911 68169 229633 68287
rect 229751 68169 229793 68287
rect 229911 68169 247633 68287
rect 247751 68169 247793 68287
rect 247911 68169 265633 68287
rect 265751 68169 265793 68287
rect 265911 68169 283633 68287
rect 283751 68169 283793 68287
rect 283911 68169 295071 68287
rect 295189 68169 295231 68287
rect 295349 68169 295365 68287
rect -3403 68153 295365 68169
rect -2443 66587 294405 66603
rect -2443 66469 -2427 66587
rect -2309 66469 -2267 66587
rect -2149 66469 11773 66587
rect 11891 66469 11933 66587
rect 12051 66469 29773 66587
rect 29891 66469 29933 66587
rect 30051 66469 47773 66587
rect 47891 66469 47933 66587
rect 48051 66469 65773 66587
rect 65891 66469 65933 66587
rect 66051 66469 83773 66587
rect 83891 66469 83933 66587
rect 84051 66469 101773 66587
rect 101891 66469 101933 66587
rect 102051 66469 119773 66587
rect 119891 66469 119933 66587
rect 120051 66469 137773 66587
rect 137891 66469 137933 66587
rect 138051 66469 155773 66587
rect 155891 66469 155933 66587
rect 156051 66469 173773 66587
rect 173891 66469 173933 66587
rect 174051 66469 191773 66587
rect 191891 66469 191933 66587
rect 192051 66469 209773 66587
rect 209891 66469 209933 66587
rect 210051 66469 227773 66587
rect 227891 66469 227933 66587
rect 228051 66469 245773 66587
rect 245891 66469 245933 66587
rect 246051 66469 263773 66587
rect 263891 66469 263933 66587
rect 264051 66469 281773 66587
rect 281891 66469 281933 66587
rect 282051 66469 294111 66587
rect 294229 66469 294271 66587
rect 294389 66469 294405 66587
rect -2443 66427 294405 66469
rect -2443 66309 -2427 66427
rect -2309 66309 -2267 66427
rect -2149 66309 11773 66427
rect 11891 66309 11933 66427
rect 12051 66309 29773 66427
rect 29891 66309 29933 66427
rect 30051 66309 47773 66427
rect 47891 66309 47933 66427
rect 48051 66309 65773 66427
rect 65891 66309 65933 66427
rect 66051 66309 83773 66427
rect 83891 66309 83933 66427
rect 84051 66309 101773 66427
rect 101891 66309 101933 66427
rect 102051 66309 119773 66427
rect 119891 66309 119933 66427
rect 120051 66309 137773 66427
rect 137891 66309 137933 66427
rect 138051 66309 155773 66427
rect 155891 66309 155933 66427
rect 156051 66309 173773 66427
rect 173891 66309 173933 66427
rect 174051 66309 191773 66427
rect 191891 66309 191933 66427
rect 192051 66309 209773 66427
rect 209891 66309 209933 66427
rect 210051 66309 227773 66427
rect 227891 66309 227933 66427
rect 228051 66309 245773 66427
rect 245891 66309 245933 66427
rect 246051 66309 263773 66427
rect 263891 66309 263933 66427
rect 264051 66309 281773 66427
rect 281891 66309 281933 66427
rect 282051 66309 294111 66427
rect 294229 66309 294271 66427
rect 294389 66309 294405 66427
rect -2443 66293 294405 66309
rect -1483 64727 293445 64743
rect -1483 64609 -1467 64727
rect -1349 64609 -1307 64727
rect -1189 64609 9913 64727
rect 10031 64609 10073 64727
rect 10191 64609 27913 64727
rect 28031 64609 28073 64727
rect 28191 64609 45913 64727
rect 46031 64609 46073 64727
rect 46191 64609 63913 64727
rect 64031 64609 64073 64727
rect 64191 64609 81913 64727
rect 82031 64609 82073 64727
rect 82191 64609 99913 64727
rect 100031 64609 100073 64727
rect 100191 64609 117913 64727
rect 118031 64609 118073 64727
rect 118191 64609 135913 64727
rect 136031 64609 136073 64727
rect 136191 64609 153913 64727
rect 154031 64609 154073 64727
rect 154191 64609 171913 64727
rect 172031 64609 172073 64727
rect 172191 64609 189913 64727
rect 190031 64609 190073 64727
rect 190191 64609 207913 64727
rect 208031 64609 208073 64727
rect 208191 64609 225913 64727
rect 226031 64609 226073 64727
rect 226191 64609 243913 64727
rect 244031 64609 244073 64727
rect 244191 64609 261913 64727
rect 262031 64609 262073 64727
rect 262191 64609 279913 64727
rect 280031 64609 280073 64727
rect 280191 64609 293151 64727
rect 293269 64609 293311 64727
rect 293429 64609 293445 64727
rect -1483 64567 293445 64609
rect -1483 64449 -1467 64567
rect -1349 64449 -1307 64567
rect -1189 64449 9913 64567
rect 10031 64449 10073 64567
rect 10191 64449 27913 64567
rect 28031 64449 28073 64567
rect 28191 64449 45913 64567
rect 46031 64449 46073 64567
rect 46191 64449 63913 64567
rect 64031 64449 64073 64567
rect 64191 64449 81913 64567
rect 82031 64449 82073 64567
rect 82191 64449 99913 64567
rect 100031 64449 100073 64567
rect 100191 64449 117913 64567
rect 118031 64449 118073 64567
rect 118191 64449 135913 64567
rect 136031 64449 136073 64567
rect 136191 64449 153913 64567
rect 154031 64449 154073 64567
rect 154191 64449 171913 64567
rect 172031 64449 172073 64567
rect 172191 64449 189913 64567
rect 190031 64449 190073 64567
rect 190191 64449 207913 64567
rect 208031 64449 208073 64567
rect 208191 64449 225913 64567
rect 226031 64449 226073 64567
rect 226191 64449 243913 64567
rect 244031 64449 244073 64567
rect 244191 64449 261913 64567
rect 262031 64449 262073 64567
rect 262191 64449 279913 64567
rect 280031 64449 280073 64567
rect 280191 64449 293151 64567
rect 293269 64449 293311 64567
rect 293429 64449 293445 64567
rect -1483 64433 293445 64449
rect -4363 61307 296325 61323
rect -4363 61189 -3867 61307
rect -3749 61189 -3707 61307
rect -3589 61189 6493 61307
rect 6611 61189 6653 61307
rect 6771 61189 24493 61307
rect 24611 61189 24653 61307
rect 24771 61189 42493 61307
rect 42611 61189 42653 61307
rect 42771 61189 60493 61307
rect 60611 61189 60653 61307
rect 60771 61189 78493 61307
rect 78611 61189 78653 61307
rect 78771 61189 96493 61307
rect 96611 61189 96653 61307
rect 96771 61189 114493 61307
rect 114611 61189 114653 61307
rect 114771 61189 132493 61307
rect 132611 61189 132653 61307
rect 132771 61189 150493 61307
rect 150611 61189 150653 61307
rect 150771 61189 168493 61307
rect 168611 61189 168653 61307
rect 168771 61189 186493 61307
rect 186611 61189 186653 61307
rect 186771 61189 204493 61307
rect 204611 61189 204653 61307
rect 204771 61189 222493 61307
rect 222611 61189 222653 61307
rect 222771 61189 240493 61307
rect 240611 61189 240653 61307
rect 240771 61189 258493 61307
rect 258611 61189 258653 61307
rect 258771 61189 276493 61307
rect 276611 61189 276653 61307
rect 276771 61189 295551 61307
rect 295669 61189 295711 61307
rect 295829 61189 296325 61307
rect -4363 61147 296325 61189
rect -4363 61029 -3867 61147
rect -3749 61029 -3707 61147
rect -3589 61029 6493 61147
rect 6611 61029 6653 61147
rect 6771 61029 24493 61147
rect 24611 61029 24653 61147
rect 24771 61029 42493 61147
rect 42611 61029 42653 61147
rect 42771 61029 60493 61147
rect 60611 61029 60653 61147
rect 60771 61029 78493 61147
rect 78611 61029 78653 61147
rect 78771 61029 96493 61147
rect 96611 61029 96653 61147
rect 96771 61029 114493 61147
rect 114611 61029 114653 61147
rect 114771 61029 132493 61147
rect 132611 61029 132653 61147
rect 132771 61029 150493 61147
rect 150611 61029 150653 61147
rect 150771 61029 168493 61147
rect 168611 61029 168653 61147
rect 168771 61029 186493 61147
rect 186611 61029 186653 61147
rect 186771 61029 204493 61147
rect 204611 61029 204653 61147
rect 204771 61029 222493 61147
rect 222611 61029 222653 61147
rect 222771 61029 240493 61147
rect 240611 61029 240653 61147
rect 240771 61029 258493 61147
rect 258611 61029 258653 61147
rect 258771 61029 276493 61147
rect 276611 61029 276653 61147
rect 276771 61029 295551 61147
rect 295669 61029 295711 61147
rect 295829 61029 296325 61147
rect -4363 61013 296325 61029
rect -3403 59447 295365 59463
rect -3403 59329 -2907 59447
rect -2789 59329 -2747 59447
rect -2629 59329 4633 59447
rect 4751 59329 4793 59447
rect 4911 59329 22633 59447
rect 22751 59329 22793 59447
rect 22911 59329 40633 59447
rect 40751 59329 40793 59447
rect 40911 59329 58633 59447
rect 58751 59329 58793 59447
rect 58911 59329 76633 59447
rect 76751 59329 76793 59447
rect 76911 59329 94633 59447
rect 94751 59329 94793 59447
rect 94911 59329 112633 59447
rect 112751 59329 112793 59447
rect 112911 59329 130633 59447
rect 130751 59329 130793 59447
rect 130911 59329 148633 59447
rect 148751 59329 148793 59447
rect 148911 59329 166633 59447
rect 166751 59329 166793 59447
rect 166911 59329 184633 59447
rect 184751 59329 184793 59447
rect 184911 59329 202633 59447
rect 202751 59329 202793 59447
rect 202911 59329 220633 59447
rect 220751 59329 220793 59447
rect 220911 59329 238633 59447
rect 238751 59329 238793 59447
rect 238911 59329 256633 59447
rect 256751 59329 256793 59447
rect 256911 59329 274633 59447
rect 274751 59329 274793 59447
rect 274911 59329 294591 59447
rect 294709 59329 294751 59447
rect 294869 59329 295365 59447
rect -3403 59287 295365 59329
rect -3403 59169 -2907 59287
rect -2789 59169 -2747 59287
rect -2629 59169 4633 59287
rect 4751 59169 4793 59287
rect 4911 59169 22633 59287
rect 22751 59169 22793 59287
rect 22911 59169 40633 59287
rect 40751 59169 40793 59287
rect 40911 59169 58633 59287
rect 58751 59169 58793 59287
rect 58911 59169 76633 59287
rect 76751 59169 76793 59287
rect 76911 59169 94633 59287
rect 94751 59169 94793 59287
rect 94911 59169 112633 59287
rect 112751 59169 112793 59287
rect 112911 59169 130633 59287
rect 130751 59169 130793 59287
rect 130911 59169 148633 59287
rect 148751 59169 148793 59287
rect 148911 59169 166633 59287
rect 166751 59169 166793 59287
rect 166911 59169 184633 59287
rect 184751 59169 184793 59287
rect 184911 59169 202633 59287
rect 202751 59169 202793 59287
rect 202911 59169 220633 59287
rect 220751 59169 220793 59287
rect 220911 59169 238633 59287
rect 238751 59169 238793 59287
rect 238911 59169 256633 59287
rect 256751 59169 256793 59287
rect 256911 59169 274633 59287
rect 274751 59169 274793 59287
rect 274911 59169 294591 59287
rect 294709 59169 294751 59287
rect 294869 59169 295365 59287
rect -3403 59153 295365 59169
rect -2443 57587 294405 57603
rect -2443 57469 -1947 57587
rect -1829 57469 -1787 57587
rect -1669 57469 2773 57587
rect 2891 57469 2933 57587
rect 3051 57469 20773 57587
rect 20891 57469 20933 57587
rect 21051 57469 38773 57587
rect 38891 57469 38933 57587
rect 39051 57469 56773 57587
rect 56891 57469 56933 57587
rect 57051 57469 74773 57587
rect 74891 57469 74933 57587
rect 75051 57469 92773 57587
rect 92891 57469 92933 57587
rect 93051 57469 110773 57587
rect 110891 57469 110933 57587
rect 111051 57469 128773 57587
rect 128891 57469 128933 57587
rect 129051 57469 146773 57587
rect 146891 57469 146933 57587
rect 147051 57469 164773 57587
rect 164891 57469 164933 57587
rect 165051 57469 182773 57587
rect 182891 57469 182933 57587
rect 183051 57469 200773 57587
rect 200891 57469 200933 57587
rect 201051 57469 218773 57587
rect 218891 57469 218933 57587
rect 219051 57469 236773 57587
rect 236891 57469 236933 57587
rect 237051 57469 254773 57587
rect 254891 57469 254933 57587
rect 255051 57469 272773 57587
rect 272891 57469 272933 57587
rect 273051 57469 290773 57587
rect 290891 57469 290933 57587
rect 291051 57469 293631 57587
rect 293749 57469 293791 57587
rect 293909 57469 294405 57587
rect -2443 57427 294405 57469
rect -2443 57309 -1947 57427
rect -1829 57309 -1787 57427
rect -1669 57309 2773 57427
rect 2891 57309 2933 57427
rect 3051 57309 20773 57427
rect 20891 57309 20933 57427
rect 21051 57309 38773 57427
rect 38891 57309 38933 57427
rect 39051 57309 56773 57427
rect 56891 57309 56933 57427
rect 57051 57309 74773 57427
rect 74891 57309 74933 57427
rect 75051 57309 92773 57427
rect 92891 57309 92933 57427
rect 93051 57309 110773 57427
rect 110891 57309 110933 57427
rect 111051 57309 128773 57427
rect 128891 57309 128933 57427
rect 129051 57309 146773 57427
rect 146891 57309 146933 57427
rect 147051 57309 164773 57427
rect 164891 57309 164933 57427
rect 165051 57309 182773 57427
rect 182891 57309 182933 57427
rect 183051 57309 200773 57427
rect 200891 57309 200933 57427
rect 201051 57309 218773 57427
rect 218891 57309 218933 57427
rect 219051 57309 236773 57427
rect 236891 57309 236933 57427
rect 237051 57309 254773 57427
rect 254891 57309 254933 57427
rect 255051 57309 272773 57427
rect 272891 57309 272933 57427
rect 273051 57309 290773 57427
rect 290891 57309 290933 57427
rect 291051 57309 293631 57427
rect 293749 57309 293791 57427
rect 293909 57309 294405 57427
rect -2443 57293 294405 57309
rect -1483 55727 293445 55743
rect -1483 55609 -987 55727
rect -869 55609 -827 55727
rect -709 55609 913 55727
rect 1031 55609 1073 55727
rect 1191 55609 18913 55727
rect 19031 55609 19073 55727
rect 19191 55609 36913 55727
rect 37031 55609 37073 55727
rect 37191 55609 54913 55727
rect 55031 55609 55073 55727
rect 55191 55609 72913 55727
rect 73031 55609 73073 55727
rect 73191 55609 90913 55727
rect 91031 55609 91073 55727
rect 91191 55609 108913 55727
rect 109031 55609 109073 55727
rect 109191 55609 126913 55727
rect 127031 55609 127073 55727
rect 127191 55609 144913 55727
rect 145031 55609 145073 55727
rect 145191 55609 162913 55727
rect 163031 55609 163073 55727
rect 163191 55609 180913 55727
rect 181031 55609 181073 55727
rect 181191 55609 198913 55727
rect 199031 55609 199073 55727
rect 199191 55609 216913 55727
rect 217031 55609 217073 55727
rect 217191 55609 234913 55727
rect 235031 55609 235073 55727
rect 235191 55609 252913 55727
rect 253031 55609 253073 55727
rect 253191 55609 270913 55727
rect 271031 55609 271073 55727
rect 271191 55609 288913 55727
rect 289031 55609 289073 55727
rect 289191 55609 292671 55727
rect 292789 55609 292831 55727
rect 292949 55609 293445 55727
rect -1483 55567 293445 55609
rect -1483 55449 -987 55567
rect -869 55449 -827 55567
rect -709 55449 913 55567
rect 1031 55449 1073 55567
rect 1191 55449 18913 55567
rect 19031 55449 19073 55567
rect 19191 55449 36913 55567
rect 37031 55449 37073 55567
rect 37191 55449 54913 55567
rect 55031 55449 55073 55567
rect 55191 55449 72913 55567
rect 73031 55449 73073 55567
rect 73191 55449 90913 55567
rect 91031 55449 91073 55567
rect 91191 55449 108913 55567
rect 109031 55449 109073 55567
rect 109191 55449 126913 55567
rect 127031 55449 127073 55567
rect 127191 55449 144913 55567
rect 145031 55449 145073 55567
rect 145191 55449 162913 55567
rect 163031 55449 163073 55567
rect 163191 55449 180913 55567
rect 181031 55449 181073 55567
rect 181191 55449 198913 55567
rect 199031 55449 199073 55567
rect 199191 55449 216913 55567
rect 217031 55449 217073 55567
rect 217191 55449 234913 55567
rect 235031 55449 235073 55567
rect 235191 55449 252913 55567
rect 253031 55449 253073 55567
rect 253191 55449 270913 55567
rect 271031 55449 271073 55567
rect 271191 55449 288913 55567
rect 289031 55449 289073 55567
rect 289191 55449 292671 55567
rect 292789 55449 292831 55567
rect 292949 55449 293445 55567
rect -1483 55433 293445 55449
rect -4363 52307 296325 52323
rect -4363 52189 -4347 52307
rect -4229 52189 -4187 52307
rect -4069 52189 15493 52307
rect 15611 52189 15653 52307
rect 15771 52189 33493 52307
rect 33611 52189 33653 52307
rect 33771 52189 51493 52307
rect 51611 52189 51653 52307
rect 51771 52189 69493 52307
rect 69611 52189 69653 52307
rect 69771 52189 87493 52307
rect 87611 52189 87653 52307
rect 87771 52189 105493 52307
rect 105611 52189 105653 52307
rect 105771 52189 123493 52307
rect 123611 52189 123653 52307
rect 123771 52189 141493 52307
rect 141611 52189 141653 52307
rect 141771 52189 159493 52307
rect 159611 52189 159653 52307
rect 159771 52189 177493 52307
rect 177611 52189 177653 52307
rect 177771 52189 195493 52307
rect 195611 52189 195653 52307
rect 195771 52189 213493 52307
rect 213611 52189 213653 52307
rect 213771 52189 231493 52307
rect 231611 52189 231653 52307
rect 231771 52189 249493 52307
rect 249611 52189 249653 52307
rect 249771 52189 267493 52307
rect 267611 52189 267653 52307
rect 267771 52189 285493 52307
rect 285611 52189 285653 52307
rect 285771 52189 296031 52307
rect 296149 52189 296191 52307
rect 296309 52189 296325 52307
rect -4363 52147 296325 52189
rect -4363 52029 -4347 52147
rect -4229 52029 -4187 52147
rect -4069 52029 15493 52147
rect 15611 52029 15653 52147
rect 15771 52029 33493 52147
rect 33611 52029 33653 52147
rect 33771 52029 51493 52147
rect 51611 52029 51653 52147
rect 51771 52029 69493 52147
rect 69611 52029 69653 52147
rect 69771 52029 87493 52147
rect 87611 52029 87653 52147
rect 87771 52029 105493 52147
rect 105611 52029 105653 52147
rect 105771 52029 123493 52147
rect 123611 52029 123653 52147
rect 123771 52029 141493 52147
rect 141611 52029 141653 52147
rect 141771 52029 159493 52147
rect 159611 52029 159653 52147
rect 159771 52029 177493 52147
rect 177611 52029 177653 52147
rect 177771 52029 195493 52147
rect 195611 52029 195653 52147
rect 195771 52029 213493 52147
rect 213611 52029 213653 52147
rect 213771 52029 231493 52147
rect 231611 52029 231653 52147
rect 231771 52029 249493 52147
rect 249611 52029 249653 52147
rect 249771 52029 267493 52147
rect 267611 52029 267653 52147
rect 267771 52029 285493 52147
rect 285611 52029 285653 52147
rect 285771 52029 296031 52147
rect 296149 52029 296191 52147
rect 296309 52029 296325 52147
rect -4363 52013 296325 52029
rect -3403 50447 295365 50463
rect -3403 50329 -3387 50447
rect -3269 50329 -3227 50447
rect -3109 50329 13633 50447
rect 13751 50329 13793 50447
rect 13911 50329 31633 50447
rect 31751 50329 31793 50447
rect 31911 50329 49633 50447
rect 49751 50329 49793 50447
rect 49911 50329 67633 50447
rect 67751 50329 67793 50447
rect 67911 50329 85633 50447
rect 85751 50329 85793 50447
rect 85911 50329 103633 50447
rect 103751 50329 103793 50447
rect 103911 50329 121633 50447
rect 121751 50329 121793 50447
rect 121911 50329 139633 50447
rect 139751 50329 139793 50447
rect 139911 50329 157633 50447
rect 157751 50329 157793 50447
rect 157911 50329 175633 50447
rect 175751 50329 175793 50447
rect 175911 50329 193633 50447
rect 193751 50329 193793 50447
rect 193911 50329 211633 50447
rect 211751 50329 211793 50447
rect 211911 50329 229633 50447
rect 229751 50329 229793 50447
rect 229911 50329 247633 50447
rect 247751 50329 247793 50447
rect 247911 50329 265633 50447
rect 265751 50329 265793 50447
rect 265911 50329 283633 50447
rect 283751 50329 283793 50447
rect 283911 50329 295071 50447
rect 295189 50329 295231 50447
rect 295349 50329 295365 50447
rect -3403 50287 295365 50329
rect -3403 50169 -3387 50287
rect -3269 50169 -3227 50287
rect -3109 50169 13633 50287
rect 13751 50169 13793 50287
rect 13911 50169 31633 50287
rect 31751 50169 31793 50287
rect 31911 50169 49633 50287
rect 49751 50169 49793 50287
rect 49911 50169 67633 50287
rect 67751 50169 67793 50287
rect 67911 50169 85633 50287
rect 85751 50169 85793 50287
rect 85911 50169 103633 50287
rect 103751 50169 103793 50287
rect 103911 50169 121633 50287
rect 121751 50169 121793 50287
rect 121911 50169 139633 50287
rect 139751 50169 139793 50287
rect 139911 50169 157633 50287
rect 157751 50169 157793 50287
rect 157911 50169 175633 50287
rect 175751 50169 175793 50287
rect 175911 50169 193633 50287
rect 193751 50169 193793 50287
rect 193911 50169 211633 50287
rect 211751 50169 211793 50287
rect 211911 50169 229633 50287
rect 229751 50169 229793 50287
rect 229911 50169 247633 50287
rect 247751 50169 247793 50287
rect 247911 50169 265633 50287
rect 265751 50169 265793 50287
rect 265911 50169 283633 50287
rect 283751 50169 283793 50287
rect 283911 50169 295071 50287
rect 295189 50169 295231 50287
rect 295349 50169 295365 50287
rect -3403 50153 295365 50169
rect -2443 48587 294405 48603
rect -2443 48469 -2427 48587
rect -2309 48469 -2267 48587
rect -2149 48469 11773 48587
rect 11891 48469 11933 48587
rect 12051 48469 29773 48587
rect 29891 48469 29933 48587
rect 30051 48469 47773 48587
rect 47891 48469 47933 48587
rect 48051 48469 65773 48587
rect 65891 48469 65933 48587
rect 66051 48469 83773 48587
rect 83891 48469 83933 48587
rect 84051 48469 101773 48587
rect 101891 48469 101933 48587
rect 102051 48469 119773 48587
rect 119891 48469 119933 48587
rect 120051 48469 137773 48587
rect 137891 48469 137933 48587
rect 138051 48469 155773 48587
rect 155891 48469 155933 48587
rect 156051 48469 173773 48587
rect 173891 48469 173933 48587
rect 174051 48469 191773 48587
rect 191891 48469 191933 48587
rect 192051 48469 209773 48587
rect 209891 48469 209933 48587
rect 210051 48469 227773 48587
rect 227891 48469 227933 48587
rect 228051 48469 245773 48587
rect 245891 48469 245933 48587
rect 246051 48469 263773 48587
rect 263891 48469 263933 48587
rect 264051 48469 281773 48587
rect 281891 48469 281933 48587
rect 282051 48469 294111 48587
rect 294229 48469 294271 48587
rect 294389 48469 294405 48587
rect -2443 48427 294405 48469
rect -2443 48309 -2427 48427
rect -2309 48309 -2267 48427
rect -2149 48309 11773 48427
rect 11891 48309 11933 48427
rect 12051 48309 29773 48427
rect 29891 48309 29933 48427
rect 30051 48309 47773 48427
rect 47891 48309 47933 48427
rect 48051 48309 65773 48427
rect 65891 48309 65933 48427
rect 66051 48309 83773 48427
rect 83891 48309 83933 48427
rect 84051 48309 101773 48427
rect 101891 48309 101933 48427
rect 102051 48309 119773 48427
rect 119891 48309 119933 48427
rect 120051 48309 137773 48427
rect 137891 48309 137933 48427
rect 138051 48309 155773 48427
rect 155891 48309 155933 48427
rect 156051 48309 173773 48427
rect 173891 48309 173933 48427
rect 174051 48309 191773 48427
rect 191891 48309 191933 48427
rect 192051 48309 209773 48427
rect 209891 48309 209933 48427
rect 210051 48309 227773 48427
rect 227891 48309 227933 48427
rect 228051 48309 245773 48427
rect 245891 48309 245933 48427
rect 246051 48309 263773 48427
rect 263891 48309 263933 48427
rect 264051 48309 281773 48427
rect 281891 48309 281933 48427
rect 282051 48309 294111 48427
rect 294229 48309 294271 48427
rect 294389 48309 294405 48427
rect -2443 48293 294405 48309
rect -1483 46727 293445 46743
rect -1483 46609 -1467 46727
rect -1349 46609 -1307 46727
rect -1189 46609 9913 46727
rect 10031 46609 10073 46727
rect 10191 46609 27913 46727
rect 28031 46609 28073 46727
rect 28191 46609 45913 46727
rect 46031 46609 46073 46727
rect 46191 46609 63913 46727
rect 64031 46609 64073 46727
rect 64191 46609 81913 46727
rect 82031 46609 82073 46727
rect 82191 46609 99913 46727
rect 100031 46609 100073 46727
rect 100191 46609 117913 46727
rect 118031 46609 118073 46727
rect 118191 46609 135913 46727
rect 136031 46609 136073 46727
rect 136191 46609 153913 46727
rect 154031 46609 154073 46727
rect 154191 46609 171913 46727
rect 172031 46609 172073 46727
rect 172191 46609 189913 46727
rect 190031 46609 190073 46727
rect 190191 46609 207913 46727
rect 208031 46609 208073 46727
rect 208191 46609 225913 46727
rect 226031 46609 226073 46727
rect 226191 46609 243913 46727
rect 244031 46609 244073 46727
rect 244191 46609 261913 46727
rect 262031 46609 262073 46727
rect 262191 46609 279913 46727
rect 280031 46609 280073 46727
rect 280191 46609 293151 46727
rect 293269 46609 293311 46727
rect 293429 46609 293445 46727
rect -1483 46567 293445 46609
rect -1483 46449 -1467 46567
rect -1349 46449 -1307 46567
rect -1189 46449 9913 46567
rect 10031 46449 10073 46567
rect 10191 46449 27913 46567
rect 28031 46449 28073 46567
rect 28191 46449 45913 46567
rect 46031 46449 46073 46567
rect 46191 46449 63913 46567
rect 64031 46449 64073 46567
rect 64191 46449 81913 46567
rect 82031 46449 82073 46567
rect 82191 46449 99913 46567
rect 100031 46449 100073 46567
rect 100191 46449 117913 46567
rect 118031 46449 118073 46567
rect 118191 46449 135913 46567
rect 136031 46449 136073 46567
rect 136191 46449 153913 46567
rect 154031 46449 154073 46567
rect 154191 46449 171913 46567
rect 172031 46449 172073 46567
rect 172191 46449 189913 46567
rect 190031 46449 190073 46567
rect 190191 46449 207913 46567
rect 208031 46449 208073 46567
rect 208191 46449 225913 46567
rect 226031 46449 226073 46567
rect 226191 46449 243913 46567
rect 244031 46449 244073 46567
rect 244191 46449 261913 46567
rect 262031 46449 262073 46567
rect 262191 46449 279913 46567
rect 280031 46449 280073 46567
rect 280191 46449 293151 46567
rect 293269 46449 293311 46567
rect 293429 46449 293445 46567
rect -1483 46433 293445 46449
rect -4363 43307 296325 43323
rect -4363 43189 -3867 43307
rect -3749 43189 -3707 43307
rect -3589 43189 6493 43307
rect 6611 43189 6653 43307
rect 6771 43189 24493 43307
rect 24611 43189 24653 43307
rect 24771 43189 42493 43307
rect 42611 43189 42653 43307
rect 42771 43189 60493 43307
rect 60611 43189 60653 43307
rect 60771 43189 78493 43307
rect 78611 43189 78653 43307
rect 78771 43189 96493 43307
rect 96611 43189 96653 43307
rect 96771 43189 114493 43307
rect 114611 43189 114653 43307
rect 114771 43189 132493 43307
rect 132611 43189 132653 43307
rect 132771 43189 150493 43307
rect 150611 43189 150653 43307
rect 150771 43189 168493 43307
rect 168611 43189 168653 43307
rect 168771 43189 186493 43307
rect 186611 43189 186653 43307
rect 186771 43189 204493 43307
rect 204611 43189 204653 43307
rect 204771 43189 222493 43307
rect 222611 43189 222653 43307
rect 222771 43189 240493 43307
rect 240611 43189 240653 43307
rect 240771 43189 258493 43307
rect 258611 43189 258653 43307
rect 258771 43189 276493 43307
rect 276611 43189 276653 43307
rect 276771 43189 295551 43307
rect 295669 43189 295711 43307
rect 295829 43189 296325 43307
rect -4363 43147 296325 43189
rect -4363 43029 -3867 43147
rect -3749 43029 -3707 43147
rect -3589 43029 6493 43147
rect 6611 43029 6653 43147
rect 6771 43029 24493 43147
rect 24611 43029 24653 43147
rect 24771 43029 42493 43147
rect 42611 43029 42653 43147
rect 42771 43029 60493 43147
rect 60611 43029 60653 43147
rect 60771 43029 78493 43147
rect 78611 43029 78653 43147
rect 78771 43029 96493 43147
rect 96611 43029 96653 43147
rect 96771 43029 114493 43147
rect 114611 43029 114653 43147
rect 114771 43029 132493 43147
rect 132611 43029 132653 43147
rect 132771 43029 150493 43147
rect 150611 43029 150653 43147
rect 150771 43029 168493 43147
rect 168611 43029 168653 43147
rect 168771 43029 186493 43147
rect 186611 43029 186653 43147
rect 186771 43029 204493 43147
rect 204611 43029 204653 43147
rect 204771 43029 222493 43147
rect 222611 43029 222653 43147
rect 222771 43029 240493 43147
rect 240611 43029 240653 43147
rect 240771 43029 258493 43147
rect 258611 43029 258653 43147
rect 258771 43029 276493 43147
rect 276611 43029 276653 43147
rect 276771 43029 295551 43147
rect 295669 43029 295711 43147
rect 295829 43029 296325 43147
rect -4363 43013 296325 43029
rect -3403 41447 295365 41463
rect -3403 41329 -2907 41447
rect -2789 41329 -2747 41447
rect -2629 41329 4633 41447
rect 4751 41329 4793 41447
rect 4911 41329 22633 41447
rect 22751 41329 22793 41447
rect 22911 41329 40633 41447
rect 40751 41329 40793 41447
rect 40911 41329 58633 41447
rect 58751 41329 58793 41447
rect 58911 41329 76633 41447
rect 76751 41329 76793 41447
rect 76911 41329 94633 41447
rect 94751 41329 94793 41447
rect 94911 41329 112633 41447
rect 112751 41329 112793 41447
rect 112911 41329 130633 41447
rect 130751 41329 130793 41447
rect 130911 41329 148633 41447
rect 148751 41329 148793 41447
rect 148911 41329 166633 41447
rect 166751 41329 166793 41447
rect 166911 41329 184633 41447
rect 184751 41329 184793 41447
rect 184911 41329 202633 41447
rect 202751 41329 202793 41447
rect 202911 41329 220633 41447
rect 220751 41329 220793 41447
rect 220911 41329 238633 41447
rect 238751 41329 238793 41447
rect 238911 41329 256633 41447
rect 256751 41329 256793 41447
rect 256911 41329 274633 41447
rect 274751 41329 274793 41447
rect 274911 41329 294591 41447
rect 294709 41329 294751 41447
rect 294869 41329 295365 41447
rect -3403 41287 295365 41329
rect -3403 41169 -2907 41287
rect -2789 41169 -2747 41287
rect -2629 41169 4633 41287
rect 4751 41169 4793 41287
rect 4911 41169 22633 41287
rect 22751 41169 22793 41287
rect 22911 41169 40633 41287
rect 40751 41169 40793 41287
rect 40911 41169 58633 41287
rect 58751 41169 58793 41287
rect 58911 41169 76633 41287
rect 76751 41169 76793 41287
rect 76911 41169 94633 41287
rect 94751 41169 94793 41287
rect 94911 41169 112633 41287
rect 112751 41169 112793 41287
rect 112911 41169 130633 41287
rect 130751 41169 130793 41287
rect 130911 41169 148633 41287
rect 148751 41169 148793 41287
rect 148911 41169 166633 41287
rect 166751 41169 166793 41287
rect 166911 41169 184633 41287
rect 184751 41169 184793 41287
rect 184911 41169 202633 41287
rect 202751 41169 202793 41287
rect 202911 41169 220633 41287
rect 220751 41169 220793 41287
rect 220911 41169 238633 41287
rect 238751 41169 238793 41287
rect 238911 41169 256633 41287
rect 256751 41169 256793 41287
rect 256911 41169 274633 41287
rect 274751 41169 274793 41287
rect 274911 41169 294591 41287
rect 294709 41169 294751 41287
rect 294869 41169 295365 41287
rect -3403 41153 295365 41169
rect -2443 39587 294405 39603
rect -2443 39469 -1947 39587
rect -1829 39469 -1787 39587
rect -1669 39469 2773 39587
rect 2891 39469 2933 39587
rect 3051 39469 20773 39587
rect 20891 39469 20933 39587
rect 21051 39469 38773 39587
rect 38891 39469 38933 39587
rect 39051 39469 56773 39587
rect 56891 39469 56933 39587
rect 57051 39469 74773 39587
rect 74891 39469 74933 39587
rect 75051 39469 92773 39587
rect 92891 39469 92933 39587
rect 93051 39469 110773 39587
rect 110891 39469 110933 39587
rect 111051 39469 128773 39587
rect 128891 39469 128933 39587
rect 129051 39469 146773 39587
rect 146891 39469 146933 39587
rect 147051 39469 164773 39587
rect 164891 39469 164933 39587
rect 165051 39469 182773 39587
rect 182891 39469 182933 39587
rect 183051 39469 200773 39587
rect 200891 39469 200933 39587
rect 201051 39469 218773 39587
rect 218891 39469 218933 39587
rect 219051 39469 236773 39587
rect 236891 39469 236933 39587
rect 237051 39469 254773 39587
rect 254891 39469 254933 39587
rect 255051 39469 272773 39587
rect 272891 39469 272933 39587
rect 273051 39469 290773 39587
rect 290891 39469 290933 39587
rect 291051 39469 293631 39587
rect 293749 39469 293791 39587
rect 293909 39469 294405 39587
rect -2443 39427 294405 39469
rect -2443 39309 -1947 39427
rect -1829 39309 -1787 39427
rect -1669 39309 2773 39427
rect 2891 39309 2933 39427
rect 3051 39309 20773 39427
rect 20891 39309 20933 39427
rect 21051 39309 38773 39427
rect 38891 39309 38933 39427
rect 39051 39309 56773 39427
rect 56891 39309 56933 39427
rect 57051 39309 74773 39427
rect 74891 39309 74933 39427
rect 75051 39309 92773 39427
rect 92891 39309 92933 39427
rect 93051 39309 110773 39427
rect 110891 39309 110933 39427
rect 111051 39309 128773 39427
rect 128891 39309 128933 39427
rect 129051 39309 146773 39427
rect 146891 39309 146933 39427
rect 147051 39309 164773 39427
rect 164891 39309 164933 39427
rect 165051 39309 182773 39427
rect 182891 39309 182933 39427
rect 183051 39309 200773 39427
rect 200891 39309 200933 39427
rect 201051 39309 218773 39427
rect 218891 39309 218933 39427
rect 219051 39309 236773 39427
rect 236891 39309 236933 39427
rect 237051 39309 254773 39427
rect 254891 39309 254933 39427
rect 255051 39309 272773 39427
rect 272891 39309 272933 39427
rect 273051 39309 290773 39427
rect 290891 39309 290933 39427
rect 291051 39309 293631 39427
rect 293749 39309 293791 39427
rect 293909 39309 294405 39427
rect -2443 39293 294405 39309
rect -1483 37727 293445 37743
rect -1483 37609 -987 37727
rect -869 37609 -827 37727
rect -709 37609 913 37727
rect 1031 37609 1073 37727
rect 1191 37609 18913 37727
rect 19031 37609 19073 37727
rect 19191 37609 36913 37727
rect 37031 37609 37073 37727
rect 37191 37609 54913 37727
rect 55031 37609 55073 37727
rect 55191 37609 72913 37727
rect 73031 37609 73073 37727
rect 73191 37609 90913 37727
rect 91031 37609 91073 37727
rect 91191 37609 108913 37727
rect 109031 37609 109073 37727
rect 109191 37609 126913 37727
rect 127031 37609 127073 37727
rect 127191 37609 144913 37727
rect 145031 37609 145073 37727
rect 145191 37609 162913 37727
rect 163031 37609 163073 37727
rect 163191 37609 180913 37727
rect 181031 37609 181073 37727
rect 181191 37609 198913 37727
rect 199031 37609 199073 37727
rect 199191 37609 216913 37727
rect 217031 37609 217073 37727
rect 217191 37609 234913 37727
rect 235031 37609 235073 37727
rect 235191 37609 252913 37727
rect 253031 37609 253073 37727
rect 253191 37609 270913 37727
rect 271031 37609 271073 37727
rect 271191 37609 288913 37727
rect 289031 37609 289073 37727
rect 289191 37609 292671 37727
rect 292789 37609 292831 37727
rect 292949 37609 293445 37727
rect -1483 37567 293445 37609
rect -1483 37449 -987 37567
rect -869 37449 -827 37567
rect -709 37449 913 37567
rect 1031 37449 1073 37567
rect 1191 37449 18913 37567
rect 19031 37449 19073 37567
rect 19191 37449 36913 37567
rect 37031 37449 37073 37567
rect 37191 37449 54913 37567
rect 55031 37449 55073 37567
rect 55191 37449 72913 37567
rect 73031 37449 73073 37567
rect 73191 37449 90913 37567
rect 91031 37449 91073 37567
rect 91191 37449 108913 37567
rect 109031 37449 109073 37567
rect 109191 37449 126913 37567
rect 127031 37449 127073 37567
rect 127191 37449 144913 37567
rect 145031 37449 145073 37567
rect 145191 37449 162913 37567
rect 163031 37449 163073 37567
rect 163191 37449 180913 37567
rect 181031 37449 181073 37567
rect 181191 37449 198913 37567
rect 199031 37449 199073 37567
rect 199191 37449 216913 37567
rect 217031 37449 217073 37567
rect 217191 37449 234913 37567
rect 235031 37449 235073 37567
rect 235191 37449 252913 37567
rect 253031 37449 253073 37567
rect 253191 37449 270913 37567
rect 271031 37449 271073 37567
rect 271191 37449 288913 37567
rect 289031 37449 289073 37567
rect 289191 37449 292671 37567
rect 292789 37449 292831 37567
rect 292949 37449 293445 37567
rect -1483 37433 293445 37449
rect -4363 34307 296325 34323
rect -4363 34189 -4347 34307
rect -4229 34189 -4187 34307
rect -4069 34189 15493 34307
rect 15611 34189 15653 34307
rect 15771 34189 33493 34307
rect 33611 34189 33653 34307
rect 33771 34189 51493 34307
rect 51611 34189 51653 34307
rect 51771 34189 69493 34307
rect 69611 34189 69653 34307
rect 69771 34189 87493 34307
rect 87611 34189 87653 34307
rect 87771 34189 105493 34307
rect 105611 34189 105653 34307
rect 105771 34189 123493 34307
rect 123611 34189 123653 34307
rect 123771 34189 141493 34307
rect 141611 34189 141653 34307
rect 141771 34189 159493 34307
rect 159611 34189 159653 34307
rect 159771 34189 177493 34307
rect 177611 34189 177653 34307
rect 177771 34189 195493 34307
rect 195611 34189 195653 34307
rect 195771 34189 213493 34307
rect 213611 34189 213653 34307
rect 213771 34189 231493 34307
rect 231611 34189 231653 34307
rect 231771 34189 249493 34307
rect 249611 34189 249653 34307
rect 249771 34189 267493 34307
rect 267611 34189 267653 34307
rect 267771 34189 285493 34307
rect 285611 34189 285653 34307
rect 285771 34189 296031 34307
rect 296149 34189 296191 34307
rect 296309 34189 296325 34307
rect -4363 34147 296325 34189
rect -4363 34029 -4347 34147
rect -4229 34029 -4187 34147
rect -4069 34029 15493 34147
rect 15611 34029 15653 34147
rect 15771 34029 33493 34147
rect 33611 34029 33653 34147
rect 33771 34029 51493 34147
rect 51611 34029 51653 34147
rect 51771 34029 69493 34147
rect 69611 34029 69653 34147
rect 69771 34029 87493 34147
rect 87611 34029 87653 34147
rect 87771 34029 105493 34147
rect 105611 34029 105653 34147
rect 105771 34029 123493 34147
rect 123611 34029 123653 34147
rect 123771 34029 141493 34147
rect 141611 34029 141653 34147
rect 141771 34029 159493 34147
rect 159611 34029 159653 34147
rect 159771 34029 177493 34147
rect 177611 34029 177653 34147
rect 177771 34029 195493 34147
rect 195611 34029 195653 34147
rect 195771 34029 213493 34147
rect 213611 34029 213653 34147
rect 213771 34029 231493 34147
rect 231611 34029 231653 34147
rect 231771 34029 249493 34147
rect 249611 34029 249653 34147
rect 249771 34029 267493 34147
rect 267611 34029 267653 34147
rect 267771 34029 285493 34147
rect 285611 34029 285653 34147
rect 285771 34029 296031 34147
rect 296149 34029 296191 34147
rect 296309 34029 296325 34147
rect -4363 34013 296325 34029
rect -3403 32447 295365 32463
rect -3403 32329 -3387 32447
rect -3269 32329 -3227 32447
rect -3109 32329 13633 32447
rect 13751 32329 13793 32447
rect 13911 32329 31633 32447
rect 31751 32329 31793 32447
rect 31911 32329 49633 32447
rect 49751 32329 49793 32447
rect 49911 32329 67633 32447
rect 67751 32329 67793 32447
rect 67911 32329 85633 32447
rect 85751 32329 85793 32447
rect 85911 32329 103633 32447
rect 103751 32329 103793 32447
rect 103911 32329 121633 32447
rect 121751 32329 121793 32447
rect 121911 32329 139633 32447
rect 139751 32329 139793 32447
rect 139911 32329 157633 32447
rect 157751 32329 157793 32447
rect 157911 32329 175633 32447
rect 175751 32329 175793 32447
rect 175911 32329 193633 32447
rect 193751 32329 193793 32447
rect 193911 32329 211633 32447
rect 211751 32329 211793 32447
rect 211911 32329 229633 32447
rect 229751 32329 229793 32447
rect 229911 32329 247633 32447
rect 247751 32329 247793 32447
rect 247911 32329 265633 32447
rect 265751 32329 265793 32447
rect 265911 32329 283633 32447
rect 283751 32329 283793 32447
rect 283911 32329 295071 32447
rect 295189 32329 295231 32447
rect 295349 32329 295365 32447
rect -3403 32287 295365 32329
rect -3403 32169 -3387 32287
rect -3269 32169 -3227 32287
rect -3109 32169 13633 32287
rect 13751 32169 13793 32287
rect 13911 32169 31633 32287
rect 31751 32169 31793 32287
rect 31911 32169 49633 32287
rect 49751 32169 49793 32287
rect 49911 32169 67633 32287
rect 67751 32169 67793 32287
rect 67911 32169 85633 32287
rect 85751 32169 85793 32287
rect 85911 32169 103633 32287
rect 103751 32169 103793 32287
rect 103911 32169 121633 32287
rect 121751 32169 121793 32287
rect 121911 32169 139633 32287
rect 139751 32169 139793 32287
rect 139911 32169 157633 32287
rect 157751 32169 157793 32287
rect 157911 32169 175633 32287
rect 175751 32169 175793 32287
rect 175911 32169 193633 32287
rect 193751 32169 193793 32287
rect 193911 32169 211633 32287
rect 211751 32169 211793 32287
rect 211911 32169 229633 32287
rect 229751 32169 229793 32287
rect 229911 32169 247633 32287
rect 247751 32169 247793 32287
rect 247911 32169 265633 32287
rect 265751 32169 265793 32287
rect 265911 32169 283633 32287
rect 283751 32169 283793 32287
rect 283911 32169 295071 32287
rect 295189 32169 295231 32287
rect 295349 32169 295365 32287
rect -3403 32153 295365 32169
rect -2443 30587 294405 30603
rect -2443 30469 -2427 30587
rect -2309 30469 -2267 30587
rect -2149 30469 11773 30587
rect 11891 30469 11933 30587
rect 12051 30469 29773 30587
rect 29891 30469 29933 30587
rect 30051 30469 47773 30587
rect 47891 30469 47933 30587
rect 48051 30469 65773 30587
rect 65891 30469 65933 30587
rect 66051 30469 83773 30587
rect 83891 30469 83933 30587
rect 84051 30469 101773 30587
rect 101891 30469 101933 30587
rect 102051 30469 119773 30587
rect 119891 30469 119933 30587
rect 120051 30469 137773 30587
rect 137891 30469 137933 30587
rect 138051 30469 155773 30587
rect 155891 30469 155933 30587
rect 156051 30469 173773 30587
rect 173891 30469 173933 30587
rect 174051 30469 191773 30587
rect 191891 30469 191933 30587
rect 192051 30469 209773 30587
rect 209891 30469 209933 30587
rect 210051 30469 227773 30587
rect 227891 30469 227933 30587
rect 228051 30469 245773 30587
rect 245891 30469 245933 30587
rect 246051 30469 263773 30587
rect 263891 30469 263933 30587
rect 264051 30469 281773 30587
rect 281891 30469 281933 30587
rect 282051 30469 294111 30587
rect 294229 30469 294271 30587
rect 294389 30469 294405 30587
rect -2443 30427 294405 30469
rect -2443 30309 -2427 30427
rect -2309 30309 -2267 30427
rect -2149 30309 11773 30427
rect 11891 30309 11933 30427
rect 12051 30309 29773 30427
rect 29891 30309 29933 30427
rect 30051 30309 47773 30427
rect 47891 30309 47933 30427
rect 48051 30309 65773 30427
rect 65891 30309 65933 30427
rect 66051 30309 83773 30427
rect 83891 30309 83933 30427
rect 84051 30309 101773 30427
rect 101891 30309 101933 30427
rect 102051 30309 119773 30427
rect 119891 30309 119933 30427
rect 120051 30309 137773 30427
rect 137891 30309 137933 30427
rect 138051 30309 155773 30427
rect 155891 30309 155933 30427
rect 156051 30309 173773 30427
rect 173891 30309 173933 30427
rect 174051 30309 191773 30427
rect 191891 30309 191933 30427
rect 192051 30309 209773 30427
rect 209891 30309 209933 30427
rect 210051 30309 227773 30427
rect 227891 30309 227933 30427
rect 228051 30309 245773 30427
rect 245891 30309 245933 30427
rect 246051 30309 263773 30427
rect 263891 30309 263933 30427
rect 264051 30309 281773 30427
rect 281891 30309 281933 30427
rect 282051 30309 294111 30427
rect 294229 30309 294271 30427
rect 294389 30309 294405 30427
rect -2443 30293 294405 30309
rect -1483 28727 293445 28743
rect -1483 28609 -1467 28727
rect -1349 28609 -1307 28727
rect -1189 28609 9913 28727
rect 10031 28609 10073 28727
rect 10191 28609 27913 28727
rect 28031 28609 28073 28727
rect 28191 28609 45913 28727
rect 46031 28609 46073 28727
rect 46191 28609 63913 28727
rect 64031 28609 64073 28727
rect 64191 28609 81913 28727
rect 82031 28609 82073 28727
rect 82191 28609 99913 28727
rect 100031 28609 100073 28727
rect 100191 28609 117913 28727
rect 118031 28609 118073 28727
rect 118191 28609 135913 28727
rect 136031 28609 136073 28727
rect 136191 28609 153913 28727
rect 154031 28609 154073 28727
rect 154191 28609 171913 28727
rect 172031 28609 172073 28727
rect 172191 28609 189913 28727
rect 190031 28609 190073 28727
rect 190191 28609 207913 28727
rect 208031 28609 208073 28727
rect 208191 28609 225913 28727
rect 226031 28609 226073 28727
rect 226191 28609 243913 28727
rect 244031 28609 244073 28727
rect 244191 28609 261913 28727
rect 262031 28609 262073 28727
rect 262191 28609 279913 28727
rect 280031 28609 280073 28727
rect 280191 28609 293151 28727
rect 293269 28609 293311 28727
rect 293429 28609 293445 28727
rect -1483 28567 293445 28609
rect -1483 28449 -1467 28567
rect -1349 28449 -1307 28567
rect -1189 28449 9913 28567
rect 10031 28449 10073 28567
rect 10191 28449 27913 28567
rect 28031 28449 28073 28567
rect 28191 28449 45913 28567
rect 46031 28449 46073 28567
rect 46191 28449 63913 28567
rect 64031 28449 64073 28567
rect 64191 28449 81913 28567
rect 82031 28449 82073 28567
rect 82191 28449 99913 28567
rect 100031 28449 100073 28567
rect 100191 28449 117913 28567
rect 118031 28449 118073 28567
rect 118191 28449 135913 28567
rect 136031 28449 136073 28567
rect 136191 28449 153913 28567
rect 154031 28449 154073 28567
rect 154191 28449 171913 28567
rect 172031 28449 172073 28567
rect 172191 28449 189913 28567
rect 190031 28449 190073 28567
rect 190191 28449 207913 28567
rect 208031 28449 208073 28567
rect 208191 28449 225913 28567
rect 226031 28449 226073 28567
rect 226191 28449 243913 28567
rect 244031 28449 244073 28567
rect 244191 28449 261913 28567
rect 262031 28449 262073 28567
rect 262191 28449 279913 28567
rect 280031 28449 280073 28567
rect 280191 28449 293151 28567
rect 293269 28449 293311 28567
rect 293429 28449 293445 28567
rect -1483 28433 293445 28449
rect -4363 25307 296325 25323
rect -4363 25189 -3867 25307
rect -3749 25189 -3707 25307
rect -3589 25189 6493 25307
rect 6611 25189 6653 25307
rect 6771 25189 24493 25307
rect 24611 25189 24653 25307
rect 24771 25189 42493 25307
rect 42611 25189 42653 25307
rect 42771 25189 60493 25307
rect 60611 25189 60653 25307
rect 60771 25189 78493 25307
rect 78611 25189 78653 25307
rect 78771 25189 96493 25307
rect 96611 25189 96653 25307
rect 96771 25189 114493 25307
rect 114611 25189 114653 25307
rect 114771 25189 132493 25307
rect 132611 25189 132653 25307
rect 132771 25189 150493 25307
rect 150611 25189 150653 25307
rect 150771 25189 168493 25307
rect 168611 25189 168653 25307
rect 168771 25189 186493 25307
rect 186611 25189 186653 25307
rect 186771 25189 204493 25307
rect 204611 25189 204653 25307
rect 204771 25189 222493 25307
rect 222611 25189 222653 25307
rect 222771 25189 240493 25307
rect 240611 25189 240653 25307
rect 240771 25189 258493 25307
rect 258611 25189 258653 25307
rect 258771 25189 276493 25307
rect 276611 25189 276653 25307
rect 276771 25189 295551 25307
rect 295669 25189 295711 25307
rect 295829 25189 296325 25307
rect -4363 25147 296325 25189
rect -4363 25029 -3867 25147
rect -3749 25029 -3707 25147
rect -3589 25029 6493 25147
rect 6611 25029 6653 25147
rect 6771 25029 24493 25147
rect 24611 25029 24653 25147
rect 24771 25029 42493 25147
rect 42611 25029 42653 25147
rect 42771 25029 60493 25147
rect 60611 25029 60653 25147
rect 60771 25029 78493 25147
rect 78611 25029 78653 25147
rect 78771 25029 96493 25147
rect 96611 25029 96653 25147
rect 96771 25029 114493 25147
rect 114611 25029 114653 25147
rect 114771 25029 132493 25147
rect 132611 25029 132653 25147
rect 132771 25029 150493 25147
rect 150611 25029 150653 25147
rect 150771 25029 168493 25147
rect 168611 25029 168653 25147
rect 168771 25029 186493 25147
rect 186611 25029 186653 25147
rect 186771 25029 204493 25147
rect 204611 25029 204653 25147
rect 204771 25029 222493 25147
rect 222611 25029 222653 25147
rect 222771 25029 240493 25147
rect 240611 25029 240653 25147
rect 240771 25029 258493 25147
rect 258611 25029 258653 25147
rect 258771 25029 276493 25147
rect 276611 25029 276653 25147
rect 276771 25029 295551 25147
rect 295669 25029 295711 25147
rect 295829 25029 296325 25147
rect -4363 25013 296325 25029
rect -3403 23447 295365 23463
rect -3403 23329 -2907 23447
rect -2789 23329 -2747 23447
rect -2629 23329 4633 23447
rect 4751 23329 4793 23447
rect 4911 23329 22633 23447
rect 22751 23329 22793 23447
rect 22911 23329 40633 23447
rect 40751 23329 40793 23447
rect 40911 23329 58633 23447
rect 58751 23329 58793 23447
rect 58911 23329 76633 23447
rect 76751 23329 76793 23447
rect 76911 23329 94633 23447
rect 94751 23329 94793 23447
rect 94911 23329 112633 23447
rect 112751 23329 112793 23447
rect 112911 23329 130633 23447
rect 130751 23329 130793 23447
rect 130911 23329 148633 23447
rect 148751 23329 148793 23447
rect 148911 23329 166633 23447
rect 166751 23329 166793 23447
rect 166911 23329 184633 23447
rect 184751 23329 184793 23447
rect 184911 23329 202633 23447
rect 202751 23329 202793 23447
rect 202911 23329 220633 23447
rect 220751 23329 220793 23447
rect 220911 23329 238633 23447
rect 238751 23329 238793 23447
rect 238911 23329 256633 23447
rect 256751 23329 256793 23447
rect 256911 23329 274633 23447
rect 274751 23329 274793 23447
rect 274911 23329 294591 23447
rect 294709 23329 294751 23447
rect 294869 23329 295365 23447
rect -3403 23287 295365 23329
rect -3403 23169 -2907 23287
rect -2789 23169 -2747 23287
rect -2629 23169 4633 23287
rect 4751 23169 4793 23287
rect 4911 23169 22633 23287
rect 22751 23169 22793 23287
rect 22911 23169 40633 23287
rect 40751 23169 40793 23287
rect 40911 23169 58633 23287
rect 58751 23169 58793 23287
rect 58911 23169 76633 23287
rect 76751 23169 76793 23287
rect 76911 23169 94633 23287
rect 94751 23169 94793 23287
rect 94911 23169 112633 23287
rect 112751 23169 112793 23287
rect 112911 23169 130633 23287
rect 130751 23169 130793 23287
rect 130911 23169 148633 23287
rect 148751 23169 148793 23287
rect 148911 23169 166633 23287
rect 166751 23169 166793 23287
rect 166911 23169 184633 23287
rect 184751 23169 184793 23287
rect 184911 23169 202633 23287
rect 202751 23169 202793 23287
rect 202911 23169 220633 23287
rect 220751 23169 220793 23287
rect 220911 23169 238633 23287
rect 238751 23169 238793 23287
rect 238911 23169 256633 23287
rect 256751 23169 256793 23287
rect 256911 23169 274633 23287
rect 274751 23169 274793 23287
rect 274911 23169 294591 23287
rect 294709 23169 294751 23287
rect 294869 23169 295365 23287
rect -3403 23153 295365 23169
rect -2443 21587 294405 21603
rect -2443 21469 -1947 21587
rect -1829 21469 -1787 21587
rect -1669 21469 2773 21587
rect 2891 21469 2933 21587
rect 3051 21469 20773 21587
rect 20891 21469 20933 21587
rect 21051 21469 38773 21587
rect 38891 21469 38933 21587
rect 39051 21469 56773 21587
rect 56891 21469 56933 21587
rect 57051 21469 74773 21587
rect 74891 21469 74933 21587
rect 75051 21469 92773 21587
rect 92891 21469 92933 21587
rect 93051 21469 110773 21587
rect 110891 21469 110933 21587
rect 111051 21469 128773 21587
rect 128891 21469 128933 21587
rect 129051 21469 146773 21587
rect 146891 21469 146933 21587
rect 147051 21469 164773 21587
rect 164891 21469 164933 21587
rect 165051 21469 182773 21587
rect 182891 21469 182933 21587
rect 183051 21469 200773 21587
rect 200891 21469 200933 21587
rect 201051 21469 218773 21587
rect 218891 21469 218933 21587
rect 219051 21469 236773 21587
rect 236891 21469 236933 21587
rect 237051 21469 254773 21587
rect 254891 21469 254933 21587
rect 255051 21469 272773 21587
rect 272891 21469 272933 21587
rect 273051 21469 290773 21587
rect 290891 21469 290933 21587
rect 291051 21469 293631 21587
rect 293749 21469 293791 21587
rect 293909 21469 294405 21587
rect -2443 21427 294405 21469
rect -2443 21309 -1947 21427
rect -1829 21309 -1787 21427
rect -1669 21309 2773 21427
rect 2891 21309 2933 21427
rect 3051 21309 20773 21427
rect 20891 21309 20933 21427
rect 21051 21309 38773 21427
rect 38891 21309 38933 21427
rect 39051 21309 56773 21427
rect 56891 21309 56933 21427
rect 57051 21309 74773 21427
rect 74891 21309 74933 21427
rect 75051 21309 92773 21427
rect 92891 21309 92933 21427
rect 93051 21309 110773 21427
rect 110891 21309 110933 21427
rect 111051 21309 128773 21427
rect 128891 21309 128933 21427
rect 129051 21309 146773 21427
rect 146891 21309 146933 21427
rect 147051 21309 164773 21427
rect 164891 21309 164933 21427
rect 165051 21309 182773 21427
rect 182891 21309 182933 21427
rect 183051 21309 200773 21427
rect 200891 21309 200933 21427
rect 201051 21309 218773 21427
rect 218891 21309 218933 21427
rect 219051 21309 236773 21427
rect 236891 21309 236933 21427
rect 237051 21309 254773 21427
rect 254891 21309 254933 21427
rect 255051 21309 272773 21427
rect 272891 21309 272933 21427
rect 273051 21309 290773 21427
rect 290891 21309 290933 21427
rect 291051 21309 293631 21427
rect 293749 21309 293791 21427
rect 293909 21309 294405 21427
rect -2443 21293 294405 21309
rect -1483 19727 293445 19743
rect -1483 19609 -987 19727
rect -869 19609 -827 19727
rect -709 19609 913 19727
rect 1031 19609 1073 19727
rect 1191 19609 18913 19727
rect 19031 19609 19073 19727
rect 19191 19609 36913 19727
rect 37031 19609 37073 19727
rect 37191 19609 54913 19727
rect 55031 19609 55073 19727
rect 55191 19609 72913 19727
rect 73031 19609 73073 19727
rect 73191 19609 90913 19727
rect 91031 19609 91073 19727
rect 91191 19609 108913 19727
rect 109031 19609 109073 19727
rect 109191 19609 126913 19727
rect 127031 19609 127073 19727
rect 127191 19609 144913 19727
rect 145031 19609 145073 19727
rect 145191 19609 162913 19727
rect 163031 19609 163073 19727
rect 163191 19609 180913 19727
rect 181031 19609 181073 19727
rect 181191 19609 198913 19727
rect 199031 19609 199073 19727
rect 199191 19609 216913 19727
rect 217031 19609 217073 19727
rect 217191 19609 234913 19727
rect 235031 19609 235073 19727
rect 235191 19609 252913 19727
rect 253031 19609 253073 19727
rect 253191 19609 270913 19727
rect 271031 19609 271073 19727
rect 271191 19609 288913 19727
rect 289031 19609 289073 19727
rect 289191 19609 292671 19727
rect 292789 19609 292831 19727
rect 292949 19609 293445 19727
rect -1483 19567 293445 19609
rect -1483 19449 -987 19567
rect -869 19449 -827 19567
rect -709 19449 913 19567
rect 1031 19449 1073 19567
rect 1191 19449 18913 19567
rect 19031 19449 19073 19567
rect 19191 19449 36913 19567
rect 37031 19449 37073 19567
rect 37191 19449 54913 19567
rect 55031 19449 55073 19567
rect 55191 19449 72913 19567
rect 73031 19449 73073 19567
rect 73191 19449 90913 19567
rect 91031 19449 91073 19567
rect 91191 19449 108913 19567
rect 109031 19449 109073 19567
rect 109191 19449 126913 19567
rect 127031 19449 127073 19567
rect 127191 19449 144913 19567
rect 145031 19449 145073 19567
rect 145191 19449 162913 19567
rect 163031 19449 163073 19567
rect 163191 19449 180913 19567
rect 181031 19449 181073 19567
rect 181191 19449 198913 19567
rect 199031 19449 199073 19567
rect 199191 19449 216913 19567
rect 217031 19449 217073 19567
rect 217191 19449 234913 19567
rect 235031 19449 235073 19567
rect 235191 19449 252913 19567
rect 253031 19449 253073 19567
rect 253191 19449 270913 19567
rect 271031 19449 271073 19567
rect 271191 19449 288913 19567
rect 289031 19449 289073 19567
rect 289191 19449 292671 19567
rect 292789 19449 292831 19567
rect 292949 19449 293445 19567
rect -1483 19433 293445 19449
rect -4363 16307 296325 16323
rect -4363 16189 -4347 16307
rect -4229 16189 -4187 16307
rect -4069 16189 15493 16307
rect 15611 16189 15653 16307
rect 15771 16189 33493 16307
rect 33611 16189 33653 16307
rect 33771 16189 51493 16307
rect 51611 16189 51653 16307
rect 51771 16189 69493 16307
rect 69611 16189 69653 16307
rect 69771 16189 87493 16307
rect 87611 16189 87653 16307
rect 87771 16189 105493 16307
rect 105611 16189 105653 16307
rect 105771 16189 123493 16307
rect 123611 16189 123653 16307
rect 123771 16189 141493 16307
rect 141611 16189 141653 16307
rect 141771 16189 159493 16307
rect 159611 16189 159653 16307
rect 159771 16189 177493 16307
rect 177611 16189 177653 16307
rect 177771 16189 195493 16307
rect 195611 16189 195653 16307
rect 195771 16189 213493 16307
rect 213611 16189 213653 16307
rect 213771 16189 231493 16307
rect 231611 16189 231653 16307
rect 231771 16189 249493 16307
rect 249611 16189 249653 16307
rect 249771 16189 267493 16307
rect 267611 16189 267653 16307
rect 267771 16189 285493 16307
rect 285611 16189 285653 16307
rect 285771 16189 296031 16307
rect 296149 16189 296191 16307
rect 296309 16189 296325 16307
rect -4363 16147 296325 16189
rect -4363 16029 -4347 16147
rect -4229 16029 -4187 16147
rect -4069 16029 15493 16147
rect 15611 16029 15653 16147
rect 15771 16029 33493 16147
rect 33611 16029 33653 16147
rect 33771 16029 51493 16147
rect 51611 16029 51653 16147
rect 51771 16029 69493 16147
rect 69611 16029 69653 16147
rect 69771 16029 87493 16147
rect 87611 16029 87653 16147
rect 87771 16029 105493 16147
rect 105611 16029 105653 16147
rect 105771 16029 123493 16147
rect 123611 16029 123653 16147
rect 123771 16029 141493 16147
rect 141611 16029 141653 16147
rect 141771 16029 159493 16147
rect 159611 16029 159653 16147
rect 159771 16029 177493 16147
rect 177611 16029 177653 16147
rect 177771 16029 195493 16147
rect 195611 16029 195653 16147
rect 195771 16029 213493 16147
rect 213611 16029 213653 16147
rect 213771 16029 231493 16147
rect 231611 16029 231653 16147
rect 231771 16029 249493 16147
rect 249611 16029 249653 16147
rect 249771 16029 267493 16147
rect 267611 16029 267653 16147
rect 267771 16029 285493 16147
rect 285611 16029 285653 16147
rect 285771 16029 296031 16147
rect 296149 16029 296191 16147
rect 296309 16029 296325 16147
rect -4363 16013 296325 16029
rect -3403 14447 295365 14463
rect -3403 14329 -3387 14447
rect -3269 14329 -3227 14447
rect -3109 14329 13633 14447
rect 13751 14329 13793 14447
rect 13911 14329 31633 14447
rect 31751 14329 31793 14447
rect 31911 14329 49633 14447
rect 49751 14329 49793 14447
rect 49911 14329 67633 14447
rect 67751 14329 67793 14447
rect 67911 14329 85633 14447
rect 85751 14329 85793 14447
rect 85911 14329 103633 14447
rect 103751 14329 103793 14447
rect 103911 14329 121633 14447
rect 121751 14329 121793 14447
rect 121911 14329 139633 14447
rect 139751 14329 139793 14447
rect 139911 14329 157633 14447
rect 157751 14329 157793 14447
rect 157911 14329 175633 14447
rect 175751 14329 175793 14447
rect 175911 14329 193633 14447
rect 193751 14329 193793 14447
rect 193911 14329 211633 14447
rect 211751 14329 211793 14447
rect 211911 14329 229633 14447
rect 229751 14329 229793 14447
rect 229911 14329 247633 14447
rect 247751 14329 247793 14447
rect 247911 14329 265633 14447
rect 265751 14329 265793 14447
rect 265911 14329 283633 14447
rect 283751 14329 283793 14447
rect 283911 14329 295071 14447
rect 295189 14329 295231 14447
rect 295349 14329 295365 14447
rect -3403 14287 295365 14329
rect -3403 14169 -3387 14287
rect -3269 14169 -3227 14287
rect -3109 14169 13633 14287
rect 13751 14169 13793 14287
rect 13911 14169 31633 14287
rect 31751 14169 31793 14287
rect 31911 14169 49633 14287
rect 49751 14169 49793 14287
rect 49911 14169 67633 14287
rect 67751 14169 67793 14287
rect 67911 14169 85633 14287
rect 85751 14169 85793 14287
rect 85911 14169 103633 14287
rect 103751 14169 103793 14287
rect 103911 14169 121633 14287
rect 121751 14169 121793 14287
rect 121911 14169 139633 14287
rect 139751 14169 139793 14287
rect 139911 14169 157633 14287
rect 157751 14169 157793 14287
rect 157911 14169 175633 14287
rect 175751 14169 175793 14287
rect 175911 14169 193633 14287
rect 193751 14169 193793 14287
rect 193911 14169 211633 14287
rect 211751 14169 211793 14287
rect 211911 14169 229633 14287
rect 229751 14169 229793 14287
rect 229911 14169 247633 14287
rect 247751 14169 247793 14287
rect 247911 14169 265633 14287
rect 265751 14169 265793 14287
rect 265911 14169 283633 14287
rect 283751 14169 283793 14287
rect 283911 14169 295071 14287
rect 295189 14169 295231 14287
rect 295349 14169 295365 14287
rect -3403 14153 295365 14169
rect -2443 12587 294405 12603
rect -2443 12469 -2427 12587
rect -2309 12469 -2267 12587
rect -2149 12469 11773 12587
rect 11891 12469 11933 12587
rect 12051 12469 29773 12587
rect 29891 12469 29933 12587
rect 30051 12469 47773 12587
rect 47891 12469 47933 12587
rect 48051 12469 65773 12587
rect 65891 12469 65933 12587
rect 66051 12469 83773 12587
rect 83891 12469 83933 12587
rect 84051 12469 101773 12587
rect 101891 12469 101933 12587
rect 102051 12469 119773 12587
rect 119891 12469 119933 12587
rect 120051 12469 137773 12587
rect 137891 12469 137933 12587
rect 138051 12469 155773 12587
rect 155891 12469 155933 12587
rect 156051 12469 173773 12587
rect 173891 12469 173933 12587
rect 174051 12469 191773 12587
rect 191891 12469 191933 12587
rect 192051 12469 209773 12587
rect 209891 12469 209933 12587
rect 210051 12469 227773 12587
rect 227891 12469 227933 12587
rect 228051 12469 245773 12587
rect 245891 12469 245933 12587
rect 246051 12469 263773 12587
rect 263891 12469 263933 12587
rect 264051 12469 281773 12587
rect 281891 12469 281933 12587
rect 282051 12469 294111 12587
rect 294229 12469 294271 12587
rect 294389 12469 294405 12587
rect -2443 12427 294405 12469
rect -2443 12309 -2427 12427
rect -2309 12309 -2267 12427
rect -2149 12309 11773 12427
rect 11891 12309 11933 12427
rect 12051 12309 29773 12427
rect 29891 12309 29933 12427
rect 30051 12309 47773 12427
rect 47891 12309 47933 12427
rect 48051 12309 65773 12427
rect 65891 12309 65933 12427
rect 66051 12309 83773 12427
rect 83891 12309 83933 12427
rect 84051 12309 101773 12427
rect 101891 12309 101933 12427
rect 102051 12309 119773 12427
rect 119891 12309 119933 12427
rect 120051 12309 137773 12427
rect 137891 12309 137933 12427
rect 138051 12309 155773 12427
rect 155891 12309 155933 12427
rect 156051 12309 173773 12427
rect 173891 12309 173933 12427
rect 174051 12309 191773 12427
rect 191891 12309 191933 12427
rect 192051 12309 209773 12427
rect 209891 12309 209933 12427
rect 210051 12309 227773 12427
rect 227891 12309 227933 12427
rect 228051 12309 245773 12427
rect 245891 12309 245933 12427
rect 246051 12309 263773 12427
rect 263891 12309 263933 12427
rect 264051 12309 281773 12427
rect 281891 12309 281933 12427
rect 282051 12309 294111 12427
rect 294229 12309 294271 12427
rect 294389 12309 294405 12427
rect -2443 12293 294405 12309
rect -1483 10727 293445 10743
rect -1483 10609 -1467 10727
rect -1349 10609 -1307 10727
rect -1189 10609 9913 10727
rect 10031 10609 10073 10727
rect 10191 10609 27913 10727
rect 28031 10609 28073 10727
rect 28191 10609 45913 10727
rect 46031 10609 46073 10727
rect 46191 10609 63913 10727
rect 64031 10609 64073 10727
rect 64191 10609 81913 10727
rect 82031 10609 82073 10727
rect 82191 10609 99913 10727
rect 100031 10609 100073 10727
rect 100191 10609 117913 10727
rect 118031 10609 118073 10727
rect 118191 10609 135913 10727
rect 136031 10609 136073 10727
rect 136191 10609 153913 10727
rect 154031 10609 154073 10727
rect 154191 10609 171913 10727
rect 172031 10609 172073 10727
rect 172191 10609 189913 10727
rect 190031 10609 190073 10727
rect 190191 10609 207913 10727
rect 208031 10609 208073 10727
rect 208191 10609 225913 10727
rect 226031 10609 226073 10727
rect 226191 10609 243913 10727
rect 244031 10609 244073 10727
rect 244191 10609 261913 10727
rect 262031 10609 262073 10727
rect 262191 10609 279913 10727
rect 280031 10609 280073 10727
rect 280191 10609 293151 10727
rect 293269 10609 293311 10727
rect 293429 10609 293445 10727
rect -1483 10567 293445 10609
rect -1483 10449 -1467 10567
rect -1349 10449 -1307 10567
rect -1189 10449 9913 10567
rect 10031 10449 10073 10567
rect 10191 10449 27913 10567
rect 28031 10449 28073 10567
rect 28191 10449 45913 10567
rect 46031 10449 46073 10567
rect 46191 10449 63913 10567
rect 64031 10449 64073 10567
rect 64191 10449 81913 10567
rect 82031 10449 82073 10567
rect 82191 10449 99913 10567
rect 100031 10449 100073 10567
rect 100191 10449 117913 10567
rect 118031 10449 118073 10567
rect 118191 10449 135913 10567
rect 136031 10449 136073 10567
rect 136191 10449 153913 10567
rect 154031 10449 154073 10567
rect 154191 10449 171913 10567
rect 172031 10449 172073 10567
rect 172191 10449 189913 10567
rect 190031 10449 190073 10567
rect 190191 10449 207913 10567
rect 208031 10449 208073 10567
rect 208191 10449 225913 10567
rect 226031 10449 226073 10567
rect 226191 10449 243913 10567
rect 244031 10449 244073 10567
rect 244191 10449 261913 10567
rect 262031 10449 262073 10567
rect 262191 10449 279913 10567
rect 280031 10449 280073 10567
rect 280191 10449 293151 10567
rect 293269 10449 293311 10567
rect 293429 10449 293445 10567
rect -1483 10433 293445 10449
rect -4363 7307 296325 7323
rect -4363 7189 -3867 7307
rect -3749 7189 -3707 7307
rect -3589 7189 6493 7307
rect 6611 7189 6653 7307
rect 6771 7189 24493 7307
rect 24611 7189 24653 7307
rect 24771 7189 42493 7307
rect 42611 7189 42653 7307
rect 42771 7189 60493 7307
rect 60611 7189 60653 7307
rect 60771 7189 78493 7307
rect 78611 7189 78653 7307
rect 78771 7189 96493 7307
rect 96611 7189 96653 7307
rect 96771 7189 114493 7307
rect 114611 7189 114653 7307
rect 114771 7189 132493 7307
rect 132611 7189 132653 7307
rect 132771 7189 150493 7307
rect 150611 7189 150653 7307
rect 150771 7189 168493 7307
rect 168611 7189 168653 7307
rect 168771 7189 186493 7307
rect 186611 7189 186653 7307
rect 186771 7189 204493 7307
rect 204611 7189 204653 7307
rect 204771 7189 222493 7307
rect 222611 7189 222653 7307
rect 222771 7189 240493 7307
rect 240611 7189 240653 7307
rect 240771 7189 258493 7307
rect 258611 7189 258653 7307
rect 258771 7189 276493 7307
rect 276611 7189 276653 7307
rect 276771 7189 295551 7307
rect 295669 7189 295711 7307
rect 295829 7189 296325 7307
rect -4363 7147 296325 7189
rect -4363 7029 -3867 7147
rect -3749 7029 -3707 7147
rect -3589 7029 6493 7147
rect 6611 7029 6653 7147
rect 6771 7029 24493 7147
rect 24611 7029 24653 7147
rect 24771 7029 42493 7147
rect 42611 7029 42653 7147
rect 42771 7029 60493 7147
rect 60611 7029 60653 7147
rect 60771 7029 78493 7147
rect 78611 7029 78653 7147
rect 78771 7029 96493 7147
rect 96611 7029 96653 7147
rect 96771 7029 114493 7147
rect 114611 7029 114653 7147
rect 114771 7029 132493 7147
rect 132611 7029 132653 7147
rect 132771 7029 150493 7147
rect 150611 7029 150653 7147
rect 150771 7029 168493 7147
rect 168611 7029 168653 7147
rect 168771 7029 186493 7147
rect 186611 7029 186653 7147
rect 186771 7029 204493 7147
rect 204611 7029 204653 7147
rect 204771 7029 222493 7147
rect 222611 7029 222653 7147
rect 222771 7029 240493 7147
rect 240611 7029 240653 7147
rect 240771 7029 258493 7147
rect 258611 7029 258653 7147
rect 258771 7029 276493 7147
rect 276611 7029 276653 7147
rect 276771 7029 295551 7147
rect 295669 7029 295711 7147
rect 295829 7029 296325 7147
rect -4363 7013 296325 7029
rect -3403 5447 295365 5463
rect -3403 5329 -2907 5447
rect -2789 5329 -2747 5447
rect -2629 5329 4633 5447
rect 4751 5329 4793 5447
rect 4911 5329 22633 5447
rect 22751 5329 22793 5447
rect 22911 5329 40633 5447
rect 40751 5329 40793 5447
rect 40911 5329 58633 5447
rect 58751 5329 58793 5447
rect 58911 5329 76633 5447
rect 76751 5329 76793 5447
rect 76911 5329 94633 5447
rect 94751 5329 94793 5447
rect 94911 5329 112633 5447
rect 112751 5329 112793 5447
rect 112911 5329 130633 5447
rect 130751 5329 130793 5447
rect 130911 5329 148633 5447
rect 148751 5329 148793 5447
rect 148911 5329 166633 5447
rect 166751 5329 166793 5447
rect 166911 5329 184633 5447
rect 184751 5329 184793 5447
rect 184911 5329 202633 5447
rect 202751 5329 202793 5447
rect 202911 5329 220633 5447
rect 220751 5329 220793 5447
rect 220911 5329 238633 5447
rect 238751 5329 238793 5447
rect 238911 5329 256633 5447
rect 256751 5329 256793 5447
rect 256911 5329 274633 5447
rect 274751 5329 274793 5447
rect 274911 5329 294591 5447
rect 294709 5329 294751 5447
rect 294869 5329 295365 5447
rect -3403 5287 295365 5329
rect -3403 5169 -2907 5287
rect -2789 5169 -2747 5287
rect -2629 5169 4633 5287
rect 4751 5169 4793 5287
rect 4911 5169 22633 5287
rect 22751 5169 22793 5287
rect 22911 5169 40633 5287
rect 40751 5169 40793 5287
rect 40911 5169 58633 5287
rect 58751 5169 58793 5287
rect 58911 5169 76633 5287
rect 76751 5169 76793 5287
rect 76911 5169 94633 5287
rect 94751 5169 94793 5287
rect 94911 5169 112633 5287
rect 112751 5169 112793 5287
rect 112911 5169 130633 5287
rect 130751 5169 130793 5287
rect 130911 5169 148633 5287
rect 148751 5169 148793 5287
rect 148911 5169 166633 5287
rect 166751 5169 166793 5287
rect 166911 5169 184633 5287
rect 184751 5169 184793 5287
rect 184911 5169 202633 5287
rect 202751 5169 202793 5287
rect 202911 5169 220633 5287
rect 220751 5169 220793 5287
rect 220911 5169 238633 5287
rect 238751 5169 238793 5287
rect 238911 5169 256633 5287
rect 256751 5169 256793 5287
rect 256911 5169 274633 5287
rect 274751 5169 274793 5287
rect 274911 5169 294591 5287
rect 294709 5169 294751 5287
rect 294869 5169 295365 5287
rect -3403 5153 295365 5169
rect -2443 3587 294405 3603
rect -2443 3469 -1947 3587
rect -1829 3469 -1787 3587
rect -1669 3469 2773 3587
rect 2891 3469 2933 3587
rect 3051 3469 20773 3587
rect 20891 3469 20933 3587
rect 21051 3469 38773 3587
rect 38891 3469 38933 3587
rect 39051 3469 56773 3587
rect 56891 3469 56933 3587
rect 57051 3469 74773 3587
rect 74891 3469 74933 3587
rect 75051 3469 92773 3587
rect 92891 3469 92933 3587
rect 93051 3469 110773 3587
rect 110891 3469 110933 3587
rect 111051 3469 128773 3587
rect 128891 3469 128933 3587
rect 129051 3469 146773 3587
rect 146891 3469 146933 3587
rect 147051 3469 164773 3587
rect 164891 3469 164933 3587
rect 165051 3469 182773 3587
rect 182891 3469 182933 3587
rect 183051 3469 200773 3587
rect 200891 3469 200933 3587
rect 201051 3469 218773 3587
rect 218891 3469 218933 3587
rect 219051 3469 236773 3587
rect 236891 3469 236933 3587
rect 237051 3469 254773 3587
rect 254891 3469 254933 3587
rect 255051 3469 272773 3587
rect 272891 3469 272933 3587
rect 273051 3469 290773 3587
rect 290891 3469 290933 3587
rect 291051 3469 293631 3587
rect 293749 3469 293791 3587
rect 293909 3469 294405 3587
rect -2443 3427 294405 3469
rect -2443 3309 -1947 3427
rect -1829 3309 -1787 3427
rect -1669 3309 2773 3427
rect 2891 3309 2933 3427
rect 3051 3309 20773 3427
rect 20891 3309 20933 3427
rect 21051 3309 38773 3427
rect 38891 3309 38933 3427
rect 39051 3309 56773 3427
rect 56891 3309 56933 3427
rect 57051 3309 74773 3427
rect 74891 3309 74933 3427
rect 75051 3309 92773 3427
rect 92891 3309 92933 3427
rect 93051 3309 110773 3427
rect 110891 3309 110933 3427
rect 111051 3309 128773 3427
rect 128891 3309 128933 3427
rect 129051 3309 146773 3427
rect 146891 3309 146933 3427
rect 147051 3309 164773 3427
rect 164891 3309 164933 3427
rect 165051 3309 182773 3427
rect 182891 3309 182933 3427
rect 183051 3309 200773 3427
rect 200891 3309 200933 3427
rect 201051 3309 218773 3427
rect 218891 3309 218933 3427
rect 219051 3309 236773 3427
rect 236891 3309 236933 3427
rect 237051 3309 254773 3427
rect 254891 3309 254933 3427
rect 255051 3309 272773 3427
rect 272891 3309 272933 3427
rect 273051 3309 290773 3427
rect 290891 3309 290933 3427
rect 291051 3309 293631 3427
rect 293749 3309 293791 3427
rect 293909 3309 294405 3427
rect -2443 3293 294405 3309
rect -1483 1727 293445 1743
rect -1483 1609 -987 1727
rect -869 1609 -827 1727
rect -709 1609 913 1727
rect 1031 1609 1073 1727
rect 1191 1609 18913 1727
rect 19031 1609 19073 1727
rect 19191 1609 36913 1727
rect 37031 1609 37073 1727
rect 37191 1609 54913 1727
rect 55031 1609 55073 1727
rect 55191 1609 72913 1727
rect 73031 1609 73073 1727
rect 73191 1609 90913 1727
rect 91031 1609 91073 1727
rect 91191 1609 108913 1727
rect 109031 1609 109073 1727
rect 109191 1609 126913 1727
rect 127031 1609 127073 1727
rect 127191 1609 144913 1727
rect 145031 1609 145073 1727
rect 145191 1609 162913 1727
rect 163031 1609 163073 1727
rect 163191 1609 180913 1727
rect 181031 1609 181073 1727
rect 181191 1609 198913 1727
rect 199031 1609 199073 1727
rect 199191 1609 216913 1727
rect 217031 1609 217073 1727
rect 217191 1609 234913 1727
rect 235031 1609 235073 1727
rect 235191 1609 252913 1727
rect 253031 1609 253073 1727
rect 253191 1609 270913 1727
rect 271031 1609 271073 1727
rect 271191 1609 288913 1727
rect 289031 1609 289073 1727
rect 289191 1609 292671 1727
rect 292789 1609 292831 1727
rect 292949 1609 293445 1727
rect -1483 1567 293445 1609
rect -1483 1449 -987 1567
rect -869 1449 -827 1567
rect -709 1449 913 1567
rect 1031 1449 1073 1567
rect 1191 1449 18913 1567
rect 19031 1449 19073 1567
rect 19191 1449 36913 1567
rect 37031 1449 37073 1567
rect 37191 1449 54913 1567
rect 55031 1449 55073 1567
rect 55191 1449 72913 1567
rect 73031 1449 73073 1567
rect 73191 1449 90913 1567
rect 91031 1449 91073 1567
rect 91191 1449 108913 1567
rect 109031 1449 109073 1567
rect 109191 1449 126913 1567
rect 127031 1449 127073 1567
rect 127191 1449 144913 1567
rect 145031 1449 145073 1567
rect 145191 1449 162913 1567
rect 163031 1449 163073 1567
rect 163191 1449 180913 1567
rect 181031 1449 181073 1567
rect 181191 1449 198913 1567
rect 199031 1449 199073 1567
rect 199191 1449 216913 1567
rect 217031 1449 217073 1567
rect 217191 1449 234913 1567
rect 235031 1449 235073 1567
rect 235191 1449 252913 1567
rect 253031 1449 253073 1567
rect 253191 1449 270913 1567
rect 271031 1449 271073 1567
rect 271191 1449 288913 1567
rect 289031 1449 289073 1567
rect 289191 1449 292671 1567
rect 292789 1449 292831 1567
rect 292949 1449 293445 1567
rect -1483 1433 293445 1449
rect -1003 -173 292965 -157
rect -1003 -291 -987 -173
rect -869 -291 -827 -173
rect -709 -291 913 -173
rect 1031 -291 1073 -173
rect 1191 -291 18913 -173
rect 19031 -291 19073 -173
rect 19191 -291 36913 -173
rect 37031 -291 37073 -173
rect 37191 -291 54913 -173
rect 55031 -291 55073 -173
rect 55191 -291 72913 -173
rect 73031 -291 73073 -173
rect 73191 -291 90913 -173
rect 91031 -291 91073 -173
rect 91191 -291 108913 -173
rect 109031 -291 109073 -173
rect 109191 -291 126913 -173
rect 127031 -291 127073 -173
rect 127191 -291 144913 -173
rect 145031 -291 145073 -173
rect 145191 -291 162913 -173
rect 163031 -291 163073 -173
rect 163191 -291 180913 -173
rect 181031 -291 181073 -173
rect 181191 -291 198913 -173
rect 199031 -291 199073 -173
rect 199191 -291 216913 -173
rect 217031 -291 217073 -173
rect 217191 -291 234913 -173
rect 235031 -291 235073 -173
rect 235191 -291 252913 -173
rect 253031 -291 253073 -173
rect 253191 -291 270913 -173
rect 271031 -291 271073 -173
rect 271191 -291 288913 -173
rect 289031 -291 289073 -173
rect 289191 -291 292671 -173
rect 292789 -291 292831 -173
rect 292949 -291 292965 -173
rect -1003 -333 292965 -291
rect -1003 -451 -987 -333
rect -869 -451 -827 -333
rect -709 -451 913 -333
rect 1031 -451 1073 -333
rect 1191 -451 18913 -333
rect 19031 -451 19073 -333
rect 19191 -451 36913 -333
rect 37031 -451 37073 -333
rect 37191 -451 54913 -333
rect 55031 -451 55073 -333
rect 55191 -451 72913 -333
rect 73031 -451 73073 -333
rect 73191 -451 90913 -333
rect 91031 -451 91073 -333
rect 91191 -451 108913 -333
rect 109031 -451 109073 -333
rect 109191 -451 126913 -333
rect 127031 -451 127073 -333
rect 127191 -451 144913 -333
rect 145031 -451 145073 -333
rect 145191 -451 162913 -333
rect 163031 -451 163073 -333
rect 163191 -451 180913 -333
rect 181031 -451 181073 -333
rect 181191 -451 198913 -333
rect 199031 -451 199073 -333
rect 199191 -451 216913 -333
rect 217031 -451 217073 -333
rect 217191 -451 234913 -333
rect 235031 -451 235073 -333
rect 235191 -451 252913 -333
rect 253031 -451 253073 -333
rect 253191 -451 270913 -333
rect 271031 -451 271073 -333
rect 271191 -451 288913 -333
rect 289031 -451 289073 -333
rect 289191 -451 292671 -333
rect 292789 -451 292831 -333
rect 292949 -451 292965 -333
rect -1003 -467 292965 -451
rect -1483 -653 293445 -637
rect -1483 -771 -1467 -653
rect -1349 -771 -1307 -653
rect -1189 -771 9913 -653
rect 10031 -771 10073 -653
rect 10191 -771 27913 -653
rect 28031 -771 28073 -653
rect 28191 -771 45913 -653
rect 46031 -771 46073 -653
rect 46191 -771 63913 -653
rect 64031 -771 64073 -653
rect 64191 -771 81913 -653
rect 82031 -771 82073 -653
rect 82191 -771 99913 -653
rect 100031 -771 100073 -653
rect 100191 -771 117913 -653
rect 118031 -771 118073 -653
rect 118191 -771 135913 -653
rect 136031 -771 136073 -653
rect 136191 -771 153913 -653
rect 154031 -771 154073 -653
rect 154191 -771 171913 -653
rect 172031 -771 172073 -653
rect 172191 -771 189913 -653
rect 190031 -771 190073 -653
rect 190191 -771 207913 -653
rect 208031 -771 208073 -653
rect 208191 -771 225913 -653
rect 226031 -771 226073 -653
rect 226191 -771 243913 -653
rect 244031 -771 244073 -653
rect 244191 -771 261913 -653
rect 262031 -771 262073 -653
rect 262191 -771 279913 -653
rect 280031 -771 280073 -653
rect 280191 -771 293151 -653
rect 293269 -771 293311 -653
rect 293429 -771 293445 -653
rect -1483 -813 293445 -771
rect -1483 -931 -1467 -813
rect -1349 -931 -1307 -813
rect -1189 -931 9913 -813
rect 10031 -931 10073 -813
rect 10191 -931 27913 -813
rect 28031 -931 28073 -813
rect 28191 -931 45913 -813
rect 46031 -931 46073 -813
rect 46191 -931 63913 -813
rect 64031 -931 64073 -813
rect 64191 -931 81913 -813
rect 82031 -931 82073 -813
rect 82191 -931 99913 -813
rect 100031 -931 100073 -813
rect 100191 -931 117913 -813
rect 118031 -931 118073 -813
rect 118191 -931 135913 -813
rect 136031 -931 136073 -813
rect 136191 -931 153913 -813
rect 154031 -931 154073 -813
rect 154191 -931 171913 -813
rect 172031 -931 172073 -813
rect 172191 -931 189913 -813
rect 190031 -931 190073 -813
rect 190191 -931 207913 -813
rect 208031 -931 208073 -813
rect 208191 -931 225913 -813
rect 226031 -931 226073 -813
rect 226191 -931 243913 -813
rect 244031 -931 244073 -813
rect 244191 -931 261913 -813
rect 262031 -931 262073 -813
rect 262191 -931 279913 -813
rect 280031 -931 280073 -813
rect 280191 -931 293151 -813
rect 293269 -931 293311 -813
rect 293429 -931 293445 -813
rect -1483 -947 293445 -931
rect -1963 -1133 293925 -1117
rect -1963 -1251 -1947 -1133
rect -1829 -1251 -1787 -1133
rect -1669 -1251 2773 -1133
rect 2891 -1251 2933 -1133
rect 3051 -1251 20773 -1133
rect 20891 -1251 20933 -1133
rect 21051 -1251 38773 -1133
rect 38891 -1251 38933 -1133
rect 39051 -1251 56773 -1133
rect 56891 -1251 56933 -1133
rect 57051 -1251 74773 -1133
rect 74891 -1251 74933 -1133
rect 75051 -1251 92773 -1133
rect 92891 -1251 92933 -1133
rect 93051 -1251 110773 -1133
rect 110891 -1251 110933 -1133
rect 111051 -1251 128773 -1133
rect 128891 -1251 128933 -1133
rect 129051 -1251 146773 -1133
rect 146891 -1251 146933 -1133
rect 147051 -1251 164773 -1133
rect 164891 -1251 164933 -1133
rect 165051 -1251 182773 -1133
rect 182891 -1251 182933 -1133
rect 183051 -1251 200773 -1133
rect 200891 -1251 200933 -1133
rect 201051 -1251 218773 -1133
rect 218891 -1251 218933 -1133
rect 219051 -1251 236773 -1133
rect 236891 -1251 236933 -1133
rect 237051 -1251 254773 -1133
rect 254891 -1251 254933 -1133
rect 255051 -1251 272773 -1133
rect 272891 -1251 272933 -1133
rect 273051 -1251 290773 -1133
rect 290891 -1251 290933 -1133
rect 291051 -1251 293631 -1133
rect 293749 -1251 293791 -1133
rect 293909 -1251 293925 -1133
rect -1963 -1293 293925 -1251
rect -1963 -1411 -1947 -1293
rect -1829 -1411 -1787 -1293
rect -1669 -1411 2773 -1293
rect 2891 -1411 2933 -1293
rect 3051 -1411 20773 -1293
rect 20891 -1411 20933 -1293
rect 21051 -1411 38773 -1293
rect 38891 -1411 38933 -1293
rect 39051 -1411 56773 -1293
rect 56891 -1411 56933 -1293
rect 57051 -1411 74773 -1293
rect 74891 -1411 74933 -1293
rect 75051 -1411 92773 -1293
rect 92891 -1411 92933 -1293
rect 93051 -1411 110773 -1293
rect 110891 -1411 110933 -1293
rect 111051 -1411 128773 -1293
rect 128891 -1411 128933 -1293
rect 129051 -1411 146773 -1293
rect 146891 -1411 146933 -1293
rect 147051 -1411 164773 -1293
rect 164891 -1411 164933 -1293
rect 165051 -1411 182773 -1293
rect 182891 -1411 182933 -1293
rect 183051 -1411 200773 -1293
rect 200891 -1411 200933 -1293
rect 201051 -1411 218773 -1293
rect 218891 -1411 218933 -1293
rect 219051 -1411 236773 -1293
rect 236891 -1411 236933 -1293
rect 237051 -1411 254773 -1293
rect 254891 -1411 254933 -1293
rect 255051 -1411 272773 -1293
rect 272891 -1411 272933 -1293
rect 273051 -1411 290773 -1293
rect 290891 -1411 290933 -1293
rect 291051 -1411 293631 -1293
rect 293749 -1411 293791 -1293
rect 293909 -1411 293925 -1293
rect -1963 -1427 293925 -1411
rect -2443 -1613 294405 -1597
rect -2443 -1731 -2427 -1613
rect -2309 -1731 -2267 -1613
rect -2149 -1731 11773 -1613
rect 11891 -1731 11933 -1613
rect 12051 -1731 29773 -1613
rect 29891 -1731 29933 -1613
rect 30051 -1731 47773 -1613
rect 47891 -1731 47933 -1613
rect 48051 -1731 65773 -1613
rect 65891 -1731 65933 -1613
rect 66051 -1731 83773 -1613
rect 83891 -1731 83933 -1613
rect 84051 -1731 101773 -1613
rect 101891 -1731 101933 -1613
rect 102051 -1731 119773 -1613
rect 119891 -1731 119933 -1613
rect 120051 -1731 137773 -1613
rect 137891 -1731 137933 -1613
rect 138051 -1731 155773 -1613
rect 155891 -1731 155933 -1613
rect 156051 -1731 173773 -1613
rect 173891 -1731 173933 -1613
rect 174051 -1731 191773 -1613
rect 191891 -1731 191933 -1613
rect 192051 -1731 209773 -1613
rect 209891 -1731 209933 -1613
rect 210051 -1731 227773 -1613
rect 227891 -1731 227933 -1613
rect 228051 -1731 245773 -1613
rect 245891 -1731 245933 -1613
rect 246051 -1731 263773 -1613
rect 263891 -1731 263933 -1613
rect 264051 -1731 281773 -1613
rect 281891 -1731 281933 -1613
rect 282051 -1731 294111 -1613
rect 294229 -1731 294271 -1613
rect 294389 -1731 294405 -1613
rect -2443 -1773 294405 -1731
rect -2443 -1891 -2427 -1773
rect -2309 -1891 -2267 -1773
rect -2149 -1891 11773 -1773
rect 11891 -1891 11933 -1773
rect 12051 -1891 29773 -1773
rect 29891 -1891 29933 -1773
rect 30051 -1891 47773 -1773
rect 47891 -1891 47933 -1773
rect 48051 -1891 65773 -1773
rect 65891 -1891 65933 -1773
rect 66051 -1891 83773 -1773
rect 83891 -1891 83933 -1773
rect 84051 -1891 101773 -1773
rect 101891 -1891 101933 -1773
rect 102051 -1891 119773 -1773
rect 119891 -1891 119933 -1773
rect 120051 -1891 137773 -1773
rect 137891 -1891 137933 -1773
rect 138051 -1891 155773 -1773
rect 155891 -1891 155933 -1773
rect 156051 -1891 173773 -1773
rect 173891 -1891 173933 -1773
rect 174051 -1891 191773 -1773
rect 191891 -1891 191933 -1773
rect 192051 -1891 209773 -1773
rect 209891 -1891 209933 -1773
rect 210051 -1891 227773 -1773
rect 227891 -1891 227933 -1773
rect 228051 -1891 245773 -1773
rect 245891 -1891 245933 -1773
rect 246051 -1891 263773 -1773
rect 263891 -1891 263933 -1773
rect 264051 -1891 281773 -1773
rect 281891 -1891 281933 -1773
rect 282051 -1891 294111 -1773
rect 294229 -1891 294271 -1773
rect 294389 -1891 294405 -1773
rect -2443 -1907 294405 -1891
rect -2923 -2093 294885 -2077
rect -2923 -2211 -2907 -2093
rect -2789 -2211 -2747 -2093
rect -2629 -2211 4633 -2093
rect 4751 -2211 4793 -2093
rect 4911 -2211 22633 -2093
rect 22751 -2211 22793 -2093
rect 22911 -2211 40633 -2093
rect 40751 -2211 40793 -2093
rect 40911 -2211 58633 -2093
rect 58751 -2211 58793 -2093
rect 58911 -2211 76633 -2093
rect 76751 -2211 76793 -2093
rect 76911 -2211 94633 -2093
rect 94751 -2211 94793 -2093
rect 94911 -2211 112633 -2093
rect 112751 -2211 112793 -2093
rect 112911 -2211 130633 -2093
rect 130751 -2211 130793 -2093
rect 130911 -2211 148633 -2093
rect 148751 -2211 148793 -2093
rect 148911 -2211 166633 -2093
rect 166751 -2211 166793 -2093
rect 166911 -2211 184633 -2093
rect 184751 -2211 184793 -2093
rect 184911 -2211 202633 -2093
rect 202751 -2211 202793 -2093
rect 202911 -2211 220633 -2093
rect 220751 -2211 220793 -2093
rect 220911 -2211 238633 -2093
rect 238751 -2211 238793 -2093
rect 238911 -2211 256633 -2093
rect 256751 -2211 256793 -2093
rect 256911 -2211 274633 -2093
rect 274751 -2211 274793 -2093
rect 274911 -2211 294591 -2093
rect 294709 -2211 294751 -2093
rect 294869 -2211 294885 -2093
rect -2923 -2253 294885 -2211
rect -2923 -2371 -2907 -2253
rect -2789 -2371 -2747 -2253
rect -2629 -2371 4633 -2253
rect 4751 -2371 4793 -2253
rect 4911 -2371 22633 -2253
rect 22751 -2371 22793 -2253
rect 22911 -2371 40633 -2253
rect 40751 -2371 40793 -2253
rect 40911 -2371 58633 -2253
rect 58751 -2371 58793 -2253
rect 58911 -2371 76633 -2253
rect 76751 -2371 76793 -2253
rect 76911 -2371 94633 -2253
rect 94751 -2371 94793 -2253
rect 94911 -2371 112633 -2253
rect 112751 -2371 112793 -2253
rect 112911 -2371 130633 -2253
rect 130751 -2371 130793 -2253
rect 130911 -2371 148633 -2253
rect 148751 -2371 148793 -2253
rect 148911 -2371 166633 -2253
rect 166751 -2371 166793 -2253
rect 166911 -2371 184633 -2253
rect 184751 -2371 184793 -2253
rect 184911 -2371 202633 -2253
rect 202751 -2371 202793 -2253
rect 202911 -2371 220633 -2253
rect 220751 -2371 220793 -2253
rect 220911 -2371 238633 -2253
rect 238751 -2371 238793 -2253
rect 238911 -2371 256633 -2253
rect 256751 -2371 256793 -2253
rect 256911 -2371 274633 -2253
rect 274751 -2371 274793 -2253
rect 274911 -2371 294591 -2253
rect 294709 -2371 294751 -2253
rect 294869 -2371 294885 -2253
rect -2923 -2387 294885 -2371
rect -3403 -2573 295365 -2557
rect -3403 -2691 -3387 -2573
rect -3269 -2691 -3227 -2573
rect -3109 -2691 13633 -2573
rect 13751 -2691 13793 -2573
rect 13911 -2691 31633 -2573
rect 31751 -2691 31793 -2573
rect 31911 -2691 49633 -2573
rect 49751 -2691 49793 -2573
rect 49911 -2691 67633 -2573
rect 67751 -2691 67793 -2573
rect 67911 -2691 85633 -2573
rect 85751 -2691 85793 -2573
rect 85911 -2691 103633 -2573
rect 103751 -2691 103793 -2573
rect 103911 -2691 121633 -2573
rect 121751 -2691 121793 -2573
rect 121911 -2691 139633 -2573
rect 139751 -2691 139793 -2573
rect 139911 -2691 157633 -2573
rect 157751 -2691 157793 -2573
rect 157911 -2691 175633 -2573
rect 175751 -2691 175793 -2573
rect 175911 -2691 193633 -2573
rect 193751 -2691 193793 -2573
rect 193911 -2691 211633 -2573
rect 211751 -2691 211793 -2573
rect 211911 -2691 229633 -2573
rect 229751 -2691 229793 -2573
rect 229911 -2691 247633 -2573
rect 247751 -2691 247793 -2573
rect 247911 -2691 265633 -2573
rect 265751 -2691 265793 -2573
rect 265911 -2691 283633 -2573
rect 283751 -2691 283793 -2573
rect 283911 -2691 295071 -2573
rect 295189 -2691 295231 -2573
rect 295349 -2691 295365 -2573
rect -3403 -2733 295365 -2691
rect -3403 -2851 -3387 -2733
rect -3269 -2851 -3227 -2733
rect -3109 -2851 13633 -2733
rect 13751 -2851 13793 -2733
rect 13911 -2851 31633 -2733
rect 31751 -2851 31793 -2733
rect 31911 -2851 49633 -2733
rect 49751 -2851 49793 -2733
rect 49911 -2851 67633 -2733
rect 67751 -2851 67793 -2733
rect 67911 -2851 85633 -2733
rect 85751 -2851 85793 -2733
rect 85911 -2851 103633 -2733
rect 103751 -2851 103793 -2733
rect 103911 -2851 121633 -2733
rect 121751 -2851 121793 -2733
rect 121911 -2851 139633 -2733
rect 139751 -2851 139793 -2733
rect 139911 -2851 157633 -2733
rect 157751 -2851 157793 -2733
rect 157911 -2851 175633 -2733
rect 175751 -2851 175793 -2733
rect 175911 -2851 193633 -2733
rect 193751 -2851 193793 -2733
rect 193911 -2851 211633 -2733
rect 211751 -2851 211793 -2733
rect 211911 -2851 229633 -2733
rect 229751 -2851 229793 -2733
rect 229911 -2851 247633 -2733
rect 247751 -2851 247793 -2733
rect 247911 -2851 265633 -2733
rect 265751 -2851 265793 -2733
rect 265911 -2851 283633 -2733
rect 283751 -2851 283793 -2733
rect 283911 -2851 295071 -2733
rect 295189 -2851 295231 -2733
rect 295349 -2851 295365 -2733
rect -3403 -2867 295365 -2851
rect -3883 -3053 295845 -3037
rect -3883 -3171 -3867 -3053
rect -3749 -3171 -3707 -3053
rect -3589 -3171 6493 -3053
rect 6611 -3171 6653 -3053
rect 6771 -3171 24493 -3053
rect 24611 -3171 24653 -3053
rect 24771 -3171 42493 -3053
rect 42611 -3171 42653 -3053
rect 42771 -3171 60493 -3053
rect 60611 -3171 60653 -3053
rect 60771 -3171 78493 -3053
rect 78611 -3171 78653 -3053
rect 78771 -3171 96493 -3053
rect 96611 -3171 96653 -3053
rect 96771 -3171 114493 -3053
rect 114611 -3171 114653 -3053
rect 114771 -3171 132493 -3053
rect 132611 -3171 132653 -3053
rect 132771 -3171 150493 -3053
rect 150611 -3171 150653 -3053
rect 150771 -3171 168493 -3053
rect 168611 -3171 168653 -3053
rect 168771 -3171 186493 -3053
rect 186611 -3171 186653 -3053
rect 186771 -3171 204493 -3053
rect 204611 -3171 204653 -3053
rect 204771 -3171 222493 -3053
rect 222611 -3171 222653 -3053
rect 222771 -3171 240493 -3053
rect 240611 -3171 240653 -3053
rect 240771 -3171 258493 -3053
rect 258611 -3171 258653 -3053
rect 258771 -3171 276493 -3053
rect 276611 -3171 276653 -3053
rect 276771 -3171 295551 -3053
rect 295669 -3171 295711 -3053
rect 295829 -3171 295845 -3053
rect -3883 -3213 295845 -3171
rect -3883 -3331 -3867 -3213
rect -3749 -3331 -3707 -3213
rect -3589 -3331 6493 -3213
rect 6611 -3331 6653 -3213
rect 6771 -3331 24493 -3213
rect 24611 -3331 24653 -3213
rect 24771 -3331 42493 -3213
rect 42611 -3331 42653 -3213
rect 42771 -3331 60493 -3213
rect 60611 -3331 60653 -3213
rect 60771 -3331 78493 -3213
rect 78611 -3331 78653 -3213
rect 78771 -3331 96493 -3213
rect 96611 -3331 96653 -3213
rect 96771 -3331 114493 -3213
rect 114611 -3331 114653 -3213
rect 114771 -3331 132493 -3213
rect 132611 -3331 132653 -3213
rect 132771 -3331 150493 -3213
rect 150611 -3331 150653 -3213
rect 150771 -3331 168493 -3213
rect 168611 -3331 168653 -3213
rect 168771 -3331 186493 -3213
rect 186611 -3331 186653 -3213
rect 186771 -3331 204493 -3213
rect 204611 -3331 204653 -3213
rect 204771 -3331 222493 -3213
rect 222611 -3331 222653 -3213
rect 222771 -3331 240493 -3213
rect 240611 -3331 240653 -3213
rect 240771 -3331 258493 -3213
rect 258611 -3331 258653 -3213
rect 258771 -3331 276493 -3213
rect 276611 -3331 276653 -3213
rect 276771 -3331 295551 -3213
rect 295669 -3331 295711 -3213
rect 295829 -3331 295845 -3213
rect -3883 -3347 295845 -3331
rect -4363 -3533 296325 -3517
rect -4363 -3651 -4347 -3533
rect -4229 -3651 -4187 -3533
rect -4069 -3651 15493 -3533
rect 15611 -3651 15653 -3533
rect 15771 -3651 33493 -3533
rect 33611 -3651 33653 -3533
rect 33771 -3651 51493 -3533
rect 51611 -3651 51653 -3533
rect 51771 -3651 69493 -3533
rect 69611 -3651 69653 -3533
rect 69771 -3651 87493 -3533
rect 87611 -3651 87653 -3533
rect 87771 -3651 105493 -3533
rect 105611 -3651 105653 -3533
rect 105771 -3651 123493 -3533
rect 123611 -3651 123653 -3533
rect 123771 -3651 141493 -3533
rect 141611 -3651 141653 -3533
rect 141771 -3651 159493 -3533
rect 159611 -3651 159653 -3533
rect 159771 -3651 177493 -3533
rect 177611 -3651 177653 -3533
rect 177771 -3651 195493 -3533
rect 195611 -3651 195653 -3533
rect 195771 -3651 213493 -3533
rect 213611 -3651 213653 -3533
rect 213771 -3651 231493 -3533
rect 231611 -3651 231653 -3533
rect 231771 -3651 249493 -3533
rect 249611 -3651 249653 -3533
rect 249771 -3651 267493 -3533
rect 267611 -3651 267653 -3533
rect 267771 -3651 285493 -3533
rect 285611 -3651 285653 -3533
rect 285771 -3651 296031 -3533
rect 296149 -3651 296191 -3533
rect 296309 -3651 296325 -3533
rect -4363 -3693 296325 -3651
rect -4363 -3811 -4347 -3693
rect -4229 -3811 -4187 -3693
rect -4069 -3811 15493 -3693
rect 15611 -3811 15653 -3693
rect 15771 -3811 33493 -3693
rect 33611 -3811 33653 -3693
rect 33771 -3811 51493 -3693
rect 51611 -3811 51653 -3693
rect 51771 -3811 69493 -3693
rect 69611 -3811 69653 -3693
rect 69771 -3811 87493 -3693
rect 87611 -3811 87653 -3693
rect 87771 -3811 105493 -3693
rect 105611 -3811 105653 -3693
rect 105771 -3811 123493 -3693
rect 123611 -3811 123653 -3693
rect 123771 -3811 141493 -3693
rect 141611 -3811 141653 -3693
rect 141771 -3811 159493 -3693
rect 159611 -3811 159653 -3693
rect 159771 -3811 177493 -3693
rect 177611 -3811 177653 -3693
rect 177771 -3811 195493 -3693
rect 195611 -3811 195653 -3693
rect 195771 -3811 213493 -3693
rect 213611 -3811 213653 -3693
rect 213771 -3811 231493 -3693
rect 231611 -3811 231653 -3693
rect 231771 -3811 249493 -3693
rect 249611 -3811 249653 -3693
rect 249771 -3811 267493 -3693
rect 267611 -3811 267653 -3693
rect 267771 -3811 285493 -3693
rect 285611 -3811 285653 -3693
rect 285771 -3811 296031 -3693
rect 296149 -3811 296191 -3693
rect 296309 -3811 296325 -3693
rect -4363 -3827 296325 -3811
<< labels >>
rlabel metal3 s 291760 142638 292480 142758 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 223049 351760 223105 352480 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 190573 351760 190629 352480 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 158143 351760 158199 352480 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 125713 351760 125769 352480 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 93237 351760 93293 352480 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 60807 351760 60863 352480 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 28377 351760 28433 352480 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -480 348610 240 348730 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -480 322498 240 322618 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -480 296454 240 296574 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 291760 169226 292480 169346 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -480 270342 240 270462 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -480 244298 240 244418 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -480 218254 240 218374 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -480 192142 240 192262 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -480 166098 240 166218 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -480 139986 240 140106 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -480 113942 240 114062 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -480 87898 240 88018 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -480 61786 240 61906 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 291760 195814 292480 195934 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 291760 222334 292480 222454 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 291760 248922 292480 249042 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 291760 275510 292480 275630 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 291760 302030 292480 302150 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 291760 328618 292480 328738 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 287909 351760 287965 352480 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 255479 351760 255535 352480 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 291760 3238 292480 3358 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 291760 228998 292480 229118 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 291760 255586 292480 255706 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 291760 282106 292480 282226 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 291760 308694 292480 308814 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 291760 335282 292480 335402 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 279813 351760 279869 352480 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 247383 351760 247439 352480 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 214907 351760 214963 352480 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 182477 351760 182533 352480 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 150047 351760 150103 352480 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 291760 23094 292480 23214 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 117571 351760 117627 352480 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 85141 351760 85197 352480 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 52711 351760 52767 352480 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 20235 351760 20291 352480 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -480 342082 240 342202 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -480 315970 240 316090 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -480 289926 240 290046 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -480 263882 240 264002 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -480 237770 240 237890 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -480 211726 240 211846 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 291760 43018 292480 43138 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -480 185614 240 185734 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -480 159570 240 159690 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -480 133526 240 133646 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -480 107414 240 107534 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -480 81370 240 81490 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -480 55258 240 55378 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -480 35742 240 35862 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -480 16158 240 16278 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 291760 62942 292480 63062 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 291760 82866 292480 82986 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 291760 102790 292480 102910 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 291760 122714 292480 122834 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 291760 149302 292480 149422 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 291760 175890 292480 176010 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 291760 202410 292480 202530 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 291760 16498 292480 16618 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 291760 242258 292480 242378 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 291760 268846 292480 268966 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 291760 295434 292480 295554 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 291760 321954 292480 322074 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 291760 348542 292480 348662 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 263575 351760 263631 352480 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 231145 351760 231201 352480 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 198715 351760 198771 352480 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 166239 351760 166295 352480 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 133809 351760 133865 352480 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 291760 36422 292480 36542 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 101379 351760 101435 352480 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 68903 351760 68959 352480 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 36473 351760 36529 352480 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 4043 351760 4099 352480 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -480 329026 240 329146 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -480 302982 240 303102 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -480 276870 240 276990 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -480 250826 240 250946 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -480 224714 240 224834 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -480 198670 240 198790 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 291760 56346 292480 56466 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -480 172626 240 172746 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -480 146514 240 146634 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -480 120470 240 120590 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -480 94358 240 94478 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -480 68314 240 68434 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -480 42270 240 42390 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -480 22686 240 22806 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -480 3170 240 3290 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 291760 76270 292480 76390 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 291760 96194 292480 96314 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 291760 116118 292480 116238 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 291760 136042 292480 136162 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 291760 162562 292480 162682 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 291760 189150 292480 189270 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 291760 215738 292480 215858 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 291760 9834 292480 9954 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 291760 235662 292480 235782 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 291760 262182 292480 262302 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 291760 288770 292480 288890 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 291760 315358 292480 315478 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 291760 341878 292480 341998 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 271717 351760 271773 352480 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 239241 351760 239297 352480 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 206811 351760 206867 352480 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 174381 351760 174437 352480 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 141905 351760 141961 352480 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 291760 29758 292480 29878 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 109475 351760 109531 352480 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 77045 351760 77101 352480 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 44569 351760 44625 352480 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 12139 351760 12195 352480 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -480 335554 240 335674 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -480 309510 240 309630 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -480 283398 240 283518 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -480 257354 240 257474 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -480 231242 240 231362 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -480 205198 240 205318 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 291760 49682 292480 49802 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -480 179154 240 179274 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -480 153042 240 153162 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -480 126998 240 127118 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -480 100886 240 101006 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -480 74842 240 74962 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -480 48730 240 48850 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -480 29214 240 29334 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -480 9630 240 9750 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 291760 69606 292480 69726 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 291760 89530 292480 89650 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 291760 109454 292480 109574 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 291760 129378 292480 129498 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 291760 155966 292480 156086 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 291760 182486 292480 182606 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 291760 209074 292480 209194 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 62923 -480 62979 240 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 240253 -480 240309 240 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 242001 -480 242057 240 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 243795 -480 243851 240 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 245543 -480 245599 240 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 247337 -480 247393 240 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 249085 -480 249141 240 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 250879 -480 250935 240 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 252673 -480 252729 240 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 254421 -480 254477 240 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 256215 -480 256271 240 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 80633 -480 80689 240 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 257963 -480 258019 240 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 259757 -480 259813 240 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 261505 -480 261561 240 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 263299 -480 263355 240 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 265047 -480 265103 240 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 266841 -480 266897 240 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 268589 -480 268645 240 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 270383 -480 270439 240 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 272177 -480 272233 240 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 273925 -480 273981 240 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 82427 -480 82483 240 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 275719 -480 275775 240 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 277467 -480 277523 240 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 279261 -480 279317 240 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 281009 -480 281065 240 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 282803 -480 282859 240 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 284551 -480 284607 240 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 286345 -480 286401 240 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 288139 -480 288195 240 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 84175 -480 84231 240 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 85969 -480 86025 240 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 87717 -480 87773 240 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 89511 -480 89567 240 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 91259 -480 91315 240 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 93053 -480 93109 240 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 94847 -480 94903 240 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 96595 -480 96651 240 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 64671 -480 64727 240 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 98389 -480 98445 240 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 100137 -480 100193 240 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 101931 -480 101987 240 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 103679 -480 103735 240 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 105473 -480 105529 240 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 107221 -480 107277 240 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 109015 -480 109071 240 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 110763 -480 110819 240 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 112557 -480 112613 240 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 114351 -480 114407 240 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 66465 -480 66521 240 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 116099 -480 116155 240 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 117893 -480 117949 240 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 119641 -480 119697 240 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 121435 -480 121491 240 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 123183 -480 123239 240 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 124977 -480 125033 240 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 126725 -480 126781 240 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 128519 -480 128575 240 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 130313 -480 130369 240 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 132061 -480 132117 240 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 68213 -480 68269 240 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 133855 -480 133911 240 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 135603 -480 135659 240 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 137397 -480 137453 240 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 139145 -480 139201 240 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 140939 -480 140995 240 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 142687 -480 142743 240 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 144481 -480 144537 240 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 146275 -480 146331 240 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 148023 -480 148079 240 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 149817 -480 149873 240 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 70007 -480 70063 240 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 151565 -480 151621 240 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 153359 -480 153415 240 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 155107 -480 155163 240 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 156901 -480 156957 240 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 158649 -480 158705 240 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 160443 -480 160499 240 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 162191 -480 162247 240 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 163985 -480 164041 240 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 165779 -480 165835 240 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 167527 -480 167583 240 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 71755 -480 71811 240 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 169321 -480 169377 240 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 171069 -480 171125 240 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 172863 -480 172919 240 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 174611 -480 174667 240 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 176405 -480 176461 240 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 178153 -480 178209 240 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 179947 -480 180003 240 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 181741 -480 181797 240 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 183489 -480 183545 240 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 185283 -480 185339 240 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 73549 -480 73605 240 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 187031 -480 187087 240 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 188825 -480 188881 240 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 190573 -480 190629 240 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 192367 -480 192423 240 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 194115 -480 194171 240 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 195909 -480 195965 240 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 197657 -480 197713 240 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 199451 -480 199507 240 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 201245 -480 201301 240 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 202993 -480 203049 240 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 75297 -480 75353 240 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 204787 -480 204843 240 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 206535 -480 206591 240 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 208329 -480 208385 240 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 210077 -480 210133 240 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 211871 -480 211927 240 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 213619 -480 213675 240 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 215413 -480 215469 240 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 217207 -480 217263 240 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 218955 -480 219011 240 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 220749 -480 220805 240 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 77091 -480 77147 240 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 222497 -480 222553 240 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 224291 -480 224347 240 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 226039 -480 226095 240 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 227833 -480 227889 240 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 229581 -480 229637 240 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 231375 -480 231431 240 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 233123 -480 233179 240 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 234917 -480 234973 240 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 236711 -480 236767 240 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 238459 -480 238515 240 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 78885 -480 78941 240 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 63475 -480 63531 240 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 240851 -480 240907 240 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 242599 -480 242655 240 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 244393 -480 244449 240 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 246141 -480 246197 240 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 247935 -480 247991 240 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 249683 -480 249739 240 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 251477 -480 251533 240 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 253225 -480 253281 240 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 255019 -480 255075 240 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 256767 -480 256823 240 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 81231 -480 81287 240 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 258561 -480 258617 240 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 260355 -480 260411 240 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 262103 -480 262159 240 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 263897 -480 263953 240 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 265645 -480 265701 240 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 267439 -480 267495 240 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 269187 -480 269243 240 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 270981 -480 271037 240 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 272729 -480 272785 240 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 274523 -480 274579 240 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 83025 -480 83081 240 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 276317 -480 276373 240 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 278065 -480 278121 240 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 279859 -480 279915 240 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 281607 -480 281663 240 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 283401 -480 283457 240 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 285149 -480 285205 240 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 286943 -480 286999 240 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 84773 -480 84829 240 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 86567 -480 86623 240 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 88315 -480 88371 240 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 90109 -480 90165 240 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 91857 -480 91913 240 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 93651 -480 93707 240 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 95399 -480 95455 240 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 97193 -480 97249 240 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 65269 -480 65325 240 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 98941 -480 98997 240 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 100735 -480 100791 240 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 102529 -480 102585 240 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 104277 -480 104333 240 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 106071 -480 106127 240 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 107819 -480 107875 240 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 109613 -480 109669 240 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 111361 -480 111417 240 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 113155 -480 113211 240 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 114903 -480 114959 240 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 67063 -480 67119 240 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 116697 -480 116753 240 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 118491 -480 118547 240 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 120239 -480 120295 240 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 122033 -480 122089 240 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 123781 -480 123837 240 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 125575 -480 125631 240 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 127323 -480 127379 240 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 129117 -480 129173 240 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 130865 -480 130921 240 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 132659 -480 132715 240 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 68811 -480 68867 240 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 134407 -480 134463 240 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 136201 -480 136257 240 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 137995 -480 138051 240 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 139743 -480 139799 240 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 141537 -480 141593 240 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 143285 -480 143341 240 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 145079 -480 145135 240 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 146827 -480 146883 240 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 148621 -480 148677 240 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 150369 -480 150425 240 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 70605 -480 70661 240 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 152163 -480 152219 240 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 153957 -480 154013 240 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 155705 -480 155761 240 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 157499 -480 157555 240 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 159247 -480 159303 240 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 161041 -480 161097 240 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 162789 -480 162845 240 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 164583 -480 164639 240 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 166331 -480 166387 240 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 168125 -480 168181 240 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 72353 -480 72409 240 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 169919 -480 169975 240 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 171667 -480 171723 240 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 173461 -480 173517 240 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 175209 -480 175265 240 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 177003 -480 177059 240 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 178751 -480 178807 240 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 180545 -480 180601 240 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 182293 -480 182349 240 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 184087 -480 184143 240 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 185835 -480 185891 240 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 74147 -480 74203 240 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 187629 -480 187685 240 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 189423 -480 189479 240 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 191171 -480 191227 240 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 192965 -480 193021 240 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 194713 -480 194769 240 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 196507 -480 196563 240 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 198255 -480 198311 240 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 200049 -480 200105 240 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 201797 -480 201853 240 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 203591 -480 203647 240 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 75895 -480 75951 240 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 205385 -480 205441 240 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 207133 -480 207189 240 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 208927 -480 208983 240 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 210675 -480 210731 240 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 212469 -480 212525 240 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 214217 -480 214273 240 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 216011 -480 216067 240 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 217759 -480 217815 240 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 219553 -480 219609 240 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 221301 -480 221357 240 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 77689 -480 77745 240 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 223095 -480 223151 240 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 224889 -480 224945 240 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 226637 -480 226693 240 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 228431 -480 228487 240 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 230179 -480 230235 240 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 231973 -480 232029 240 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 233721 -480 233777 240 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 235515 -480 235571 240 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 237263 -480 237319 240 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 239057 -480 239113 240 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 79437 -480 79493 240 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 64073 -480 64129 240 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 241403 -480 241459 240 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 243197 -480 243253 240 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 244945 -480 245001 240 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 246739 -480 246795 240 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 248533 -480 248589 240 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 250281 -480 250337 240 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 252075 -480 252131 240 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 253823 -480 253879 240 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 255617 -480 255673 240 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 257365 -480 257421 240 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 81829 -480 81885 240 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 259159 -480 259215 240 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 260907 -480 260963 240 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 262701 -480 262757 240 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 264495 -480 264551 240 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 266243 -480 266299 240 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 268037 -480 268093 240 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 269785 -480 269841 240 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 271579 -480 271635 240 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 273327 -480 273383 240 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 275121 -480 275177 240 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 83577 -480 83633 240 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 276869 -480 276925 240 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 278663 -480 278719 240 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 280411 -480 280467 240 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 282205 -480 282261 240 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 283999 -480 284055 240 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 285747 -480 285803 240 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 287541 -480 287597 240 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 289289 -480 289345 240 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 85371 -480 85427 240 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 87119 -480 87175 240 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 88913 -480 88969 240 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 90707 -480 90763 240 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 92455 -480 92511 240 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 94249 -480 94305 240 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 95997 -480 96053 240 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 97791 -480 97847 240 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 65867 -480 65923 240 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 99539 -480 99595 240 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 101333 -480 101389 240 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 103081 -480 103137 240 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 104875 -480 104931 240 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 106669 -480 106725 240 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 108417 -480 108473 240 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 110211 -480 110267 240 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 111959 -480 112015 240 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 113753 -480 113809 240 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 115501 -480 115557 240 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 67615 -480 67671 240 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 117295 -480 117351 240 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 119043 -480 119099 240 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 120837 -480 120893 240 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 122585 -480 122641 240 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 124379 -480 124435 240 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 126173 -480 126229 240 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 127921 -480 127977 240 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 129715 -480 129771 240 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 131463 -480 131519 240 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 133257 -480 133313 240 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 69409 -480 69465 240 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 135005 -480 135061 240 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 136799 -480 136855 240 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 138547 -480 138603 240 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 140341 -480 140397 240 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 142135 -480 142191 240 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 143883 -480 143939 240 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 145677 -480 145733 240 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 147425 -480 147481 240 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 149219 -480 149275 240 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 150967 -480 151023 240 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 71203 -480 71259 240 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 152761 -480 152817 240 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 154509 -480 154565 240 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 156303 -480 156359 240 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 158097 -480 158153 240 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 159845 -480 159901 240 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 161639 -480 161695 240 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 163387 -480 163443 240 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 165181 -480 165237 240 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 166929 -480 166985 240 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 168723 -480 168779 240 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 72951 -480 73007 240 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 170471 -480 170527 240 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 172265 -480 172321 240 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 174013 -480 174069 240 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 175807 -480 175863 240 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 177601 -480 177657 240 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 179349 -480 179405 240 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 181143 -480 181199 240 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 182891 -480 182947 240 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 184685 -480 184741 240 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 186433 -480 186489 240 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 74745 -480 74801 240 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 188227 -480 188283 240 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 189975 -480 190031 240 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 191769 -480 191825 240 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 193563 -480 193619 240 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 195311 -480 195367 240 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 197105 -480 197161 240 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 198853 -480 198909 240 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 200647 -480 200703 240 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 202395 -480 202451 240 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 204189 -480 204245 240 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 76493 -480 76549 240 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 205937 -480 205993 240 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 207731 -480 207787 240 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 209479 -480 209535 240 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 211273 -480 211329 240 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 213067 -480 213123 240 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 214815 -480 214871 240 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 216609 -480 216665 240 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 218357 -480 218413 240 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 220151 -480 220207 240 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 221899 -480 221955 240 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 78287 -480 78343 240 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 223693 -480 223749 240 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 225441 -480 225497 240 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 227235 -480 227291 240 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 229029 -480 229085 240 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 230777 -480 230833 240 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 232571 -480 232627 240 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 234319 -480 234375 240 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 236113 -480 236169 240 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 237861 -480 237917 240 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 239655 -480 239711 240 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 80035 -480 80091 240 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 289887 -480 289943 240 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 290485 -480 290541 240 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 291083 -480 291139 240 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 291681 -480 291737 240 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -1003 -467 292965 -157 8 vccd1
port 531 nsew power input
rlabel metal5 s -1483 1433 293445 1743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 19433 293445 19743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 37433 293445 37743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 55433 293445 55743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 73433 293445 73743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 91433 293445 91743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 109433 293445 109743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 127433 293445 127743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 145433 293445 145743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 163433 293445 163743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 181433 293445 181743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 199433 293445 199743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 217433 293445 217743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 235433 293445 235743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 253433 293445 253743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 271433 293445 271743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 289433 293445 289743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 307433 293445 307743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 325433 293445 325743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1483 343433 293445 343743 6 vccd1
port 531 nsew power input
rlabel metal5 s -1003 352125 292965 352435 6 vccd1
port 531 nsew power input
rlabel metal4 s -1003 -467 -693 352435 4 vccd1
port 531 nsew power input
rlabel metal4 s 292655 -467 292965 352435 6 vccd1
port 531 nsew power input
rlabel metal4 s 897 -947 1207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 18897 -947 19207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 36897 -947 37207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 54897 -947 55207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 72897 -947 73207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 90897 -947 91207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 108897 -947 109207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 126897 -947 127207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 144897 -947 145207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 162897 -947 163207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 180897 -947 181207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 198897 -947 199207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 216897 -947 217207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 234897 -947 235207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 252897 -947 253207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 270897 -947 271207 352915 6 vccd1
port 531 nsew power input
rlabel metal4 s 288897 -947 289207 352915 6 vccd1
port 531 nsew power input
rlabel metal5 s -1963 -1427 293925 -1117 8 vccd2
port 532 nsew power input
rlabel metal5 s -2443 3293 294405 3603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 21293 294405 21603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 39293 294405 39603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 57293 294405 57603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 75293 294405 75603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 93293 294405 93603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 111293 294405 111603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 129293 294405 129603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 147293 294405 147603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 165293 294405 165603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 183293 294405 183603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 201293 294405 201603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 219293 294405 219603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 237293 294405 237603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 255293 294405 255603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 273293 294405 273603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 291293 294405 291603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 309293 294405 309603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 327293 294405 327603 6 vccd2
port 532 nsew power input
rlabel metal5 s -2443 345293 294405 345603 6 vccd2
port 532 nsew power input
rlabel metal5 s -1963 353085 293925 353395 6 vccd2
port 532 nsew power input
rlabel metal4 s -1963 -1427 -1653 353395 4 vccd2
port 532 nsew power input
rlabel metal4 s 293615 -1427 293925 353395 6 vccd2
port 532 nsew power input
rlabel metal4 s 2757 -1907 3067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 20757 -1907 21067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 38757 -1907 39067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 56757 -1907 57067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 74757 -1907 75067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 92757 -1907 93067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 110757 -1907 111067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 128757 -1907 129067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 146757 -1907 147067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 164757 -1907 165067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 182757 -1907 183067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 200757 -1907 201067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 218757 -1907 219067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 236757 -1907 237067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 254757 -1907 255067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 272757 -1907 273067 353875 6 vccd2
port 532 nsew power input
rlabel metal4 s 290757 -1907 291067 353875 6 vccd2
port 532 nsew power input
rlabel metal5 s -2923 -2387 294885 -2077 8 vdda1
port 533 nsew power input
rlabel metal5 s -3403 5153 295365 5463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 23153 295365 23463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 41153 295365 41463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 59153 295365 59463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 77153 295365 77463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 95153 295365 95463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 113153 295365 113463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 131153 295365 131463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 149153 295365 149463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 167153 295365 167463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 185153 295365 185463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 203153 295365 203463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 221153 295365 221463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 239153 295365 239463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 257153 295365 257463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 275153 295365 275463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 293153 295365 293463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 311153 295365 311463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 329153 295365 329463 6 vdda1
port 533 nsew power input
rlabel metal5 s -3403 347153 295365 347463 6 vdda1
port 533 nsew power input
rlabel metal5 s -2923 354045 294885 354355 6 vdda1
port 533 nsew power input
rlabel metal4 s -2923 -2387 -2613 354355 4 vdda1
port 533 nsew power input
rlabel metal4 s 294575 -2387 294885 354355 6 vdda1
port 533 nsew power input
rlabel metal4 s 4617 -2867 4927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 22617 -2867 22927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 40617 -2867 40927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 58617 -2867 58927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 76617 -2867 76927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 94617 -2867 94927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 112617 -2867 112927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 130617 -2867 130927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 148617 -2867 148927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 166617 -2867 166927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 184617 -2867 184927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 202617 -2867 202927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 220617 -2867 220927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 238617 -2867 238927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 256617 -2867 256927 354835 6 vdda1
port 533 nsew power input
rlabel metal4 s 274617 -2867 274927 354835 6 vdda1
port 533 nsew power input
rlabel metal5 s -3883 -3347 295845 -3037 8 vdda2
port 534 nsew power input
rlabel metal5 s -4363 7013 296325 7323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 25013 296325 25323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 43013 296325 43323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 61013 296325 61323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 79013 296325 79323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 97013 296325 97323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 115013 296325 115323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 133013 296325 133323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 151013 296325 151323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 169013 296325 169323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 187013 296325 187323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 205013 296325 205323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 223013 296325 223323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 241013 296325 241323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 259013 296325 259323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 277013 296325 277323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 295013 296325 295323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 313013 296325 313323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 331013 296325 331323 6 vdda2
port 534 nsew power input
rlabel metal5 s -4363 349013 296325 349323 6 vdda2
port 534 nsew power input
rlabel metal5 s -3883 355005 295845 355315 6 vdda2
port 534 nsew power input
rlabel metal4 s -3883 -3347 -3573 355315 4 vdda2
port 534 nsew power input
rlabel metal4 s 295535 -3347 295845 355315 6 vdda2
port 534 nsew power input
rlabel metal4 s 6477 -3827 6787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 24477 -3827 24787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 42477 -3827 42787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 60477 -3827 60787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 78477 -3827 78787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 96477 -3827 96787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 114477 -3827 114787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 132477 -3827 132787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 150477 -3827 150787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 168477 -3827 168787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 186477 -3827 186787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 204477 -3827 204787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 222477 -3827 222787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 240477 -3827 240787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 258477 -3827 258787 355795 6 vdda2
port 534 nsew power input
rlabel metal4 s 276477 -3827 276787 355795 6 vdda2
port 534 nsew power input
rlabel metal5 s -3403 -2867 295365 -2557 8 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 14153 295365 14463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 32153 295365 32463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 50153 295365 50463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 68153 295365 68463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 86153 295365 86463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 104153 295365 104463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 122153 295365 122463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 140153 295365 140463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 158153 295365 158463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 176153 295365 176463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 194153 295365 194463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 212153 295365 212463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 230153 295365 230463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 248153 295365 248463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 266153 295365 266463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 284153 295365 284463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 302153 295365 302463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 320153 295365 320463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 338153 295365 338463 6 vssa1
port 535 nsew ground input
rlabel metal5 s -3403 354525 295365 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s -3403 -2867 -3093 354835 4 vssa1
port 535 nsew ground input
rlabel metal4 s 13617 -2867 13927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 31617 -2867 31927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 49617 -2867 49927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 67617 -2867 67927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 85617 -2867 85927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 103617 -2867 103927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 121617 -2867 121927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 139617 -2867 139927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 157617 -2867 157927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 175617 -2867 175927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 193617 -2867 193927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 211617 -2867 211927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 229617 -2867 229927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 247617 -2867 247927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 265617 -2867 265927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 283617 -2867 283927 354835 6 vssa1
port 535 nsew ground input
rlabel metal4 s 295055 -2867 295365 354835 6 vssa1
port 535 nsew ground input
rlabel metal5 s -4363 -3827 296325 -3517 8 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 16013 296325 16323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 34013 296325 34323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 52013 296325 52323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 70013 296325 70323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 88013 296325 88323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 106013 296325 106323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 124013 296325 124323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 142013 296325 142323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 160013 296325 160323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 178013 296325 178323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 196013 296325 196323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 214013 296325 214323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 232013 296325 232323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 250013 296325 250323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 268013 296325 268323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 286013 296325 286323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 304013 296325 304323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 322013 296325 322323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 340013 296325 340323 6 vssa2
port 536 nsew ground input
rlabel metal5 s -4363 355485 296325 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s -4363 -3827 -4053 355795 4 vssa2
port 536 nsew ground input
rlabel metal4 s 15477 -3827 15787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 33477 -3827 33787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 51477 -3827 51787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 69477 -3827 69787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 87477 -3827 87787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 105477 -3827 105787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 123477 -3827 123787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 141477 -3827 141787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 159477 -3827 159787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 177477 -3827 177787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 195477 -3827 195787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 213477 -3827 213787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 231477 -3827 231787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 249477 -3827 249787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 267477 -3827 267787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 285477 -3827 285787 355795 6 vssa2
port 536 nsew ground input
rlabel metal4 s 296015 -3827 296325 355795 6 vssa2
port 536 nsew ground input
rlabel metal5 s -1483 -947 293445 -637 8 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 10433 293445 10743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 28433 293445 28743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 46433 293445 46743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 64433 293445 64743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 82433 293445 82743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 100433 293445 100743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 118433 293445 118743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 136433 293445 136743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 154433 293445 154743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 172433 293445 172743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 190433 293445 190743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 208433 293445 208743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 226433 293445 226743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 244433 293445 244743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 262433 293445 262743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 280433 293445 280743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 298433 293445 298743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 316433 293445 316743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 334433 293445 334743 6 vssd1
port 537 nsew ground input
rlabel metal5 s -1483 352605 293445 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s -1483 -947 -1173 352915 4 vssd1
port 537 nsew ground input
rlabel metal4 s 9897 -947 10207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 27897 -947 28207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 45897 -947 46207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 63897 -947 64207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 81897 -947 82207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 99897 -947 100207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 117897 -947 118207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 135897 -947 136207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 153897 -947 154207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 171897 -947 172207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 189897 -947 190207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 207897 -947 208207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 225897 -947 226207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 243897 -947 244207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 261897 -947 262207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 279897 -947 280207 352915 6 vssd1
port 537 nsew ground input
rlabel metal4 s 293135 -947 293445 352915 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2443 -1907 294405 -1597 8 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 12293 294405 12603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 30293 294405 30603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 48293 294405 48603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 66293 294405 66603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 84293 294405 84603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 102293 294405 102603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 120293 294405 120603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 138293 294405 138603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 156293 294405 156603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 174293 294405 174603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 192293 294405 192603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 210293 294405 210603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 228293 294405 228603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 246293 294405 246603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 264293 294405 264603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 282293 294405 282603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 300293 294405 300603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 318293 294405 318603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 336293 294405 336603 6 vssd2
port 538 nsew ground input
rlabel metal5 s -2443 353565 294405 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s -2443 -1907 -2133 353875 4 vssd2
port 538 nsew ground input
rlabel metal4 s 11757 -1907 12067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 29757 -1907 30067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 47757 -1907 48067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 65757 -1907 66067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 83757 -1907 84067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 101757 -1907 102067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 119757 -1907 120067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 137757 -1907 138067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 155757 -1907 156067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 173757 -1907 174067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 191757 -1907 192067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 209757 -1907 210067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 227757 -1907 228067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 245757 -1907 246067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 263757 -1907 264067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 281757 -1907 282067 353875 6 vssd2
port 538 nsew ground input
rlabel metal4 s 294095 -1907 294405 353875 6 vssd2
port 538 nsew ground input
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 23915 -480 23971 240 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 25663 -480 25719 240 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 27457 -480 27513 240 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 29205 -480 29261 240 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 30999 -480 31055 240 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 32747 -480 32803 240 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 34541 -480 34597 240 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 36289 -480 36345 240 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 38083 -480 38139 240 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 39831 -480 39887 240 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 6159 -480 6215 240 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 41625 -480 41681 240 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 43419 -480 43475 240 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 45167 -480 45223 240 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 46961 -480 47017 240 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 48709 -480 48765 240 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 50503 -480 50559 240 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 52251 -480 52307 240 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 54045 -480 54101 240 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 55793 -480 55849 240 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 57587 -480 57643 240 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 8505 -480 8561 240 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 59381 -480 59437 240 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 61129 -480 61185 240 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 10897 -480 10953 240 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 13243 -480 13299 240 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 15037 -480 15093 240 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 16785 -480 16841 240 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 18579 -480 18635 240 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 20327 -480 20383 240 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 22121 -480 22177 240 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 4365 -480 4421 240 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 24467 -480 24523 240 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 26261 -480 26317 240 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 28009 -480 28065 240 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 29803 -480 29859 240 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 31597 -480 31653 240 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 33345 -480 33401 240 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 35139 -480 35195 240 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 36887 -480 36943 240 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 38681 -480 38737 240 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 40429 -480 40485 240 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 6757 -480 6813 240 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 42223 -480 42279 240 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 43971 -480 44027 240 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 45765 -480 45821 240 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 47559 -480 47615 240 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 49307 -480 49363 240 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 51101 -480 51157 240 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 52849 -480 52905 240 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 54643 -480 54699 240 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 56391 -480 56447 240 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 58185 -480 58241 240 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 9103 -480 9159 240 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 59933 -480 59989 240 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 61727 -480 61783 240 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 11495 -480 11551 240 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 13841 -480 13897 240 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 15635 -480 15691 240 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 17383 -480 17439 240 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 19177 -480 19233 240 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 20925 -480 20981 240 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 22719 -480 22775 240 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 4963 -480 5019 240 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 25065 -480 25121 240 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 26859 -480 26915 240 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 28607 -480 28663 240 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 30401 -480 30457 240 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 32149 -480 32205 240 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 33943 -480 33999 240 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 35737 -480 35793 240 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 37485 -480 37541 240 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 39279 -480 39335 240 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 41027 -480 41083 240 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 7355 -480 7411 240 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 42821 -480 42877 240 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 44569 -480 44625 240 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 46363 -480 46419 240 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 48111 -480 48167 240 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 49905 -480 49961 240 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 51653 -480 51709 240 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 53447 -480 53503 240 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 55241 -480 55297 240 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 56989 -480 57045 240 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 58783 -480 58839 240 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 9701 -480 9757 240 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 60531 -480 60587 240 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 62325 -480 62381 240 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 12093 -480 12149 240 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 14439 -480 14495 240 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 16187 -480 16243 240 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 17981 -480 18037 240 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 19775 -480 19831 240 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 21523 -480 21579 240 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 23317 -480 23373 240 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 5561 -480 5617 240 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 7953 -480 8009 240 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 10299 -480 10355 240 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 12645 -480 12701 240 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
