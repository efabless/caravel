magic
tech sky130A
magscale 36 1
timestamp 1598787136
<< metal5 >>
rect 0 75 15 90
rect 30 75 45 105
rect 0 60 45 75
rect 30 0 45 60
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
