magic
tech sky130A
magscale 1 2
timestamp 1636146659
<< viali >>
rect 4721 833 4755 867
rect 949 765 983 799
rect 1501 765 1535 799
rect 1777 765 1811 799
rect 2053 765 2087 799
rect 2513 765 2547 799
rect 2973 765 3007 799
rect 3433 765 3467 799
rect 3893 765 3927 799
rect 4353 765 4387 799
rect 5273 765 5307 799
rect 1225 629 1259 663
rect 4813 629 4847 663
<< metal1 >>
rect 0 2202 5980 2224
rect 0 2150 78 2202
rect 130 2150 142 2202
rect 194 2150 206 2202
rect 258 2150 270 2202
rect 322 2150 1478 2202
rect 1530 2150 1542 2202
rect 1594 2150 1606 2202
rect 1658 2150 1670 2202
rect 1722 2150 2878 2202
rect 2930 2150 2942 2202
rect 2994 2150 3006 2202
rect 3058 2150 3070 2202
rect 3122 2150 4278 2202
rect 4330 2150 4342 2202
rect 4394 2150 4406 2202
rect 4458 2150 4470 2202
rect 4522 2150 5980 2202
rect 0 2128 5980 2150
rect 0 1658 5980 1680
rect 0 1606 778 1658
rect 830 1606 842 1658
rect 894 1606 906 1658
rect 958 1606 970 1658
rect 1022 1606 2178 1658
rect 2230 1606 2242 1658
rect 2294 1606 2306 1658
rect 2358 1606 2370 1658
rect 2422 1606 3578 1658
rect 3630 1606 3642 1658
rect 3694 1606 3706 1658
rect 3758 1606 3770 1658
rect 3822 1606 4978 1658
rect 5030 1606 5042 1658
rect 5094 1606 5106 1658
rect 5158 1606 5170 1658
rect 5222 1606 5980 1658
rect 0 1584 5980 1606
rect 0 1114 5980 1136
rect 0 1062 78 1114
rect 130 1062 142 1114
rect 194 1062 206 1114
rect 258 1062 270 1114
rect 322 1062 1478 1114
rect 1530 1062 1542 1114
rect 1594 1062 1606 1114
rect 1658 1062 1670 1114
rect 1722 1062 2878 1114
rect 2930 1062 2942 1114
rect 2994 1062 3006 1114
rect 3058 1062 3070 1114
rect 3122 1062 4278 1114
rect 4330 1062 4342 1114
rect 4394 1062 4406 1114
rect 4458 1062 4470 1114
rect 4522 1062 5980 1114
rect 0 1040 5980 1062
rect 4709 867 4767 873
rect 4709 833 4721 867
rect 4755 864 4767 867
rect 5718 864 5724 876
rect 4755 836 5724 864
rect 4755 833 4767 836
rect 4709 827 4767 833
rect 5718 824 5724 836
rect 5776 824 5782 876
rect 198 756 204 808
rect 256 796 262 808
rect 937 799 995 805
rect 937 796 949 799
rect 256 768 949 796
rect 256 756 262 768
rect 937 765 949 768
rect 983 765 995 799
rect 937 759 995 765
rect 1118 756 1124 808
rect 1176 796 1182 808
rect 1489 799 1547 805
rect 1489 796 1501 799
rect 1176 768 1501 796
rect 1176 756 1182 768
rect 1489 765 1501 768
rect 1535 765 1547 799
rect 1489 759 1547 765
rect 1578 756 1584 808
rect 1636 796 1642 808
rect 1765 799 1823 805
rect 1765 796 1777 799
rect 1636 768 1777 796
rect 1636 756 1642 768
rect 1765 765 1777 768
rect 1811 765 1823 799
rect 2038 796 2044 808
rect 1999 768 2044 796
rect 1765 759 1823 765
rect 2038 756 2044 768
rect 2096 756 2102 808
rect 2498 796 2504 808
rect 2459 768 2504 796
rect 2498 756 2504 768
rect 2556 756 2562 808
rect 2958 796 2964 808
rect 2919 768 2964 796
rect 2958 756 2964 768
rect 3016 756 3022 808
rect 3418 796 3424 808
rect 3379 768 3424 796
rect 3418 756 3424 768
rect 3476 756 3482 808
rect 3878 796 3884 808
rect 3839 768 3884 796
rect 3878 756 3884 768
rect 3936 756 3942 808
rect 4338 796 4344 808
rect 4299 768 4344 796
rect 4338 756 4344 768
rect 4396 756 4402 808
rect 5258 796 5264 808
rect 5219 768 5264 796
rect 5258 756 5264 768
rect 5316 756 5322 808
rect 658 620 664 672
rect 716 660 722 672
rect 1213 663 1271 669
rect 1213 660 1225 663
rect 716 632 1225 660
rect 716 620 722 632
rect 1213 629 1225 632
rect 1259 629 1271 663
rect 4798 660 4804 672
rect 4759 632 4804 660
rect 1213 623 1271 629
rect 4798 620 4804 632
rect 4856 620 4862 672
rect 0 570 5980 592
rect 0 518 778 570
rect 830 518 842 570
rect 894 518 906 570
rect 958 518 970 570
rect 1022 518 2178 570
rect 2230 518 2242 570
rect 2294 518 2306 570
rect 2358 518 2370 570
rect 2422 518 3578 570
rect 3630 518 3642 570
rect 3694 518 3706 570
rect 3758 518 3770 570
rect 3822 518 4978 570
rect 5030 518 5042 570
rect 5094 518 5106 570
rect 5158 518 5170 570
rect 5222 518 5980 570
rect 0 496 5980 518
<< via1 >>
rect 78 2150 130 2202
rect 142 2150 194 2202
rect 206 2150 258 2202
rect 270 2150 322 2202
rect 1478 2150 1530 2202
rect 1542 2150 1594 2202
rect 1606 2150 1658 2202
rect 1670 2150 1722 2202
rect 2878 2150 2930 2202
rect 2942 2150 2994 2202
rect 3006 2150 3058 2202
rect 3070 2150 3122 2202
rect 4278 2150 4330 2202
rect 4342 2150 4394 2202
rect 4406 2150 4458 2202
rect 4470 2150 4522 2202
rect 778 1606 830 1658
rect 842 1606 894 1658
rect 906 1606 958 1658
rect 970 1606 1022 1658
rect 2178 1606 2230 1658
rect 2242 1606 2294 1658
rect 2306 1606 2358 1658
rect 2370 1606 2422 1658
rect 3578 1606 3630 1658
rect 3642 1606 3694 1658
rect 3706 1606 3758 1658
rect 3770 1606 3822 1658
rect 4978 1606 5030 1658
rect 5042 1606 5094 1658
rect 5106 1606 5158 1658
rect 5170 1606 5222 1658
rect 78 1062 130 1114
rect 142 1062 194 1114
rect 206 1062 258 1114
rect 270 1062 322 1114
rect 1478 1062 1530 1114
rect 1542 1062 1594 1114
rect 1606 1062 1658 1114
rect 1670 1062 1722 1114
rect 2878 1062 2930 1114
rect 2942 1062 2994 1114
rect 3006 1062 3058 1114
rect 3070 1062 3122 1114
rect 4278 1062 4330 1114
rect 4342 1062 4394 1114
rect 4406 1062 4458 1114
rect 4470 1062 4522 1114
rect 5724 824 5776 876
rect 204 756 256 808
rect 1124 756 1176 808
rect 1584 756 1636 808
rect 2044 799 2096 808
rect 2044 765 2053 799
rect 2053 765 2087 799
rect 2087 765 2096 799
rect 2044 756 2096 765
rect 2504 799 2556 808
rect 2504 765 2513 799
rect 2513 765 2547 799
rect 2547 765 2556 799
rect 2504 756 2556 765
rect 2964 799 3016 808
rect 2964 765 2973 799
rect 2973 765 3007 799
rect 3007 765 3016 799
rect 2964 756 3016 765
rect 3424 799 3476 808
rect 3424 765 3433 799
rect 3433 765 3467 799
rect 3467 765 3476 799
rect 3424 756 3476 765
rect 3884 799 3936 808
rect 3884 765 3893 799
rect 3893 765 3927 799
rect 3927 765 3936 799
rect 3884 756 3936 765
rect 4344 799 4396 808
rect 4344 765 4353 799
rect 4353 765 4387 799
rect 4387 765 4396 799
rect 4344 756 4396 765
rect 5264 799 5316 808
rect 5264 765 5273 799
rect 5273 765 5307 799
rect 5307 765 5316 799
rect 5264 756 5316 765
rect 664 620 716 672
rect 4804 663 4856 672
rect 4804 629 4813 663
rect 4813 629 4847 663
rect 4847 629 4856 663
rect 4804 620 4856 629
rect 778 518 830 570
rect 842 518 894 570
rect 906 518 958 570
rect 970 518 1022 570
rect 2178 518 2230 570
rect 2242 518 2294 570
rect 2306 518 2358 570
rect 2370 518 2422 570
rect 3578 518 3630 570
rect 3642 518 3694 570
rect 3706 518 3758 570
rect 3770 518 3822 570
rect 4978 518 5030 570
rect 5042 518 5094 570
rect 5106 518 5158 570
rect 5170 518 5222 570
<< metal2 >>
rect 78 2204 322 2224
rect 78 2202 92 2204
rect 148 2202 172 2204
rect 228 2202 252 2204
rect 308 2202 322 2204
rect 78 2148 92 2150
rect 148 2148 172 2150
rect 228 2148 252 2150
rect 308 2148 322 2150
rect 78 2128 322 2148
rect 1478 2204 1722 2224
rect 1478 2202 1492 2204
rect 1548 2202 1572 2204
rect 1628 2202 1652 2204
rect 1708 2202 1722 2204
rect 1478 2148 1492 2150
rect 1548 2148 1572 2150
rect 1628 2148 1652 2150
rect 1708 2148 1722 2150
rect 1478 2128 1722 2148
rect 2878 2204 3122 2224
rect 2878 2202 2892 2204
rect 2948 2202 2972 2204
rect 3028 2202 3052 2204
rect 3108 2202 3122 2204
rect 2878 2148 2892 2150
rect 2948 2148 2972 2150
rect 3028 2148 3052 2150
rect 3108 2148 3122 2150
rect 2878 2128 3122 2148
rect 4278 2204 4522 2224
rect 4278 2202 4292 2204
rect 4348 2202 4372 2204
rect 4428 2202 4452 2204
rect 4508 2202 4522 2204
rect 4278 2148 4292 2150
rect 4348 2148 4372 2150
rect 4428 2148 4452 2150
rect 4508 2148 4522 2150
rect 4278 2128 4522 2148
rect 778 1660 1022 1680
rect 778 1658 792 1660
rect 848 1658 872 1660
rect 928 1658 952 1660
rect 1008 1658 1022 1660
rect 778 1604 792 1606
rect 848 1604 872 1606
rect 928 1604 952 1606
rect 1008 1604 1022 1606
rect 778 1584 1022 1604
rect 2178 1660 2422 1680
rect 2178 1658 2192 1660
rect 2248 1658 2272 1660
rect 2328 1658 2352 1660
rect 2408 1658 2422 1660
rect 2178 1604 2192 1606
rect 2248 1604 2272 1606
rect 2328 1604 2352 1606
rect 2408 1604 2422 1606
rect 2178 1584 2422 1604
rect 3578 1660 3822 1680
rect 3578 1658 3592 1660
rect 3648 1658 3672 1660
rect 3728 1658 3752 1660
rect 3808 1658 3822 1660
rect 3578 1604 3592 1606
rect 3648 1604 3672 1606
rect 3728 1604 3752 1606
rect 3808 1604 3822 1606
rect 3578 1584 3822 1604
rect 4978 1660 5222 1680
rect 4978 1658 4992 1660
rect 5048 1658 5072 1660
rect 5128 1658 5152 1660
rect 5208 1658 5222 1660
rect 4978 1604 4992 1606
rect 5048 1604 5072 1606
rect 5128 1604 5152 1606
rect 5208 1604 5222 1606
rect 4978 1584 5222 1604
rect 78 1116 322 1136
rect 78 1114 92 1116
rect 148 1114 172 1116
rect 228 1114 252 1116
rect 308 1114 322 1116
rect 78 1060 92 1062
rect 148 1060 172 1062
rect 228 1060 252 1062
rect 308 1060 322 1062
rect 78 1040 322 1060
rect 1478 1116 1722 1136
rect 1478 1114 1492 1116
rect 1548 1114 1572 1116
rect 1628 1114 1652 1116
rect 1708 1114 1722 1116
rect 1478 1060 1492 1062
rect 1548 1060 1572 1062
rect 1628 1060 1652 1062
rect 1708 1060 1722 1062
rect 1478 1040 1722 1060
rect 2878 1116 3122 1136
rect 2878 1114 2892 1116
rect 2948 1114 2972 1116
rect 3028 1114 3052 1116
rect 3108 1114 3122 1116
rect 2878 1060 2892 1062
rect 2948 1060 2972 1062
rect 3028 1060 3052 1062
rect 3108 1060 3122 1062
rect 2878 1040 3122 1060
rect 4278 1116 4522 1136
rect 4278 1114 4292 1116
rect 4348 1114 4372 1116
rect 4428 1114 4452 1116
rect 4508 1114 4522 1116
rect 4278 1060 4292 1062
rect 4348 1060 4372 1062
rect 4428 1060 4452 1062
rect 4508 1060 4522 1062
rect 4278 1040 4522 1060
rect 5724 876 5776 882
rect 5724 818 5776 824
rect 204 808 256 814
rect 204 750 256 756
rect 1124 808 1176 814
rect 1124 750 1176 756
rect 1584 808 1636 814
rect 1584 750 1636 756
rect 2044 808 2096 814
rect 2044 750 2096 756
rect 2504 808 2556 814
rect 2504 750 2556 756
rect 2964 808 3016 814
rect 2964 750 3016 756
rect 3424 808 3476 814
rect 3424 750 3476 756
rect 3884 808 3936 814
rect 3884 750 3936 756
rect 4344 808 4396 814
rect 4344 750 4396 756
rect 5264 808 5316 814
rect 5264 750 5316 756
rect 216 400 244 750
rect 664 672 716 678
rect 664 614 716 620
rect 676 400 704 614
rect 778 572 1022 592
rect 778 570 792 572
rect 848 570 872 572
rect 928 570 952 572
rect 1008 570 1022 572
rect 778 516 792 518
rect 848 516 872 518
rect 928 516 952 518
rect 1008 516 1022 518
rect 778 496 1022 516
rect 1136 400 1164 750
rect 1596 400 1624 750
rect 2056 400 2084 750
rect 2178 572 2422 592
rect 2178 570 2192 572
rect 2248 570 2272 572
rect 2328 570 2352 572
rect 2408 570 2422 572
rect 2178 516 2192 518
rect 2248 516 2272 518
rect 2328 516 2352 518
rect 2408 516 2422 518
rect 2178 496 2422 516
rect 2516 400 2544 750
rect 2976 400 3004 750
rect 3436 400 3464 750
rect 3578 572 3822 592
rect 3578 570 3592 572
rect 3648 570 3672 572
rect 3728 570 3752 572
rect 3808 570 3822 572
rect 3578 516 3592 518
rect 3648 516 3672 518
rect 3728 516 3752 518
rect 3808 516 3822 518
rect 3578 496 3822 516
rect 3896 400 3924 750
rect 4356 400 4384 750
rect 4804 672 4856 678
rect 4804 614 4856 620
rect 4816 400 4844 614
rect 4978 572 5222 592
rect 4978 570 4992 572
rect 5048 570 5072 572
rect 5128 570 5152 572
rect 5208 570 5222 572
rect 4978 516 4992 518
rect 5048 516 5072 518
rect 5128 516 5152 518
rect 5208 516 5222 518
rect 4978 496 5222 516
rect 5276 400 5304 750
rect 5736 400 5764 818
rect 202 0 258 400
rect 662 0 718 400
rect 1122 0 1178 400
rect 1582 0 1638 400
rect 2042 0 2098 400
rect 2502 0 2558 400
rect 2962 0 3018 400
rect 3422 0 3478 400
rect 3882 0 3938 400
rect 4342 0 4398 400
rect 4802 0 4858 400
rect 5262 0 5318 400
rect 5722 0 5778 400
<< via2 >>
rect 92 2202 148 2204
rect 172 2202 228 2204
rect 252 2202 308 2204
rect 92 2150 130 2202
rect 130 2150 142 2202
rect 142 2150 148 2202
rect 172 2150 194 2202
rect 194 2150 206 2202
rect 206 2150 228 2202
rect 252 2150 258 2202
rect 258 2150 270 2202
rect 270 2150 308 2202
rect 92 2148 148 2150
rect 172 2148 228 2150
rect 252 2148 308 2150
rect 1492 2202 1548 2204
rect 1572 2202 1628 2204
rect 1652 2202 1708 2204
rect 1492 2150 1530 2202
rect 1530 2150 1542 2202
rect 1542 2150 1548 2202
rect 1572 2150 1594 2202
rect 1594 2150 1606 2202
rect 1606 2150 1628 2202
rect 1652 2150 1658 2202
rect 1658 2150 1670 2202
rect 1670 2150 1708 2202
rect 1492 2148 1548 2150
rect 1572 2148 1628 2150
rect 1652 2148 1708 2150
rect 2892 2202 2948 2204
rect 2972 2202 3028 2204
rect 3052 2202 3108 2204
rect 2892 2150 2930 2202
rect 2930 2150 2942 2202
rect 2942 2150 2948 2202
rect 2972 2150 2994 2202
rect 2994 2150 3006 2202
rect 3006 2150 3028 2202
rect 3052 2150 3058 2202
rect 3058 2150 3070 2202
rect 3070 2150 3108 2202
rect 2892 2148 2948 2150
rect 2972 2148 3028 2150
rect 3052 2148 3108 2150
rect 4292 2202 4348 2204
rect 4372 2202 4428 2204
rect 4452 2202 4508 2204
rect 4292 2150 4330 2202
rect 4330 2150 4342 2202
rect 4342 2150 4348 2202
rect 4372 2150 4394 2202
rect 4394 2150 4406 2202
rect 4406 2150 4428 2202
rect 4452 2150 4458 2202
rect 4458 2150 4470 2202
rect 4470 2150 4508 2202
rect 4292 2148 4348 2150
rect 4372 2148 4428 2150
rect 4452 2148 4508 2150
rect 792 1658 848 1660
rect 872 1658 928 1660
rect 952 1658 1008 1660
rect 792 1606 830 1658
rect 830 1606 842 1658
rect 842 1606 848 1658
rect 872 1606 894 1658
rect 894 1606 906 1658
rect 906 1606 928 1658
rect 952 1606 958 1658
rect 958 1606 970 1658
rect 970 1606 1008 1658
rect 792 1604 848 1606
rect 872 1604 928 1606
rect 952 1604 1008 1606
rect 2192 1658 2248 1660
rect 2272 1658 2328 1660
rect 2352 1658 2408 1660
rect 2192 1606 2230 1658
rect 2230 1606 2242 1658
rect 2242 1606 2248 1658
rect 2272 1606 2294 1658
rect 2294 1606 2306 1658
rect 2306 1606 2328 1658
rect 2352 1606 2358 1658
rect 2358 1606 2370 1658
rect 2370 1606 2408 1658
rect 2192 1604 2248 1606
rect 2272 1604 2328 1606
rect 2352 1604 2408 1606
rect 3592 1658 3648 1660
rect 3672 1658 3728 1660
rect 3752 1658 3808 1660
rect 3592 1606 3630 1658
rect 3630 1606 3642 1658
rect 3642 1606 3648 1658
rect 3672 1606 3694 1658
rect 3694 1606 3706 1658
rect 3706 1606 3728 1658
rect 3752 1606 3758 1658
rect 3758 1606 3770 1658
rect 3770 1606 3808 1658
rect 3592 1604 3648 1606
rect 3672 1604 3728 1606
rect 3752 1604 3808 1606
rect 4992 1658 5048 1660
rect 5072 1658 5128 1660
rect 5152 1658 5208 1660
rect 4992 1606 5030 1658
rect 5030 1606 5042 1658
rect 5042 1606 5048 1658
rect 5072 1606 5094 1658
rect 5094 1606 5106 1658
rect 5106 1606 5128 1658
rect 5152 1606 5158 1658
rect 5158 1606 5170 1658
rect 5170 1606 5208 1658
rect 4992 1604 5048 1606
rect 5072 1604 5128 1606
rect 5152 1604 5208 1606
rect 92 1114 148 1116
rect 172 1114 228 1116
rect 252 1114 308 1116
rect 92 1062 130 1114
rect 130 1062 142 1114
rect 142 1062 148 1114
rect 172 1062 194 1114
rect 194 1062 206 1114
rect 206 1062 228 1114
rect 252 1062 258 1114
rect 258 1062 270 1114
rect 270 1062 308 1114
rect 92 1060 148 1062
rect 172 1060 228 1062
rect 252 1060 308 1062
rect 1492 1114 1548 1116
rect 1572 1114 1628 1116
rect 1652 1114 1708 1116
rect 1492 1062 1530 1114
rect 1530 1062 1542 1114
rect 1542 1062 1548 1114
rect 1572 1062 1594 1114
rect 1594 1062 1606 1114
rect 1606 1062 1628 1114
rect 1652 1062 1658 1114
rect 1658 1062 1670 1114
rect 1670 1062 1708 1114
rect 1492 1060 1548 1062
rect 1572 1060 1628 1062
rect 1652 1060 1708 1062
rect 2892 1114 2948 1116
rect 2972 1114 3028 1116
rect 3052 1114 3108 1116
rect 2892 1062 2930 1114
rect 2930 1062 2942 1114
rect 2942 1062 2948 1114
rect 2972 1062 2994 1114
rect 2994 1062 3006 1114
rect 3006 1062 3028 1114
rect 3052 1062 3058 1114
rect 3058 1062 3070 1114
rect 3070 1062 3108 1114
rect 2892 1060 2948 1062
rect 2972 1060 3028 1062
rect 3052 1060 3108 1062
rect 4292 1114 4348 1116
rect 4372 1114 4428 1116
rect 4452 1114 4508 1116
rect 4292 1062 4330 1114
rect 4330 1062 4342 1114
rect 4342 1062 4348 1114
rect 4372 1062 4394 1114
rect 4394 1062 4406 1114
rect 4406 1062 4428 1114
rect 4452 1062 4458 1114
rect 4458 1062 4470 1114
rect 4470 1062 4508 1114
rect 4292 1060 4348 1062
rect 4372 1060 4428 1062
rect 4452 1060 4508 1062
rect 792 570 848 572
rect 872 570 928 572
rect 952 570 1008 572
rect 792 518 830 570
rect 830 518 842 570
rect 842 518 848 570
rect 872 518 894 570
rect 894 518 906 570
rect 906 518 928 570
rect 952 518 958 570
rect 958 518 970 570
rect 970 518 1008 570
rect 792 516 848 518
rect 872 516 928 518
rect 952 516 1008 518
rect 2192 570 2248 572
rect 2272 570 2328 572
rect 2352 570 2408 572
rect 2192 518 2230 570
rect 2230 518 2242 570
rect 2242 518 2248 570
rect 2272 518 2294 570
rect 2294 518 2306 570
rect 2306 518 2328 570
rect 2352 518 2358 570
rect 2358 518 2370 570
rect 2370 518 2408 570
rect 2192 516 2248 518
rect 2272 516 2328 518
rect 2352 516 2408 518
rect 3592 570 3648 572
rect 3672 570 3728 572
rect 3752 570 3808 572
rect 3592 518 3630 570
rect 3630 518 3642 570
rect 3642 518 3648 570
rect 3672 518 3694 570
rect 3694 518 3706 570
rect 3706 518 3728 570
rect 3752 518 3758 570
rect 3758 518 3770 570
rect 3770 518 3808 570
rect 3592 516 3648 518
rect 3672 516 3728 518
rect 3752 516 3808 518
rect 4992 570 5048 572
rect 5072 570 5128 572
rect 5152 570 5208 572
rect 4992 518 5030 570
rect 5030 518 5042 570
rect 5042 518 5048 570
rect 5072 518 5094 570
rect 5094 518 5106 570
rect 5106 518 5128 570
rect 5152 518 5158 570
rect 5158 518 5170 570
rect 5170 518 5208 570
rect 4992 516 5048 518
rect 5072 516 5128 518
rect 5152 516 5208 518
<< metal3 >>
rect 60 2208 340 2209
rect 60 2144 88 2208
rect 152 2144 168 2208
rect 232 2144 248 2208
rect 312 2144 340 2208
rect 60 2143 340 2144
rect 1460 2208 1740 2209
rect 1460 2144 1488 2208
rect 1552 2144 1568 2208
rect 1632 2144 1648 2208
rect 1712 2144 1740 2208
rect 1460 2143 1740 2144
rect 2860 2208 3140 2209
rect 2860 2144 2888 2208
rect 2952 2144 2968 2208
rect 3032 2144 3048 2208
rect 3112 2144 3140 2208
rect 2860 2143 3140 2144
rect 4260 2208 4540 2209
rect 4260 2144 4288 2208
rect 4352 2144 4368 2208
rect 4432 2144 4448 2208
rect 4512 2144 4540 2208
rect 4260 2143 4540 2144
rect 760 1664 1040 1665
rect 760 1600 788 1664
rect 852 1600 868 1664
rect 932 1600 948 1664
rect 1012 1600 1040 1664
rect 760 1599 1040 1600
rect 2160 1664 2440 1665
rect 2160 1600 2188 1664
rect 2252 1600 2268 1664
rect 2332 1600 2348 1664
rect 2412 1600 2440 1664
rect 2160 1599 2440 1600
rect 3560 1664 3840 1665
rect 3560 1600 3588 1664
rect 3652 1600 3668 1664
rect 3732 1600 3748 1664
rect 3812 1600 3840 1664
rect 3560 1599 3840 1600
rect 4960 1664 5240 1665
rect 4960 1600 4988 1664
rect 5052 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5240 1664
rect 4960 1599 5240 1600
rect 60 1120 340 1121
rect 60 1056 88 1120
rect 152 1056 168 1120
rect 232 1056 248 1120
rect 312 1056 340 1120
rect 60 1055 340 1056
rect 1460 1120 1740 1121
rect 1460 1056 1488 1120
rect 1552 1056 1568 1120
rect 1632 1056 1648 1120
rect 1712 1056 1740 1120
rect 1460 1055 1740 1056
rect 2860 1120 3140 1121
rect 2860 1056 2888 1120
rect 2952 1056 2968 1120
rect 3032 1056 3048 1120
rect 3112 1056 3140 1120
rect 2860 1055 3140 1056
rect 4260 1120 4540 1121
rect 4260 1056 4288 1120
rect 4352 1056 4368 1120
rect 4432 1056 4448 1120
rect 4512 1056 4540 1120
rect 4260 1055 4540 1056
rect 760 576 1040 577
rect 760 512 788 576
rect 852 512 868 576
rect 932 512 948 576
rect 1012 512 1040 576
rect 760 511 1040 512
rect 2160 576 2440 577
rect 2160 512 2188 576
rect 2252 512 2268 576
rect 2332 512 2348 576
rect 2412 512 2440 576
rect 2160 511 2440 512
rect 3560 576 3840 577
rect 3560 512 3588 576
rect 3652 512 3668 576
rect 3732 512 3748 576
rect 3812 512 3840 576
rect 3560 511 3840 512
rect 4960 576 5240 577
rect 4960 512 4988 576
rect 5052 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5240 576
rect 4960 511 5240 512
<< via3 >>
rect 88 2204 152 2208
rect 88 2148 92 2204
rect 92 2148 148 2204
rect 148 2148 152 2204
rect 88 2144 152 2148
rect 168 2204 232 2208
rect 168 2148 172 2204
rect 172 2148 228 2204
rect 228 2148 232 2204
rect 168 2144 232 2148
rect 248 2204 312 2208
rect 248 2148 252 2204
rect 252 2148 308 2204
rect 308 2148 312 2204
rect 248 2144 312 2148
rect 1488 2204 1552 2208
rect 1488 2148 1492 2204
rect 1492 2148 1548 2204
rect 1548 2148 1552 2204
rect 1488 2144 1552 2148
rect 1568 2204 1632 2208
rect 1568 2148 1572 2204
rect 1572 2148 1628 2204
rect 1628 2148 1632 2204
rect 1568 2144 1632 2148
rect 1648 2204 1712 2208
rect 1648 2148 1652 2204
rect 1652 2148 1708 2204
rect 1708 2148 1712 2204
rect 1648 2144 1712 2148
rect 2888 2204 2952 2208
rect 2888 2148 2892 2204
rect 2892 2148 2948 2204
rect 2948 2148 2952 2204
rect 2888 2144 2952 2148
rect 2968 2204 3032 2208
rect 2968 2148 2972 2204
rect 2972 2148 3028 2204
rect 3028 2148 3032 2204
rect 2968 2144 3032 2148
rect 3048 2204 3112 2208
rect 3048 2148 3052 2204
rect 3052 2148 3108 2204
rect 3108 2148 3112 2204
rect 3048 2144 3112 2148
rect 4288 2204 4352 2208
rect 4288 2148 4292 2204
rect 4292 2148 4348 2204
rect 4348 2148 4352 2204
rect 4288 2144 4352 2148
rect 4368 2204 4432 2208
rect 4368 2148 4372 2204
rect 4372 2148 4428 2204
rect 4428 2148 4432 2204
rect 4368 2144 4432 2148
rect 4448 2204 4512 2208
rect 4448 2148 4452 2204
rect 4452 2148 4508 2204
rect 4508 2148 4512 2204
rect 4448 2144 4512 2148
rect 788 1660 852 1664
rect 788 1604 792 1660
rect 792 1604 848 1660
rect 848 1604 852 1660
rect 788 1600 852 1604
rect 868 1660 932 1664
rect 868 1604 872 1660
rect 872 1604 928 1660
rect 928 1604 932 1660
rect 868 1600 932 1604
rect 948 1660 1012 1664
rect 948 1604 952 1660
rect 952 1604 1008 1660
rect 1008 1604 1012 1660
rect 948 1600 1012 1604
rect 2188 1660 2252 1664
rect 2188 1604 2192 1660
rect 2192 1604 2248 1660
rect 2248 1604 2252 1660
rect 2188 1600 2252 1604
rect 2268 1660 2332 1664
rect 2268 1604 2272 1660
rect 2272 1604 2328 1660
rect 2328 1604 2332 1660
rect 2268 1600 2332 1604
rect 2348 1660 2412 1664
rect 2348 1604 2352 1660
rect 2352 1604 2408 1660
rect 2408 1604 2412 1660
rect 2348 1600 2412 1604
rect 3588 1660 3652 1664
rect 3588 1604 3592 1660
rect 3592 1604 3648 1660
rect 3648 1604 3652 1660
rect 3588 1600 3652 1604
rect 3668 1660 3732 1664
rect 3668 1604 3672 1660
rect 3672 1604 3728 1660
rect 3728 1604 3732 1660
rect 3668 1600 3732 1604
rect 3748 1660 3812 1664
rect 3748 1604 3752 1660
rect 3752 1604 3808 1660
rect 3808 1604 3812 1660
rect 3748 1600 3812 1604
rect 4988 1660 5052 1664
rect 4988 1604 4992 1660
rect 4992 1604 5048 1660
rect 5048 1604 5052 1660
rect 4988 1600 5052 1604
rect 5068 1660 5132 1664
rect 5068 1604 5072 1660
rect 5072 1604 5128 1660
rect 5128 1604 5132 1660
rect 5068 1600 5132 1604
rect 5148 1660 5212 1664
rect 5148 1604 5152 1660
rect 5152 1604 5208 1660
rect 5208 1604 5212 1660
rect 5148 1600 5212 1604
rect 88 1116 152 1120
rect 88 1060 92 1116
rect 92 1060 148 1116
rect 148 1060 152 1116
rect 88 1056 152 1060
rect 168 1116 232 1120
rect 168 1060 172 1116
rect 172 1060 228 1116
rect 228 1060 232 1116
rect 168 1056 232 1060
rect 248 1116 312 1120
rect 248 1060 252 1116
rect 252 1060 308 1116
rect 308 1060 312 1116
rect 248 1056 312 1060
rect 1488 1116 1552 1120
rect 1488 1060 1492 1116
rect 1492 1060 1548 1116
rect 1548 1060 1552 1116
rect 1488 1056 1552 1060
rect 1568 1116 1632 1120
rect 1568 1060 1572 1116
rect 1572 1060 1628 1116
rect 1628 1060 1632 1116
rect 1568 1056 1632 1060
rect 1648 1116 1712 1120
rect 1648 1060 1652 1116
rect 1652 1060 1708 1116
rect 1708 1060 1712 1116
rect 1648 1056 1712 1060
rect 2888 1116 2952 1120
rect 2888 1060 2892 1116
rect 2892 1060 2948 1116
rect 2948 1060 2952 1116
rect 2888 1056 2952 1060
rect 2968 1116 3032 1120
rect 2968 1060 2972 1116
rect 2972 1060 3028 1116
rect 3028 1060 3032 1116
rect 2968 1056 3032 1060
rect 3048 1116 3112 1120
rect 3048 1060 3052 1116
rect 3052 1060 3108 1116
rect 3108 1060 3112 1116
rect 3048 1056 3112 1060
rect 4288 1116 4352 1120
rect 4288 1060 4292 1116
rect 4292 1060 4348 1116
rect 4348 1060 4352 1116
rect 4288 1056 4352 1060
rect 4368 1116 4432 1120
rect 4368 1060 4372 1116
rect 4372 1060 4428 1116
rect 4428 1060 4432 1116
rect 4368 1056 4432 1060
rect 4448 1116 4512 1120
rect 4448 1060 4452 1116
rect 4452 1060 4508 1116
rect 4508 1060 4512 1116
rect 4448 1056 4512 1060
rect 788 572 852 576
rect 788 516 792 572
rect 792 516 848 572
rect 848 516 852 572
rect 788 512 852 516
rect 868 572 932 576
rect 868 516 872 572
rect 872 516 928 572
rect 928 516 932 572
rect 868 512 932 516
rect 948 572 1012 576
rect 948 516 952 572
rect 952 516 1008 572
rect 1008 516 1012 572
rect 948 512 1012 516
rect 2188 572 2252 576
rect 2188 516 2192 572
rect 2192 516 2248 572
rect 2248 516 2252 572
rect 2188 512 2252 516
rect 2268 572 2332 576
rect 2268 516 2272 572
rect 2272 516 2328 572
rect 2328 516 2332 572
rect 2268 512 2332 516
rect 2348 572 2412 576
rect 2348 516 2352 572
rect 2352 516 2408 572
rect 2408 516 2412 572
rect 2348 512 2412 516
rect 3588 572 3652 576
rect 3588 516 3592 572
rect 3592 516 3648 572
rect 3648 516 3652 572
rect 3588 512 3652 516
rect 3668 572 3732 576
rect 3668 516 3672 572
rect 3672 516 3728 572
rect 3728 516 3732 572
rect 3668 512 3732 516
rect 3748 572 3812 576
rect 3748 516 3752 572
rect 3752 516 3808 572
rect 3808 516 3812 572
rect 3748 512 3812 516
rect 4988 572 5052 576
rect 4988 516 4992 572
rect 4992 516 5048 572
rect 5048 516 5052 572
rect 4988 512 5052 516
rect 5068 572 5132 576
rect 5068 516 5072 572
rect 5072 516 5128 572
rect 5128 516 5132 572
rect 5068 512 5132 516
rect 5148 572 5212 576
rect 5148 516 5152 572
rect 5152 516 5208 572
rect 5208 516 5212 572
rect 5148 512 5212 516
<< metal4 >>
rect 60 2208 340 2224
rect 60 2144 88 2208
rect 152 2144 168 2208
rect 232 2144 248 2208
rect 312 2144 340 2208
rect 60 1120 340 2144
rect 60 1056 88 1120
rect 152 1056 168 1120
rect 232 1056 248 1120
rect 312 1056 340 1120
rect 60 1014 340 1056
rect 60 778 82 1014
rect 318 778 340 1014
rect 60 496 340 778
rect 760 1714 1040 2224
rect 760 1478 782 1714
rect 1018 1478 1040 1714
rect 760 576 1040 1478
rect 760 512 788 576
rect 852 512 868 576
rect 932 512 948 576
rect 1012 512 1040 576
rect 760 496 1040 512
rect 1460 2208 1740 2224
rect 1460 2144 1488 2208
rect 1552 2144 1568 2208
rect 1632 2144 1648 2208
rect 1712 2144 1740 2208
rect 1460 1120 1740 2144
rect 1460 1056 1488 1120
rect 1552 1056 1568 1120
rect 1632 1056 1648 1120
rect 1712 1056 1740 1120
rect 1460 1014 1740 1056
rect 1460 778 1482 1014
rect 1718 778 1740 1014
rect 1460 496 1740 778
rect 2160 1714 2440 2224
rect 2160 1478 2182 1714
rect 2418 1478 2440 1714
rect 2160 576 2440 1478
rect 2160 512 2188 576
rect 2252 512 2268 576
rect 2332 512 2348 576
rect 2412 512 2440 576
rect 2160 496 2440 512
rect 2860 2208 3140 2224
rect 2860 2144 2888 2208
rect 2952 2144 2968 2208
rect 3032 2144 3048 2208
rect 3112 2144 3140 2208
rect 2860 1120 3140 2144
rect 2860 1056 2888 1120
rect 2952 1056 2968 1120
rect 3032 1056 3048 1120
rect 3112 1056 3140 1120
rect 2860 1014 3140 1056
rect 2860 778 2882 1014
rect 3118 778 3140 1014
rect 2860 496 3140 778
rect 3560 1714 3840 2224
rect 3560 1478 3582 1714
rect 3818 1478 3840 1714
rect 3560 576 3840 1478
rect 3560 512 3588 576
rect 3652 512 3668 576
rect 3732 512 3748 576
rect 3812 512 3840 576
rect 3560 496 3840 512
rect 4260 2208 4540 2224
rect 4260 2144 4288 2208
rect 4352 2144 4368 2208
rect 4432 2144 4448 2208
rect 4512 2144 4540 2208
rect 4260 1120 4540 2144
rect 4260 1056 4288 1120
rect 4352 1056 4368 1120
rect 4432 1056 4448 1120
rect 4512 1056 4540 1120
rect 4260 1014 4540 1056
rect 4260 778 4282 1014
rect 4518 778 4540 1014
rect 4260 496 4540 778
rect 4960 1714 5240 2224
rect 4960 1478 4982 1714
rect 5218 1478 5240 1714
rect 4960 576 5240 1478
rect 4960 512 4988 576
rect 5052 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5240 576
rect 4960 496 5240 512
<< via4 >>
rect 82 778 318 1014
rect 782 1664 1018 1714
rect 782 1600 788 1664
rect 788 1600 852 1664
rect 852 1600 868 1664
rect 868 1600 932 1664
rect 932 1600 948 1664
rect 948 1600 1012 1664
rect 1012 1600 1018 1664
rect 782 1478 1018 1600
rect 1482 778 1718 1014
rect 2182 1664 2418 1714
rect 2182 1600 2188 1664
rect 2188 1600 2252 1664
rect 2252 1600 2268 1664
rect 2268 1600 2332 1664
rect 2332 1600 2348 1664
rect 2348 1600 2412 1664
rect 2412 1600 2418 1664
rect 2182 1478 2418 1600
rect 2882 778 3118 1014
rect 3582 1664 3818 1714
rect 3582 1600 3588 1664
rect 3588 1600 3652 1664
rect 3652 1600 3668 1664
rect 3668 1600 3732 1664
rect 3732 1600 3748 1664
rect 3748 1600 3812 1664
rect 3812 1600 3818 1664
rect 3582 1478 3818 1600
rect 4282 778 4518 1014
rect 4982 1664 5218 1714
rect 4982 1600 4988 1664
rect 4988 1600 5052 1664
rect 5052 1600 5068 1664
rect 5068 1600 5132 1664
rect 5132 1600 5148 1664
rect 5148 1600 5212 1664
rect 5212 1600 5218 1664
rect 4982 1478 5218 1600
<< metal5 >>
rect 0 1714 5980 1756
rect 0 1478 782 1714
rect 1018 1478 2182 1714
rect 2418 1478 3582 1714
rect 3818 1478 4982 1714
rect 5218 1478 5980 1714
rect 0 1436 5980 1478
rect 0 1014 5980 1056
rect 0 778 82 1014
rect 318 778 1482 1014
rect 1718 778 2882 1014
rect 3118 778 4282 1014
rect 4518 778 5980 1014
rect 0 736 5980 778
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 276 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 276 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 0 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 0 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 1196 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1635271187
transform 1 0 1380 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[1\]
timestamp 1635271187
transform 1 0 1196 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[2\]
timestamp 1635271187
transform -1 0 1748 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[3\]
timestamp 1635271187
transform -1 0 2024 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[4\]
timestamp 1635271187
transform -1 0 2300 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[5\]
timestamp 1635271187
transform 1 0 2300 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1635271187
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3036 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1635271187
transform 1 0 3496 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1635271187
transform 1 0 2484 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[6\]
timestamp 1635271187
transform 1 0 2760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[7\]
timestamp 1635271187
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1635271187
transform 1 0 3956 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48
timestamp 1635271187
transform 1 0 4416 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1635271187
transform 1 0 3588 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4692 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[12\]
timestamp 1635271187
transform 1 0 4508 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[8\]
timestamp 1635271187
transform 1 0 3680 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[9\]
timestamp 1635271187
transform 1 0 4140 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[10\]
timestamp 1635271187
transform 1 0 4784 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1635271187
transform 1 0 5152 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_7
timestamp 1635271187
transform 1 0 5152 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1635271187
transform 1 0 5060 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1635271187
transform 1 0 5060 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[11\]
timestamp 1635271187
transform -1 0 5520 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1635271187
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1635271187
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1635271187
transform 1 0 5520 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 5980 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 5980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1635271187
transform 1 0 276 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635271187
transform 1 0 0 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1635271187
transform 1 0 1380 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635271187
transform 1 0 2484 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635271187
transform 1 0 2668 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1635271187
transform 1 0 2576 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635271187
transform 1 0 3772 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp 1635271187
transform 1 0 4876 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1635271187
transform 1 0 5244 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1635271187
transform 1 0 5612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 5980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1635271187
transform 1 0 5152 0 1 1632
box -38 -48 130 592
<< labels >>
rlabel metal5 s 0 1436 5980 1756 6 VGND
port 0 nsew ground input
rlabel metal4 s 760 496 1040 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 2160 496 2440 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 3560 496 3840 2224 6 VGND
port 0 nsew ground input
rlabel metal4 s 4960 496 5240 2224 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 736 5980 1056 6 VPWR
port 1 nsew power input
rlabel metal4 s 60 496 340 2224 6 VPWR
port 1 nsew power input
rlabel metal4 s 1460 496 1740 2224 6 VPWR
port 1 nsew power input
rlabel metal4 s 2860 496 3140 2224 6 VPWR
port 1 nsew power input
rlabel metal4 s 4260 496 4540 2224 6 VPWR
port 1 nsew power input
rlabel metal2 s 202 0 258 400 6 gpio_defaults[0]
port 2 nsew signal tristate
rlabel metal2 s 4802 0 4858 400 6 gpio_defaults[10]
port 3 nsew signal tristate
rlabel metal2 s 5262 0 5318 400 6 gpio_defaults[11]
port 4 nsew signal tristate
rlabel metal2 s 5722 0 5778 400 6 gpio_defaults[12]
port 5 nsew signal tristate
rlabel metal2 s 662 0 718 400 6 gpio_defaults[1]
port 6 nsew signal tristate
rlabel metal2 s 1122 0 1178 400 6 gpio_defaults[2]
port 7 nsew signal tristate
rlabel metal2 s 1582 0 1638 400 6 gpio_defaults[3]
port 8 nsew signal tristate
rlabel metal2 s 2042 0 2098 400 6 gpio_defaults[4]
port 9 nsew signal tristate
rlabel metal2 s 2502 0 2558 400 6 gpio_defaults[5]
port 10 nsew signal tristate
rlabel metal2 s 2962 0 3018 400 6 gpio_defaults[6]
port 11 nsew signal tristate
rlabel metal2 s 3422 0 3478 400 6 gpio_defaults[7]
port 12 nsew signal tristate
rlabel metal2 s 3882 0 3938 400 6 gpio_defaults[8]
port 13 nsew signal tristate
rlabel metal2 s 4342 0 4398 400 6 gpio_defaults[9]
port 14 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 6000 2200
<< end >>
