magic
tech sky130A
magscale 1 2
timestamp 1675162490
<< obsli1 >>
rect 460 1071 3220 4369
<< obsm1 >>
rect 460 1040 3220 4400
<< metal2 >>
rect 754 5000 810 6200
rect 1122 5000 1178 6200
rect 800 1040 1080 4400
rect 2680 1040 2960 4400
rect 754 -600 810 600
rect 1122 -600 1178 600
<< obsm2 >>
rect 572 4944 698 5114
rect 866 4944 1066 5114
rect 1234 4944 1452 5114
rect 572 4456 1452 4944
rect 572 984 744 4456
rect 1136 984 1452 4456
rect 572 656 1452 984
rect 572 462 698 656
rect 866 462 1066 656
rect 1234 462 1452 656
<< metal3 >>
rect -600 4224 600 4344
rect -600 3952 600 4072
rect -600 3680 600 3800
rect 412 3268 3268 3548
rect -600 2864 600 2984
rect -600 2592 600 2712
rect -600 2320 600 2440
rect 412 1788 3268 2068
rect -600 1504 600 1624
rect -600 1232 600 1352
rect -600 960 600 1080
<< obsm3 >>
rect 680 3628 1367 4317
rect 600 3064 1367 3188
rect 680 2240 1367 3064
rect 600 2148 1367 2240
rect 600 1704 1367 1708
rect 680 990 1367 1704
<< labels >>
rlabel metal2 s 2680 1040 2960 4400 6 VGND
port 1 nsew ground bidirectional
rlabel metal3 s 412 3268 3268 3548 6 VGND
port 1 nsew ground bidirectional
rlabel metal2 s 800 1040 1080 4400 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 412 1788 3268 2068 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 754 5000 810 6200 6 gpio_defaults[0]
port 3 nsew signal output
rlabel metal3 s -600 4224 600 4344 4 gpio_defaults[10]
port 4 nsew signal output
rlabel metal2 s 754 -600 810 600 8 gpio_defaults[11]
port 5 nsew signal output
rlabel metal2 s 1122 -600 1178 600 8 gpio_defaults[12]
port 6 nsew signal output
rlabel metal2 s 1122 5000 1178 6200 6 gpio_defaults[1]
port 7 nsew signal output
rlabel metal3 s -600 960 600 1080 4 gpio_defaults[2]
port 8 nsew signal output
rlabel metal3 s -600 1232 600 1352 4 gpio_defaults[3]
port 9 nsew signal output
rlabel metal3 s -600 1504 600 1624 4 gpio_defaults[4]
port 10 nsew signal output
rlabel metal3 s -600 2320 600 2440 4 gpio_defaults[5]
port 11 nsew signal output
rlabel metal3 s -600 2592 600 2712 4 gpio_defaults[6]
port 12 nsew signal output
rlabel metal3 s -600 2864 600 2984 4 gpio_defaults[7]
port 13 nsew signal output
rlabel metal3 s -600 3680 600 3800 4 gpio_defaults[8]
port 14 nsew signal output
rlabel metal3 s -600 3952 600 4072 4 gpio_defaults[9]
port 15 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3400 5600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44334
string GDS_FILE /home/hosni/caravel_sky130/caravel/openlane/gpio_defaults_block/runs/23_01_31_02_54/results/signoff/gpio_defaults_block.magic.gds
string GDS_START 19988
<< end >>

