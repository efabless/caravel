module empty_macro_1 ();
endmodule
